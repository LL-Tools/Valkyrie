

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810;

  NAND2_X2 U5011 ( .A1(n7936), .A2(n7935), .ZN(n9797) );
  INV_X1 U5012 ( .A(n7601), .ZN(n7605) );
  INV_X4 U5013 ( .A(n8500), .ZN(n8506) );
  AND2_X1 U5014 ( .A1(n6600), .A2(n6599), .ZN(n8054) );
  CLKBUF_X1 U5015 ( .A(n5771), .Z(n6089) );
  OR2_X1 U5016 ( .A1(n7290), .A2(n10687), .ZN(n7465) );
  OR2_X1 U5017 ( .A1(n7572), .A2(n5146), .ZN(n5143) );
  NAND2_X1 U5018 ( .A1(n8512), .A2(n8515), .ZN(n7098) );
  INV_X2 U5019 ( .A(n9376), .ZN(n4948) );
  INV_X1 U5020 ( .A(n7394), .ZN(n8043) );
  INV_X1 U5021 ( .A(n8693), .ZN(n8890) );
  INV_X2 U5022 ( .A(n5861), .ZN(n8307) );
  INV_X1 U5023 ( .A(n9370), .ZN(n9307) );
  INV_X1 U5024 ( .A(n9376), .ZN(n9309) );
  CLKBUF_X2 U5026 ( .A(n5558), .Z(n8071) );
  INV_X1 U5027 ( .A(n8079), .ZN(n10578) );
  XNOR2_X1 U5028 ( .A(n6252), .B(n6997), .ZN(n6990) );
  INV_X1 U5029 ( .A(n6264), .ZN(n8516) );
  INV_X1 U5030 ( .A(n6941), .ZN(n6983) );
  XNOR2_X1 U5031 ( .A(n6017), .B(n6018), .ZN(n8044) );
  CLKBUF_X3 U5032 ( .A(n7890), .Z(n5056) );
  AND2_X1 U5033 ( .A1(n5336), .A2(n5686), .ZN(n4947) );
  XNOR2_X2 U5034 ( .A(n5689), .B(n5688), .ZN(n6363) );
  INV_X1 U5035 ( .A(n5700), .ZN(n9149) );
  NAND2_X2 U5036 ( .A1(n5413), .A2(n5592), .ZN(n5872) );
  AND2_X2 U5037 ( .A1(n5401), .A2(n5400), .ZN(n6252) );
  OAI21_X2 U5038 ( .B1(n7469), .B2(n5170), .A(n6155), .ZN(n7336) );
  NOR2_X2 U5039 ( .A1(n7157), .A2(n6280), .ZN(n6281) );
  AOI211_X2 U5040 ( .C1(n8415), .C2(n8409), .A(n8408), .B(n8407), .ZN(n8410)
         );
  OAI21_X2 U5041 ( .B1(n5925), .B2(n5613), .A(n5612), .ZN(n5941) );
  OAI22_X2 U5042 ( .A1(n8543), .A2(n8695), .B1(n7866), .B2(n7865), .ZN(n8602)
         );
  XNOR2_X2 U5043 ( .A(n7865), .B(n7866), .ZN(n8543) );
  NOR2_X2 U5044 ( .A1(n6253), .A2(n6989), .ZN(n7156) );
  AOI22_X2 U5045 ( .A1(n8602), .A2(n8603), .B1(n8901), .B2(n7867), .ZN(n8577)
         );
  OR2_X1 U5046 ( .A1(n9227), .A2(n5376), .ZN(n5375) );
  INV_X1 U5047 ( .A(n8692), .ZN(n8880) );
  NAND2_X1 U5048 ( .A1(n8092), .A2(n8030), .ZN(n7077) );
  INV_X1 U5049 ( .A(n8958), .ZN(n8989) );
  AND2_X1 U5050 ( .A1(n8302), .A2(n10130), .ZN(n7206) );
  CLKBUF_X2 U5051 ( .A(n6102), .Z(n6119) );
  CLKBUF_X2 U5052 ( .A(n5772), .Z(n6102) );
  NAND2_X1 U5053 ( .A1(n7392), .A2(n5057), .ZN(n7394) );
  CLKBUF_X2 U5054 ( .A(n5873), .Z(n6113) );
  INV_X2 U5055 ( .A(n9674), .ZN(n9671) );
  AOI21_X1 U5056 ( .B1(n6480), .B2(P1_IR_REG_28__SCAN_IN), .A(n5296), .ZN(
        n5295) );
  NOR2_X2 U5057 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6419) );
  NOR2_X1 U5058 ( .A1(n9747), .A2(n9746), .ZN(n9748) );
  NAND2_X1 U5059 ( .A1(n8609), .A2(n7859), .ZN(n8560) );
  OR2_X1 U5060 ( .A1(n9829), .A2(n10015), .ZN(n9810) );
  AND2_X1 U5061 ( .A1(n9773), .A2(n8172), .ZN(n9791) );
  NAND2_X1 U5062 ( .A1(n7955), .A2(n7954), .ZN(n9831) );
  NAND2_X1 U5063 ( .A1(n5410), .A2(n5409), .ZN(n5408) );
  NAND2_X1 U5064 ( .A1(n7827), .A2(n8646), .ZN(n8651) );
  OR2_X1 U5065 ( .A1(n8732), .A2(n6287), .ZN(n5240) );
  AND2_X1 U5066 ( .A1(n5042), .A2(n8647), .ZN(n7768) );
  OAI211_X1 U5067 ( .C1(n8434), .C2(n8433), .A(n8432), .B(n8431), .ZN(n8435)
         );
  MUX2_X1 U5068 ( .A(n8428), .B(n8427), .S(n8506), .Z(n8434) );
  OR2_X1 U5069 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  NAND2_X1 U5070 ( .A1(n5896), .A2(n5895), .ZN(n10724) );
  NAND2_X1 U5071 ( .A1(n5875), .A2(n5438), .ZN(n10705) );
  NAND2_X1 U5072 ( .A1(n6983), .A2(n8079), .ZN(n8232) );
  OAI21_X1 U5073 ( .B1(n8379), .B2(n8378), .A(n8377), .ZN(n8390) );
  XNOR2_X1 U5074 ( .A(n5857), .B(n5856), .ZN(n7346) );
  NAND4_X1 U5075 ( .A1(n7049), .A2(n7048), .A3(n7047), .A4(n7046), .ZN(n9560)
         );
  NAND4_X1 U5076 ( .A1(n6604), .A2(n6603), .A3(n6602), .A4(n6601), .ZN(n6799)
         );
  CLKBUF_X3 U5077 ( .A(n7206), .Z(n8072) );
  NOR2_X2 U5078 ( .A1(n6779), .A2(n8506), .ZN(n6190) );
  NAND3_X1 U5079 ( .A1(n5150), .A2(n5149), .A3(n5016), .ZN(n6250) );
  INV_X1 U5080 ( .A(n6599), .ZN(n10130) );
  NAND2_X1 U5081 ( .A1(n8365), .A2(n8367), .ZN(n6138) );
  OR2_X1 U5082 ( .A1(n10486), .A2(n5816), .ZN(n6277) );
  NAND4_X2 U5083 ( .A1(n5802), .A2(n5801), .A3(n5800), .A4(n5799), .ZN(n10636)
         );
  NAND4_X2 U5084 ( .A1(n5790), .A2(n5789), .A3(n5788), .A4(n5787), .ZN(n10592)
         );
  OR2_X1 U5085 ( .A1(n8709), .A2(n6773), .ZN(n8363) );
  AND2_X1 U5086 ( .A1(n6598), .A2(n5554), .ZN(n6599) );
  OR2_X2 U5087 ( .A1(n10454), .A2(n6315), .ZN(n5151) );
  AND2_X2 U5088 ( .A1(n5487), .A2(n8520), .ZN(n8500) );
  MUX2_X1 U5089 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6597), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n6598) );
  INV_X1 U5090 ( .A(n8362), .ZN(n5487) );
  INV_X1 U5091 ( .A(n7138), .ZN(n10571) );
  NAND4_X2 U5092 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n8708)
         );
  CLKBUF_X3 U5093 ( .A(n5786), .Z(n8314) );
  NAND3_X1 U5094 ( .A1(n6453), .A2(n6403), .A3(n6402), .ZN(n6969) );
  NAND2_X1 U5095 ( .A1(n8231), .A2(n7546), .ZN(n10556) );
  NAND2_X2 U5096 ( .A1(n5295), .A2(n5294), .ZN(n7392) );
  INV_X4 U5097 ( .A(n8310), .ZN(n5828) );
  OR2_X1 U5098 ( .A1(n10449), .A2(n6316), .ZN(n5230) );
  NAND2_X1 U5099 ( .A1(n6240), .A2(n5056), .ZN(n5858) );
  INV_X2 U5100 ( .A(n6240), .ZN(n6036) );
  NAND2_X1 U5101 ( .A1(n5113), .A2(n5110), .ZN(n5294) );
  NAND2_X2 U5102 ( .A1(n6363), .A2(n6358), .ZN(n6240) );
  INV_X1 U5103 ( .A(n5701), .ZN(n9154) );
  NAND2_X1 U5104 ( .A1(n6135), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U5105 ( .A1(n9146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5697) );
  NAND2_X2 U5106 ( .A1(n5057), .A2(P1_U3086), .ZN(n10138) );
  BUF_X4 U5107 ( .A(n5617), .Z(n5057) );
  AND2_X1 U5108 ( .A1(n5020), .A2(n6391), .ZN(n5541) );
  NOR2_X1 U5109 ( .A1(n5844), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5862) );
  NOR2_X2 U5110 ( .A1(n5782), .A2(n5888), .ZN(n10433) );
  NAND2_X1 U5111 ( .A1(n5759), .A2(n5760), .ZN(n6675) );
  AND2_X1 U5112 ( .A1(n5780), .A2(n5781), .ZN(n5888) );
  CLKBUF_X1 U5113 ( .A(n5780), .Z(n6268) );
  AND3_X1 U5114 ( .A1(n5094), .A2(n6181), .A3(n5093), .ZN(n5685) );
  AND2_X1 U5115 ( .A1(n5683), .A2(n5682), .ZN(n6020) );
  AND4_X1 U5116 ( .A1(n5886), .A2(n5885), .A3(n5678), .A4(n5677), .ZN(n4952)
         );
  NAND2_X1 U5117 ( .A1(n6381), .A2(n5526), .ZN(n5525) );
  NOR2_X1 U5118 ( .A1(n10124), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5110) );
  INV_X4 U5119 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U5120 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6384) );
  NOR2_X1 U5121 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6385) );
  NOR2_X1 U5122 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6386) );
  NOR2_X1 U5123 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5683) );
  NOR2_X1 U5124 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5682) );
  INV_X4 U5125 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5126 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5696) );
  NAND4_X2 U5127 ( .A1(n5709), .A2(n5708), .A3(n5707), .A4(n5706), .ZN(n8843)
         );
  NOR2_X2 U5128 ( .A1(n5977), .A2(n8760), .ZN(n8759) );
  OAI211_X2 U5129 ( .C1(n5861), .C2(n6435), .A(n5860), .B(n5859), .ZN(n10687)
         );
  NOR4_X2 U5130 ( .A1(n8840), .A2(n8351), .A3(n8350), .A4(n8349), .ZN(n8352)
         );
  OAI21_X2 U5131 ( .B1(n9846), .B2(n5299), .A(n5297), .ZN(n9792) );
  AND2_X1 U5132 ( .A1(n9796), .A2(n5122), .ZN(n9731) );
  NOR2_X2 U5133 ( .A1(n9810), .A2(n9797), .ZN(n9796) );
  AOI21_X2 U5134 ( .B1(n9925), .B2(n5306), .A(n5303), .ZN(n9891) );
  AND2_X1 U5135 ( .A1(n5646), .A2(n5645), .ZN(n6048) );
  NAND2_X1 U5136 ( .A1(n6766), .A2(n6767), .ZN(n6769) );
  INV_X1 U5137 ( .A(n5520), .ZN(n5518) );
  OR2_X1 U5138 ( .A1(n8795), .A2(n9083), .ZN(n5128) );
  NAND2_X1 U5139 ( .A1(n5187), .A2(n8135), .ZN(n8140) );
  NAND2_X1 U5140 ( .A1(n8124), .A2(n8123), .ZN(n5189) );
  INV_X1 U5141 ( .A(n8458), .ZN(n5224) );
  MUX2_X1 U5142 ( .A(n8454), .B(n8453), .S(n8506), .Z(n8458) );
  AOI21_X1 U5143 ( .B1(n5180), .B2(n9700), .A(n5179), .ZN(n5178) );
  NOR2_X1 U5144 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5885) );
  NOR2_X1 U5145 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5886) );
  INV_X1 U5146 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6391) );
  INV_X1 U5147 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6381) );
  OAI21_X1 U5148 ( .B1(n8495), .B2(n8494), .A(n8493), .ZN(n8496) );
  NAND2_X1 U5149 ( .A1(n8495), .A2(n8494), .ZN(n5052) );
  INV_X1 U5150 ( .A(n8325), .ZN(n5492) );
  OAI21_X1 U5151 ( .B1(n8850), .B2(n8840), .A(n8323), .ZN(n8325) );
  OR2_X1 U5152 ( .A1(n6675), .A2(n6269), .ZN(n5228) );
  OR2_X1 U5153 ( .A1(n6234), .A2(n5746), .ZN(n8499) );
  OR2_X1 U5154 ( .A1(n8839), .A2(n8854), .ZN(n6126) );
  OAI21_X1 U5155 ( .B1(n5423), .B2(n5419), .A(n4994), .ZN(n5418) );
  INV_X1 U5156 ( .A(n5555), .ZN(n5419) );
  NAND2_X1 U5157 ( .A1(n8882), .A2(n8486), .ZN(n5483) );
  AND2_X1 U5158 ( .A1(n5470), .A2(n5098), .ZN(n5097) );
  NAND2_X1 U5159 ( .A1(n8456), .A2(n5099), .ZN(n5098) );
  INV_X1 U5160 ( .A(n6015), .ZN(n5099) );
  OR2_X1 U5161 ( .A1(n9010), .A2(n8988), .ZN(n8448) );
  AND2_X1 U5162 ( .A1(n5431), .A2(n6162), .ZN(n5430) );
  OR2_X1 U5163 ( .A1(n5432), .A2(n7589), .ZN(n5431) );
  NAND2_X1 U5164 ( .A1(n7590), .A2(n7588), .ZN(n6160) );
  AND2_X1 U5165 ( .A1(n5354), .A2(n6444), .ZN(n6767) );
  AND2_X1 U5166 ( .A1(n6211), .A2(n5356), .ZN(n5355) );
  NAND2_X1 U5167 ( .A1(n5160), .A2(n4947), .ZN(n6203) );
  AND4_X1 U5168 ( .A1(n5162), .A2(n5161), .A3(n4952), .A4(n4983), .ZN(n5160)
         );
  OR2_X1 U5169 ( .A1(n5888), .A2(n5807), .ZN(n5806) );
  INV_X1 U5170 ( .A(n9536), .ZN(n5380) );
  INV_X1 U5171 ( .A(n9537), .ZN(n5379) );
  OR2_X1 U5172 ( .A1(n9991), .A2(n10369), .ZN(n8213) );
  AND2_X1 U5173 ( .A1(n5004), .A2(n5505), .ZN(n5503) );
  AND2_X1 U5174 ( .A1(n9721), .A2(n4974), .ZN(n5508) );
  OR2_X1 U5175 ( .A1(n9765), .A2(n9780), .ZN(n9745) );
  OAI21_X1 U5176 ( .B1(n7884), .B2(n10266), .A(n7883), .ZN(n8067) );
  XNOR2_X1 U5177 ( .A(n7882), .B(n7881), .ZN(n7884) );
  NAND2_X1 U5178 ( .A1(n5723), .A2(n5722), .ZN(n5734) );
  INV_X1 U5179 ( .A(n6437), .ZN(n6390) );
  NAND2_X1 U5180 ( .A1(n6390), .A2(n5328), .ZN(n6606) );
  AND2_X1 U5181 ( .A1(n5541), .A2(n6389), .ZN(n5328) );
  OAI21_X1 U5182 ( .B1(n6072), .B2(n5277), .A(n5275), .ZN(n6097) );
  AOI21_X1 U5183 ( .B1(n6071), .B2(n5278), .A(n5276), .ZN(n5275) );
  INV_X1 U5184 ( .A(n5278), .ZN(n5277) );
  INV_X1 U5185 ( .A(n5659), .ZN(n5276) );
  AND2_X1 U5186 ( .A1(n5663), .A2(n5662), .ZN(n6096) );
  NAND2_X1 U5187 ( .A1(n5959), .A2(n5958), .ZN(n8357) );
  NAND2_X1 U5188 ( .A1(n5364), .A2(n4980), .ZN(n7454) );
  INV_X1 U5189 ( .A(n5567), .ZN(n5363) );
  NAND2_X1 U5190 ( .A1(n8635), .A2(n7864), .ZN(n7865) );
  OR2_X1 U5191 ( .A1(n6771), .A2(n10591), .ZN(n6775) );
  NAND2_X1 U5192 ( .A1(n9149), .A2(n9154), .ZN(n5786) );
  OAI21_X1 U5193 ( .B1(n7376), .B2(n5444), .A(n5443), .ZN(n7673) );
  NAND2_X1 U5194 ( .A1(n5447), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5444) );
  INV_X1 U5195 ( .A(n7674), .ZN(n5447) );
  NAND2_X1 U5196 ( .A1(n5049), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U5197 ( .A1(n5238), .A2(n5237), .ZN(n5442) );
  INV_X1 U5198 ( .A(n8711), .ZN(n5237) );
  NOR2_X1 U5199 ( .A1(n8733), .A2(n5950), .ZN(n8732) );
  NAND2_X1 U5200 ( .A1(n5129), .A2(n5130), .ZN(n5410) );
  INV_X1 U5201 ( .A(n5131), .ZN(n5130) );
  OAI21_X1 U5202 ( .B1(n6258), .B2(P2_REG1_REG_13__SCAN_IN), .A(n5134), .ZN(
        n5131) );
  NAND2_X1 U5203 ( .A1(n5240), .A2(n5239), .ZN(n5440) );
  INV_X1 U5204 ( .A(n8743), .ZN(n5239) );
  INV_X1 U5205 ( .A(n6190), .ZN(n9005) );
  NAND2_X1 U5206 ( .A1(n9991), .A2(n10369), .ZN(n8281) );
  NOR2_X1 U5207 ( .A1(n6388), .A2(n6437), .ZN(n6392) );
  AND2_X1 U5208 ( .A1(n5551), .A2(n9727), .ZN(n5546) );
  NOR2_X1 U5209 ( .A1(n9754), .A2(n5549), .ZN(n5548) );
  INV_X1 U5210 ( .A(n9725), .ZN(n5549) );
  NAND2_X1 U5211 ( .A1(n5515), .A2(n5517), .ZN(n5514) );
  INV_X1 U5212 ( .A(n5521), .ZN(n5515) );
  INV_X1 U5213 ( .A(n7392), .ZN(n8045) );
  INV_X1 U5214 ( .A(n6943), .ZN(n8046) );
  NAND2_X1 U5215 ( .A1(n7897), .A2(n7896), .ZN(n9682) );
  INV_X1 U5216 ( .A(n6468), .ZN(n6640) );
  INV_X1 U5217 ( .A(n5113), .ZN(n6476) );
  INV_X1 U5218 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U5219 ( .A1(n5250), .A2(n5255), .ZN(n6049) );
  NAND2_X1 U5220 ( .A1(n6017), .A2(n5257), .ZN(n5250) );
  INV_X2 U5221 ( .A(P2_U3893), .ZN(n8812) );
  OR2_X1 U5222 ( .A1(n8728), .A2(n5946), .ZN(n5133) );
  XOR2_X1 U5223 ( .A(n5050), .B(n6257), .Z(n8728) );
  AND2_X1 U5224 ( .A1(n4973), .A2(n5128), .ZN(n8808) );
  INV_X1 U5225 ( .A(n5396), .ZN(n6262) );
  NAND2_X1 U5226 ( .A1(n8105), .A2(n8250), .ZN(n8120) );
  MUX2_X1 U5227 ( .A(n8095), .B(n8094), .S(n8181), .Z(n8103) );
  INV_X1 U5228 ( .A(n8120), .ZN(n8116) );
  AND2_X1 U5229 ( .A1(n8264), .A2(n8174), .ZN(n5191) );
  NAND2_X1 U5230 ( .A1(n8147), .A2(n8148), .ZN(n5195) );
  OR3_X1 U5231 ( .A1(n8146), .A2(n8174), .A3(n8256), .ZN(n8147) );
  NOR2_X1 U5232 ( .A1(n8174), .A2(n5194), .ZN(n5193) );
  INV_X1 U5233 ( .A(n8259), .ZN(n5194) );
  NAND2_X1 U5234 ( .A1(n5224), .A2(n5221), .ZN(n5220) );
  NAND2_X1 U5235 ( .A1(n8450), .A2(n5222), .ZN(n5221) );
  INV_X1 U5236 ( .A(n8455), .ZN(n5222) );
  AOI21_X1 U5237 ( .B1(n5223), .B2(n5219), .A(n5218), .ZN(n5217) );
  INV_X1 U5238 ( .A(n8450), .ZN(n5219) );
  INV_X1 U5239 ( .A(n8457), .ZN(n5218) );
  OR2_X1 U5240 ( .A1(n5216), .A2(n8451), .ZN(n5213) );
  OAI21_X1 U5241 ( .B1(n8154), .B2(n8193), .A(n5204), .ZN(n5203) );
  AND2_X1 U5242 ( .A1(n9889), .A2(n8262), .ZN(n5204) );
  NAND2_X1 U5243 ( .A1(n9855), .A2(n5198), .ZN(n5197) );
  NAND2_X1 U5244 ( .A1(n5199), .A2(n8174), .ZN(n5198) );
  NOR2_X1 U5245 ( .A1(n5202), .A2(n5201), .ZN(n5200) );
  NAND2_X1 U5246 ( .A1(n8267), .A2(n8174), .ZN(n5201) );
  AND2_X1 U5247 ( .A1(n5182), .A2(n5181), .ZN(n5180) );
  NAND2_X1 U5248 ( .A1(n9773), .A2(n4970), .ZN(n5181) );
  INV_X1 U5249 ( .A(n8171), .ZN(n5182) );
  AND2_X1 U5250 ( .A1(n8484), .A2(n8483), .ZN(n5208) );
  AOI21_X1 U5251 ( .B1(n5174), .B2(n5177), .A(n4975), .ZN(n5173) );
  INV_X1 U5252 ( .A(SI_11_), .ZN(n10185) );
  NOR2_X1 U5253 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5887) );
  NAND2_X1 U5254 ( .A1(n5119), .A2(n10106), .ZN(n5118) );
  NOR2_X1 U5255 ( .A1(n9932), .A2(n9952), .ZN(n5119) );
  AOI21_X1 U5256 ( .B1(n5255), .B2(n5253), .A(n5252), .ZN(n5251) );
  INV_X1 U5257 ( .A(n6048), .ZN(n5252) );
  INV_X1 U5258 ( .A(n5257), .ZN(n5253) );
  INV_X1 U5259 ( .A(n5255), .ZN(n5254) );
  INV_X1 U5260 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6383) );
  INV_X1 U5261 ( .A(n5910), .ZN(n5263) );
  INV_X1 U5262 ( .A(n5601), .ZN(n5267) );
  INV_X1 U5263 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5526) );
  AOI21_X1 U5264 ( .B1(n5352), .B2(n5350), .A(n4996), .ZN(n5349) );
  INV_X1 U5265 ( .A(n8668), .ZN(n5350) );
  NAND2_X1 U5266 ( .A1(n9094), .A2(n8828), .ZN(n5491) );
  NOR2_X1 U5267 ( .A1(n5226), .A2(n5751), .ZN(n5225) );
  INV_X1 U5268 ( .A(n6270), .ZN(n5226) );
  NAND2_X1 U5269 ( .A1(n10435), .A2(n6246), .ZN(n6247) );
  NAND2_X1 U5270 ( .A1(n10521), .A2(n5448), .ZN(n5231) );
  NAND2_X1 U5271 ( .A1(n10512), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U5272 ( .A1(n5422), .A2(n5555), .ZN(n5421) );
  INV_X1 U5273 ( .A(n5424), .ZN(n5422) );
  NOR2_X1 U5274 ( .A1(n5484), .A2(n5482), .ZN(n5481) );
  INV_X1 U5275 ( .A(n8485), .ZN(n5482) );
  INV_X1 U5276 ( .A(n5025), .ZN(n5484) );
  NAND2_X1 U5277 ( .A1(n5003), .A2(n4956), .ZN(n5423) );
  NAND2_X1 U5278 ( .A1(n6126), .A2(n6125), .ZN(n8840) );
  NAND2_X1 U5279 ( .A1(n5459), .A2(n6108), .ZN(n5458) );
  NAND2_X1 U5280 ( .A1(n5460), .A2(n5462), .ZN(n5459) );
  INV_X1 U5281 ( .A(n6172), .ZN(n5165) );
  OR2_X1 U5282 ( .A1(n8655), .A2(n8989), .ZN(n8964) );
  INV_X1 U5283 ( .A(n5108), .ZN(n5107) );
  NOR2_X1 U5284 ( .A1(n5109), .A2(n8341), .ZN(n5108) );
  INV_X1 U5285 ( .A(n5969), .ZN(n5109) );
  NOR2_X1 U5286 ( .A1(n8438), .A2(n5479), .ZN(n5478) );
  INV_X1 U5287 ( .A(n5955), .ZN(n5479) );
  AND2_X1 U5288 ( .A1(n6240), .A2(n5057), .ZN(n5779) );
  NAND2_X1 U5289 ( .A1(n5495), .A2(n6207), .ZN(n5493) );
  AND3_X1 U5290 ( .A1(n5780), .A2(n5887), .A3(n5679), .ZN(n5336) );
  INV_X1 U5291 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5679) );
  NOR2_X1 U5292 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5677) );
  AND2_X1 U5293 ( .A1(n5336), .A2(n4952), .ZN(n5681) );
  INV_X1 U5294 ( .A(n9447), .ZN(n5387) );
  INV_X1 U5295 ( .A(n5391), .ZN(n5386) );
  NOR2_X1 U5296 ( .A1(n9447), .A2(n9343), .ZN(n5388) );
  NOR2_X1 U5297 ( .A1(n5070), .A2(n5067), .ZN(n5066) );
  INV_X1 U5298 ( .A(n9364), .ZN(n5067) );
  INV_X1 U5299 ( .A(n5368), .ZN(n5070) );
  NOR2_X1 U5300 ( .A1(n5372), .A2(n5369), .ZN(n5368) );
  INV_X1 U5301 ( .A(n9403), .ZN(n5372) );
  INV_X1 U5302 ( .A(n9469), .ZN(n5369) );
  NAND2_X1 U5303 ( .A1(n9403), .A2(n5371), .ZN(n5370) );
  NOR2_X1 U5304 ( .A1(n8183), .A2(n8231), .ZN(n5271) );
  OAI21_X1 U5305 ( .B1(n5184), .B2(n5183), .A(n4995), .ZN(n8180) );
  NOR2_X1 U5306 ( .A1(n10005), .A2(n9765), .ZN(n5126) );
  INV_X1 U5307 ( .A(n9696), .ZN(n5300) );
  OR2_X1 U5308 ( .A1(n10015), .A2(n9794), .ZN(n9699) );
  NOR2_X1 U5309 ( .A1(n9717), .A2(n5517), .ZN(n5513) );
  OR2_X1 U5310 ( .A1(n9932), .A2(n9950), .ZN(n8263) );
  NAND2_X1 U5311 ( .A1(n5310), .A2(n5309), .ZN(n5308) );
  INV_X1 U5312 ( .A(n9925), .ZN(n5310) );
  AOI21_X1 U5313 ( .B1(n5317), .B2(n5319), .A(n5316), .ZN(n5315) );
  INV_X1 U5314 ( .A(n9959), .ZN(n5316) );
  INV_X1 U5315 ( .A(n7721), .ZN(n5317) );
  NOR2_X1 U5316 ( .A1(n8141), .A2(n5320), .ZN(n5319) );
  INV_X1 U5317 ( .A(n8142), .ZN(n5320) );
  OR2_X1 U5318 ( .A1(n10778), .A2(n9509), .ZN(n8139) );
  OR2_X1 U5319 ( .A1(n7323), .A2(n8098), .ZN(n5314) );
  NAND2_X1 U5320 ( .A1(n7272), .A2(n10618), .ZN(n8096) );
  NOR2_X2 U5321 ( .A1(n9896), .A2(n9881), .ZN(n9880) );
  NOR2_X1 U5322 ( .A1(n9968), .A2(n9952), .ZN(n9951) );
  NAND2_X1 U5323 ( .A1(n6473), .A2(n5112), .ZN(n5111) );
  INV_X1 U5324 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6473) );
  INV_X1 U5325 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5112) );
  OAI21_X1 U5326 ( .B1(n5664), .B2(n5032), .A(n5288), .ZN(n5721) );
  INV_X1 U5327 ( .A(n5289), .ZN(n5288) );
  OAI21_X1 U5328 ( .B1(n5292), .B2(n5032), .A(n5672), .ZN(n5289) );
  INV_X1 U5329 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6394) );
  INV_X1 U5330 ( .A(n6393), .ZN(n5542) );
  INV_X1 U5331 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6404) );
  OAI21_X1 U5332 ( .B1(n5971), .B2(n5625), .A(n5624), .ZN(n5986) );
  OAI21_X1 U5333 ( .B1(n5941), .B2(n5283), .A(n5281), .ZN(n5971) );
  AOI21_X1 U5334 ( .B1(n5940), .B2(n5284), .A(n5282), .ZN(n5281) );
  INV_X1 U5335 ( .A(n5284), .ZN(n5283) );
  INV_X1 U5336 ( .A(n5622), .ZN(n5282) );
  NOR2_X1 U5337 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6380) );
  OAI21_X1 U5338 ( .B1(n7890), .B2(n5044), .A(n5043), .ZN(n5571) );
  NAND2_X1 U5339 ( .A1(n7890), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5043) );
  INV_X1 U5340 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5244) );
  INV_X1 U5341 ( .A(n5349), .ZN(n5347) );
  INV_X1 U5342 ( .A(n6888), .ZN(n6889) );
  NOR2_X1 U5343 ( .A1(n7257), .A2(n5366), .ZN(n5365) );
  INV_X1 U5344 ( .A(n7254), .ZN(n5366) );
  NAND2_X1 U5345 ( .A1(n7837), .A2(n8533), .ZN(n8535) );
  OAI21_X1 U5346 ( .B1(n5489), .B2(n5486), .A(n5485), .ZN(n8514) );
  NAND2_X1 U5347 ( .A1(n5488), .A2(n5487), .ZN(n5486) );
  NAND2_X1 U5348 ( .A1(n8355), .A2(n8362), .ZN(n5485) );
  NOR3_X1 U5349 ( .A1(n5492), .A2(n8510), .A3(n5490), .ZN(n5489) );
  NAND2_X1 U5350 ( .A1(n5681), .A2(n5680), .ZN(n6019) );
  INV_X1 U5351 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5680) );
  XNOR2_X1 U5352 ( .A(n10433), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n10437) );
  NAND2_X1 U5353 ( .A1(n10436), .A2(n10437), .ZN(n10435) );
  OR2_X1 U5354 ( .A1(n5151), .A2(n10470), .ZN(n5150) );
  OR2_X1 U5355 ( .A1(n10470), .A2(n5412), .ZN(n5149) );
  NAND2_X1 U5356 ( .A1(n10522), .A2(n10523), .ZN(n10521) );
  NOR2_X1 U5357 ( .A1(n10488), .A2(n6251), .ZN(n10510) );
  OR2_X1 U5358 ( .A1(n10510), .A2(n10509), .ZN(n5401) );
  XNOR2_X1 U5359 ( .A(n5231), .B(n6436), .ZN(n6992) );
  XNOR2_X1 U5360 ( .A(n6281), .B(n7381), .ZN(n7376) );
  NOR2_X1 U5361 ( .A1(n6339), .A2(n7161), .ZN(n7379) );
  NOR2_X1 U5362 ( .A1(n7381), .A2(n6281), .ZN(n6282) );
  OR2_X1 U5363 ( .A1(n7376), .A2(n5879), .ZN(n5446) );
  AOI21_X1 U5364 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6472), .A(n7662), .ZN(
        n6255) );
  AND3_X1 U5365 ( .A1(n5144), .A2(n5143), .A3(n5037), .ZN(n6257) );
  NAND2_X1 U5366 ( .A1(n5397), .A2(n5039), .ZN(n5396) );
  NOR2_X1 U5367 ( .A1(n6128), .A2(n5103), .ZN(n5102) );
  OR2_X1 U5368 ( .A1(n6124), .A2(n5104), .ZN(n5103) );
  INV_X1 U5369 ( .A(n8488), .ZN(n5104) );
  AOI211_X1 U5370 ( .C1(n8320), .C2(n6125), .A(n5749), .B(n5748), .ZN(n8323)
         );
  INV_X1 U5371 ( .A(n8843), .ZN(n8868) );
  INV_X1 U5372 ( .A(n8943), .ZN(n8913) );
  AOI21_X1 U5373 ( .B1(n5470), .B2(n5474), .A(n5469), .ZN(n5468) );
  NAND2_X1 U5374 ( .A1(n5097), .A2(n5100), .ZN(n5095) );
  NOR2_X1 U5375 ( .A1(n4992), .A2(n5416), .ZN(n5415) );
  INV_X1 U5376 ( .A(n6167), .ZN(n5416) );
  NAND2_X1 U5377 ( .A1(n8986), .A2(n8990), .ZN(n6168) );
  AND2_X1 U5378 ( .A1(n8964), .A2(n8456), .ZN(n8978) );
  AND4_X1 U5379 ( .A1(n6000), .A2(n5999), .A3(n5998), .A4(n5997), .ZN(n8988)
         );
  INV_X1 U5380 ( .A(n8696), .ZN(n9004) );
  NAND2_X1 U5381 ( .A1(n7745), .A2(n5108), .ZN(n9007) );
  AOI21_X1 U5382 ( .B1(n5430), .B2(n5429), .A(n5428), .ZN(n5427) );
  NOR2_X1 U5383 ( .A1(n6163), .A2(n6161), .ZN(n5429) );
  NAND2_X1 U5384 ( .A1(n7681), .A2(n8432), .ZN(n5480) );
  NAND2_X1 U5385 ( .A1(n5480), .A2(n5478), .ZN(n7745) );
  NAND2_X1 U5386 ( .A1(n10705), .A2(n5437), .ZN(n8404) );
  NAND2_X1 U5387 ( .A1(n7466), .A2(n8418), .ZN(n5465) );
  NAND2_X1 U5388 ( .A1(n5434), .A2(n5171), .ZN(n5170) );
  NAND2_X1 U5389 ( .A1(n7097), .A2(n7096), .ZN(n9021) );
  NAND2_X1 U5390 ( .A1(n5741), .A2(n5740), .ZN(n6234) );
  NAND2_X1 U5391 ( .A1(n6074), .A2(n6073), .ZN(n8347) );
  INV_X1 U5392 ( .A(n10720), .ZN(n10801) );
  NAND2_X1 U5393 ( .A1(n6210), .A2(n6211), .ZN(n6443) );
  XNOR2_X1 U5394 ( .A(n5699), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5701) );
  OR2_X1 U5395 ( .A1(n5698), .A2(n5807), .ZN(n5699) );
  INV_X1 U5396 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U5397 ( .A1(n5159), .A2(n4947), .ZN(n6205) );
  NAND2_X1 U5398 ( .A1(n5808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5824) );
  INV_X1 U5399 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5823) );
  INV_X1 U5400 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6408) );
  OR2_X1 U5401 ( .A1(n4957), .A2(n5018), .ZN(n5376) );
  NOR2_X1 U5402 ( .A1(n9219), .A2(n5090), .ZN(n5089) );
  INV_X1 U5403 ( .A(n5091), .ZN(n5090) );
  INV_X1 U5404 ( .A(n5376), .ZN(n5086) );
  INV_X1 U5405 ( .A(n6858), .ZN(n5064) );
  NAND3_X1 U5406 ( .A1(n9455), .A2(n9389), .A3(n9176), .ZN(n5395) );
  NAND2_X1 U5407 ( .A1(n5064), .A2(n6856), .ZN(n6977) );
  INV_X1 U5408 ( .A(n5548), .ZN(n5544) );
  AND2_X1 U5409 ( .A1(n5123), .A2(n5124), .ZN(n5122) );
  XNOR2_X1 U5410 ( .A(n9704), .B(n9729), .ZN(n5327) );
  NAND2_X1 U5411 ( .A1(n9775), .A2(n9702), .ZN(n9759) );
  AOI21_X1 U5412 ( .B1(n5508), .B2(n5506), .A(n4987), .ZN(n5505) );
  INV_X1 U5413 ( .A(n5508), .ZN(n5507) );
  OR2_X1 U5414 ( .A1(n9881), .A2(n9893), .ZN(n9718) );
  NOR2_X1 U5415 ( .A1(n9713), .A2(n5522), .ZN(n5521) );
  INV_X1 U5416 ( .A(n5560), .ZN(n5522) );
  OR2_X1 U5417 ( .A1(n9932), .A2(n9911), .ZN(n5520) );
  OR2_X1 U5418 ( .A1(n10114), .A2(n9712), .ZN(n5560) );
  OR2_X1 U5419 ( .A1(n9971), .A2(n9948), .ZN(n9944) );
  AND2_X1 U5420 ( .A1(n9708), .A2(n9965), .ZN(n9709) );
  AOI21_X1 U5421 ( .B1(n5534), .B2(n5539), .A(n4961), .ZN(n5531) );
  INV_X1 U5422 ( .A(n7702), .ZN(n5538) );
  NOR2_X1 U5423 ( .A1(n9510), .A2(n9415), .ZN(n5535) );
  NAND2_X1 U5424 ( .A1(n5313), .A2(n5311), .ZN(n7523) );
  AND2_X1 U5425 ( .A1(n8244), .A2(n5312), .ZN(n5311) );
  OR2_X1 U5426 ( .A1(n10556), .A2(n6836), .ZN(n9915) );
  NOR2_X1 U5427 ( .A1(n5074), .A2(n5073), .ZN(n5072) );
  OR2_X1 U5428 ( .A1(n6605), .A2(n5076), .ZN(n5075) );
  NOR2_X1 U5429 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5073) );
  NAND2_X1 U5430 ( .A1(n7964), .A2(n7963), .ZN(n10024) );
  NAND2_X1 U5431 ( .A1(n7974), .A2(n7973), .ZN(n10030) );
  NAND2_X1 U5432 ( .A1(n8048), .A2(n8047), .ZN(n9917) );
  AND2_X1 U5433 ( .A1(n6817), .A2(n6829), .ZN(n6822) );
  NAND2_X1 U5434 ( .A1(n6452), .A2(n6453), .ZN(n6468) );
  XNOR2_X1 U5435 ( .A(n7894), .B(n7893), .ZN(n9145) );
  OAI21_X1 U5436 ( .B1(n8067), .B2(n8066), .A(n7889), .ZN(n7894) );
  XNOR2_X1 U5437 ( .A(n6595), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U5438 ( .A1(n5554), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6595) );
  INV_X1 U5439 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6593) );
  XNOR2_X1 U5440 ( .A(n6395), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U5441 ( .A1(n4965), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U5442 ( .A1(n5291), .A2(n5668), .ZN(n5710) );
  NAND2_X1 U5443 ( .A1(n5664), .A2(n5292), .ZN(n5291) );
  NAND2_X1 U5444 ( .A1(n6606), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U5445 ( .A1(n5280), .A2(n5278), .ZN(n6086) );
  NAND2_X1 U5446 ( .A1(n5280), .A2(n5653), .ZN(n6084) );
  NAND2_X1 U5447 ( .A1(n5286), .A2(n5616), .ZN(n5957) );
  INV_X1 U5448 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6459) );
  INV_X1 U5449 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6382) );
  XNOR2_X1 U5450 ( .A(n5872), .B(n5871), .ZN(n7395) );
  NAND2_X1 U5451 ( .A1(n5414), .A2(n5589), .ZN(n5857) );
  INV_X1 U5452 ( .A(n8695), .ZN(n8912) );
  NOR2_X1 U5453 ( .A1(n5340), .A2(n8676), .ZN(n5338) );
  NOR2_X1 U5454 ( .A1(n5343), .A2(n5346), .ZN(n5340) );
  NOR2_X1 U5455 ( .A1(n5347), .A2(n7875), .ZN(n5346) );
  NAND2_X1 U5456 ( .A1(n5342), .A2(n5348), .ZN(n5341) );
  NAND2_X1 U5457 ( .A1(n5352), .A2(n7875), .ZN(n5348) );
  INV_X1 U5458 ( .A(n5343), .ZN(n5342) );
  NAND2_X1 U5459 ( .A1(n5725), .A2(n5724), .ZN(n8839) );
  AND2_X1 U5460 ( .A1(n6775), .A2(n6772), .ZN(n6788) );
  NAND2_X1 U5461 ( .A1(n6009), .A2(n6008), .ZN(n8599) );
  NAND2_X1 U5462 ( .A1(n6762), .A2(n10650), .ZN(n8673) );
  MUX2_X1 U5463 ( .A(n6299), .B(n8812), .S(n8517), .Z(n10511) );
  NAND2_X1 U5464 ( .A1(n5140), .A2(n6464), .ZN(n5138) );
  NAND2_X1 U5465 ( .A1(n7156), .A2(n4954), .ZN(n5136) );
  NAND2_X1 U5466 ( .A1(n5054), .A2(n4968), .ZN(n5238) );
  NAND2_X1 U5467 ( .A1(n5144), .A2(n5143), .ZN(n8719) );
  INV_X1 U5468 ( .A(n5442), .ZN(n8710) );
  INV_X1 U5469 ( .A(n5051), .ZN(n6286) );
  INV_X1 U5470 ( .A(n5410), .ZN(n8751) );
  INV_X1 U5471 ( .A(n5440), .ZN(n8742) );
  INV_X1 U5472 ( .A(n5408), .ZN(n6260) );
  NAND2_X1 U5473 ( .A1(n5048), .A2(n5046), .ZN(n5045) );
  NOR3_X1 U5474 ( .A1(n5033), .A2(n8802), .A3(n5047), .ZN(n5046) );
  NAND2_X1 U5475 ( .A1(n8803), .A2(n10519), .ZN(n5048) );
  INV_X1 U5476 ( .A(n8801), .ZN(n5047) );
  XNOR2_X1 U5477 ( .A(n5396), .B(n8799), .ZN(n8795) );
  XNOR2_X1 U5478 ( .A(n5236), .B(n5235), .ZN(n5234) );
  INV_X1 U5479 ( .A(n8816), .ZN(n5235) );
  NOR2_X1 U5480 ( .A1(n8814), .A2(n8815), .ZN(n5236) );
  NAND2_X1 U5481 ( .A1(n5453), .A2(n8553), .ZN(n5452) );
  NAND2_X1 U5482 ( .A1(n10516), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U5483 ( .A1(n5038), .A2(n5404), .ZN(n5403) );
  OR2_X1 U5484 ( .A1(n6364), .A2(n10464), .ZN(n6365) );
  XNOR2_X1 U5485 ( .A(n5455), .B(n6360), .ZN(n5454) );
  NAND2_X1 U5486 ( .A1(n5000), .A2(n5456), .ZN(n5455) );
  OR2_X1 U5487 ( .A1(n6186), .A2(n9000), .ZN(n6199) );
  INV_X1 U5488 ( .A(n5157), .ZN(n5156) );
  OAI22_X1 U5489 ( .A1(n8854), .A2(n9005), .B1(n9003), .B2(n8880), .ZN(n5157)
         );
  NAND2_X1 U5490 ( .A1(n8870), .A2(n8488), .ZN(n8856) );
  NAND2_X1 U5491 ( .A1(n5471), .A2(n5472), .ZN(n8923) );
  INV_X1 U5492 ( .A(n5466), .ZN(n5472) );
  OR2_X1 U5493 ( .A1(n8965), .A2(n5474), .ZN(n5471) );
  NAND2_X1 U5494 ( .A1(n6063), .A2(n6062), .ZN(n9062) );
  NAND2_X1 U5495 ( .A1(n5477), .A2(n5475), .ZN(n8937) );
  AND2_X1 U5496 ( .A1(n5477), .A2(n6045), .ZN(n8935) );
  NAND2_X1 U5497 ( .A1(n6051), .A2(n6050), .ZN(n8950) );
  NAND2_X1 U5498 ( .A1(n8362), .A2(n7545), .ZN(n10799) );
  NOR2_X1 U5499 ( .A1(n7091), .A2(n6377), .ZN(n10748) );
  NOR2_X1 U5500 ( .A1(n8831), .A2(n6200), .ZN(n6378) );
  AND2_X1 U5501 ( .A1(n8833), .A2(n10739), .ZN(n6200) );
  INV_X1 U5502 ( .A(n6211), .ZN(n7825) );
  INV_X1 U5503 ( .A(n9826), .ZN(n9862) );
  INV_X1 U5504 ( .A(n9562), .ZN(n7119) );
  INV_X1 U5505 ( .A(n9964), .ZN(n9712) );
  NAND2_X1 U5506 ( .A1(n5547), .A2(n5546), .ZN(n9737) );
  NOR2_X1 U5507 ( .A1(n8122), .A2(n4971), .ZN(n5188) );
  OAI21_X1 U5508 ( .B1(n8103), .B2(n8102), .A(n8101), .ZN(n8111) );
  NAND2_X1 U5509 ( .A1(n8140), .A2(n5186), .ZN(n8143) );
  AND2_X1 U5510 ( .A1(n8138), .A2(n8139), .ZN(n5186) );
  OR2_X1 U5511 ( .A1(n5224), .A2(n5223), .ZN(n5212) );
  NAND2_X1 U5512 ( .A1(n5192), .A2(n5190), .ZN(n8152) );
  OAI21_X1 U5513 ( .B1(n5195), .B2(n8149), .A(n5193), .ZN(n5192) );
  OAI21_X1 U5514 ( .B1(n5195), .B2(n8151), .A(n5191), .ZN(n5190) );
  AOI21_X1 U5515 ( .B1(n4999), .B2(n8966), .A(n8462), .ZN(n5214) );
  AND2_X1 U5516 ( .A1(n8086), .A2(n8085), .ZN(n8091) );
  OAI21_X1 U5517 ( .B1(n8159), .B2(n8174), .A(n5196), .ZN(n8160) );
  AOI21_X1 U5518 ( .B1(n5203), .B2(n5200), .A(n5197), .ZN(n5196) );
  INV_X1 U5519 ( .A(n5178), .ZN(n5177) );
  INV_X1 U5520 ( .A(n5180), .ZN(n5176) );
  INV_X1 U5521 ( .A(SI_19_), .ZN(n10277) );
  INV_X1 U5522 ( .A(SI_16_), .ZN(n10250) );
  INV_X1 U5523 ( .A(SI_14_), .ZN(n10286) );
  INV_X1 U5524 ( .A(SI_8_), .ZN(n10298) );
  NAND2_X1 U5525 ( .A1(n5361), .A2(n5359), .ZN(n5358) );
  INV_X1 U5526 ( .A(n8533), .ZN(n5359) );
  INV_X1 U5527 ( .A(n8492), .ZN(n5205) );
  INV_X1 U5528 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5494) );
  INV_X1 U5529 ( .A(n9279), .ZN(n5371) );
  AOI21_X1 U5530 ( .B1(n8176), .B2(n4978), .A(n5185), .ZN(n5184) );
  NAND2_X1 U5531 ( .A1(n9729), .A2(n8177), .ZN(n5185) );
  NAND2_X1 U5532 ( .A1(n5739), .A2(n5738), .ZN(n7882) );
  INV_X1 U5533 ( .A(n5668), .ZN(n5290) );
  NAND2_X1 U5534 ( .A1(n6615), .A2(n6616), .ZN(n6393) );
  NOR2_X1 U5535 ( .A1(n5956), .A2(n5285), .ZN(n5284) );
  INV_X1 U5536 ( .A(n5616), .ZN(n5285) );
  INV_X1 U5537 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5618) );
  INV_X1 U5538 ( .A(n5361), .ZN(n5360) );
  NAND2_X1 U5539 ( .A1(n8326), .A2(n8327), .ZN(n5488) );
  OAI21_X1 U5540 ( .B1(n6675), .B2(n6243), .A(n6244), .ZN(n6679) );
  AND2_X1 U5541 ( .A1(n5440), .A2(n5439), .ZN(n6289) );
  NAND2_X1 U5542 ( .A1(n8750), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5439) );
  AOI21_X1 U5543 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8784), .A(n8785), .ZN(
        n6292) );
  AOI21_X1 U5544 ( .B1(n6354), .B2(n6353), .A(n6352), .ZN(n6356) );
  OR2_X1 U5545 ( .A1(n6353), .A2(n6292), .ZN(n6295) );
  NAND2_X1 U5546 ( .A1(n4956), .A2(n5565), .ZN(n5424) );
  INV_X1 U5547 ( .A(n8456), .ZN(n5100) );
  NOR2_X1 U5548 ( .A1(n5466), .A2(n6070), .ZN(n5470) );
  INV_X1 U5549 ( .A(n8468), .ZN(n5469) );
  OR2_X1 U5550 ( .A1(n9062), .A2(n8913), .ZN(n8467) );
  INV_X1 U5551 ( .A(n7468), .ZN(n5171) );
  NAND2_X1 U5552 ( .A1(n7465), .A2(n8405), .ZN(n6151) );
  INV_X1 U5553 ( .A(n6767), .ZN(n7095) );
  AND2_X1 U5554 ( .A1(n8512), .A2(n7176), .ZN(n6373) );
  OR2_X1 U5555 ( .A1(n6443), .A2(n6223), .ZN(n6368) );
  OR2_X1 U5556 ( .A1(n8506), .A2(n6373), .ZN(n6743) );
  NAND2_X1 U5557 ( .A1(n6143), .A2(n6142), .ZN(n7099) );
  OR2_X1 U5558 ( .A1(n5912), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5913) );
  INV_X1 U5559 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5853) );
  INV_X1 U5560 ( .A(n7192), .ZN(n5078) );
  NOR2_X1 U5561 ( .A1(n5382), .A2(n7219), .ZN(n5082) );
  NOR2_X1 U5562 ( .A1(n4991), .A2(n5080), .ZN(n5079) );
  NOR2_X1 U5563 ( .A1(n7202), .A2(n5081), .ZN(n5080) );
  INV_X1 U5564 ( .A(n7219), .ZN(n5081) );
  NAND2_X1 U5565 ( .A1(n7193), .A2(n7192), .ZN(n5083) );
  NAND3_X1 U5566 ( .A1(n8185), .A2(n6807), .A3(n10556), .ZN(n5059) );
  OR2_X1 U5567 ( .A1(n9995), .A2(n9728), .ZN(n8212) );
  NAND2_X1 U5568 ( .A1(n5287), .A2(n9550), .ZN(n8217) );
  INV_X1 U5569 ( .A(n8288), .ZN(n5287) );
  NAND2_X1 U5570 ( .A1(n6392), .A2(n6391), .ZN(n6614) );
  NOR2_X1 U5571 ( .A1(n9995), .A2(n5125), .ZN(n5124) );
  INV_X1 U5572 ( .A(n5126), .ZN(n5125) );
  OR2_X1 U5573 ( .A1(n10030), .A2(n9848), .ZN(n8198) );
  INV_X1 U5574 ( .A(n8263), .ZN(n5307) );
  AND2_X1 U5575 ( .A1(n7491), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7527) );
  NOR2_X1 U5576 ( .A1(n7733), .A2(n10778), .ZN(n7734) );
  OR2_X1 U5577 ( .A1(n7630), .A2(n9197), .ZN(n7733) );
  NAND2_X1 U5578 ( .A1(n4966), .A2(n8098), .ZN(n5312) );
  OR2_X1 U5579 ( .A1(n9188), .A2(n7515), .ZN(n8250) );
  INV_X1 U5580 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7352) );
  OR2_X1 U5581 ( .A1(n7353), .A2(n7352), .ZN(n7404) );
  AOI22_X1 U5582 ( .A1(n5558), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n8054), .ZN(n6736) );
  NAND2_X1 U5583 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n5076) );
  INV_X1 U5584 ( .A(n6606), .ZN(n5074) );
  AND2_X1 U5585 ( .A1(n6613), .A2(n6831), .ZN(n8223) );
  NAND3_X1 U5586 ( .A1(n9759), .A2(n9744), .A3(n9745), .ZN(n9743) );
  OR2_X1 U5587 ( .A1(n9839), .A2(n9831), .ZN(n9829) );
  NAND2_X1 U5588 ( .A1(n5116), .A2(n5120), .ZN(n5115) );
  INV_X1 U5589 ( .A(n5118), .ZN(n5116) );
  NOR2_X1 U5590 ( .A1(n9968), .A2(n5117), .ZN(n9930) );
  INV_X1 U5591 ( .A(n5119), .ZN(n5117) );
  AND2_X1 U5592 ( .A1(n7734), .A2(n9488), .ZN(n7796) );
  XNOR2_X1 U5593 ( .A(n6798), .B(n6938), .ZN(n6800) );
  NAND2_X1 U5594 ( .A1(n5113), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6480) );
  AND2_X1 U5595 ( .A1(n5722), .A2(n5676), .ZN(n5720) );
  NOR2_X1 U5596 ( .A1(n5665), .A2(n5293), .ZN(n5292) );
  INV_X1 U5597 ( .A(n5663), .ZN(n5293) );
  NOR2_X1 U5598 ( .A1(n6083), .A2(n5279), .ZN(n5278) );
  INV_X1 U5599 ( .A(n5653), .ZN(n5279) );
  NAND2_X1 U5600 ( .A1(n5249), .A2(n5247), .ZN(n6061) );
  AOI21_X1 U5601 ( .B1(n5251), .B2(n5254), .A(n5248), .ZN(n5247) );
  INV_X1 U5602 ( .A(n5646), .ZN(n5248) );
  NOR2_X1 U5603 ( .A1(n6032), .A2(n5258), .ZN(n5257) );
  INV_X1 U5604 ( .A(n5637), .ZN(n5258) );
  AOI21_X1 U5605 ( .B1(n5259), .B2(n5257), .A(n5256), .ZN(n5255) );
  INV_X1 U5606 ( .A(n5641), .ZN(n5256) );
  INV_X1 U5607 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6615) );
  INV_X1 U5608 ( .A(n6018), .ZN(n5259) );
  OAI21_X1 U5609 ( .B1(n5986), .B2(n5985), .A(n5629), .ZN(n6005) );
  AND2_X1 U5610 ( .A1(n5633), .A2(n5632), .ZN(n6004) );
  AOI21_X1 U5611 ( .B1(n4950), .B2(n5268), .A(n5262), .ZN(n5261) );
  INV_X1 U5612 ( .A(n5609), .ZN(n5262) );
  AOI21_X1 U5613 ( .B1(n5266), .B2(n5898), .A(n4998), .ZN(n5265) );
  NOR2_X1 U5614 ( .A1(n5561), .A2(n5267), .ZN(n5266) );
  INV_X1 U5615 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6457) );
  AND2_X1 U5616 ( .A1(n5524), .A2(n5523), .ZN(n6433) );
  NOR2_X1 U5617 ( .A1(n5525), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5523) );
  AOI22_X1 U5618 ( .A1(n5349), .A2(n5344), .B1(n5347), .B2(n5345), .ZN(n5343)
         );
  NAND2_X1 U5619 ( .A1(n5351), .A2(n5345), .ZN(n5344) );
  INV_X1 U5620 ( .A(n7875), .ZN(n5345) );
  NAND2_X1 U5621 ( .A1(n7655), .A2(n7654), .ZN(n7764) );
  NAND2_X1 U5622 ( .A1(n8651), .A2(n4982), .ZN(n8623) );
  NAND2_X1 U5623 ( .A1(n7764), .A2(n5367), .ZN(n8647) );
  AND2_X1 U5624 ( .A1(n7765), .A2(n7763), .ZN(n5367) );
  CLKBUF_X1 U5625 ( .A(n7826), .Z(n8649) );
  XNOR2_X1 U5626 ( .A(n6770), .B(n7874), .ZN(n6882) );
  NOR2_X1 U5627 ( .A1(n8677), .A2(n5362), .ZN(n5361) );
  INV_X1 U5628 ( .A(n7839), .ZN(n5362) );
  NAND2_X1 U5629 ( .A1(n5557), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6134) );
  OR2_X1 U5630 ( .A1(n8314), .A2(n5796), .ZN(n5801) );
  NAND2_X1 U5631 ( .A1(n5398), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6681) );
  INV_X1 U5632 ( .A(n6679), .ZN(n5398) );
  NAND2_X1 U5633 ( .A1(n5228), .A2(n6270), .ZN(n5227) );
  NAND2_X1 U5634 ( .A1(n5135), .A2(n6323), .ZN(n5411) );
  INV_X1 U5635 ( .A(n6277), .ZN(n10485) );
  NAND2_X1 U5636 ( .A1(n6277), .A2(n6276), .ZN(n10522) );
  NOR2_X1 U5637 ( .A1(n6333), .A2(n6332), .ZN(n6995) );
  INV_X1 U5638 ( .A(n5231), .ZN(n6278) );
  NAND2_X1 U5639 ( .A1(n10512), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U5640 ( .A1(n7155), .A2(n4954), .ZN(n5137) );
  NAND2_X1 U5641 ( .A1(n5399), .A2(n6464), .ZN(n5139) );
  AOI21_X1 U5642 ( .B1(n7381), .B2(n6341), .A(n7378), .ZN(n7669) );
  INV_X1 U5643 ( .A(n5054), .ZN(n7573) );
  AOI21_X1 U5644 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n6472), .A(n7673), .ZN(
        n6284) );
  OR2_X1 U5645 ( .A1(n7572), .A2(n5916), .ZN(n5148) );
  OR2_X1 U5646 ( .A1(n8720), .A2(n5916), .ZN(n5146) );
  NAND2_X1 U5647 ( .A1(n6256), .A2(n5145), .ZN(n5144) );
  INV_X1 U5648 ( .A(n8720), .ZN(n5145) );
  XNOR2_X1 U5649 ( .A(n5051), .B(n5050), .ZN(n8733) );
  NAND2_X1 U5650 ( .A1(n5442), .A2(n5441), .ZN(n5051) );
  NAND2_X1 U5651 ( .A1(n8718), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5441) );
  INV_X1 U5652 ( .A(n6258), .ZN(n5132) );
  NAND2_X1 U5653 ( .A1(n8750), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5409) );
  AOI21_X1 U5654 ( .B1(n5406), .B2(n8807), .A(n5405), .ZN(n5404) );
  NOR2_X1 U5655 ( .A1(n6263), .A2(n6357), .ZN(n5405) );
  AND2_X1 U5656 ( .A1(n6497), .A2(n8516), .ZN(n10492) );
  NAND2_X1 U5657 ( .A1(n8815), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U5658 ( .A1(n5420), .A2(n5417), .ZN(n6180) );
  INV_X1 U5659 ( .A(n5418), .ZN(n5417) );
  AND2_X1 U5660 ( .A1(n8322), .A2(n8321), .ZN(n8850) );
  AND2_X1 U5661 ( .A1(n8488), .A2(n8855), .ZN(n8869) );
  INV_X1 U5662 ( .A(n8477), .ZN(n5462) );
  INV_X1 U5663 ( .A(n5461), .ZN(n5460) );
  OAI21_X1 U5664 ( .B1(n5462), .B2(n8472), .A(n8476), .ZN(n5461) );
  NOR2_X1 U5665 ( .A1(n6174), .A2(n5165), .ZN(n5164) );
  INV_X1 U5666 ( .A(n8694), .ZN(n8901) );
  INV_X1 U5667 ( .A(n6090), .ZN(n6076) );
  NOR2_X1 U5668 ( .A1(n6065), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6075) );
  INV_X1 U5669 ( .A(n5475), .ZN(n5474) );
  NAND2_X1 U5670 ( .A1(n8979), .A2(n8456), .ZN(n8965) );
  OAI21_X1 U5671 ( .B1(n6046), .B2(n5467), .A(n8464), .ZN(n5466) );
  NAND2_X1 U5672 ( .A1(n8938), .A2(n5473), .ZN(n5467) );
  INV_X1 U5673 ( .A(n6047), .ZN(n5473) );
  NOR2_X1 U5674 ( .A1(n6046), .A2(n5476), .ZN(n5475) );
  NAND2_X1 U5675 ( .A1(n8965), .A2(n6047), .ZN(n5477) );
  NOR2_X1 U5676 ( .A1(n6039), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U5677 ( .A1(n10144), .A2(n6025), .ZN(n6039) );
  NAND2_X1 U5678 ( .A1(n6016), .A2(n6015), .ZN(n8979) );
  NOR2_X1 U5679 ( .A1(n6010), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6025) );
  OAI21_X1 U5680 ( .B1(n5480), .B2(n5107), .A(n5105), .ZN(n6003) );
  INV_X1 U5681 ( .A(n5106), .ZN(n5105) );
  OAI21_X1 U5682 ( .B1(n5478), .B2(n5107), .A(n6002), .ZN(n5106) );
  NOR2_X1 U5683 ( .A1(n5978), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5995) );
  OR2_X1 U5684 ( .A1(n5961), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5978) );
  AND2_X1 U5685 ( .A1(n5968), .A2(n8444), .ZN(n8438) );
  OAI21_X1 U5686 ( .B1(n6160), .B2(n5432), .A(n5430), .ZN(n7746) );
  NAND2_X1 U5687 ( .A1(n5945), .A2(n5944), .ZN(n8361) );
  NAND2_X1 U5688 ( .A1(n6160), .A2(n7589), .ZN(n7682) );
  NOR2_X1 U5689 ( .A1(n5933), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U5690 ( .A1(n6159), .A2(n6158), .ZN(n7590) );
  OR2_X1 U5691 ( .A1(n5917), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5933) );
  OAI21_X1 U5692 ( .B1(n7551), .B2(n8413), .A(n8420), .ZN(n7564) );
  NAND2_X1 U5693 ( .A1(n5877), .A2(n5876), .ZN(n5904) );
  NAND2_X1 U5694 ( .A1(n10721), .A2(n8417), .ZN(n7551) );
  AND4_X1 U5695 ( .A1(n5909), .A2(n5908), .A3(n5907), .A4(n5906), .ZN(n8641)
         );
  INV_X1 U5696 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7164) );
  AND2_X1 U5697 ( .A1(n5862), .A2(n7164), .ZN(n5877) );
  INV_X1 U5698 ( .A(n6151), .ZN(n8403) );
  OR2_X1 U5699 ( .A1(n5829), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5844) );
  AND4_X1 U5700 ( .A1(n5849), .A2(n5848), .A3(n5847), .A4(n5846), .ZN(n7290)
         );
  AND2_X1 U5701 ( .A1(n8388), .A2(n8382), .ZN(n8329) );
  INV_X1 U5702 ( .A(n8371), .ZN(n10587) );
  OR2_X1 U5703 ( .A1(n6240), .A2(n6675), .ZN(n5761) );
  NAND2_X1 U5704 ( .A1(n5779), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5762) );
  AND2_X1 U5705 ( .A1(n6779), .A2(n8500), .ZN(n10637) );
  AND2_X1 U5706 ( .A1(n8500), .A2(n6373), .ZN(n9022) );
  OR2_X1 U5707 ( .A1(n8500), .A2(n6372), .ZN(n7094) );
  OR2_X1 U5708 ( .A1(n6443), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U5709 ( .A1(n8309), .A2(n8308), .ZN(n8828) );
  NAND2_X1 U5710 ( .A1(n8044), .A2(n6113), .ZN(n6024) );
  NAND2_X1 U5711 ( .A1(n5692), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U5712 ( .A1(n6203), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5690) );
  AND2_X1 U5713 ( .A1(n6204), .A2(n6203), .ZN(n6211) );
  OR2_X1 U5714 ( .A1(n6205), .A2(n5493), .ZN(n6201) );
  XNOR2_X1 U5715 ( .A(n6233), .B(n5686), .ZN(n7561) );
  INV_X1 U5716 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5972) );
  XNOR2_X1 U5717 ( .A(n5806), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6323) );
  OR2_X1 U5718 ( .A1(n9505), .A2(n9504), .ZN(n5091) );
  NAND2_X1 U5719 ( .A1(n5084), .A2(n5024), .ZN(n5092) );
  INV_X1 U5720 ( .A(n9503), .ZN(n5084) );
  AND2_X1 U5721 ( .A1(n5385), .A2(n9445), .ZN(n5384) );
  NAND2_X1 U5722 ( .A1(n5387), .A2(n5386), .ZN(n5385) );
  NAND2_X1 U5723 ( .A1(n9293), .A2(n9294), .ZN(n5391) );
  NAND2_X1 U5724 ( .A1(n5389), .A2(n9490), .ZN(n5392) );
  AND2_X1 U5725 ( .A1(n5563), .A2(n5390), .ZN(n5389) );
  INV_X1 U5726 ( .A(n6976), .ZN(n5062) );
  OR2_X1 U5727 ( .A1(n7712), .A2(n7711), .ZN(n7725) );
  AOI21_X1 U5728 ( .B1(n5368), .B2(n5069), .A(n5001), .ZN(n5068) );
  INV_X1 U5729 ( .A(n9271), .ZN(n5069) );
  AND2_X1 U5730 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n7965), .ZN(n7967) );
  NOR2_X1 U5731 ( .A1(n9191), .A2(n5394), .ZN(n5393) );
  INV_X1 U5732 ( .A(n9184), .ZN(n5394) );
  AND2_X1 U5733 ( .A1(n9258), .A2(n9257), .ZN(n9517) );
  NOR2_X1 U5734 ( .A1(n9250), .A2(n5378), .ZN(n5374) );
  AND2_X1 U5735 ( .A1(n8004), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U5736 ( .A1(n5083), .A2(n7202), .ZN(n7220) );
  OR2_X1 U5737 ( .A1(n5083), .A2(n7202), .ZN(n7221) );
  OR2_X1 U5738 ( .A1(n8076), .A2(n9705), .ZN(n8288) );
  AND2_X1 U5739 ( .A1(n8227), .A2(n9674), .ZN(n6650) );
  NAND2_X1 U5740 ( .A1(n9671), .A2(n8231), .ZN(n8185) );
  NAND2_X1 U5741 ( .A1(n5274), .A2(n6831), .ZN(n5272) );
  AOI21_X1 U5742 ( .B1(n5271), .B2(n5274), .A(n8227), .ZN(n5270) );
  AND2_X1 U5743 ( .A1(n9745), .A2(n8189), .ZN(n9754) );
  NOR2_X1 U5744 ( .A1(n7937), .A2(n7929), .ZN(n7928) );
  NAND2_X1 U5745 ( .A1(n9774), .A2(n9701), .ZN(n9775) );
  NAND2_X1 U5746 ( .A1(n5502), .A2(n5501), .ZN(n9790) );
  AOI21_X1 U5747 ( .B1(n5503), .B2(n5507), .A(n4990), .ZN(n5501) );
  AND2_X1 U5748 ( .A1(n5298), .A2(n9699), .ZN(n5297) );
  AND2_X1 U5749 ( .A1(n7957), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7947) );
  INV_X1 U5750 ( .A(n9723), .ZN(n9809) );
  NAND2_X1 U5751 ( .A1(n9850), .A2(n9696), .ZN(n9822) );
  INV_X1 U5752 ( .A(n9722), .ZN(n9847) );
  NAND2_X1 U5753 ( .A1(n5302), .A2(n5506), .ZN(n9850) );
  INV_X1 U5754 ( .A(n9846), .ZN(n5302) );
  AND2_X1 U5755 ( .A1(n9880), .A2(n9868), .ZN(n9863) );
  NOR2_X1 U5756 ( .A1(n7995), .A2(n7985), .ZN(n7984) );
  AOI21_X1 U5757 ( .B1(n5513), .B2(n4951), .A(n5512), .ZN(n5511) );
  INV_X1 U5758 ( .A(n9716), .ZN(n5512) );
  INV_X1 U5759 ( .A(n5304), .ZN(n5303) );
  AOI21_X1 U5760 ( .B1(n4949), .B2(n5306), .A(n5305), .ZN(n5304) );
  INV_X1 U5761 ( .A(n8266), .ZN(n5305) );
  NAND2_X1 U5762 ( .A1(n5308), .A2(n8263), .ZN(n9906) );
  NAND2_X1 U5763 ( .A1(n5308), .A2(n5306), .ZN(n9908) );
  INV_X1 U5764 ( .A(n9911), .ZN(n9950) );
  INV_X1 U5765 ( .A(n5319), .ZN(n5318) );
  OAI21_X1 U5766 ( .B1(n7702), .B2(n5530), .A(n5528), .ZN(n9711) );
  NAND2_X1 U5767 ( .A1(n5531), .A2(n4969), .ZN(n5530) );
  AND2_X1 U5768 ( .A1(n5529), .A2(n5559), .ZN(n5528) );
  NAND2_X1 U5769 ( .A1(n7784), .A2(n5319), .ZN(n9961) );
  NAND2_X1 U5770 ( .A1(n10753), .A2(n7721), .ZN(n7784) );
  OR2_X1 U5771 ( .A1(n7615), .A2(n7614), .ZN(n7712) );
  AND2_X1 U5772 ( .A1(n8130), .A2(n8128), .ZN(n8038) );
  NAND2_X1 U5773 ( .A1(n7524), .A2(n7525), .ZN(n7621) );
  NAND2_X1 U5774 ( .A1(n5127), .A2(n4955), .ZN(n7537) );
  AOI21_X1 U5775 ( .B1(n7361), .B2(n5500), .A(n4989), .ZN(n5499) );
  INV_X1 U5776 ( .A(n7344), .ZN(n5500) );
  NAND2_X1 U5777 ( .A1(n5314), .A2(n4966), .ZN(n7519) );
  NAND2_X1 U5778 ( .A1(n5127), .A2(n7605), .ZN(n7416) );
  NAND2_X1 U5779 ( .A1(n7265), .A2(n8087), .ZN(n7323) );
  OR2_X1 U5780 ( .A1(n7264), .A2(n7263), .ZN(n7265) );
  AND2_X1 U5781 ( .A1(n7327), .A2(n10662), .ZN(n7325) );
  NOR2_X1 U5782 ( .A1(n7125), .A2(n10618), .ZN(n7327) );
  NAND2_X1 U5783 ( .A1(n6958), .A2(n8031), .ZN(n7123) );
  INV_X1 U5784 ( .A(n9561), .ZN(n7272) );
  NAND2_X1 U5785 ( .A1(n6956), .A2(n6955), .ZN(n8092) );
  INV_X1 U5786 ( .A(n10551), .ZN(n10756) );
  NOR2_X1 U5787 ( .A1(n6726), .A2(n10567), .ZN(n7085) );
  AND2_X1 U5788 ( .A1(n6816), .A2(n6815), .ZN(n6829) );
  NAND2_X1 U5789 ( .A1(n10135), .A2(n8223), .ZN(n10551) );
  NAND2_X1 U5790 ( .A1(n9152), .A2(n8043), .ZN(n7903) );
  NAND2_X1 U5791 ( .A1(n7919), .A2(n7918), .ZN(n9765) );
  NAND2_X1 U5792 ( .A1(n7945), .A2(n7944), .ZN(n10015) );
  NAND2_X1 U5793 ( .A1(n8025), .A2(n8024), .ZN(n9971) );
  NAND2_X1 U5794 ( .A1(n7710), .A2(n7709), .ZN(n9212) );
  AND2_X1 U5795 ( .A1(n5127), .A2(n4958), .ZN(n7538) );
  NAND2_X1 U5796 ( .A1(n7351), .A2(n7361), .ZN(n7391) );
  NAND2_X1 U5797 ( .A1(n7345), .A2(n7344), .ZN(n7351) );
  OR2_X1 U5798 ( .A1(n7394), .A2(n6716), .ZN(n6717) );
  INV_X1 U5799 ( .A(n10765), .ZN(n10619) );
  INV_X1 U5800 ( .A(n10767), .ZN(n10623) );
  XNOR2_X1 U5801 ( .A(n8067), .B(n8066), .ZN(n8306) );
  XNOR2_X1 U5802 ( .A(n7884), .B(SI_29_), .ZN(n9152) );
  XNOR2_X1 U5803 ( .A(n5734), .B(n5733), .ZN(n9155) );
  NAND2_X1 U5804 ( .A1(n5329), .A2(n6390), .ZN(n6396) );
  AND3_X1 U5805 ( .A1(n5541), .A2(n6389), .A3(n5019), .ZN(n5329) );
  NAND2_X1 U5806 ( .A1(n6405), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6482) );
  INV_X1 U5807 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6616) );
  OR2_X1 U5808 ( .A1(n6697), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6698) );
  OR2_X1 U5809 ( .A1(n6574), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6697) );
  AND2_X1 U5810 ( .A1(n6570), .A2(n6574), .ZN(n7704) );
  XNOR2_X1 U5811 ( .A(n5925), .B(n5924), .ZN(n7703) );
  NAND2_X1 U5812 ( .A1(n5264), .A2(n5601), .ZN(n5899) );
  NAND2_X1 U5813 ( .A1(n5884), .A2(n5561), .ZN(n5264) );
  NAND2_X1 U5814 ( .A1(n5587), .A2(n5586), .ZN(n5836) );
  AND2_X1 U5815 ( .A1(n6424), .A2(n6423), .ZN(n6528) );
  NAND2_X1 U5816 ( .A1(n5581), .A2(n5580), .ZN(n5803) );
  XNOR2_X1 U5817 ( .A(n5571), .B(n5568), .ZN(n5757) );
  NAND3_X1 U5818 ( .A1(n5242), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5241) );
  INV_X1 U5819 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5242) );
  NOR2_X1 U5820 ( .A1(n7288), .A2(n5567), .ZN(n7294) );
  NAND2_X1 U5821 ( .A1(n5694), .A2(n5693), .ZN(n8859) );
  AND4_X1 U5822 ( .A1(n5954), .A2(n5953), .A3(n5952), .A4(n5951), .ZN(n8566)
         );
  NAND2_X1 U5823 ( .A1(n6088), .A2(n6087), .ZN(n8904) );
  NAND2_X1 U5824 ( .A1(n6890), .A2(n6889), .ZN(n6903) );
  AND2_X1 U5825 ( .A1(n7131), .A2(n6774), .ZN(n6789) );
  NAND2_X1 U5826 ( .A1(n8651), .A2(n7830), .ZN(n8571) );
  NAND2_X1 U5827 ( .A1(n5994), .A2(n5993), .ZN(n9010) );
  OAI21_X1 U5828 ( .B1(n6890), .B2(n5335), .A(n5331), .ZN(n7018) );
  NOR2_X1 U5829 ( .A1(n6889), .A2(n5334), .ZN(n5333) );
  NAND2_X1 U5830 ( .A1(n6099), .A2(n6098), .ZN(n8891) );
  INV_X1 U5831 ( .A(n9019), .ZN(n6773) );
  NAND2_X1 U5832 ( .A1(n7862), .A2(n4979), .ZN(n8635) );
  INV_X1 U5833 ( .A(n7861), .ZN(n5357) );
  NAND2_X1 U5834 ( .A1(n7862), .A2(n7861), .ZN(n8634) );
  XNOR2_X1 U5835 ( .A(n6882), .B(n8708), .ZN(n6777) );
  OR2_X1 U5836 ( .A1(n8657), .A2(n8656), .ZN(n8658) );
  INV_X1 U5837 ( .A(n8680), .ZN(n8663) );
  INV_X1 U5838 ( .A(n5364), .ZN(n7288) );
  NAND2_X1 U5839 ( .A1(n7255), .A2(n7254), .ZN(n7256) );
  NAND2_X1 U5840 ( .A1(n5713), .A2(n5712), .ZN(n8871) );
  NAND2_X1 U5841 ( .A1(n8535), .A2(n5361), .ZN(n5556) );
  NAND2_X1 U5842 ( .A1(n8535), .A2(n7839), .ZN(n8678) );
  AND2_X1 U5843 ( .A1(n6780), .A2(n6757), .ZN(n8686) );
  NAND2_X1 U5844 ( .A1(n8514), .A2(n8513), .ZN(n5210) );
  XNOR2_X1 U5845 ( .A(n6137), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8520) );
  OR2_X1 U5846 ( .A1(n5010), .A2(n6019), .ZN(n6136) );
  NAND4_X1 U5847 ( .A1(n5719), .A2(n5718), .A3(n5717), .A4(n5716), .ZN(n8692)
         );
  INV_X1 U5848 ( .A(n8566), .ZN(n8700) );
  OR2_X1 U5849 ( .A1(n5786), .A2(n5751), .ZN(n5752) );
  NAND2_X1 U5850 ( .A1(n5150), .A2(n5149), .ZN(n10469) );
  NOR2_X1 U5851 ( .A1(n10479), .A2(n10478), .ZN(n10477) );
  AND2_X1 U5852 ( .A1(n5230), .A2(n4953), .ZN(n10479) );
  AOI21_X1 U5853 ( .B1(n6323), .B2(n6322), .A(n10461), .ZN(n10476) );
  INV_X1 U5854 ( .A(n5401), .ZN(n10508) );
  INV_X1 U5855 ( .A(n5446), .ZN(n7375) );
  NOR2_X1 U5856 ( .A1(n6254), .A2(n7373), .ZN(n7664) );
  INV_X1 U5857 ( .A(n6282), .ZN(n5445) );
  AOI21_X1 U5858 ( .B1(n6133), .B2(n6132), .A(n6131), .ZN(n8833) );
  NAND2_X1 U5859 ( .A1(n6115), .A2(n6114), .ZN(n9045) );
  NAND2_X1 U5860 ( .A1(n6082), .A2(n8472), .ZN(n8902) );
  NAND2_X1 U5861 ( .A1(n6173), .A2(n6172), .ZN(n5166) );
  NAND2_X1 U5862 ( .A1(n6168), .A2(n6167), .ZN(n8975) );
  NAND2_X1 U5863 ( .A1(n7745), .A2(n5969), .ZN(n7812) );
  NAND2_X1 U5864 ( .A1(n5976), .A2(n5975), .ZN(n8356) );
  NAND2_X1 U5865 ( .A1(n5465), .A2(n5463), .ZN(n10721) );
  NOR2_X1 U5866 ( .A1(n8334), .A2(n5464), .ZN(n5463) );
  INV_X1 U5867 ( .A(n8404), .ZN(n5464) );
  NAND2_X1 U5868 ( .A1(n5465), .A2(n8404), .ZN(n7339) );
  AND2_X1 U5869 ( .A1(n5874), .A2(n5007), .ZN(n5438) );
  OR2_X1 U5870 ( .A1(n7346), .A2(n5858), .ZN(n5859) );
  OR2_X1 U5871 ( .A1(n9021), .A2(n10598), .ZN(n10653) );
  AND2_X1 U5872 ( .A1(n10709), .A2(n10700), .ZN(n9015) );
  AND2_X1 U5873 ( .A1(n8305), .A2(n8304), .ZN(n9094) );
  INV_X1 U5874 ( .A(n8828), .ZN(n9098) );
  INV_X1 U5875 ( .A(n8839), .ZN(n9102) );
  INV_X1 U5876 ( .A(n8859), .ZN(n9105) );
  AND2_X1 U5877 ( .A1(n10720), .A2(n9038), .ZN(n5155) );
  OR2_X1 U5878 ( .A1(n9066), .A2(n9065), .ZN(n9126) );
  OR2_X1 U5879 ( .A1(n9070), .A2(n9069), .ZN(n9127) );
  INV_X1 U5880 ( .A(n8655), .ZN(n9135) );
  NAND2_X1 U5881 ( .A1(n6758), .A2(n6443), .ZN(n6450) );
  XNOR2_X1 U5882 ( .A(n6208), .B(n6207), .ZN(n7741) );
  XNOR2_X1 U5883 ( .A(n6206), .B(n5495), .ZN(n7698) );
  INV_X1 U5884 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7174) );
  INV_X1 U5885 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6913) );
  INV_X1 U5886 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6899) );
  INV_X1 U5887 ( .A(n6301), .ZN(n8784) );
  INV_X1 U5888 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6694) );
  INV_X1 U5889 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6493) );
  INV_X1 U5890 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6470) );
  INV_X1 U5891 ( .A(n7678), .ZN(n6472) );
  INV_X1 U5892 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6463) );
  INV_X1 U5893 ( .A(n6323), .ZN(n10459) );
  OAI21_X1 U5894 ( .B1(n5780), .B2(n5450), .A(n5449), .ZN(n5782) );
  NAND2_X1 U5895 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5450) );
  NAND2_X1 U5896 ( .A1(n5807), .A2(n5781), .ZN(n5449) );
  NAND2_X1 U5897 ( .A1(n7783), .A2(n7782), .ZN(n9708) );
  NAND2_X1 U5898 ( .A1(n9490), .A2(n5563), .ZN(n9489) );
  NAND2_X1 U5899 ( .A1(n6977), .A2(n6976), .ZN(n7029) );
  AND3_X1 U5900 ( .A1(n9528), .A2(n9320), .A3(n9321), .ZN(n9379) );
  BUF_X1 U5901 ( .A(n6797), .Z(n6726) );
  NAND2_X1 U5902 ( .A1(n5373), .A2(n9279), .ZN(n9404) );
  NAND2_X1 U5903 ( .A1(n9468), .A2(n9469), .ZN(n5373) );
  INV_X1 U5904 ( .A(n9825), .ZN(n9794) );
  INV_X1 U5905 ( .A(n9553), .ZN(n9948) );
  INV_X1 U5906 ( .A(n5088), .ZN(n5087) );
  NAND2_X1 U5907 ( .A1(n5086), .A2(n5024), .ZN(n5085) );
  OAI21_X1 U5908 ( .B1(n5376), .B2(n5089), .A(n5377), .ZN(n5088) );
  NAND2_X1 U5909 ( .A1(n8013), .A2(n8012), .ZN(n9952) );
  AND2_X1 U5910 ( .A1(n5392), .A2(n5391), .ZN(n9449) );
  NAND2_X1 U5911 ( .A1(n5071), .A2(n9271), .ZN(n9468) );
  NAND2_X1 U5912 ( .A1(n9363), .A2(n9364), .ZN(n5071) );
  NAND2_X1 U5913 ( .A1(n7983), .A2(n7982), .ZN(n9881) );
  INV_X1 U5914 ( .A(n9542), .ZN(n9496) );
  OAI211_X1 U5915 ( .C1(n7392), .C2(n6847), .A(n6846), .B(n6845), .ZN(n8079)
         );
  NAND2_X1 U5916 ( .A1(n5381), .A2(n7221), .ZN(n7423) );
  NAND2_X1 U5917 ( .A1(n7220), .A2(n7219), .ZN(n5381) );
  NAND3_X1 U5918 ( .A1(n9527), .A2(n9530), .A3(n9526), .ZN(n9528) );
  AND2_X1 U5919 ( .A1(n6644), .A2(n6642), .ZN(n9529) );
  INV_X1 U5920 ( .A(n9529), .ZN(n9548) );
  INV_X1 U5921 ( .A(n7546), .ZN(n6613) );
  AND4_X1 U5922 ( .A1(n7907), .A2(n7906), .A3(n7905), .A4(n7904), .ZN(n10369)
         );
  NAND4_X1 U5923 ( .A1(n6864), .A2(n6863), .A3(n6862), .A4(n6861), .ZN(n9562)
         );
  NAND2_X1 U5924 ( .A1(n7898), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6864) );
  NAND2_X1 U5925 ( .A1(n7206), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6862) );
  INV_X1 U5926 ( .A(n6392), .ZN(n6914) );
  OR2_X1 U5927 ( .A1(n9658), .A2(n9657), .ZN(n9673) );
  NOR2_X1 U5928 ( .A1(n9683), .A2(n9915), .ZN(n9982) );
  INV_X1 U5929 ( .A(n5546), .ZN(n5545) );
  AOI21_X1 U5930 ( .B1(n5546), .B2(n5544), .A(n4962), .ZN(n5543) );
  INV_X1 U5931 ( .A(n5325), .ZN(n5324) );
  NAND2_X1 U5932 ( .A1(n5327), .A2(n10752), .ZN(n5326) );
  OAI22_X1 U5933 ( .A1(n9728), .A2(n9949), .B1(n9706), .B2(n9705), .ZN(n5325)
         );
  NAND2_X1 U5934 ( .A1(n5504), .A2(n5505), .ZN(n9804) );
  OR2_X1 U5935 ( .A1(n9838), .A2(n5507), .ZN(n5504) );
  AND2_X1 U5936 ( .A1(n5509), .A2(n4974), .ZN(n9818) );
  NAND2_X1 U5937 ( .A1(n9838), .A2(n9845), .ZN(n5509) );
  OAI21_X1 U5938 ( .B1(n9939), .B2(n5516), .A(n4951), .ZN(n9888) );
  NAND2_X1 U5939 ( .A1(n5519), .A2(n5520), .ZN(n9904) );
  NAND2_X1 U5940 ( .A1(n9939), .A2(n5521), .ZN(n5519) );
  NAND2_X1 U5941 ( .A1(n9939), .A2(n5560), .ZN(n9924) );
  NAND2_X1 U5942 ( .A1(n5527), .A2(n5531), .ZN(n7779) );
  NAND2_X1 U5943 ( .A1(n7702), .A2(n5534), .ZN(n5527) );
  INV_X1 U5944 ( .A(n5535), .ZN(n5533) );
  NAND2_X1 U5945 ( .A1(n5538), .A2(n5537), .ZN(n5536) );
  INV_X1 U5946 ( .A(n9188), .ZN(n10729) );
  INV_X1 U5947 ( .A(n10618), .ZN(n7271) );
  NAND2_X1 U5948 ( .A1(n7635), .A2(n7083), .ZN(n10781) );
  NAND2_X1 U5949 ( .A1(n6646), .A2(n10553), .ZN(n7126) );
  AND2_X1 U5950 ( .A1(n8227), .A2(n9671), .ZN(n10553) );
  AND2_X2 U5951 ( .A1(n6822), .A2(n6821), .ZN(n10770) );
  INV_X1 U5952 ( .A(n9682), .ZN(n10073) );
  INV_X1 U5953 ( .A(n8076), .ZN(n10077) );
  NAND2_X1 U5954 ( .A1(n5002), .A2(n5321), .ZN(n10078) );
  NOR2_X1 U5955 ( .A1(n9990), .A2(n5322), .ZN(n5321) );
  NAND2_X1 U5956 ( .A1(n9992), .A2(n5323), .ZN(n5322) );
  NAND2_X1 U5957 ( .A1(n9991), .A2(n10619), .ZN(n5323) );
  INV_X1 U5958 ( .A(n9765), .ZN(n10083) );
  INV_X1 U5959 ( .A(n9797), .ZN(n10088) );
  INV_X1 U5960 ( .A(n9831), .ZN(n10093) );
  INV_X1 U5961 ( .A(n9952), .ZN(n10114) );
  INV_X1 U5962 ( .A(n9971), .ZN(n10118) );
  INV_X1 U5963 ( .A(n9212), .ZN(n9488) );
  NAND2_X1 U5964 ( .A1(n10774), .A2(n10619), .ZN(n10122) );
  AOI21_X1 U5965 ( .B1(n6640), .B2(n6456), .A(n6454), .ZN(n6827) );
  NAND2_X1 U5966 ( .A1(n6651), .A2(n6468), .ZN(n10141) );
  AND2_X1 U5967 ( .A1(n5017), .A2(n6481), .ZN(n5552) );
  INV_X1 U5968 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5553) );
  XNOR2_X1 U5969 ( .A(n6401), .B(P1_IR_REG_24__SCAN_IN), .ZN(n7700) );
  XNOR2_X1 U5970 ( .A(n6482), .B(n6406), .ZN(n7546) );
  INV_X1 U5971 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7173) );
  INV_X1 U5972 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6898) );
  AND2_X1 U5973 ( .A1(n6490), .A2(n6461), .ZN(n7512) );
  NOR2_X1 U5974 ( .A1(n6744), .A2(n6242), .ZN(P2_U3893) );
  NAND2_X1 U5975 ( .A1(n5341), .A2(n8624), .ZN(n5339) );
  INV_X1 U5976 ( .A(n5238), .ZN(n8712) );
  INV_X1 U5977 ( .A(n5133), .ZN(n8727) );
  INV_X1 U5978 ( .A(n5240), .ZN(n8744) );
  INV_X1 U5979 ( .A(n5397), .ZN(n8776) );
  AOI21_X1 U5980 ( .B1(n4960), .B2(n10525), .A(n5045), .ZN(n8804) );
  INV_X1 U5981 ( .A(n5128), .ZN(n8794) );
  AOI21_X1 U5982 ( .B1(n5234), .B2(n10525), .A(n5232), .ZN(n8822) );
  AOI21_X1 U5983 ( .B1(n5454), .B2(n10525), .A(n5451), .ZN(n6366) );
  AND2_X1 U5984 ( .A1(n6367), .A2(n6365), .ZN(n5055) );
  OR2_X1 U5985 ( .A1(n5452), .A2(n6300), .ZN(n5451) );
  OAI21_X1 U5986 ( .B1(n6378), .B2(n10805), .A(n5435), .ZN(P2_U3488) );
  NOR2_X1 U5987 ( .A1(n5436), .A2(n5027), .ZN(n5435) );
  NOR2_X1 U5988 ( .A1(n10806), .A2(n6379), .ZN(n5436) );
  OAI21_X1 U5989 ( .B1(n6378), .B2(n10807), .A(n6238), .ZN(P2_U3456) );
  OAI21_X1 U5990 ( .B1(n8834), .B2(n9143), .A(n6236), .ZN(n6237) );
  NAND2_X1 U5991 ( .A1(n5154), .A2(n5152), .ZN(P2_U3454) );
  INV_X1 U5992 ( .A(n5153), .ZN(n5152) );
  OR2_X1 U5993 ( .A1(n9103), .A2(n10807), .ZN(n5154) );
  OAI22_X1 U5994 ( .A1(n9105), .A2(n9143), .B1(n10810), .B2(n9104), .ZN(n5153)
         );
  AOI211_X1 U5995 ( .C1(n9994), .C2(n9972), .A(n9752), .B(n9751), .ZN(n9753)
         );
  INV_X1 U5996 ( .A(n9845), .ZN(n5506) );
  NAND2_X1 U5997 ( .A1(n8263), .A2(n8153), .ZN(n4949) );
  AND2_X1 U5998 ( .A1(n5265), .A2(n5263), .ZN(n4950) );
  AND2_X1 U5999 ( .A1(n4993), .A2(n5514), .ZN(n4951) );
  NAND2_X1 U6000 ( .A1(n6273), .A2(n10459), .ZN(n4953) );
  AND2_X1 U6001 ( .A1(n5141), .A2(n7381), .ZN(n4954) );
  AND2_X1 U6002 ( .A1(n10691), .A2(n7605), .ZN(n4955) );
  OR2_X1 U6003 ( .A1(n8859), .A2(n8843), .ZN(n4956) );
  OR2_X1 U6004 ( .A1(n9797), .A2(n9809), .ZN(n9773) );
  INV_X1 U6005 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10124) );
  NAND2_X1 U6006 ( .A1(n7613), .A2(n7612), .ZN(n9197) );
  NOR2_X1 U6007 ( .A1(n9226), .A2(n9225), .ZN(n4957) );
  AND2_X1 U6008 ( .A1(n4955), .A2(n10713), .ZN(n4958) );
  INV_X1 U6009 ( .A(n8209), .ZN(n5179) );
  NAND2_X1 U6010 ( .A1(n7909), .A2(n7908), .ZN(n9995) );
  XOR2_X1 U6011 ( .A(n8853), .B(n8857), .Z(n4959) );
  OR2_X1 U6012 ( .A1(n8814), .A2(n4967), .ZN(n4960) );
  AND2_X1 U6013 ( .A1(n5540), .A2(n9509), .ZN(n4961) );
  AND2_X1 U6014 ( .A1(n9995), .A2(n5550), .ZN(n4962) );
  AND2_X1 U6015 ( .A1(n7845), .A2(n4984), .ZN(n4963) );
  AND2_X1 U6016 ( .A1(n8859), .A2(n8843), .ZN(n4964) );
  NAND2_X1 U6017 ( .A1(n6903), .A2(n5330), .ZN(n7016) );
  INV_X1 U6018 ( .A(n5779), .ZN(n5861) );
  INV_X1 U6019 ( .A(n8705), .ZN(n5437) );
  OR2_X1 U6020 ( .A1(n6396), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4965) );
  AND2_X1 U6021 ( .A1(n8238), .A2(n8239), .ZN(n4966) );
  AND2_X1 U6022 ( .A1(n8800), .A2(n8993), .ZN(n4967) );
  OR2_X1 U6023 ( .A1(n6344), .A2(n6284), .ZN(n4968) );
  OR2_X1 U6024 ( .A1(n9212), .A2(n10757), .ZN(n4969) );
  AND2_X1 U6025 ( .A1(n8169), .A2(n8174), .ZN(n4970) );
  AND2_X1 U6026 ( .A1(n8129), .A2(n8174), .ZN(n4971) );
  OR3_X1 U6027 ( .A1(n8819), .A2(n8821), .A3(n10464), .ZN(n4972) );
  XNOR2_X1 U6028 ( .A(n5870), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7165) );
  INV_X1 U6029 ( .A(n8196), .ZN(n5202) );
  OR2_X1 U6030 ( .A1(n6353), .A2(n6262), .ZN(n4973) );
  INV_X1 U6031 ( .A(n8938), .ZN(n5476) );
  AND2_X1 U6032 ( .A1(n8213), .A2(n8281), .ZN(n9729) );
  INV_X1 U6033 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5495) );
  INV_X1 U6034 ( .A(n9756), .ZN(n5175) );
  INV_X1 U6035 ( .A(n6997), .ZN(n6436) );
  AND2_X1 U6036 ( .A1(n5869), .A2(n5855), .ZN(n6997) );
  INV_X1 U6037 ( .A(n8444), .ZN(n5428) );
  NOR2_X1 U6038 ( .A1(n6614), .A2(n6393), .ZN(n6605) );
  NAND2_X1 U6039 ( .A1(n5524), .A2(n6381), .ZN(n6420) );
  OR2_X1 U6040 ( .A1(n10024), .A2(n9826), .ZN(n4974) );
  AND2_X1 U6041 ( .A1(n8273), .A2(n8181), .ZN(n4975) );
  INV_X1 U6042 ( .A(n7155), .ZN(n5140) );
  OR2_X1 U6043 ( .A1(n6396), .A2(n5111), .ZN(n5113) );
  INV_X1 U6044 ( .A(n7890), .ZN(n5617) );
  NOR2_X1 U6045 ( .A1(n9905), .A2(n5307), .ZN(n5306) );
  OR2_X1 U6046 ( .A1(n8219), .A2(n8181), .ZN(n4976) );
  NAND2_X1 U6047 ( .A1(n8499), .A2(n8498), .ZN(n8328) );
  INV_X1 U6048 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5807) );
  AND2_X1 U6049 ( .A1(n5547), .A2(n9727), .ZN(n4977) );
  INV_X1 U6050 ( .A(n9932), .ZN(n10110) );
  NAND2_X1 U6051 ( .A1(n8003), .A2(n8002), .ZN(n9932) );
  AND2_X1 U6052 ( .A1(n8175), .A2(n9744), .ZN(n4978) );
  NOR2_X1 U6053 ( .A1(n8633), .A2(n5357), .ZN(n4979) );
  INV_X1 U6054 ( .A(n9343), .ZN(n5390) );
  INV_X1 U6055 ( .A(n5539), .ZN(n5537) );
  NOR2_X1 U6056 ( .A1(n9197), .A2(n10758), .ZN(n5539) );
  INV_X1 U6057 ( .A(n10005), .ZN(n9787) );
  NAND2_X1 U6058 ( .A1(n7927), .A2(n7926), .ZN(n10005) );
  AND2_X1 U6059 ( .A1(n7293), .A2(n5363), .ZN(n4980) );
  AND2_X1 U6060 ( .A1(n4983), .A2(n5687), .ZN(n4981) );
  AND2_X1 U6061 ( .A1(n7831), .A2(n7830), .ZN(n4982) );
  AND3_X1 U6062 ( .A1(n6207), .A2(n5495), .A3(n5494), .ZN(n4983) );
  OR2_X1 U6063 ( .A1(n7846), .A2(n5358), .ZN(n4984) );
  INV_X1 U6064 ( .A(n5517), .ZN(n5516) );
  NOR2_X1 U6065 ( .A1(n9715), .A2(n5518), .ZN(n5517) );
  AND2_X1 U6066 ( .A1(n5133), .A2(n5132), .ZN(n4985) );
  INV_X1 U6067 ( .A(n6388), .ZN(n6389) );
  AND2_X1 U6068 ( .A1(n5142), .A2(n5141), .ZN(n4986) );
  AND2_X1 U6069 ( .A1(n9831), .A2(n9722), .ZN(n4987) );
  NOR2_X1 U6070 ( .A1(n8707), .A2(n7013), .ZN(n4988) );
  INV_X1 U6071 ( .A(n5565), .ZN(n5426) );
  AND2_X1 U6072 ( .A1(n7390), .A2(n7605), .ZN(n4989) );
  AND2_X1 U6073 ( .A1(n9815), .A2(n9794), .ZN(n4990) );
  INV_X1 U6074 ( .A(n5378), .ZN(n5377) );
  NOR2_X1 U6075 ( .A1(n5380), .A2(n5379), .ZN(n5378) );
  AND2_X1 U6076 ( .A1(n7424), .A2(n7425), .ZN(n4991) );
  AND2_X1 U6077 ( .A1(n8655), .A2(n8958), .ZN(n4992) );
  OR2_X1 U6078 ( .A1(n10106), .A2(n9714), .ZN(n4993) );
  INV_X1 U6079 ( .A(n6161), .ZN(n5432) );
  NAND2_X1 U6080 ( .A1(n6419), .A2(n6380), .ZN(n6412) );
  NAND2_X1 U6081 ( .A1(n8839), .A2(n8691), .ZN(n4994) );
  AND2_X1 U6082 ( .A1(n4976), .A2(n8218), .ZN(n4995) );
  INV_X1 U6083 ( .A(n5564), .ZN(n5425) );
  AND2_X1 U6084 ( .A1(n7873), .A2(n8843), .ZN(n4996) );
  OR2_X1 U6085 ( .A1(n6205), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n4997) );
  AND2_X1 U6086 ( .A1(n5604), .A2(SI_10_), .ZN(n4998) );
  NAND2_X1 U6087 ( .A1(n5220), .A2(n5217), .ZN(n4999) );
  AND2_X1 U6088 ( .A1(n6297), .A2(n6296), .ZN(n5000) );
  NAND2_X1 U6089 ( .A1(n5370), .A2(n9287), .ZN(n5001) );
  INV_X1 U6090 ( .A(n5399), .ZN(n5141) );
  NOR2_X1 U6091 ( .A1(n7165), .A2(n6310), .ZN(n5399) );
  INV_X1 U6092 ( .A(n4949), .ZN(n5309) );
  AND2_X1 U6093 ( .A1(n5326), .A2(n5324), .ZN(n5002) );
  INV_X1 U6094 ( .A(n5352), .ZN(n5351) );
  AND2_X1 U6095 ( .A1(n8524), .A2(n5353), .ZN(n5352) );
  OR2_X1 U6096 ( .A1(n4964), .A2(n5564), .ZN(n5003) );
  OR2_X1 U6097 ( .A1(n9815), .A2(n9794), .ZN(n5004) );
  AND2_X1 U6098 ( .A1(n8486), .A2(n8485), .ZN(n5005) );
  NOR2_X1 U6099 ( .A1(n8704), .A2(n10724), .ZN(n5006) );
  OR2_X1 U6100 ( .A1(n6442), .A2(n6240), .ZN(n5007) );
  NOR2_X1 U6101 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5008) );
  NOR2_X1 U6102 ( .A1(n5082), .A2(n5078), .ZN(n5009) );
  NAND3_X1 U6103 ( .A1(n6020), .A2(n5685), .A3(n5684), .ZN(n5010) );
  OR2_X1 U6104 ( .A1(n9125), .A2(n8900), .ZN(n5011) );
  AND2_X1 U6105 ( .A1(n8857), .A2(n8489), .ZN(n5012) );
  AND2_X1 U6106 ( .A1(n5430), .A2(n5968), .ZN(n5013) );
  AND2_X1 U6107 ( .A1(n4951), .A2(n8000), .ZN(n5014) );
  NAND2_X1 U6108 ( .A1(n7027), .A2(n7026), .ZN(n5015) );
  NAND2_X1 U6109 ( .A1(n10471), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5016) );
  AND2_X1 U6110 ( .A1(n6593), .A2(n5553), .ZN(n5017) );
  AND2_X1 U6111 ( .A1(n5380), .A2(n5379), .ZN(n5018) );
  NOR2_X1 U6112 ( .A1(n6399), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5019) );
  AND2_X1 U6113 ( .A1(n5542), .A2(n6394), .ZN(n5020) );
  OR2_X1 U6114 ( .A1(n7846), .A2(n5360), .ZN(n5021) );
  INV_X1 U6115 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5093) );
  NAND2_X1 U6116 ( .A1(n10471), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5022) );
  AND2_X1 U6117 ( .A1(n5137), .A2(n5139), .ZN(n5023) );
  NAND2_X1 U6118 ( .A1(n5898), .A2(n5601), .ZN(n5268) );
  INV_X1 U6119 ( .A(n6608), .ZN(n9376) );
  INV_X1 U6120 ( .A(n8054), .ZN(n7993) );
  INV_X2 U6121 ( .A(n7993), .ZN(n7948) );
  NAND2_X1 U6122 ( .A1(n9505), .A2(n9504), .ZN(n5024) );
  NAND2_X1 U6123 ( .A1(n5092), .A2(n5091), .ZN(n9327) );
  INV_X1 U6124 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U6125 ( .A1(n5536), .A2(n5533), .ZN(n10751) );
  INV_X1 U6126 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6406) );
  INV_X1 U6127 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5094) );
  INV_X1 U6128 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5892) );
  OR2_X1 U6129 ( .A1(n9881), .A2(n9861), .ZN(n9857) );
  INV_X1 U6130 ( .A(n9857), .ZN(n5199) );
  AND4_X1 U6131 ( .A1(n7917), .A2(n7916), .A3(n7915), .A4(n7914), .ZN(n9728)
         );
  INV_X1 U6132 ( .A(n9728), .ZN(n5550) );
  NAND2_X1 U6133 ( .A1(n7903), .A2(n7902), .ZN(n9991) );
  INV_X1 U6134 ( .A(n9991), .ZN(n5123) );
  NOR2_X1 U6135 ( .A1(n9968), .A2(n5115), .ZN(n5114) );
  AND2_X1 U6136 ( .A1(n8490), .A2(n8855), .ZN(n5025) );
  AND2_X1 U6137 ( .A1(n5480), .A2(n5955), .ZN(n5026) );
  NOR2_X1 U6138 ( .A1(n8834), .A2(n9089), .ZN(n5027) );
  INV_X1 U6139 ( .A(n5121), .ZN(n9914) );
  NOR2_X1 U6140 ( .A1(n9968), .A2(n5118), .ZN(n5121) );
  AND2_X1 U6141 ( .A1(n7784), .A2(n8142), .ZN(n5028) );
  AND2_X1 U6142 ( .A1(n8212), .A2(n9703), .ZN(n9744) );
  INV_X1 U6143 ( .A(n9744), .ZN(n5551) );
  AND2_X1 U6144 ( .A1(n5314), .A2(n8239), .ZN(n5029) );
  INV_X1 U6145 ( .A(n8667), .ZN(n5353) );
  NOR2_X1 U6146 ( .A1(n9227), .A2(n4957), .ZN(n5030) );
  AND2_X1 U6147 ( .A1(n5148), .A2(n5147), .ZN(n5031) );
  NAND2_X2 U6148 ( .A1(n9021), .A2(n10650), .ZN(n10709) );
  INV_X1 U6149 ( .A(n7367), .ZN(n5127) );
  NAND2_X1 U6150 ( .A1(n7992), .A2(n7991), .ZN(n9897) );
  INV_X1 U6151 ( .A(n9897), .ZN(n5120) );
  NAND2_X1 U6152 ( .A1(n7706), .A2(n7705), .ZN(n10778) );
  INV_X1 U6153 ( .A(n10778), .ZN(n5540) );
  OR2_X1 U6154 ( .A1(n5711), .A2(n5290), .ZN(n5032) );
  AND2_X1 U6155 ( .A1(n10516), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n5033) );
  INV_X1 U6156 ( .A(n10805), .ZN(n10806) );
  INV_X1 U6157 ( .A(n10748), .ZN(n10805) );
  AND2_X1 U6158 ( .A1(n5008), .A2(n6020), .ZN(n5162) );
  INV_X1 U6159 ( .A(n5534), .ZN(n5532) );
  NOR2_X1 U6160 ( .A1(n10755), .A2(n5535), .ZN(n5534) );
  AND2_X1 U6161 ( .A1(n5446), .A2(n5445), .ZN(n5034) );
  AND2_X1 U6162 ( .A1(n6476), .A2(n6481), .ZN(n6594) );
  NAND4_X1 U6163 ( .A1(n5162), .A2(n5161), .A3(n4952), .A4(n5336), .ZN(n5035)
         );
  AND2_X1 U6164 ( .A1(n6903), .A2(n6902), .ZN(n5036) );
  OR2_X1 U6165 ( .A1(n6308), .A2(n5932), .ZN(n5037) );
  INV_X1 U6166 ( .A(n6307), .ZN(n5050) );
  AND2_X1 U6167 ( .A1(n6185), .A2(n6224), .ZN(n9000) );
  INV_X1 U6168 ( .A(n9000), .ZN(n10641) );
  AND2_X1 U6169 ( .A1(n8186), .A2(n6807), .ZN(n10563) );
  INV_X1 U6170 ( .A(n10563), .ZN(n10752) );
  OR2_X1 U6171 ( .A1(n8807), .A2(n6357), .ZN(n5038) );
  INV_X1 U6172 ( .A(n6800), .ZN(n8029) );
  NAND2_X1 U6173 ( .A1(n8784), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5039) );
  INV_X1 U6174 ( .A(n5407), .ZN(n5406) );
  NAND2_X1 U6175 ( .A1(n6263), .A2(n6357), .ZN(n5407) );
  AND2_X1 U6176 ( .A1(n5404), .A2(n5407), .ZN(n5040) );
  AND2_X1 U6177 ( .A1(n5151), .A2(n5412), .ZN(n5041) );
  INV_X1 U6178 ( .A(n6831), .ZN(n8231) );
  XNOR2_X1 U6179 ( .A(n6483), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6831) );
  XNOR2_X1 U6180 ( .A(n6134), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8515) );
  INV_X1 U6181 ( .A(n8515), .ZN(n7176) );
  NAND2_X1 U6182 ( .A1(n5075), .A2(n5072), .ZN(n8227) );
  INV_X1 U6183 ( .A(n8227), .ZN(n6836) );
  INV_X1 U6184 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5246) );
  INV_X1 U6185 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6186 ( .A1(n7767), .A2(n7766), .ZN(n5042) );
  NAND2_X1 U6187 ( .A1(n8611), .A2(n8610), .ZN(n8609) );
  INV_X1 U6188 ( .A(n6247), .ZN(n5135) );
  NAND2_X1 U6189 ( .A1(n5412), .A2(n5411), .ZN(n10454) );
  NOR2_X1 U6190 ( .A1(n10487), .A2(n5812), .ZN(n10488) );
  NAND2_X1 U6191 ( .A1(n6366), .A2(n5055), .ZN(P2_U3201) );
  OAI21_X2 U6192 ( .B1(n8898), .B2(n6175), .A(n6176), .ZN(n8888) );
  NAND2_X1 U6193 ( .A1(n8925), .A2(n8924), .ZN(n6173) );
  NAND2_X1 U6194 ( .A1(n6164), .A2(n8440), .ZN(n8999) );
  NAND2_X1 U6195 ( .A1(n5167), .A2(n5427), .ZN(n7815) );
  NAND2_X1 U6196 ( .A1(n5058), .A2(n5476), .ZN(n8941) );
  NAND2_X1 U6197 ( .A1(n5158), .A2(n5156), .ZN(n9037) );
  OAI21_X1 U6198 ( .B1(n8866), .B2(n5426), .A(n5425), .ZN(n5168) );
  AOI21_X1 U6199 ( .B1(n7336), .B2(n8334), .A(n5006), .ZN(n5433) );
  MUX2_X1 U6200 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7890), .Z(n5575) );
  AND2_X2 U6201 ( .A1(n5243), .A2(n5241), .ZN(n7890) );
  INV_X1 U6202 ( .A(n10705), .ZN(n7477) );
  NAND2_X1 U6203 ( .A1(n6160), .A2(n5013), .ZN(n5167) );
  NAND2_X1 U6204 ( .A1(n7815), .A2(n8341), .ZN(n6164) );
  NAND2_X1 U6205 ( .A1(n4959), .A2(n10641), .ZN(n5158) );
  NOR2_X1 U6206 ( .A1(n9037), .A2(n5155), .ZN(n9103) );
  INV_X1 U6207 ( .A(n5433), .ZN(n7552) );
  INV_X1 U6208 ( .A(n8939), .ZN(n5058) );
  NAND2_X1 U6209 ( .A1(n8954), .A2(n6169), .ZN(n8955) );
  INV_X1 U6210 ( .A(n5168), .ZN(n8853) );
  INV_X1 U6211 ( .A(n6154), .ZN(n5434) );
  OAI21_X1 U6212 ( .B1(n8866), .B2(n5424), .A(n5423), .ZN(n8841) );
  NOR2_X1 U6213 ( .A1(n6992), .A2(n6313), .ZN(n6991) );
  INV_X1 U6214 ( .A(n7574), .ZN(n5049) );
  NOR2_X1 U6215 ( .A1(n7813), .A2(n8762), .ZN(n8761) );
  NOR2_X1 U6216 ( .A1(n5053), .A2(n5229), .ZN(n6275) );
  XNOR2_X1 U6217 ( .A(n6275), .B(n6326), .ZN(n10486) );
  NOR2_X1 U6218 ( .A1(n5230), .A2(n10478), .ZN(n5053) );
  NOR2_X1 U6219 ( .A1(n6279), .A2(n6991), .ZN(n7159) );
  OAI22_X1 U6220 ( .A1(n8412), .A2(n8411), .B1(n8410), .B2(n8506), .ZN(n8422)
         );
  AOI211_X1 U6221 ( .C1(n10800), .C2(n8443), .A(n8442), .B(n8441), .ZN(n8452)
         );
  NAND3_X2 U6222 ( .A1(n5159), .A2(n4947), .A3(n4981), .ZN(n5692) );
  AOI21_X1 U6223 ( .B1(n8505), .B2(n8503), .A(n8502), .ZN(n8504) );
  OR2_X1 U6224 ( .A1(n10592), .A2(n10605), .ZN(n8388) );
  NAND2_X1 U6225 ( .A1(n5211), .A2(n5210), .ZN(n5209) );
  NAND3_X1 U6226 ( .A1(n8496), .A2(n6128), .A3(n5052), .ZN(n8505) );
  NAND2_X1 U6227 ( .A1(n5260), .A2(n5261), .ZN(n5925) );
  XNOR2_X1 U6228 ( .A(n5209), .B(n8515), .ZN(n8523) );
  NAND2_X1 U6229 ( .A1(n5212), .A2(n8966), .ZN(n5216) );
  AOI21_X1 U6230 ( .B1(n5206), .B2(n5012), .A(n5205), .ZN(n8495) );
  OAI21_X1 U6231 ( .B1(n8511), .B2(n8510), .A(n8512), .ZN(n5211) );
  OAI21_X1 U6232 ( .B1(n8482), .B2(n5208), .A(n5005), .ZN(n5207) );
  NAND2_X1 U6233 ( .A1(n10429), .A2(n6272), .ZN(n6273) );
  NAND2_X1 U6234 ( .A1(n10430), .A2(n10431), .ZN(n10429) );
  NAND2_X1 U6235 ( .A1(n8814), .A2(n8816), .ZN(n5456) );
  NAND2_X1 U6236 ( .A1(n8820), .A2(n8821), .ZN(n5233) );
  NAND2_X1 U6237 ( .A1(n5163), .A2(n5011), .ZN(n8898) );
  NAND2_X1 U6238 ( .A1(n8878), .A2(n6178), .ZN(n5169) );
  XNOR2_X1 U6239 ( .A(n6289), .B(n6303), .ZN(n8762) );
  NAND2_X1 U6240 ( .A1(n6282), .A2(n5447), .ZN(n5443) );
  INV_X1 U6241 ( .A(n5395), .ZN(n9456) );
  NAND2_X2 U6242 ( .A1(n9314), .A2(n9370), .ZN(n6725) );
  NAND2_X4 U6243 ( .A1(n5059), .A2(n6969), .ZN(n9314) );
  NAND2_X1 U6244 ( .A1(n6836), .A2(n6831), .ZN(n6807) );
  NAND2_X1 U6245 ( .A1(n7028), .A2(n5062), .ZN(n5060) );
  NAND2_X1 U6246 ( .A1(n5060), .A2(n5015), .ZN(n5061) );
  AOI21_X2 U6247 ( .B1(n5064), .B2(n5063), .A(n5061), .ZN(n7040) );
  AND2_X1 U6248 ( .A1(n6856), .A2(n7028), .ZN(n5063) );
  NAND2_X1 U6249 ( .A1(n9363), .A2(n5066), .ZN(n5065) );
  NAND2_X1 U6250 ( .A1(n5065), .A2(n5068), .ZN(n9292) );
  NAND2_X1 U6251 ( .A1(n5077), .A2(n5079), .ZN(n7429) );
  NAND2_X1 U6252 ( .A1(n7193), .A2(n5009), .ZN(n5077) );
  OAI21_X1 U6253 ( .B1(n9503), .B2(n5085), .A(n5087), .ZN(n9426) );
  AND2_X1 U6254 ( .A1(n5092), .A2(n5089), .ZN(n9227) );
  NAND2_X1 U6255 ( .A1(n6016), .A2(n5097), .ZN(n5096) );
  NAND3_X1 U6256 ( .A1(n5096), .A2(n5468), .A3(n5095), .ZN(n8915) );
  NAND2_X1 U6257 ( .A1(n8870), .A2(n5102), .ZN(n5101) );
  NAND2_X1 U6258 ( .A1(n6130), .A2(n5101), .ZN(n6131) );
  NAND3_X1 U6259 ( .A1(n6199), .A2(n6197), .A3(n6198), .ZN(n8831) );
  INV_X1 U6260 ( .A(n5114), .ZN(n9896) );
  AND2_X1 U6261 ( .A1(n9796), .A2(n5126), .ZN(n9764) );
  NAND2_X1 U6262 ( .A1(n9796), .A2(n5124), .ZN(n9738) );
  NAND2_X1 U6263 ( .A1(n9796), .A2(n9787), .ZN(n9781) );
  NAND3_X1 U6264 ( .A1(n5127), .A2(n10729), .A3(n4958), .ZN(n7630) );
  NAND2_X1 U6265 ( .A1(n8728), .A2(n5132), .ZN(n5129) );
  INV_X1 U6266 ( .A(n8752), .ZN(n5134) );
  NAND2_X1 U6267 ( .A1(n6681), .A2(n6244), .ZN(n10436) );
  OAI211_X1 U6268 ( .C1(n7156), .C2(n5138), .A(n5136), .B(n5023), .ZN(n7374)
         );
  NOR2_X1 U6269 ( .A1(n7374), .A2(n10725), .ZN(n7373) );
  OR2_X1 U6270 ( .A1(n7156), .A2(n7155), .ZN(n5142) );
  INV_X1 U6271 ( .A(n5142), .ZN(n7154) );
  INV_X1 U6272 ( .A(n5148), .ZN(n7571) );
  INV_X1 U6273 ( .A(n6256), .ZN(n5147) );
  INV_X1 U6274 ( .A(n5151), .ZN(n10456) );
  NAND2_X2 U6275 ( .A1(n5691), .A2(n5692), .ZN(n6358) );
  AND3_X1 U6276 ( .A1(n5162), .A2(n5161), .A3(n4952), .ZN(n5159) );
  AND2_X2 U6277 ( .A1(n5685), .A2(n5684), .ZN(n5161) );
  NAND2_X1 U6278 ( .A1(n6173), .A2(n5164), .ZN(n5163) );
  XNOR2_X1 U6279 ( .A(n5166), .B(n8914), .ZN(n8911) );
  NAND2_X2 U6280 ( .A1(n5169), .A2(n6179), .ZN(n8866) );
  NAND2_X1 U6281 ( .A1(n5172), .A2(n5173), .ZN(n8173) );
  NAND2_X1 U6282 ( .A1(n8170), .A2(n5174), .ZN(n5172) );
  AOI21_X1 U6283 ( .B1(n5178), .B2(n5176), .A(n5175), .ZN(n5174) );
  NAND3_X1 U6284 ( .A1(n8178), .A2(n8217), .A3(n8219), .ZN(n5183) );
  NAND3_X1 U6285 ( .A1(n5189), .A2(n8127), .A3(n5188), .ZN(n5187) );
  OAI21_X2 U6286 ( .B1(n5872), .B2(n5871), .A(n5597), .ZN(n5884) );
  NAND3_X1 U6287 ( .A1(n5207), .A2(n8869), .A3(n8487), .ZN(n5206) );
  OR2_X1 U6288 ( .A1(n8452), .A2(n5213), .ZN(n5215) );
  AND2_X1 U6289 ( .A1(n5215), .A2(n5214), .ZN(n8466) );
  AND2_X1 U6290 ( .A1(n8978), .A2(n8455), .ZN(n5223) );
  NAND2_X1 U6291 ( .A1(n5228), .A2(n5225), .ZN(n6677) );
  NAND2_X1 U6292 ( .A1(n5227), .A2(n5751), .ZN(n6676) );
  OAI21_X1 U6293 ( .B1(n10478), .B2(n4953), .A(n5022), .ZN(n5229) );
  INV_X1 U6294 ( .A(n5230), .ZN(n10448) );
  NAND4_X1 U6295 ( .A1(n5233), .A2(n8818), .A3(n4972), .A4(n8817), .ZN(n5232)
         );
  NAND3_X1 U6296 ( .A1(n5246), .A2(n5245), .A3(n5244), .ZN(n5243) );
  NAND2_X1 U6297 ( .A1(n6017), .A2(n5251), .ZN(n5249) );
  OAI21_X1 U6298 ( .B1(n6017), .B2(n5259), .A(n5637), .ZN(n6033) );
  NAND2_X1 U6299 ( .A1(n5884), .A2(n4950), .ZN(n5260) );
  OAI21_X1 U6300 ( .B1(n5884), .B2(n5268), .A(n5265), .ZN(n5911) );
  OR2_X1 U6301 ( .A1(n8228), .A2(n5269), .ZN(n5273) );
  OAI21_X1 U6302 ( .B1(n8184), .B2(n5272), .A(n5270), .ZN(n5269) );
  AOI21_X1 U6303 ( .B1(n8184), .B2(n8183), .A(n8231), .ZN(n8187) );
  AOI21_X1 U6304 ( .B1(n8285), .B2(n9671), .A(n6613), .ZN(n5274) );
  NOR2_X1 U6305 ( .A1(n5273), .A2(n8229), .ZN(n8301) );
  NAND2_X1 U6306 ( .A1(n6072), .A2(n5651), .ZN(n5280) );
  NAND2_X1 U6307 ( .A1(n5941), .A2(n5614), .ZN(n5286) );
  NAND2_X1 U6308 ( .A1(n5664), .A2(n5663), .ZN(n6112) );
  NOR2_X1 U6309 ( .A1(n6481), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5296) );
  NAND3_X1 U6310 ( .A1(n5301), .A2(n9698), .A3(n5300), .ZN(n5298) );
  NAND2_X1 U6311 ( .A1(n5301), .A2(n9698), .ZN(n5299) );
  NAND2_X1 U6312 ( .A1(n9696), .A2(n9845), .ZN(n5301) );
  NAND2_X1 U6313 ( .A1(n7323), .A2(n4966), .ZN(n5313) );
  OAI21_X1 U6314 ( .B1(n10753), .B2(n5318), .A(n5315), .ZN(n8191) );
  NAND2_X1 U6315 ( .A1(n6594), .A2(n6593), .ZN(n6596) );
  NAND2_X1 U6316 ( .A1(n6433), .A2(n6382), .ZN(n6437) );
  INV_X1 U6317 ( .A(n6061), .ZN(n5647) );
  NAND2_X1 U6318 ( .A1(n6776), .A2(n6777), .ZN(n6885) );
  INV_X4 U6319 ( .A(n7870), .ZN(n7874) );
  INV_X1 U6320 ( .A(n5335), .ZN(n5330) );
  AOI21_X1 U6321 ( .B1(n6907), .B2(n5333), .A(n5332), .ZN(n5331) );
  INV_X1 U6322 ( .A(n7015), .ZN(n5332) );
  INV_X1 U6323 ( .A(n6902), .ZN(n5334) );
  NAND2_X1 U6324 ( .A1(n6907), .A2(n6902), .ZN(n5335) );
  AND2_X1 U6325 ( .A1(n6020), .A2(n5684), .ZN(n6034) );
  INV_X1 U6326 ( .A(n5681), .ZN(n5942) );
  NAND2_X1 U6327 ( .A1(n8666), .A2(n5338), .ZN(n5337) );
  AOI21_X1 U6328 ( .B1(n8666), .B2(n8668), .A(n8667), .ZN(n8525) );
  OAI211_X1 U6329 ( .C1(n8666), .C2(n5339), .A(n5337), .B(n7880), .ZN(P2_U3160) );
  NAND2_X1 U6330 ( .A1(n5355), .A2(n6210), .ZN(n5354) );
  INV_X1 U6331 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5356) );
  OAI21_X1 U6332 ( .B1(n7837), .B2(n5021), .A(n4963), .ZN(n7849) );
  NAND2_X1 U6333 ( .A1(n7255), .A2(n5365), .ZN(n5364) );
  NAND2_X1 U6334 ( .A1(n7764), .A2(n7763), .ZN(n7767) );
  NAND2_X1 U6335 ( .A1(n5375), .A2(n5374), .ZN(n9258) );
  INV_X1 U6336 ( .A(n7202), .ZN(n5382) );
  NAND2_X1 U6337 ( .A1(n5383), .A2(n5384), .ZN(n9419) );
  NAND3_X1 U6338 ( .A1(n9490), .A2(n5563), .A3(n5388), .ZN(n5383) );
  INV_X1 U6339 ( .A(n5392), .ZN(n9342) );
  NAND2_X1 U6340 ( .A1(n5395), .A2(n9184), .ZN(n9192) );
  NAND2_X1 U6341 ( .A1(n5395), .A2(n5393), .ZN(n9350) );
  OR2_X2 U6342 ( .A1(n8778), .A2(n8777), .ZN(n5397) );
  NAND2_X1 U6343 ( .A1(n8808), .A2(n5040), .ZN(n5402) );
  OAI211_X1 U6344 ( .C1(n8808), .C2(n5403), .A(n5402), .B(n10492), .ZN(n6367)
         );
  NOR2_X1 U6345 ( .A1(n8808), .A2(n8807), .ZN(n8806) );
  XNOR2_X2 U6346 ( .A(n5408), .B(n8766), .ZN(n8760) );
  NAND2_X1 U6347 ( .A1(n6247), .A2(n10459), .ZN(n5412) );
  NAND2_X1 U6348 ( .A1(n5857), .A2(n5856), .ZN(n5413) );
  NAND2_X1 U6349 ( .A1(n5836), .A2(n5835), .ZN(n5414) );
  NAND2_X1 U6350 ( .A1(n6168), .A2(n5415), .ZN(n8954) );
  OR2_X1 U6351 ( .A1(n8866), .A2(n5421), .ZN(n5420) );
  NAND2_X1 U6352 ( .A1(n8398), .A2(n8404), .ZN(n8333) );
  NOR2_X2 U6353 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5780) );
  OAI21_X1 U6354 ( .B1(n6082), .B2(n5462), .A(n5460), .ZN(n8895) );
  INV_X1 U6355 ( .A(n5457), .ZN(n6110) );
  AOI21_X1 U6356 ( .B1(n6082), .B2(n5460), .A(n5458), .ZN(n5457) );
  NAND2_X1 U6357 ( .A1(n5483), .A2(n8485), .ZN(n8870) );
  NAND2_X1 U6358 ( .A1(n5483), .A2(n5481), .ZN(n8322) );
  NAND3_X1 U6359 ( .A1(n5491), .A2(n8498), .A3(n8508), .ZN(n5490) );
  OAI21_X1 U6360 ( .B1(n7345), .B2(n5497), .A(n5499), .ZN(n7398) );
  NAND3_X1 U6361 ( .A1(n5498), .A2(n7401), .A3(n5496), .ZN(n7504) );
  NAND2_X1 U6362 ( .A1(n5499), .A2(n5497), .ZN(n5496) );
  INV_X1 U6363 ( .A(n7361), .ZN(n5497) );
  NAND2_X1 U6364 ( .A1(n7345), .A2(n5499), .ZN(n5498) );
  NAND2_X1 U6365 ( .A1(n9838), .A2(n5503), .ZN(n5502) );
  NAND2_X1 U6366 ( .A1(n9939), .A2(n5014), .ZN(n5510) );
  NAND2_X1 U6367 ( .A1(n5510), .A2(n5511), .ZN(n9871) );
  NOR2_X1 U6368 ( .A1(n6412), .A2(n5525), .ZN(n6422) );
  INV_X1 U6369 ( .A(n6412), .ZN(n5524) );
  NAND3_X1 U6370 ( .A1(n5531), .A2(n5532), .A3(n4969), .ZN(n5529) );
  OAI21_X1 U6371 ( .B1(n9726), .B2(n5545), .A(n5543), .ZN(n9730) );
  NAND2_X1 U6372 ( .A1(n9726), .A2(n5548), .ZN(n5547) );
  NAND2_X1 U6373 ( .A1(n9726), .A2(n9725), .ZN(n9755) );
  NAND2_X1 U6374 ( .A1(n6476), .A2(n5552), .ZN(n5554) );
  NAND2_X1 U6375 ( .A1(n6128), .A2(n6127), .ZN(n6129) );
  NAND2_X1 U6376 ( .A1(n5785), .A2(n8373), .ZN(n7109) );
  INV_X1 U6377 ( .A(n9764), .ZN(n9740) );
  INV_X1 U6378 ( .A(n6797), .ZN(n6938) );
  NAND2_X1 U6379 ( .A1(n8373), .A2(n8374), .ZN(n8371) );
  OR2_X1 U6380 ( .A1(n8322), .A2(n6129), .ZN(n6130) );
  NAND4_X2 U6381 ( .A1(n5766), .A2(n5765), .A3(n5764), .A4(n5763), .ZN(n8709)
         );
  NAND4_X2 U6382 ( .A1(n5755), .A2(n5754), .A3(n5753), .A4(n5752), .ZN(n10591)
         );
  OR2_X1 U6383 ( .A1(n6102), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5787) );
  INV_X1 U6384 ( .A(n6798), .ZN(n10552) );
  OR2_X1 U6385 ( .A1(n8839), .A2(n8691), .ZN(n5555) );
  INV_X1 U6386 ( .A(n8840), .ZN(n6127) );
  NAND2_X1 U6387 ( .A1(n6035), .A2(n6034), .ZN(n5557) );
  AND2_X2 U6388 ( .A1(n6600), .A2(n10130), .ZN(n5558) );
  OR2_X1 U6389 ( .A1(n9488), .A2(n7778), .ZN(n5559) );
  AND2_X2 U6390 ( .A1(n6410), .A2(n7559), .ZN(P1_U3973) );
  INV_X1 U6391 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5686) );
  INV_X1 U6392 ( .A(n7381), .ZN(n6464) );
  AND2_X1 U6393 ( .A1(n5894), .A2(n5912), .ZN(n7381) );
  INV_X1 U6394 ( .A(n7165), .ZN(n6442) );
  AND2_X1 U6395 ( .A1(n5601), .A2(n5600), .ZN(n5561) );
  INV_X1 U6396 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5947) );
  INV_X1 U6397 ( .A(n9915), .ZN(n10762) );
  NAND2_X2 U6398 ( .A1(n9090), .A2(n6761), .ZN(n10650) );
  XOR2_X1 U6399 ( .A(n9249), .B(n9373), .Z(n5562) );
  AND4_X1 U6400 ( .A1(n5732), .A2(n5731), .A3(n5730), .A4(n5729), .ZN(n8854)
         );
  INV_X1 U6401 ( .A(n8854), .ZN(n8691) );
  INV_X1 U6402 ( .A(n5858), .ZN(n5873) );
  INV_X1 U6403 ( .A(n8328), .ZN(n6128) );
  OR2_X1 U6404 ( .A1(n9292), .A2(n9291), .ZN(n5563) );
  AND2_X2 U6405 ( .A1(n9091), .A2(n6758), .ZN(n10810) );
  AND2_X1 U6406 ( .A1(n8871), .A2(n8692), .ZN(n5564) );
  OR2_X1 U6407 ( .A1(n8871), .A2(n8692), .ZN(n5565) );
  NOR2_X1 U6408 ( .A1(n7851), .A2(n8551), .ZN(n5566) );
  AND2_X1 U6409 ( .A1(n7287), .A2(n10635), .ZN(n5567) );
  NAND2_X1 U6410 ( .A1(n6294), .A2(n7010), .ZN(n6297) );
  INV_X1 U6411 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5684) );
  OR4_X1 U6412 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6635) );
  NOR2_X1 U6413 ( .A1(n7165), .A2(n6311), .ZN(n6280) );
  INV_X1 U6414 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5687) );
  INV_X1 U6415 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n5642) );
  INV_X1 U6416 ( .A(n7658), .ZN(n7654) );
  INV_X1 U6417 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5876) );
  OAI21_X1 U6418 ( .B1(n7143), .B2(n8392), .A(n5842), .ZN(n5843) );
  INV_X1 U6419 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10144) );
  INV_X1 U6420 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7403) );
  INV_X1 U6421 ( .A(SI_27_), .ZN(n10256) );
  INV_X1 U6422 ( .A(SI_23_), .ZN(n10255) );
  INV_X1 U6423 ( .A(SI_17_), .ZN(n10251) );
  INV_X1 U6424 ( .A(SI_9_), .ZN(n10248) );
  NAND2_X1 U6425 ( .A1(n7768), .A2(n8641), .ZN(n7826) );
  INV_X1 U6426 ( .A(n8572), .ZN(n7831) );
  INV_X1 U6427 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10340) );
  OR2_X1 U6428 ( .A1(n5715), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5727) );
  OR2_X1 U6429 ( .A1(n6116), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U6430 ( .A1(n5702), .A2(n6076), .ZN(n6100) );
  NAND2_X1 U6431 ( .A1(n10146), .A2(n6053), .ZN(n6065) );
  OR2_X1 U6432 ( .A1(n5904), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U6433 ( .A1(n6212), .A2(n6446), .ZN(n7093) );
  INV_X1 U6434 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5695) );
  AND2_X1 U6435 ( .A1(n5889), .A2(n5888), .ZN(n5893) );
  NOR2_X1 U6436 ( .A1(n8017), .A2(n8005), .ZN(n8004) );
  INV_X1 U6437 ( .A(n7975), .ZN(n7965) );
  NAND2_X1 U6438 ( .A1(n7392), .A2(n5056), .ZN(n6943) );
  NOR2_X1 U6439 ( .A1(n7725), .A2(n7724), .ZN(n7786) );
  OR2_X1 U6440 ( .A1(n8015), .A2(n8014), .ZN(n8017) );
  OR2_X1 U6441 ( .A1(n7882), .A2(n7881), .ZN(n7883) );
  INV_X1 U6442 ( .A(SI_21_), .ZN(n10253) );
  INV_X1 U6443 ( .A(SI_18_), .ZN(n5635) );
  INV_X1 U6444 ( .A(SI_15_), .ZN(n10283) );
  INV_X1 U6445 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6568) );
  INV_X1 U6446 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5814) );
  INV_X1 U6447 ( .A(n8686), .ZN(n8660) );
  INV_X1 U6448 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5688) );
  INV_X1 U6449 ( .A(n6358), .ZN(n6264) );
  AND2_X1 U6450 ( .A1(n5727), .A2(n5705), .ZN(n8860) );
  INV_X1 U6451 ( .A(n8698), .ZN(n9002) );
  NOR2_X1 U6452 ( .A1(n7095), .A2(n7093), .ZN(n6370) );
  AND2_X1 U6453 ( .A1(n7550), .A2(n7549), .ZN(n8335) );
  INV_X1 U6454 ( .A(n10637), .ZN(n9003) );
  NOR2_X1 U6455 ( .A1(n9022), .A2(n6188), .ZN(n10634) );
  AND2_X1 U6456 ( .A1(n7967), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7957) );
  INV_X1 U6457 ( .A(n9927), .ZN(n9714) );
  INV_X1 U6458 ( .A(n9965), .ZN(n9707) );
  AND2_X1 U6459 ( .A1(n9199), .A2(n9198), .ZN(n9504) );
  INV_X1 U6460 ( .A(n9539), .ZN(n9498) );
  NAND2_X1 U6461 ( .A1(n6653), .A2(n10135), .ZN(n9542) );
  AND2_X1 U6462 ( .A1(n8223), .A2(n6650), .ZN(n10555) );
  INV_X1 U6463 ( .A(n9995), .ZN(n9742) );
  INV_X1 U6464 ( .A(n9552), .ZN(n9780) );
  INV_X1 U6465 ( .A(n10015), .ZN(n9815) );
  INV_X1 U6466 ( .A(n10024), .ZN(n9844) );
  NAND2_X1 U6467 ( .A1(n8069), .A2(n8068), .ZN(n8076) );
  AND2_X1 U6468 ( .A1(n8139), .A2(n8136), .ZN(n10755) );
  OR2_X1 U6469 ( .A1(n10135), .A2(n6805), .ZN(n9949) );
  OR2_X1 U6470 ( .A1(n10556), .A2(n6650), .ZN(n10765) );
  OR2_X1 U6471 ( .A1(n6812), .A2(n6613), .ZN(n7316) );
  INV_X1 U6472 ( .A(n8676), .ZN(n8624) );
  OR2_X1 U6473 ( .A1(n6119), .A2(n8824), .ZN(n8318) );
  OR2_X1 U6474 ( .A1(n6119), .A2(n8883), .ZN(n6121) );
  AND4_X1 U6475 ( .A1(n6043), .A2(n6042), .A3(n6041), .A4(n6040), .ZN(n8977)
         );
  AND2_X1 U6476 ( .A1(n9156), .A2(n6298), .ZN(n6497) );
  INV_X1 U6477 ( .A(n10506), .ZN(n10516) );
  NOR2_X1 U6478 ( .A1(n6261), .A2(n8759), .ZN(n8778) );
  INV_X1 U6479 ( .A(n10464), .ZN(n10519) );
  AND2_X1 U6480 ( .A1(n8425), .A2(n8423), .ZN(n8339) );
  AND2_X1 U6481 ( .A1(n8385), .A2(n8393), .ZN(n8331) );
  INV_X1 U6482 ( .A(n10650), .ZN(n10706) );
  NAND2_X1 U6483 ( .A1(n6376), .A2(n6375), .ZN(n6377) );
  INV_X1 U6484 ( .A(n6760), .ZN(n9090) );
  INV_X1 U6485 ( .A(n10643), .ZN(n10739) );
  INV_X1 U6486 ( .A(n10799), .ZN(n10747) );
  OR2_X1 U6487 ( .A1(n10634), .A2(n10739), .ZN(n10720) );
  AND2_X1 U6488 ( .A1(n6744), .A2(n6448), .ZN(n6758) );
  INV_X1 U6489 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6181) );
  AND2_X1 U6490 ( .A1(n7913), .A2(n7912), .ZN(n9749) );
  INV_X1 U6491 ( .A(n9543), .ZN(n9473) );
  INV_X1 U6492 ( .A(n7446), .ZN(n9546) );
  AND3_X1 U6493 ( .A1(n7901), .A2(n7900), .A3(n7899), .ZN(n9686) );
  OR2_X1 U6494 ( .A1(n6487), .A2(n6486), .ZN(n9669) );
  NOR2_X1 U6495 ( .A1(n6516), .A2(n8295), .ZN(n10538) );
  NAND2_X1 U6496 ( .A1(n8209), .A2(n9756), .ZN(n9778) );
  OAI21_X1 U6497 ( .B1(n10030), .B2(n9876), .A(n9720), .ZN(n9838) );
  INV_X1 U6498 ( .A(n9976), .ZN(n10777) );
  INV_X1 U6499 ( .A(n9949), .ZN(n10759) );
  INV_X1 U6500 ( .A(n7629), .ZN(n7400) );
  AOI21_X1 U6501 ( .B1(n6640), .B2(n6629), .A(n6628), .ZN(n6821) );
  NAND2_X1 U6502 ( .A1(n7629), .A2(n7316), .ZN(n10767) );
  INV_X1 U6503 ( .A(n10556), .ZN(n10566) );
  AND2_X1 U6504 ( .A1(n6575), .A2(n6697), .ZN(n7708) );
  OR2_X1 U6505 ( .A1(n7825), .A2(n6232), .ZN(n6744) );
  NAND2_X1 U6506 ( .A1(n6754), .A2(n6758), .ZN(n8676) );
  INV_X1 U6507 ( .A(n8673), .ZN(n8689) );
  INV_X1 U6508 ( .A(n8988), .ZN(n8697) );
  INV_X1 U6509 ( .A(n8641), .ZN(n8703) );
  OR2_X1 U6510 ( .A1(P2_U3150), .A2(n6266), .ZN(n10506) );
  OR2_X1 U6511 ( .A1(n6267), .A2(n8516), .ZN(n10496) );
  INV_X1 U6512 ( .A(n10492), .ZN(n10514) );
  INV_X1 U6513 ( .A(n10709), .ZN(n9017) );
  INV_X1 U6514 ( .A(n9015), .ZN(n8968) );
  NAND2_X1 U6515 ( .A1(n10806), .A2(n10747), .ZN(n9089) );
  INV_X1 U6516 ( .A(n8347), .ZN(n9125) );
  INV_X1 U6517 ( .A(n10810), .ZN(n10807) );
  AND2_X1 U6518 ( .A1(n7561), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6448) );
  INV_X1 U6519 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7314) );
  INV_X1 U6520 ( .A(n6308), .ZN(n8718) );
  INV_X1 U6521 ( .A(n6326), .ZN(n10498) );
  XNOR2_X1 U6522 ( .A(n6409), .B(n6408), .ZN(n7559) );
  AND2_X1 U6523 ( .A1(n6647), .A2(n7126), .ZN(n9543) );
  INV_X1 U6524 ( .A(n10552), .ZN(n9564) );
  NAND2_X1 U6525 ( .A1(n6513), .A2(n10139), .ZN(n10546) );
  AND2_X1 U6526 ( .A1(n7415), .A2(n7414), .ZN(n10696) );
  INV_X1 U6527 ( .A(n10781), .ZN(n9979) );
  NAND2_X2 U6528 ( .A1(n6830), .A2(n7126), .ZN(n10560) );
  NAND2_X1 U6529 ( .A1(n10770), .A2(n10619), .ZN(n10069) );
  INV_X1 U6530 ( .A(n10770), .ZN(n10768) );
  INV_X1 U6531 ( .A(n9917), .ZN(n10106) );
  INV_X1 U6532 ( .A(n9708), .ZN(n10123) );
  INV_X1 U6533 ( .A(n10774), .ZN(n10771) );
  AND2_X2 U6534 ( .A1(n6822), .A2(n6828), .ZN(n10774) );
  AND3_X1 U6535 ( .A1(n6969), .A2(P1_STATE_REG_SCAN_IN), .A3(n7559), .ZN(n6651) );
  XNOR2_X1 U6536 ( .A(n6475), .B(n6593), .ZN(n10135) );
  INV_X1 U6537 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6916) );
  INV_X1 U6538 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6467) );
  INV_X1 U6539 ( .A(SI_1_), .ZN(n5568) );
  AND2_X1 U6540 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U6541 ( .A1(n5617), .A2(n5569), .ZN(n6611) );
  AND2_X1 U6542 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U6543 ( .A1(n5056), .A2(n5570), .ZN(n5769) );
  NAND2_X1 U6544 ( .A1(n6611), .A2(n5769), .ZN(n5756) );
  NAND2_X1 U6545 ( .A1(n5757), .A2(n5756), .ZN(n5573) );
  NAND2_X1 U6546 ( .A1(n5571), .A2(SI_1_), .ZN(n5572) );
  NAND2_X1 U6547 ( .A1(n5573), .A2(n5572), .ZN(n5778) );
  INV_X1 U6548 ( .A(SI_2_), .ZN(n5574) );
  XNOR2_X1 U6549 ( .A(n5575), .B(n5574), .ZN(n5777) );
  NAND2_X1 U6550 ( .A1(n5778), .A2(n5777), .ZN(n5577) );
  NAND2_X1 U6551 ( .A1(n5575), .A2(SI_2_), .ZN(n5576) );
  NAND2_X1 U6552 ( .A1(n5577), .A2(n5576), .ZN(n5791) );
  MUX2_X1 U6553 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5617), .Z(n5579) );
  INV_X1 U6554 ( .A(SI_3_), .ZN(n5578) );
  XNOR2_X1 U6555 ( .A(n5579), .B(n5578), .ZN(n5792) );
  NAND2_X1 U6556 ( .A1(n5791), .A2(n5792), .ZN(n5581) );
  NAND2_X1 U6557 ( .A1(n5579), .A2(SI_3_), .ZN(n5580) );
  MUX2_X1 U6558 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5617), .Z(n5582) );
  INV_X1 U6559 ( .A(SI_4_), .ZN(n10195) );
  XNOR2_X1 U6560 ( .A(n5582), .B(n10195), .ZN(n5804) );
  NAND2_X1 U6561 ( .A1(n5803), .A2(n5804), .ZN(n5584) );
  NAND2_X1 U6562 ( .A1(n5582), .A2(SI_4_), .ZN(n5583) );
  NAND2_X1 U6563 ( .A1(n5584), .A2(n5583), .ZN(n5821) );
  MUX2_X1 U6564 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5057), .Z(n5585) );
  INV_X1 U6565 ( .A(SI_5_), .ZN(n10246) );
  XNOR2_X1 U6566 ( .A(n5585), .B(n10246), .ZN(n5822) );
  NAND2_X1 U6567 ( .A1(n5821), .A2(n5822), .ZN(n5587) );
  NAND2_X1 U6568 ( .A1(n5585), .A2(SI_5_), .ZN(n5586) );
  MUX2_X1 U6569 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5057), .Z(n5588) );
  INV_X1 U6570 ( .A(SI_6_), .ZN(n10151) );
  XNOR2_X1 U6571 ( .A(n5588), .B(n10151), .ZN(n5835) );
  NAND2_X1 U6572 ( .A1(n5588), .A2(SI_6_), .ZN(n5589) );
  MUX2_X1 U6573 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5057), .Z(n5591) );
  INV_X1 U6574 ( .A(SI_7_), .ZN(n5590) );
  XNOR2_X1 U6575 ( .A(n5591), .B(n5590), .ZN(n5856) );
  NAND2_X1 U6576 ( .A1(n5591), .A2(SI_7_), .ZN(n5592) );
  INV_X1 U6577 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6440) );
  INV_X1 U6578 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5593) );
  MUX2_X1 U6579 ( .A(n6440), .B(n5593), .S(n5057), .Z(n5594) );
  NAND2_X1 U6580 ( .A1(n5594), .A2(n10298), .ZN(n5597) );
  INV_X1 U6581 ( .A(n5594), .ZN(n5595) );
  NAND2_X1 U6582 ( .A1(n5595), .A2(SI_8_), .ZN(n5596) );
  NAND2_X1 U6583 ( .A1(n5597), .A2(n5596), .ZN(n5871) );
  MUX2_X1 U6584 ( .A(n6463), .B(n6467), .S(n5057), .Z(n5598) );
  NAND2_X1 U6585 ( .A1(n5598), .A2(n10248), .ZN(n5601) );
  INV_X1 U6586 ( .A(n5598), .ZN(n5599) );
  NAND2_X1 U6587 ( .A1(n5599), .A2(SI_9_), .ZN(n5600) );
  INV_X1 U6588 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5602) );
  MUX2_X1 U6589 ( .A(n6470), .B(n5602), .S(n5057), .Z(n5603) );
  XNOR2_X1 U6590 ( .A(n5603), .B(SI_10_), .ZN(n5898) );
  INV_X1 U6591 ( .A(n5603), .ZN(n5604) );
  INV_X1 U6592 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5605) );
  MUX2_X1 U6593 ( .A(n6493), .B(n5605), .S(n5057), .Z(n5606) );
  NAND2_X1 U6594 ( .A1(n5606), .A2(n10185), .ZN(n5609) );
  INV_X1 U6595 ( .A(n5606), .ZN(n5607) );
  NAND2_X1 U6596 ( .A1(n5607), .A2(SI_11_), .ZN(n5608) );
  NAND2_X1 U6597 ( .A1(n5609), .A2(n5608), .ZN(n5910) );
  MUX2_X1 U6598 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n5057), .Z(n5611) );
  INV_X1 U6599 ( .A(SI_12_), .ZN(n5610) );
  XNOR2_X1 U6600 ( .A(n5611), .B(n5610), .ZN(n5924) );
  INV_X1 U6601 ( .A(n5924), .ZN(n5613) );
  NAND2_X1 U6602 ( .A1(n5611), .A2(SI_12_), .ZN(n5612) );
  MUX2_X1 U6603 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5057), .Z(n5615) );
  XNOR2_X1 U6604 ( .A(n5615), .B(SI_13_), .ZN(n5940) );
  INV_X1 U6605 ( .A(n5940), .ZN(n5614) );
  NAND2_X1 U6606 ( .A1(n5615), .A2(SI_13_), .ZN(n5616) );
  MUX2_X1 U6607 ( .A(n6694), .B(n5618), .S(n5057), .Z(n5619) );
  NAND2_X1 U6608 ( .A1(n5619), .A2(n10286), .ZN(n5622) );
  INV_X1 U6609 ( .A(n5619), .ZN(n5620) );
  NAND2_X1 U6610 ( .A1(n5620), .A2(SI_14_), .ZN(n5621) );
  NAND2_X1 U6611 ( .A1(n5622), .A2(n5621), .ZN(n5956) );
  MUX2_X1 U6612 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5057), .Z(n5623) );
  XNOR2_X1 U6613 ( .A(n5623), .B(n10283), .ZN(n5970) );
  INV_X1 U6614 ( .A(n5970), .ZN(n5625) );
  NAND2_X1 U6615 ( .A1(n5623), .A2(SI_15_), .ZN(n5624) );
  MUX2_X1 U6616 ( .A(n6899), .B(n6898), .S(n5057), .Z(n5626) );
  NAND2_X1 U6617 ( .A1(n5626), .A2(n10250), .ZN(n5629) );
  INV_X1 U6618 ( .A(n5626), .ZN(n5627) );
  NAND2_X1 U6619 ( .A1(n5627), .A2(SI_16_), .ZN(n5628) );
  NAND2_X1 U6620 ( .A1(n5629), .A2(n5628), .ZN(n5985) );
  MUX2_X1 U6621 ( .A(n6913), .B(n6916), .S(n5057), .Z(n5630) );
  NAND2_X1 U6622 ( .A1(n5630), .A2(n10251), .ZN(n5633) );
  INV_X1 U6623 ( .A(n5630), .ZN(n5631) );
  NAND2_X1 U6624 ( .A1(n5631), .A2(SI_17_), .ZN(n5632) );
  NAND2_X1 U6625 ( .A1(n6005), .A2(n6004), .ZN(n5634) );
  NAND2_X2 U6626 ( .A1(n5634), .A2(n5633), .ZN(n6017) );
  MUX2_X1 U6627 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5057), .Z(n5636) );
  XNOR2_X1 U6628 ( .A(n5636), .B(n5635), .ZN(n6018) );
  NAND2_X1 U6629 ( .A1(n5636), .A2(SI_18_), .ZN(n5637) );
  MUX2_X1 U6630 ( .A(n7174), .B(n7173), .S(n5057), .Z(n5638) );
  NAND2_X1 U6631 ( .A1(n5638), .A2(n10277), .ZN(n5641) );
  INV_X1 U6632 ( .A(n5638), .ZN(n5639) );
  NAND2_X1 U6633 ( .A1(n5639), .A2(SI_19_), .ZN(n5640) );
  NAND2_X1 U6634 ( .A1(n5641), .A2(n5640), .ZN(n6032) );
  MUX2_X1 U6635 ( .A(n7314), .B(n5642), .S(n5057), .Z(n5643) );
  INV_X1 U6636 ( .A(SI_20_), .ZN(n10155) );
  NAND2_X1 U6637 ( .A1(n5643), .A2(n10155), .ZN(n5646) );
  INV_X1 U6638 ( .A(n5643), .ZN(n5644) );
  NAND2_X1 U6639 ( .A1(n5644), .A2(SI_20_), .ZN(n5645) );
  MUX2_X1 U6640 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5057), .Z(n5648) );
  XNOR2_X1 U6641 ( .A(n5648), .B(n10253), .ZN(n6060) );
  NAND2_X1 U6642 ( .A1(n5647), .A2(n6060), .ZN(n5650) );
  NAND2_X1 U6643 ( .A1(n5648), .A2(SI_21_), .ZN(n5649) );
  NAND2_X1 U6644 ( .A1(n5650), .A2(n5649), .ZN(n6072) );
  MUX2_X1 U6645 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n5057), .Z(n5652) );
  XNOR2_X1 U6646 ( .A(n5652), .B(SI_22_), .ZN(n6071) );
  INV_X1 U6647 ( .A(n6071), .ZN(n5651) );
  NAND2_X1 U6648 ( .A1(n5652), .A2(SI_22_), .ZN(n5653) );
  INV_X1 U6649 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5655) );
  INV_X1 U6650 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5654) );
  MUX2_X1 U6651 ( .A(n5655), .B(n5654), .S(n5057), .Z(n5656) );
  NAND2_X1 U6652 ( .A1(n5656), .A2(n10255), .ZN(n5659) );
  INV_X1 U6653 ( .A(n5656), .ZN(n5657) );
  NAND2_X1 U6654 ( .A1(n5657), .A2(SI_23_), .ZN(n5658) );
  NAND2_X1 U6655 ( .A1(n5659), .A2(n5658), .ZN(n6083) );
  INV_X1 U6656 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7697) );
  INV_X1 U6657 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7701) );
  MUX2_X1 U6658 ( .A(n7697), .B(n7701), .S(n5057), .Z(n5660) );
  INV_X1 U6659 ( .A(SI_24_), .ZN(n10163) );
  NAND2_X1 U6660 ( .A1(n5660), .A2(n10163), .ZN(n5663) );
  INV_X1 U6661 ( .A(n5660), .ZN(n5661) );
  NAND2_X1 U6662 ( .A1(n5661), .A2(SI_24_), .ZN(n5662) );
  NAND2_X1 U6663 ( .A1(n6097), .A2(n6096), .ZN(n5664) );
  INV_X1 U6664 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7740) );
  INV_X1 U6665 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7742) );
  MUX2_X1 U6666 ( .A(n7740), .B(n7742), .S(n5057), .Z(n5666) );
  XNOR2_X1 U6667 ( .A(n5666), .B(SI_25_), .ZN(n6111) );
  INV_X1 U6668 ( .A(n6111), .ZN(n5665) );
  INV_X1 U6669 ( .A(n5666), .ZN(n5667) );
  NAND2_X1 U6670 ( .A1(n5667), .A2(SI_25_), .ZN(n5668) );
  INV_X1 U6671 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7823) );
  INV_X1 U6672 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7822) );
  MUX2_X1 U6673 ( .A(n7823), .B(n7822), .S(n5057), .Z(n5669) );
  INV_X1 U6674 ( .A(SI_26_), .ZN(n10165) );
  NAND2_X1 U6675 ( .A1(n5669), .A2(n10165), .ZN(n5672) );
  INV_X1 U6676 ( .A(n5669), .ZN(n5670) );
  NAND2_X1 U6677 ( .A1(n5670), .A2(SI_26_), .ZN(n5671) );
  NAND2_X1 U6678 ( .A1(n5672), .A2(n5671), .ZN(n5711) );
  INV_X1 U6679 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5673) );
  INV_X1 U6680 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10136) );
  MUX2_X1 U6681 ( .A(n5673), .B(n10136), .S(n5057), .Z(n5674) );
  NAND2_X1 U6682 ( .A1(n5674), .A2(n10256), .ZN(n5722) );
  INV_X1 U6683 ( .A(n5674), .ZN(n5675) );
  NAND2_X1 U6684 ( .A1(n5675), .A2(SI_27_), .ZN(n5676) );
  XNOR2_X1 U6685 ( .A(n5721), .B(n5720), .ZN(n9158) );
  NOR2_X1 U6686 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5678) );
  MUX2_X1 U6687 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5690), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5691) );
  NAND2_X1 U6688 ( .A1(n9158), .A2(n6113), .ZN(n5694) );
  NAND2_X1 U6689 ( .A1(n8307), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5693) );
  NOR2_X2 U6690 ( .A1(n5692), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U6691 ( .A1(n5698), .A2(n5695), .ZN(n9146) );
  XNOR2_X2 U6692 ( .A(n5697), .B(n5696), .ZN(n5700) );
  NAND2_X2 U6693 ( .A1(n5700), .A2(n9154), .ZN(n8312) );
  INV_X2 U6694 ( .A(n8312), .ZN(n5771) );
  NAND2_X1 U6695 ( .A1(n6089), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5709) );
  AND2_X4 U6696 ( .A1(n5700), .A2(n5701), .ZN(n8310) );
  INV_X1 U6697 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9039) );
  OR2_X1 U6698 ( .A1(n5828), .A2(n9039), .ZN(n5708) );
  NAND2_X1 U6699 ( .A1(n9149), .A2(n5701), .ZN(n5772) );
  INV_X1 U6700 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5702) );
  INV_X1 U6701 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10235) );
  INV_X1 U6702 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10146) );
  NOR2_X1 U6703 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5813) );
  NAND2_X1 U6704 ( .A1(n5813), .A2(n5814), .ZN(n5829) );
  NAND2_X1 U6705 ( .A1(n5948), .A2(n5947), .ZN(n5961) );
  NAND2_X1 U6706 ( .A1(n10340), .A2(n5995), .ZN(n6010) );
  NAND2_X1 U6707 ( .A1(n10235), .A2(n6075), .ZN(n6090) );
  INV_X1 U6708 ( .A(n6100), .ZN(n5703) );
  INV_X1 U6709 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10346) );
  NAND2_X1 U6710 ( .A1(n5703), .A2(n10346), .ZN(n6116) );
  INV_X1 U6711 ( .A(n6118), .ZN(n5704) );
  INV_X1 U6712 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10364) );
  NAND2_X1 U6713 ( .A1(n5704), .A2(n10364), .ZN(n5715) );
  NAND2_X1 U6714 ( .A1(n5715), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5705) );
  OR2_X2 U6715 ( .A1(n6119), .A2(n8860), .ZN(n5707) );
  INV_X1 U6716 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8861) );
  OR2_X1 U6717 ( .A1(n8314), .A2(n8861), .ZN(n5706) );
  NAND2_X1 U6718 ( .A1(n8859), .A2(n8868), .ZN(n8490) );
  XNOR2_X1 U6719 ( .A(n5710), .B(n5711), .ZN(n7925) );
  NAND2_X1 U6720 ( .A1(n7925), .A2(n6113), .ZN(n5713) );
  NAND2_X1 U6721 ( .A1(n8307), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U6722 ( .A1(n6089), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5719) );
  INV_X1 U6723 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9043) );
  OR2_X1 U6724 ( .A1(n5828), .A2(n9043), .ZN(n5718) );
  NAND2_X1 U6725 ( .A1(n6118), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5714) );
  AND2_X1 U6726 ( .A1(n5715), .A2(n5714), .ZN(n8872) );
  OR2_X1 U6727 ( .A1(n6102), .A2(n8872), .ZN(n5717) );
  INV_X1 U6728 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8873) );
  OR2_X1 U6729 ( .A1(n8314), .A2(n8873), .ZN(n5716) );
  NAND2_X1 U6730 ( .A1(n8871), .A2(n8880), .ZN(n8855) );
  NAND2_X1 U6731 ( .A1(n5721), .A2(n5720), .ZN(n5723) );
  MUX2_X1 U6732 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n5056), .Z(n5735) );
  INV_X1 U6733 ( .A(SI_28_), .ZN(n5736) );
  XNOR2_X1 U6734 ( .A(n5735), .B(n5736), .ZN(n5733) );
  NAND2_X1 U6735 ( .A1(n9155), .A2(n6113), .ZN(n5725) );
  NAND2_X1 U6736 ( .A1(n8307), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U6737 ( .A1(n8310), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5732) );
  INV_X1 U6738 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9100) );
  OR2_X1 U6739 ( .A1(n8312), .A2(n9100), .ZN(n5731) );
  INV_X1 U6740 ( .A(n5727), .ZN(n5726) );
  INV_X1 U6741 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10325) );
  NAND2_X1 U6742 ( .A1(n5726), .A2(n10325), .ZN(n8824) );
  NAND2_X1 U6743 ( .A1(n5727), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8848) );
  AND2_X1 U6744 ( .A1(n8824), .A2(n8848), .ZN(n7878) );
  OR2_X1 U6745 ( .A1(n6102), .A2(n7878), .ZN(n5730) );
  INV_X1 U6746 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5728) );
  OR2_X1 U6747 ( .A1(n8314), .A2(n5728), .ZN(n5729) );
  OR2_X2 U6748 ( .A1(n8859), .A2(n8868), .ZN(n8491) );
  NAND2_X1 U6749 ( .A1(n6126), .A2(n8491), .ZN(n6124) );
  NAND2_X1 U6750 ( .A1(n5734), .A2(n5733), .ZN(n5739) );
  INV_X1 U6751 ( .A(n5735), .ZN(n5737) );
  NAND2_X1 U6752 ( .A1(n5737), .A2(n5736), .ZN(n5738) );
  INV_X1 U6753 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10131) );
  INV_X1 U6754 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10370) );
  MUX2_X1 U6755 ( .A(n10131), .B(n10370), .S(n5056), .Z(n7881) );
  NAND2_X1 U6756 ( .A1(n9152), .A2(n6113), .ZN(n5741) );
  NAND2_X1 U6757 ( .A1(n8307), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U6758 ( .A1(n8310), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5745) );
  INV_X1 U6759 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5742) );
  OR2_X1 U6760 ( .A1(n8314), .A2(n5742), .ZN(n5744) );
  INV_X1 U6761 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6235) );
  OR2_X1 U6762 ( .A1(n8312), .A2(n6235), .ZN(n5743) );
  NAND4_X1 U6763 ( .A1(n8318), .A2(n5745), .A3(n5744), .A4(n5743), .ZN(n8844)
         );
  INV_X1 U6764 ( .A(n8844), .ZN(n5746) );
  NAND2_X1 U6765 ( .A1(n6234), .A2(n5746), .ZN(n8498) );
  NAND2_X1 U6766 ( .A1(n8839), .A2(n8854), .ZN(n6125) );
  OAI211_X1 U6767 ( .C1(n5025), .C2(n6124), .A(n8328), .B(n6125), .ZN(n6133)
         );
  OR2_X2 U6768 ( .A1(n8871), .A2(n8880), .ZN(n8488) );
  NAND2_X1 U6769 ( .A1(n8491), .A2(n8488), .ZN(n5747) );
  AND2_X1 U6770 ( .A1(n5747), .A2(n8490), .ZN(n8320) );
  INV_X1 U6771 ( .A(n6126), .ZN(n5749) );
  INV_X1 U6772 ( .A(n8499), .ZN(n5748) );
  NAND2_X1 U6773 ( .A1(n8323), .A2(n8498), .ZN(n6132) );
  INV_X1 U6774 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6795) );
  OR2_X1 U6775 ( .A1(n5772), .A2(n6795), .ZN(n5755) );
  INV_X1 U6776 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5750) );
  OR2_X1 U6777 ( .A1(n8312), .A2(n5750), .ZN(n5754) );
  NAND2_X1 U6778 ( .A1(n8310), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5753) );
  INV_X1 U6779 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5751) );
  XNOR2_X1 U6780 ( .A(n5757), .B(n5756), .ZN(n6716) );
  NAND2_X1 U6781 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5758) );
  MUX2_X1 U6782 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5758), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5760) );
  INV_X1 U6783 ( .A(n6268), .ZN(n5759) );
  OAI211_X2 U6784 ( .C1(n5858), .C2(n6716), .A(n5762), .B(n5761), .ZN(n7138)
         );
  OR2_X2 U6785 ( .A1(n10591), .A2(n10571), .ZN(n8365) );
  NAND2_X1 U6786 ( .A1(n10591), .A2(n10571), .ZN(n8367) );
  INV_X1 U6787 ( .A(n6138), .ZN(n7137) );
  NAND2_X1 U6788 ( .A1(n5771), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5766) );
  INV_X1 U6789 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6317) );
  OR2_X1 U6790 ( .A1(n5828), .A2(n6317), .ZN(n5765) );
  INV_X1 U6791 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6318) );
  OR2_X1 U6792 ( .A1(n5786), .A2(n6318), .ZN(n5764) );
  INV_X1 U6793 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6765) );
  OR2_X1 U6794 ( .A1(n5772), .A2(n6765), .ZN(n5763) );
  NAND2_X1 U6795 ( .A1(n5056), .A2(SI_0_), .ZN(n5768) );
  INV_X1 U6796 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U6797 ( .A1(n5768), .A2(n5767), .ZN(n5770) );
  AND2_X1 U6798 ( .A1(n5770), .A2(n5769), .ZN(n9163) );
  MUX2_X1 U6799 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9163), .S(n6240), .Z(n9019) );
  INV_X1 U6800 ( .A(n8363), .ZN(n7136) );
  NAND2_X1 U6801 ( .A1(n7137), .A2(n7136), .ZN(n7135) );
  NAND2_X1 U6802 ( .A1(n7135), .A2(n8365), .ZN(n10585) );
  NAND2_X1 U6803 ( .A1(n5771), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5776) );
  INV_X1 U6804 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6245) );
  OR2_X1 U6805 ( .A1(n5828), .A2(n6245), .ZN(n5775) );
  INV_X1 U6806 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6271) );
  OR2_X1 U6807 ( .A1(n5786), .A2(n6271), .ZN(n5774) );
  INV_X1 U6808 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10597) );
  OR2_X1 U6809 ( .A1(n5772), .A2(n10597), .ZN(n5773) );
  XNOR2_X1 U6810 ( .A(n5778), .B(n5777), .ZN(n6843) );
  NAND2_X1 U6811 ( .A1(n5779), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5784) );
  INV_X1 U6812 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U6813 ( .A1(n6036), .A2(n10433), .ZN(n5783) );
  OAI211_X1 U6814 ( .C1(n5858), .C2(n6843), .A(n5784), .B(n5783), .ZN(n6770)
         );
  INV_X1 U6815 ( .A(n6770), .ZN(n10599) );
  OR2_X1 U6816 ( .A1(n8708), .A2(n10599), .ZN(n8373) );
  NAND2_X1 U6817 ( .A1(n8708), .A2(n10599), .ZN(n8374) );
  NAND2_X1 U6818 ( .A1(n10585), .A2(n10587), .ZN(n5785) );
  NAND2_X1 U6819 ( .A1(n5771), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5790) );
  INV_X1 U6820 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6315) );
  OR2_X1 U6821 ( .A1(n5828), .A2(n6315), .ZN(n5789) );
  INV_X1 U6822 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6316) );
  OR2_X1 U6823 ( .A1(n5786), .A2(n6316), .ZN(n5788) );
  XNOR2_X1 U6824 ( .A(n5791), .B(n5792), .ZN(n6942) );
  NAND2_X1 U6825 ( .A1(n5779), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U6826 ( .A1(n6036), .A2(n6323), .ZN(n5793) );
  OAI211_X1 U6827 ( .C1(n5858), .C2(n6942), .A(n5794), .B(n5793), .ZN(n6886)
         );
  INV_X1 U6828 ( .A(n6886), .ZN(n10605) );
  NAND2_X1 U6829 ( .A1(n10592), .A2(n10605), .ZN(n8382) );
  NAND2_X1 U6830 ( .A1(n7109), .A2(n8329), .ZN(n5795) );
  NAND2_X1 U6831 ( .A1(n5795), .A2(n8388), .ZN(n7090) );
  NAND2_X1 U6832 ( .A1(n8310), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5802) );
  INV_X1 U6833 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5796) );
  AND2_X1 U6834 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5797) );
  NOR2_X1 U6835 ( .A1(n5813), .A2(n5797), .ZN(n7103) );
  OR2_X1 U6836 ( .A1(n6102), .A2(n7103), .ZN(n5800) );
  INV_X1 U6837 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5798) );
  OR2_X1 U6838 ( .A1(n8312), .A2(n5798), .ZN(n5799) );
  XNOR2_X1 U6839 ( .A(n5803), .B(n5804), .ZN(n7030) );
  NAND2_X1 U6840 ( .A1(n8307), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5810) );
  INV_X1 U6841 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U6842 ( .A1(n5806), .A2(n5805), .ZN(n5808) );
  XNOR2_X2 U6843 ( .A(n5824), .B(n5823), .ZN(n10471) );
  INV_X1 U6844 ( .A(n10471), .ZN(n6325) );
  NAND2_X1 U6845 ( .A1(n6036), .A2(n6325), .ZN(n5809) );
  OAI211_X1 U6846 ( .C1(n5858), .C2(n7030), .A(n5810), .B(n5809), .ZN(n6904)
         );
  NAND2_X1 U6847 ( .A1(n10636), .A2(n6904), .ZN(n10628) );
  OR2_X1 U6848 ( .A1(n10636), .A2(n6904), .ZN(n5811) );
  NAND2_X1 U6849 ( .A1(n10628), .A2(n5811), .ZN(n8377) );
  NAND2_X1 U6850 ( .A1(n7090), .A2(n8377), .ZN(n7143) );
  NAND2_X1 U6851 ( .A1(n6089), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5820) );
  INV_X1 U6852 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5812) );
  OR2_X1 U6853 ( .A1(n5828), .A2(n5812), .ZN(n5819) );
  OR2_X1 U6854 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  AND2_X1 U6855 ( .A1(n5829), .A2(n5815), .ZN(n10651) );
  OR2_X1 U6856 ( .A1(n6119), .A2(n10651), .ZN(n5818) );
  INV_X1 U6857 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5816) );
  OR2_X1 U6858 ( .A1(n8314), .A2(n5816), .ZN(n5817) );
  NAND4_X1 U6859 ( .A1(n5820), .A2(n5819), .A3(n5818), .A4(n5817), .ZN(n8707)
         );
  XNOR2_X1 U6860 ( .A(n5821), .B(n5822), .ZN(n7194) );
  NAND2_X1 U6861 ( .A1(n8307), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U6862 ( .A1(n5824), .A2(n5823), .ZN(n5825) );
  NAND2_X1 U6863 ( .A1(n5825), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5838) );
  XNOR2_X1 U6864 ( .A(n5838), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U6865 ( .A1(n6036), .A2(n6326), .ZN(n5826) );
  OAI211_X1 U6866 ( .C1(n5858), .C2(n7194), .A(n5827), .B(n5826), .ZN(n7013)
         );
  INV_X1 U6867 ( .A(n7013), .ZN(n10652) );
  NAND2_X1 U6868 ( .A1(n8707), .A2(n10652), .ZN(n8384) );
  INV_X1 U6869 ( .A(n8384), .ZN(n8392) );
  INV_X1 U6870 ( .A(n6904), .ZN(n10612) );
  NOR2_X1 U6871 ( .A1(n10636), .A2(n10612), .ZN(n8380) );
  OR2_X1 U6872 ( .A1(n8707), .A2(n10652), .ZN(n7145) );
  NAND2_X1 U6873 ( .A1(n5771), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5834) );
  INV_X1 U6874 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6314) );
  OR2_X1 U6875 ( .A1(n5828), .A2(n6314), .ZN(n5833) );
  NAND2_X1 U6876 ( .A1(n5829), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5830) );
  AND2_X1 U6877 ( .A1(n5844), .A2(n5830), .ZN(n7251) );
  OR2_X1 U6878 ( .A1(n6102), .A2(n7251), .ZN(n5832) );
  INV_X1 U6879 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7151) );
  OR2_X1 U6880 ( .A1(n8314), .A2(n7151), .ZN(n5831) );
  NAND4_X1 U6881 ( .A1(n5834), .A2(n5833), .A3(n5832), .A4(n5831), .ZN(n10635)
         );
  XNOR2_X1 U6882 ( .A(n5836), .B(n5835), .ZN(n7222) );
  NAND2_X1 U6883 ( .A1(n8307), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5841) );
  INV_X1 U6884 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U6885 ( .A1(n5838), .A2(n5837), .ZN(n5839) );
  NAND2_X1 U6886 ( .A1(n5839), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5851) );
  XNOR2_X1 U6887 ( .A(n5851), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U6888 ( .A1(n6036), .A2(n6329), .ZN(n5840) );
  OAI211_X1 U6889 ( .C1(n5858), .C2(n7222), .A(n5841), .B(n5840), .ZN(n7260)
         );
  INV_X1 U6890 ( .A(n7260), .ZN(n10668) );
  OR2_X1 U6891 ( .A1(n10635), .A2(n10668), .ZN(n8385) );
  NAND2_X1 U6892 ( .A1(n7145), .A2(n8385), .ZN(n8394) );
  AOI21_X1 U6893 ( .B1(n8380), .B2(n8384), .A(n8394), .ZN(n5842) );
  NAND2_X1 U6894 ( .A1(n10635), .A2(n10668), .ZN(n8393) );
  NAND2_X1 U6895 ( .A1(n5843), .A2(n8393), .ZN(n7309) );
  NAND2_X1 U6896 ( .A1(n6089), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5849) );
  INV_X1 U6897 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6312) );
  OR2_X1 U6898 ( .A1(n5828), .A2(n6312), .ZN(n5848) );
  AND2_X1 U6899 ( .A1(n5844), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5845) );
  NOR2_X1 U6900 ( .A1(n5862), .A2(n5845), .ZN(n7308) );
  OR2_X1 U6901 ( .A1(n6102), .A2(n7308), .ZN(n5847) );
  INV_X1 U6902 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6313) );
  OR2_X1 U6903 ( .A1(n8314), .A2(n6313), .ZN(n5846) );
  INV_X1 U6904 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6435) );
  INV_X1 U6905 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U6906 ( .A1(n5851), .A2(n5850), .ZN(n5852) );
  NAND2_X1 U6907 ( .A1(n5852), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U6908 ( .A1(n5854), .A2(n5853), .ZN(n5869) );
  OR2_X1 U6909 ( .A1(n5854), .A2(n5853), .ZN(n5855) );
  NAND2_X1 U6910 ( .A1(n6036), .A2(n6997), .ZN(n5860) );
  NAND2_X1 U6911 ( .A1(n7290), .A2(n10687), .ZN(n8405) );
  NAND2_X1 U6912 ( .A1(n7309), .A2(n8403), .ZN(n7466) );
  NAND2_X1 U6913 ( .A1(n5771), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5868) );
  INV_X1 U6914 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6310) );
  OR2_X1 U6915 ( .A1(n5828), .A2(n6310), .ZN(n5867) );
  NOR2_X1 U6916 ( .A1(n5862), .A2(n7164), .ZN(n5863) );
  OR2_X1 U6917 ( .A1(n5877), .A2(n5863), .ZN(n10707) );
  INV_X1 U6918 ( .A(n10707), .ZN(n5864) );
  OR2_X1 U6919 ( .A1(n6102), .A2(n5864), .ZN(n5866) );
  INV_X1 U6920 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6311) );
  OR2_X1 U6921 ( .A1(n8314), .A2(n6311), .ZN(n5865) );
  NAND4_X1 U6922 ( .A1(n5868), .A2(n5867), .A3(n5866), .A4(n5865), .ZN(n8705)
         );
  NAND2_X1 U6923 ( .A1(n5869), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U6924 ( .A1(n7395), .A2(n5873), .ZN(n5875) );
  NAND2_X1 U6925 ( .A1(n8307), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U6926 ( .A1(n8705), .A2(n7477), .ZN(n8398) );
  AND2_X1 U6927 ( .A1(n7465), .A2(n8398), .ZN(n8418) );
  NAND2_X1 U6928 ( .A1(n6089), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5883) );
  OR2_X1 U6929 ( .A1(n5828), .A2(n10725), .ZN(n5882) );
  OR2_X1 U6930 ( .A1(n5877), .A2(n5876), .ZN(n5878) );
  AND2_X1 U6931 ( .A1(n5904), .A2(n5878), .ZN(n7650) );
  OR2_X1 U6932 ( .A1(n6119), .A2(n7650), .ZN(n5881) );
  INV_X1 U6933 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5879) );
  OR2_X1 U6934 ( .A1(n8314), .A2(n5879), .ZN(n5880) );
  NAND4_X1 U6935 ( .A1(n5883), .A2(n5882), .A3(n5881), .A4(n5880), .ZN(n8704)
         );
  INV_X1 U6936 ( .A(n8704), .ZN(n7461) );
  XNOR2_X1 U6937 ( .A(n5884), .B(n5561), .ZN(n7483) );
  NAND2_X1 U6938 ( .A1(n7483), .A2(n6113), .ZN(n5896) );
  AND3_X1 U6939 ( .A1(n5887), .A2(n5886), .A3(n5885), .ZN(n5889) );
  NOR2_X1 U6940 ( .A1(n5893), .A2(n5807), .ZN(n5890) );
  MUX2_X1 U6941 ( .A(n5807), .B(n5890), .S(P2_IR_REG_9__SCAN_IN), .Z(n5891) );
  INV_X1 U6942 ( .A(n5891), .ZN(n5894) );
  NAND2_X1 U6943 ( .A1(n5893), .A2(n5892), .ZN(n5912) );
  AOI22_X1 U6944 ( .A1(n8307), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6036), .B2(
        n7381), .ZN(n5895) );
  NAND2_X1 U6945 ( .A1(n7461), .A2(n10724), .ZN(n8406) );
  INV_X1 U6946 ( .A(n10724), .ZN(n5897) );
  NAND2_X1 U6947 ( .A1(n5897), .A2(n8704), .ZN(n8417) );
  NAND2_X1 U6948 ( .A1(n8406), .A2(n8417), .ZN(n8334) );
  XNOR2_X1 U6949 ( .A(n5899), .B(n5898), .ZN(n7511) );
  NAND2_X1 U6950 ( .A1(n7511), .A2(n6113), .ZN(n5902) );
  NAND2_X1 U6951 ( .A1(n5912), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5900) );
  XNOR2_X1 U6952 ( .A(n5900), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7678) );
  AOI22_X1 U6953 ( .A1(n8307), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6036), .B2(
        n7678), .ZN(n5901) );
  NAND2_X1 U6954 ( .A1(n5902), .A2(n5901), .ZN(n10735) );
  NAND2_X1 U6955 ( .A1(n5771), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5909) );
  INV_X1 U6956 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5903) );
  OR2_X1 U6957 ( .A1(n5828), .A2(n5903), .ZN(n5908) );
  NAND2_X1 U6958 ( .A1(n5904), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5905) );
  AND2_X1 U6959 ( .A1(n5917), .A2(n5905), .ZN(n7774) );
  OR2_X1 U6960 ( .A1(n6102), .A2(n7774), .ZN(n5907) );
  INV_X1 U6961 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6283) );
  OR2_X1 U6962 ( .A1(n8314), .A2(n6283), .ZN(n5906) );
  NOR2_X1 U6963 ( .A1(n10735), .A2(n8641), .ZN(n8413) );
  NAND2_X1 U6964 ( .A1(n10735), .A2(n8641), .ZN(n8420) );
  XNOR2_X1 U6965 ( .A(n5911), .B(n5910), .ZN(n7610) );
  NAND2_X1 U6966 ( .A1(n7610), .A2(n6113), .ZN(n5915) );
  NAND2_X1 U6967 ( .A1(n5913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5927) );
  INV_X1 U6968 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5926) );
  XNOR2_X1 U6969 ( .A(n5927), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6344) );
  AOI22_X1 U6970 ( .A1(n8307), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6036), .B2(
        n6344), .ZN(n5914) );
  NAND2_X1 U6971 ( .A1(n5915), .A2(n5914), .ZN(n10746) );
  NAND2_X1 U6972 ( .A1(n6089), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5922) );
  INV_X1 U6973 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5916) );
  OR2_X1 U6974 ( .A1(n5828), .A2(n5916), .ZN(n5921) );
  INV_X1 U6975 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7567) );
  OR2_X1 U6976 ( .A1(n8314), .A2(n7567), .ZN(n5920) );
  NAND2_X1 U6977 ( .A1(n5917), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5918) );
  AND2_X1 U6978 ( .A1(n5933), .A2(n5918), .ZN(n8645) );
  OR2_X1 U6979 ( .A1(n6119), .A2(n8645), .ZN(n5919) );
  NAND4_X1 U6980 ( .A1(n5922), .A2(n5921), .A3(n5920), .A4(n5919), .ZN(n8702)
         );
  INV_X1 U6981 ( .A(n8702), .ZN(n7828) );
  OR2_X1 U6982 ( .A1(n10746), .A2(n7828), .ZN(n8425) );
  NAND2_X1 U6983 ( .A1(n10746), .A2(n7828), .ZN(n8423) );
  NAND2_X1 U6984 ( .A1(n7564), .A2(n8339), .ZN(n5923) );
  NAND2_X1 U6985 ( .A1(n5923), .A2(n8423), .ZN(n7595) );
  NAND2_X1 U6986 ( .A1(n7703), .A2(n6113), .ZN(n5931) );
  NAND2_X1 U6987 ( .A1(n5927), .A2(n5926), .ZN(n5928) );
  NAND2_X1 U6988 ( .A1(n5928), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5929) );
  XNOR2_X1 U6989 ( .A(n5929), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6308) );
  AOI22_X1 U6990 ( .A1(n8307), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6036), .B2(
        n6308), .ZN(n5930) );
  NAND2_X1 U6991 ( .A1(n5931), .A2(n5930), .ZN(n8575) );
  NAND2_X1 U6992 ( .A1(n5771), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5938) );
  INV_X1 U6993 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5932) );
  OR2_X1 U6994 ( .A1(n5828), .A2(n5932), .ZN(n5937) );
  AND2_X1 U6995 ( .A1(n5933), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5934) );
  NOR2_X1 U6996 ( .A1(n5948), .A2(n5934), .ZN(n8569) );
  OR2_X1 U6997 ( .A1(n6119), .A2(n8569), .ZN(n5936) );
  INV_X1 U6998 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6285) );
  OR2_X1 U6999 ( .A1(n8314), .A2(n6285), .ZN(n5935) );
  NAND4_X1 U7000 ( .A1(n5938), .A2(n5937), .A3(n5936), .A4(n5935), .ZN(n8701)
         );
  INV_X1 U7001 ( .A(n8701), .ZN(n8627) );
  OR2_X1 U7002 ( .A1(n8575), .A2(n8627), .ZN(n8429) );
  NAND2_X1 U7003 ( .A1(n7595), .A2(n8429), .ZN(n5939) );
  NAND2_X1 U7004 ( .A1(n8575), .A2(n8627), .ZN(n8430) );
  NAND2_X1 U7005 ( .A1(n5939), .A2(n8430), .ZN(n7681) );
  XNOR2_X1 U7006 ( .A(n5941), .B(n5940), .ZN(n7707) );
  NAND2_X1 U7007 ( .A1(n7707), .A2(n6113), .ZN(n5945) );
  NAND2_X1 U7008 ( .A1(n5942), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5943) );
  XNOR2_X1 U7009 ( .A(n5943), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6307) );
  AOI22_X1 U7010 ( .A1(n8307), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6036), .B2(
        n6307), .ZN(n5944) );
  NAND2_X1 U7011 ( .A1(n6089), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5954) );
  INV_X1 U7012 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5946) );
  OR2_X1 U7013 ( .A1(n5828), .A2(n5946), .ZN(n5953) );
  OR2_X1 U7014 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  AND2_X1 U7015 ( .A1(n5949), .A2(n5961), .ZN(n8628) );
  OR2_X1 U7016 ( .A1(n6119), .A2(n8628), .ZN(n5952) );
  INV_X1 U7017 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5950) );
  OR2_X1 U7018 ( .A1(n8314), .A2(n5950), .ZN(n5951) );
  XNOR2_X1 U7019 ( .A(n8361), .B(n8700), .ZN(n8432) );
  NAND2_X1 U7020 ( .A1(n8361), .A2(n8566), .ZN(n5955) );
  XNOR2_X1 U7021 ( .A(n5957), .B(n5956), .ZN(n7780) );
  NAND2_X1 U7022 ( .A1(n7780), .A2(n6113), .ZN(n5959) );
  NAND2_X1 U7023 ( .A1(n6019), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5973) );
  XNOR2_X1 U7024 ( .A(n5973), .B(n5972), .ZN(n8750) );
  INV_X1 U7025 ( .A(n8750), .ZN(n6305) );
  AOI22_X1 U7026 ( .A1(n8307), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6036), .B2(
        n6305), .ZN(n5958) );
  NAND2_X1 U7027 ( .A1(n5771), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5967) );
  INV_X1 U7028 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5960) );
  OR2_X1 U7029 ( .A1(n5828), .A2(n5960), .ZN(n5966) );
  NAND2_X1 U7030 ( .A1(n5961), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5962) );
  AND2_X1 U7031 ( .A1(n5978), .A2(n5962), .ZN(n8538) );
  OR2_X1 U7032 ( .A1(n6119), .A2(n8538), .ZN(n5965) );
  INV_X1 U7033 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5963) );
  OR2_X1 U7034 ( .A1(n8314), .A2(n5963), .ZN(n5964) );
  NAND4_X1 U7035 ( .A1(n5967), .A2(n5966), .A3(n5965), .A4(n5964), .ZN(n8699)
         );
  NOR2_X1 U7036 ( .A1(n8357), .A2(n8699), .ZN(n6163) );
  INV_X1 U7037 ( .A(n6163), .ZN(n5968) );
  NAND2_X1 U7038 ( .A1(n8357), .A2(n8699), .ZN(n8444) );
  INV_X1 U7039 ( .A(n8699), .ZN(n8681) );
  OR2_X1 U7040 ( .A1(n8357), .A2(n8681), .ZN(n5969) );
  XNOR2_X1 U7041 ( .A(n5971), .B(n5970), .ZN(n8022) );
  NAND2_X1 U7042 ( .A1(n8022), .A2(n6113), .ZN(n5976) );
  NAND2_X1 U7043 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  NAND2_X1 U7044 ( .A1(n5974), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5988) );
  XNOR2_X1 U7045 ( .A(n5988), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6303) );
  AOI22_X1 U7046 ( .A1(n8307), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6036), .B2(
        n6303), .ZN(n5975) );
  NAND2_X1 U7047 ( .A1(n6089), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5983) );
  INV_X1 U7048 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5977) );
  OR2_X1 U7049 ( .A1(n5828), .A2(n5977), .ZN(n5982) );
  AND2_X1 U7050 ( .A1(n5978), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5979) );
  NOR2_X1 U7051 ( .A1(n5995), .A2(n5979), .ZN(n8682) );
  OR2_X1 U7052 ( .A1(n6119), .A2(n8682), .ZN(n5981) );
  INV_X1 U7053 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7813) );
  OR2_X1 U7054 ( .A1(n8314), .A2(n7813), .ZN(n5980) );
  NAND4_X1 U7055 ( .A1(n5983), .A2(n5982), .A3(n5981), .A4(n5980), .ZN(n8698)
         );
  NAND2_X1 U7056 ( .A1(n8356), .A2(n9002), .ZN(n9006) );
  OR2_X1 U7057 ( .A1(n8356), .A2(n9002), .ZN(n5984) );
  NAND2_X1 U7058 ( .A1(n9006), .A2(n5984), .ZN(n8341) );
  XNOR2_X1 U7059 ( .A(n5986), .B(n5985), .ZN(n8011) );
  NAND2_X1 U7060 ( .A1(n8011), .A2(n6113), .ZN(n5994) );
  INV_X1 U7061 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7062 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  NAND2_X1 U7063 ( .A1(n5989), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5991) );
  INV_X1 U7064 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7065 ( .A1(n5991), .A2(n5990), .ZN(n6006) );
  OR2_X1 U7066 ( .A1(n5991), .A2(n5990), .ZN(n5992) );
  AND2_X1 U7067 ( .A1(n6006), .A2(n5992), .ZN(n6301) );
  AOI22_X1 U7068 ( .A1(n8307), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6036), .B2(
        n6301), .ZN(n5993) );
  NAND2_X1 U7069 ( .A1(n6089), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6000) );
  INV_X1 U7070 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9087) );
  OR2_X1 U7071 ( .A1(n5828), .A2(n9087), .ZN(n5999) );
  OR2_X1 U7072 ( .A1(n5995), .A2(n10340), .ZN(n5996) );
  AND2_X1 U7073 ( .A1(n5996), .A2(n6010), .ZN(n9011) );
  OR2_X1 U7074 ( .A1(n6119), .A2(n9011), .ZN(n5998) );
  INV_X1 U7075 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9012) );
  OR2_X1 U7076 ( .A1(n8314), .A2(n9012), .ZN(n5997) );
  NAND2_X1 U7077 ( .A1(n9010), .A2(n8988), .ZN(n8449) );
  NAND2_X1 U7078 ( .A1(n8448), .A2(n8449), .ZN(n8998) );
  INV_X1 U7079 ( .A(n9006), .ZN(n6001) );
  NOR2_X1 U7080 ( .A1(n8998), .A2(n6001), .ZN(n6002) );
  NAND2_X1 U7081 ( .A1(n6003), .A2(n8448), .ZN(n8991) );
  XNOR2_X1 U7082 ( .A(n6005), .B(n6004), .ZN(n8001) );
  NAND2_X1 U7083 ( .A1(n8001), .A2(n6113), .ZN(n6009) );
  NAND2_X1 U7084 ( .A1(n6006), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6007) );
  XNOR2_X1 U7085 ( .A(n6007), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6353) );
  AOI22_X1 U7086 ( .A1(n8307), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6036), .B2(
        n6353), .ZN(n6008) );
  NAND2_X1 U7087 ( .A1(n5771), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6014) );
  INV_X1 U7088 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9083) );
  OR2_X1 U7089 ( .A1(n5828), .A2(n9083), .ZN(n6013) );
  INV_X1 U7090 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8993) );
  OR2_X1 U7091 ( .A1(n8314), .A2(n8993), .ZN(n6012) );
  AOI21_X1 U7092 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(n6010), .A(n6025), .ZN(
        n8992) );
  OR2_X1 U7093 ( .A1(n6119), .A2(n8992), .ZN(n6011) );
  NAND4_X1 U7094 ( .A1(n6014), .A2(n6013), .A3(n6012), .A4(n6011), .ZN(n8696)
         );
  XNOR2_X1 U7095 ( .A(n8599), .B(n9004), .ZN(n8990) );
  INV_X1 U7096 ( .A(n8990), .ZN(n8344) );
  NAND2_X1 U7097 ( .A1(n8991), .A2(n8344), .ZN(n6016) );
  OR2_X1 U7098 ( .A1(n8599), .A2(n9004), .ZN(n6015) );
  INV_X1 U7099 ( .A(n6019), .ZN(n6035) );
  NAND2_X1 U7100 ( .A1(n6035), .A2(n6020), .ZN(n6021) );
  NAND2_X1 U7101 ( .A1(n6021), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6022) );
  XNOR2_X1 U7102 ( .A(n6022), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8821) );
  AOI22_X1 U7103 ( .A1(n8307), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6036), .B2(
        n8821), .ZN(n6023) );
  NAND2_X2 U7104 ( .A1(n6024), .A2(n6023), .ZN(n8655) );
  NAND2_X1 U7105 ( .A1(n8310), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6031) );
  INV_X1 U7106 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8981) );
  OR2_X1 U7107 ( .A1(n8314), .A2(n8981), .ZN(n6030) );
  INV_X1 U7108 ( .A(n6025), .ZN(n6027) );
  INV_X1 U7109 ( .A(n6039), .ZN(n6026) );
  AOI21_X1 U7110 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(n6027), .A(n6026), .ZN(
        n8980) );
  OR2_X1 U7111 ( .A1(n6102), .A2(n8980), .ZN(n6029) );
  INV_X1 U7112 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9133) );
  OR2_X1 U7113 ( .A1(n8312), .A2(n9133), .ZN(n6028) );
  NAND4_X1 U7114 ( .A1(n6031), .A2(n6030), .A3(n6029), .A4(n6028), .ZN(n8958)
         );
  NAND2_X1 U7115 ( .A1(n8655), .A2(n8989), .ZN(n8456) );
  XNOR2_X1 U7116 ( .A(n6033), .B(n6032), .ZN(n7990) );
  NAND2_X1 U7117 ( .A1(n7990), .A2(n6113), .ZN(n6038) );
  AOI22_X1 U7118 ( .A1(n8307), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8515), .B2(
        n6036), .ZN(n6037) );
  NAND2_X1 U7119 ( .A1(n6038), .A2(n6037), .ZN(n8972) );
  NAND2_X1 U7120 ( .A1(n5771), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6043) );
  INV_X1 U7121 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9075) );
  OR2_X1 U7122 ( .A1(n5828), .A2(n9075), .ZN(n6042) );
  AOI21_X1 U7123 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(n6039), .A(n6053), .ZN(
        n8962) );
  OR2_X1 U7124 ( .A1(n6119), .A2(n8962), .ZN(n6041) );
  INV_X1 U7125 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8963) );
  OR2_X1 U7126 ( .A1(n8314), .A2(n8963), .ZN(n6040) );
  OR2_X1 U7127 ( .A1(n8972), .A2(n8977), .ZN(n6044) );
  AND2_X1 U7128 ( .A1(n8964), .A2(n6044), .ZN(n6047) );
  INV_X1 U7129 ( .A(n6044), .ZN(n8460) );
  NAND2_X1 U7130 ( .A1(n8972), .A2(n8977), .ZN(n8459) );
  NAND2_X1 U7131 ( .A1(n6044), .A2(n8459), .ZN(n8956) );
  INV_X1 U7132 ( .A(n8956), .ZN(n8966) );
  OR2_X1 U7133 ( .A1(n8460), .A2(n8966), .ZN(n6045) );
  INV_X1 U7134 ( .A(n6045), .ZN(n6046) );
  XNOR2_X1 U7135 ( .A(n6049), .B(n6048), .ZN(n7981) );
  NAND2_X1 U7136 ( .A1(n7981), .A2(n6113), .ZN(n6051) );
  NAND2_X1 U7137 ( .A1(n8307), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7138 ( .A1(n6089), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6059) );
  INV_X1 U7139 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n6052) );
  OR2_X1 U7140 ( .A1(n5828), .A2(n6052), .ZN(n6058) );
  INV_X1 U7141 ( .A(n6053), .ZN(n6055) );
  INV_X1 U7142 ( .A(n6065), .ZN(n6054) );
  AOI21_X1 U7143 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(n6055), .A(n6054), .ZN(
        n8947) );
  OR2_X1 U7144 ( .A1(n6102), .A2(n8947), .ZN(n6057) );
  INV_X1 U7145 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8948) );
  OR2_X1 U7146 ( .A1(n8314), .A2(n8948), .ZN(n6056) );
  NAND4_X1 U7147 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(n8959)
         );
  XNOR2_X1 U7148 ( .A(n8950), .B(n8959), .ZN(n8938) );
  INV_X1 U7149 ( .A(n8959), .ZN(n8554) );
  OR2_X1 U7150 ( .A1(n8950), .A2(n8554), .ZN(n8464) );
  XNOR2_X1 U7151 ( .A(n6061), .B(n6060), .ZN(n7972) );
  NAND2_X1 U7152 ( .A1(n7972), .A2(n6113), .ZN(n6063) );
  NAND2_X1 U7153 ( .A1(n8307), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7154 ( .A1(n5771), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6069) );
  INV_X1 U7155 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6064) );
  OR2_X1 U7156 ( .A1(n5828), .A2(n6064), .ZN(n6068) );
  AOI21_X1 U7157 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(n6065), .A(n6075), .ZN(
        n8930) );
  OR2_X1 U7158 ( .A1(n6119), .A2(n8930), .ZN(n6067) );
  INV_X1 U7159 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8931) );
  OR2_X1 U7160 ( .A1(n8314), .A2(n8931), .ZN(n6066) );
  NAND4_X1 U7161 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n8943)
         );
  INV_X1 U7162 ( .A(n8467), .ZN(n6070) );
  NAND2_X1 U7163 ( .A1(n9062), .A2(n8913), .ZN(n8468) );
  XNOR2_X1 U7164 ( .A(n6072), .B(n6071), .ZN(n7962) );
  NAND2_X1 U7165 ( .A1(n7962), .A2(n6113), .ZN(n6074) );
  NAND2_X1 U7166 ( .A1(n8307), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7167 ( .A1(n8310), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6081) );
  INV_X1 U7168 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8917) );
  OR2_X1 U7169 ( .A1(n8314), .A2(n8917), .ZN(n6080) );
  INV_X1 U7170 ( .A(n6075), .ZN(n6077) );
  AOI21_X1 U7171 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n6077), .A(n6076), .ZN(
        n8916) );
  OR2_X1 U7172 ( .A1(n6102), .A2(n8916), .ZN(n6079) );
  INV_X1 U7173 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9123) );
  OR2_X1 U7174 ( .A1(n8312), .A2(n9123), .ZN(n6078) );
  NAND4_X1 U7175 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6078), .ZN(n8927)
         );
  INV_X1 U7176 ( .A(n8927), .ZN(n8900) );
  OR2_X1 U7177 ( .A1(n8347), .A2(n8900), .ZN(n8471) );
  NAND2_X1 U7178 ( .A1(n8915), .A2(n8471), .ZN(n6082) );
  NAND2_X1 U7179 ( .A1(n8347), .A2(n8900), .ZN(n8472) );
  NAND2_X1 U7180 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  NAND2_X1 U7181 ( .A1(n6086), .A2(n6085), .ZN(n7953) );
  NAND2_X1 U7182 ( .A1(n7953), .A2(n6113), .ZN(n6088) );
  NAND2_X1 U7183 ( .A1(n8307), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7184 ( .A1(n6089), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6095) );
  INV_X1 U7185 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9056) );
  OR2_X1 U7186 ( .A1(n5828), .A2(n9056), .ZN(n6094) );
  NAND2_X1 U7187 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(n6090), .ZN(n6091) );
  AND2_X1 U7188 ( .A1(n6100), .A2(n6091), .ZN(n8905) );
  OR2_X1 U7189 ( .A1(n6119), .A2(n8905), .ZN(n6093) );
  INV_X1 U7190 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8906) );
  OR2_X1 U7191 ( .A1(n8314), .A2(n8906), .ZN(n6092) );
  NAND4_X1 U7192 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n8695)
         );
  OR2_X1 U7193 ( .A1(n8904), .A2(n8912), .ZN(n8477) );
  NAND2_X1 U7194 ( .A1(n8904), .A2(n8912), .ZN(n8476) );
  XNOR2_X1 U7195 ( .A(n6097), .B(n6096), .ZN(n7943) );
  NAND2_X1 U7196 ( .A1(n7943), .A2(n6113), .ZN(n6099) );
  NAND2_X1 U7197 ( .A1(n8307), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7198 ( .A1(n5771), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6107) );
  INV_X1 U7199 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9052) );
  OR2_X1 U7200 ( .A1(n5828), .A2(n9052), .ZN(n6106) );
  NAND2_X1 U7201 ( .A1(n6100), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6101) );
  AND2_X1 U7202 ( .A1(n6116), .A2(n6101), .ZN(n8892) );
  OR2_X1 U7203 ( .A1(n6102), .A2(n8892), .ZN(n6105) );
  INV_X1 U7204 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6103) );
  OR2_X1 U7205 ( .A1(n8314), .A2(n6103), .ZN(n6104) );
  NAND4_X1 U7206 ( .A1(n6107), .A2(n6106), .A3(n6105), .A4(n6104), .ZN(n8694)
         );
  OR2_X1 U7207 ( .A1(n8891), .A2(n8901), .ZN(n6108) );
  NAND2_X1 U7208 ( .A1(n8891), .A2(n8901), .ZN(n6109) );
  NAND2_X1 U7209 ( .A1(n6110), .A2(n6109), .ZN(n8882) );
  XNOR2_X1 U7210 ( .A(n6112), .B(n6111), .ZN(n7934) );
  NAND2_X1 U7211 ( .A1(n7934), .A2(n6113), .ZN(n6115) );
  NAND2_X1 U7212 ( .A1(n8307), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7213 ( .A1(n5771), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6123) );
  INV_X1 U7214 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9048) );
  OR2_X1 U7215 ( .A1(n5828), .A2(n9048), .ZN(n6122) );
  NAND2_X1 U7216 ( .A1(n6116), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6117) );
  AND2_X1 U7217 ( .A1(n6118), .A2(n6117), .ZN(n8883) );
  INV_X1 U7218 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8884) );
  OR2_X1 U7219 ( .A1(n8314), .A2(n8884), .ZN(n6120) );
  NAND4_X1 U7220 ( .A1(n6123), .A2(n6122), .A3(n6121), .A4(n6120), .ZN(n8693)
         );
  OR2_X1 U7221 ( .A1(n9045), .A2(n8890), .ZN(n8486) );
  NAND2_X1 U7222 ( .A1(n9045), .A2(n8890), .ZN(n8485) );
  NAND2_X1 U7223 ( .A1(n6134), .A2(n5093), .ZN(n6135) );
  XNOR2_X2 U7224 ( .A(n6182), .B(n6181), .ZN(n8512) );
  NAND2_X1 U7225 ( .A1(n6136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6137) );
  OR2_X1 U7226 ( .A1(n7098), .A2(n8520), .ZN(n10643) );
  NAND2_X1 U7227 ( .A1(n8709), .A2(n9019), .ZN(n7131) );
  NAND2_X1 U7228 ( .A1(n6138), .A2(n7131), .ZN(n10588) );
  OR2_X1 U7229 ( .A1(n10591), .A2(n7138), .ZN(n10586) );
  NAND2_X1 U7230 ( .A1(n10588), .A2(n10586), .ZN(n6139) );
  NAND2_X1 U7231 ( .A1(n6139), .A2(n8371), .ZN(n10590) );
  OR2_X1 U7232 ( .A1(n8708), .A2(n6770), .ZN(n6140) );
  NAND2_X1 U7233 ( .A1(n10590), .A2(n6140), .ZN(n7111) );
  NAND2_X1 U7234 ( .A1(n10592), .A2(n6886), .ZN(n6141) );
  NAND2_X1 U7235 ( .A1(n7111), .A2(n6141), .ZN(n6143) );
  OR2_X1 U7236 ( .A1(n10592), .A2(n6886), .ZN(n6142) );
  INV_X1 U7237 ( .A(n7099), .ZN(n6145) );
  INV_X1 U7238 ( .A(n8377), .ZN(n6144) );
  NAND2_X1 U7239 ( .A1(n6145), .A2(n6144), .ZN(n10629) );
  NAND2_X1 U7240 ( .A1(n8707), .A2(n7013), .ZN(n6146) );
  AND2_X1 U7241 ( .A1(n10628), .A2(n6146), .ZN(n6147) );
  AOI21_X2 U7242 ( .B1(n10629), .B2(n6147), .A(n4988), .ZN(n7469) );
  NAND2_X1 U7243 ( .A1(n10635), .A2(n7260), .ZN(n6148) );
  NAND2_X1 U7244 ( .A1(n6151), .A2(n6148), .ZN(n7468) );
  OR2_X1 U7245 ( .A1(n8705), .A2(n10705), .ZN(n6152) );
  INV_X1 U7246 ( .A(n6152), .ZN(n6149) );
  NOR2_X1 U7247 ( .A1(n6149), .A2(n8333), .ZN(n6154) );
  NOR2_X1 U7248 ( .A1(n10635), .A2(n7260), .ZN(n6150) );
  INV_X1 U7249 ( .A(n10687), .ZN(n7302) );
  AOI22_X1 U7250 ( .A1(n6151), .A2(n6150), .B1(n7290), .B2(n7302), .ZN(n7470)
         );
  AND2_X1 U7251 ( .A1(n7470), .A2(n6152), .ZN(n6153) );
  NAND2_X1 U7252 ( .A1(n8703), .A2(n10735), .ZN(n7549) );
  NAND2_X1 U7253 ( .A1(n7552), .A2(n7549), .ZN(n6156) );
  OR2_X1 U7254 ( .A1(n8703), .A2(n10735), .ZN(n7550) );
  NAND2_X1 U7255 ( .A1(n6156), .A2(n7550), .ZN(n7565) );
  NAND2_X1 U7256 ( .A1(n10746), .A2(n8702), .ZN(n6157) );
  NAND2_X1 U7257 ( .A1(n7565), .A2(n6157), .ZN(n6159) );
  OR2_X1 U7258 ( .A1(n10746), .A2(n8702), .ZN(n6158) );
  NAND2_X1 U7259 ( .A1(n8575), .A2(n8701), .ZN(n7588) );
  OR2_X1 U7260 ( .A1(n8575), .A2(n8701), .ZN(n7589) );
  NAND2_X1 U7261 ( .A1(n8361), .A2(n8700), .ZN(n6161) );
  OR2_X1 U7262 ( .A1(n8361), .A2(n8700), .ZN(n6162) );
  NAND2_X1 U7263 ( .A1(n8356), .A2(n8698), .ZN(n8440) );
  NAND2_X1 U7264 ( .A1(n8999), .A2(n8998), .ZN(n6166) );
  NAND2_X1 U7265 ( .A1(n9010), .A2(n8697), .ZN(n6165) );
  NAND2_X1 U7266 ( .A1(n6166), .A2(n6165), .ZN(n8986) );
  NAND2_X1 U7267 ( .A1(n8599), .A2(n8696), .ZN(n6167) );
  OR2_X1 U7268 ( .A1(n8655), .A2(n8958), .ZN(n8953) );
  AND2_X1 U7269 ( .A1(n8956), .A2(n8953), .ZN(n6169) );
  INV_X1 U7270 ( .A(n8977), .ZN(n8944) );
  NAND2_X1 U7271 ( .A1(n8972), .A2(n8944), .ZN(n6170) );
  NAND2_X1 U7272 ( .A1(n8955), .A2(n6170), .ZN(n8939) );
  OR2_X1 U7273 ( .A1(n8950), .A2(n8959), .ZN(n6171) );
  NAND2_X1 U7274 ( .A1(n8941), .A2(n6171), .ZN(n8925) );
  NAND2_X1 U7275 ( .A1(n8467), .A2(n8468), .ZN(n8924) );
  OR2_X1 U7276 ( .A1(n9062), .A2(n8943), .ZN(n6172) );
  NOR2_X1 U7277 ( .A1(n8347), .A2(n8927), .ZN(n6174) );
  AND2_X1 U7278 ( .A1(n8904), .A2(n8695), .ZN(n6175) );
  OR2_X1 U7279 ( .A1(n8904), .A2(n8695), .ZN(n6176) );
  NAND2_X1 U7280 ( .A1(n8891), .A2(n8694), .ZN(n8479) );
  NAND2_X1 U7281 ( .A1(n8888), .A2(n8479), .ZN(n6177) );
  OR2_X1 U7282 ( .A1(n8891), .A2(n8694), .ZN(n8483) );
  NAND2_X1 U7283 ( .A1(n6177), .A2(n8483), .ZN(n8878) );
  NAND2_X1 U7284 ( .A1(n9045), .A2(n8693), .ZN(n6178) );
  OR2_X1 U7285 ( .A1(n9045), .A2(n8693), .ZN(n6179) );
  XNOR2_X1 U7286 ( .A(n6180), .B(n8328), .ZN(n6186) );
  NAND2_X1 U7287 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  NAND2_X1 U7288 ( .A1(n6183), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6184) );
  XNOR2_X2 U7289 ( .A(n6184), .B(n5094), .ZN(n8362) );
  OR2_X1 U7290 ( .A1(n8362), .A2(n8512), .ZN(n6185) );
  NAND2_X1 U7291 ( .A1(n8520), .A2(n8515), .ZN(n6224) );
  NAND2_X1 U7292 ( .A1(n8520), .A2(n7176), .ZN(n6371) );
  INV_X1 U7293 ( .A(n6371), .ZN(n6187) );
  INV_X1 U7294 ( .A(n8520), .ZN(n7545) );
  OAI21_X1 U7295 ( .B1(n6373), .B2(n6187), .A(n10799), .ZN(n6188) );
  NAND2_X1 U7296 ( .A1(n8833), .A2(n10634), .ZN(n6198) );
  INV_X1 U7297 ( .A(n6363), .ZN(n8517) );
  NAND2_X1 U7298 ( .A1(n8517), .A2(n6264), .ZN(n6189) );
  AND2_X1 U7299 ( .A1(n6240), .A2(n6189), .ZN(n6779) );
  NAND2_X1 U7300 ( .A1(n6240), .A2(P2_B_REG_SCAN_IN), .ZN(n6191) );
  AND2_X1 U7301 ( .A1(n6190), .A2(n6191), .ZN(n8825) );
  NAND2_X1 U7302 ( .A1(n8310), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6196) );
  INV_X1 U7303 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6192) );
  OR2_X1 U7304 ( .A1(n8312), .A2(n6192), .ZN(n6195) );
  INV_X1 U7305 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6193) );
  OR2_X1 U7306 ( .A1(n8314), .A2(n6193), .ZN(n6194) );
  NAND4_X1 U7307 ( .A1(n8318), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(n8690)
         );
  AOI22_X1 U7308 ( .A1(n8691), .A2(n10637), .B1(n8825), .B2(n8690), .ZN(n6197)
         );
  NAND2_X1 U7309 ( .A1(n6201), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6202) );
  MUX2_X1 U7310 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6202), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6204) );
  NAND2_X1 U7311 ( .A1(n6205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6206) );
  XNOR2_X1 U7312 ( .A(n7698), .B(P2_B_REG_SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7313 ( .A1(n4997), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7314 ( .A1(n6209), .A2(n7741), .ZN(n6210) );
  NAND2_X1 U7315 ( .A1(n7825), .A2(n7698), .ZN(n6444) );
  NAND2_X1 U7316 ( .A1(n7825), .A2(n7741), .ZN(n6446) );
  NOR2_X1 U7317 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6216) );
  NOR4_X1 U7318 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6215) );
  NOR4_X1 U7319 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6214) );
  NOR4_X1 U7320 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6213) );
  NAND4_X1 U7321 ( .A1(n6216), .A2(n6215), .A3(n6214), .A4(n6213), .ZN(n6222)
         );
  NOR4_X1 U7322 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6220) );
  NOR4_X1 U7323 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6219) );
  NOR4_X1 U7324 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6218) );
  NOR4_X1 U7325 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6217) );
  NAND4_X1 U7326 ( .A1(n6220), .A2(n6219), .A3(n6218), .A4(n6217), .ZN(n6221)
         );
  NOR2_X1 U7327 ( .A1(n6222), .A2(n6221), .ZN(n6223) );
  NAND2_X1 U7328 ( .A1(n6370), .A2(n6368), .ZN(n6759) );
  OR2_X1 U7329 ( .A1(n6224), .A2(n8512), .ZN(n6226) );
  NOR2_X1 U7330 ( .A1(n6226), .A2(n5487), .ZN(n6751) );
  NOR2_X1 U7331 ( .A1(n9022), .A2(n6751), .ZN(n6225) );
  OR2_X1 U7332 ( .A1(n6759), .A2(n6225), .ZN(n6229) );
  NAND3_X1 U7333 ( .A1(n7095), .A2(n7093), .A3(n6368), .ZN(n6756) );
  INV_X1 U7334 ( .A(n6756), .ZN(n6227) );
  NAND3_X1 U7335 ( .A1(n8506), .A2(n10799), .A3(n6226), .ZN(n6753) );
  INV_X1 U7336 ( .A(n7098), .ZN(n6761) );
  OR2_X1 U7337 ( .A1(n10799), .A2(n6761), .ZN(n10598) );
  NAND2_X1 U7338 ( .A1(n6753), .A2(n10598), .ZN(n6742) );
  NAND2_X1 U7339 ( .A1(n6227), .A2(n6742), .ZN(n6228) );
  NAND2_X1 U7340 ( .A1(n6229), .A2(n6228), .ZN(n9091) );
  INV_X1 U7341 ( .A(n7741), .ZN(n6231) );
  INV_X1 U7342 ( .A(n7698), .ZN(n6230) );
  NAND2_X1 U7343 ( .A1(n6231), .A2(n6230), .ZN(n6232) );
  NAND2_X1 U7344 ( .A1(n5035), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6233) );
  INV_X1 U7345 ( .A(n6234), .ZN(n8834) );
  NAND2_X1 U7346 ( .A1(n10810), .A2(n10747), .ZN(n9143) );
  OR2_X1 U7347 ( .A1(n10810), .A2(n6235), .ZN(n6236) );
  INV_X1 U7348 ( .A(n6237), .ZN(n6238) );
  NAND2_X1 U7349 ( .A1(n6744), .A2(n8506), .ZN(n6239) );
  NAND2_X1 U7350 ( .A1(n6239), .A2(n7561), .ZN(n6298) );
  NAND2_X1 U7351 ( .A1(n6240), .A2(n6298), .ZN(n6241) );
  NAND2_X1 U7352 ( .A1(n6241), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7353 ( .A(n6448), .ZN(n6242) );
  INV_X1 U7354 ( .A(n6329), .ZN(n10512) );
  MUX2_X1 U7355 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6314), .S(n6329), .Z(n10509)
         );
  NOR2_X1 U7356 ( .A1(n6317), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7357 ( .A1(n6268), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6244) );
  INV_X1 U7358 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10575) );
  OR2_X1 U7359 ( .A1(n10433), .A2(n6245), .ZN(n6246) );
  NAND2_X1 U7360 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n10471), .ZN(n6248) );
  OAI21_X1 U7361 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n10471), .A(n6248), .ZN(
        n10470) );
  NAND2_X1 U7362 ( .A1(n6250), .A2(n10498), .ZN(n6249) );
  INV_X1 U7363 ( .A(n6249), .ZN(n6251) );
  OAI21_X1 U7364 ( .B1(n6250), .B2(n10498), .A(n6249), .ZN(n10487) );
  NOR2_X1 U7365 ( .A1(n6997), .A2(n6252), .ZN(n6253) );
  NOR2_X1 U7366 ( .A1(n6312), .A2(n6990), .ZN(n6989) );
  AOI22_X1 U7367 ( .A1(n7165), .A2(P2_REG1_REG_8__SCAN_IN), .B1(n6310), .B2(
        n6442), .ZN(n7155) );
  NOR2_X1 U7368 ( .A1(n7381), .A2(n4986), .ZN(n6254) );
  INV_X1 U7369 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U7370 ( .A1(n7678), .A2(P2_REG1_REG_10__SCAN_IN), .B1(n5903), .B2(
        n6472), .ZN(n7663) );
  NOR2_X1 U7371 ( .A1(n7664), .A2(n7663), .ZN(n7662) );
  NOR2_X1 U7372 ( .A1(n6344), .A2(n6255), .ZN(n6256) );
  XNOR2_X1 U7373 ( .A(n6255), .B(n6344), .ZN(n7572) );
  AOI22_X1 U7374 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6308), .B1(n8718), .B2(
        n5932), .ZN(n8720) );
  NOR2_X1 U7375 ( .A1(n6307), .A2(n6257), .ZN(n6258) );
  NAND2_X1 U7376 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8750), .ZN(n6259) );
  OAI21_X1 U7377 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8750), .A(n6259), .ZN(
        n8752) );
  NOR2_X1 U7378 ( .A1(n6303), .A2(n6260), .ZN(n6261) );
  INV_X1 U7379 ( .A(n6303), .ZN(n8766) );
  AOI22_X1 U7380 ( .A1(n6301), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n9087), .B2(
        n8784), .ZN(n8777) );
  INV_X1 U7381 ( .A(n6353), .ZN(n8799) );
  INV_X1 U7382 ( .A(n8821), .ZN(n7010) );
  NAND2_X1 U7383 ( .A1(n7010), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6263) );
  OAI21_X1 U7384 ( .B1(n7010), .B2(P2_REG1_REG_18__SCAN_IN), .A(n6263), .ZN(
        n8807) );
  XNOR2_X1 U7385 ( .A(n8515), .B(n9075), .ZN(n6357) );
  NOR2_X1 U7386 ( .A1(n6363), .A2(P2_U3151), .ZN(n9156) );
  INV_X1 U7387 ( .A(n7561), .ZN(n6265) );
  NOR2_X1 U7388 ( .A1(n6744), .A2(n6265), .ZN(n6266) );
  INV_X1 U7389 ( .A(n6497), .ZN(n6267) );
  XNOR2_X1 U7390 ( .A(n10433), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n10431) );
  NOR2_X1 U7391 ( .A1(n6318), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7392 ( .A1(n6268), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7393 ( .A1(n6677), .A2(n6270), .ZN(n10430) );
  OR2_X1 U7394 ( .A1(n10433), .A2(n6271), .ZN(n6272) );
  XNOR2_X1 U7395 ( .A(n6273), .B(n10459), .ZN(n10449) );
  NAND2_X1 U7396 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n10471), .ZN(n6274) );
  OAI21_X1 U7397 ( .B1(n10471), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6274), .ZN(
        n10478) );
  OR2_X1 U7398 ( .A1(n6275), .A2(n6326), .ZN(n6276) );
  MUX2_X1 U7399 ( .A(n7151), .B(P2_REG2_REG_6__SCAN_IN), .S(n6329), .Z(n10523)
         );
  NOR2_X1 U7400 ( .A1(n6997), .A2(n6278), .ZN(n6279) );
  AOI22_X1 U7401 ( .A1(n7165), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n6311), .B2(
        n6442), .ZN(n7158) );
  NOR2_X1 U7402 ( .A1(n7159), .A2(n7158), .ZN(n7157) );
  MUX2_X1 U7403 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n6283), .S(n7678), .Z(n7674)
         );
  XNOR2_X1 U7404 ( .A(n6344), .B(n6284), .ZN(n7574) );
  MUX2_X1 U7405 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6285), .S(n6308), .Z(n8711)
         );
  NOR2_X1 U7406 ( .A1(n6307), .A2(n6286), .ZN(n6287) );
  NAND2_X1 U7407 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8750), .ZN(n6288) );
  OAI21_X1 U7408 ( .B1(n8750), .B2(P2_REG2_REG_14__SCAN_IN), .A(n6288), .ZN(
        n8743) );
  NOR2_X1 U7409 ( .A1(n6303), .A2(n6289), .ZN(n6290) );
  NOR2_X1 U7410 ( .A1(n8761), .A2(n6290), .ZN(n8787) );
  NOR2_X1 U7411 ( .A1(n8784), .A2(n9012), .ZN(n6291) );
  AOI21_X1 U7412 ( .B1(n9012), .B2(n8784), .A(n6291), .ZN(n8786) );
  NOR2_X1 U7413 ( .A1(n8787), .A2(n8786), .ZN(n8785) );
  NAND2_X1 U7414 ( .A1(n6353), .A2(n6292), .ZN(n6293) );
  NAND2_X1 U7415 ( .A1(n6295), .A2(n6293), .ZN(n8800) );
  NOR2_X2 U7416 ( .A1(n8800), .A2(n8993), .ZN(n8814) );
  XNOR2_X1 U7417 ( .A(n8821), .B(P2_REG2_REG_18__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U7418 ( .A1(n6295), .A2(n8981), .ZN(n6294) );
  INV_X1 U7419 ( .A(n6295), .ZN(n8815) );
  XNOR2_X1 U7420 ( .A(n8515), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U7421 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8553) );
  NOR2_X1 U7422 ( .A1(n6358), .A2(P2_U3151), .ZN(n9159) );
  NAND2_X1 U7423 ( .A1(n9159), .A2(n6298), .ZN(n6299) );
  NOR2_X1 U7424 ( .A1(n10511), .A2(n7176), .ZN(n6300) );
  MUX2_X1 U7425 ( .A(n8993), .B(n9083), .S(n8516), .Z(n6354) );
  XNOR2_X1 U7426 ( .A(n6354), .B(n8799), .ZN(n8798) );
  MUX2_X1 U7427 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6358), .Z(n6302) );
  OR2_X1 U7428 ( .A1(n6302), .A2(n8784), .ZN(n6351) );
  XNOR2_X1 U7429 ( .A(n6302), .B(n6301), .ZN(n8781) );
  MUX2_X1 U7430 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8516), .Z(n6304) );
  OR2_X1 U7431 ( .A1(n6304), .A2(n8766), .ZN(n6350) );
  XNOR2_X1 U7432 ( .A(n6304), .B(n6303), .ZN(n8771) );
  MUX2_X1 U7433 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8516), .Z(n6306) );
  OR2_X1 U7434 ( .A1(n6306), .A2(n8750), .ZN(n6349) );
  XNOR2_X1 U7435 ( .A(n6306), .B(n6305), .ZN(n8746) );
  MUX2_X1 U7436 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8516), .Z(n6348) );
  XNOR2_X1 U7437 ( .A(n6348), .B(n6307), .ZN(n8731) );
  MUX2_X1 U7438 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6358), .Z(n6309) );
  OR2_X1 U7439 ( .A1(n6309), .A2(n8718), .ZN(n6347) );
  XNOR2_X1 U7440 ( .A(n6309), .B(n6308), .ZN(n8715) );
  MUX2_X1 U7441 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8516), .Z(n6345) );
  INV_X1 U7442 ( .A(n6344), .ZN(n7578) );
  OR2_X1 U7443 ( .A1(n6345), .A2(n7578), .ZN(n6346) );
  MUX2_X1 U7444 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8516), .Z(n6340) );
  INV_X1 U7445 ( .A(n6340), .ZN(n6341) );
  MUX2_X1 U7446 ( .A(n6311), .B(n6310), .S(n6358), .Z(n6338) );
  NAND2_X1 U7447 ( .A1(n6338), .A2(n7165), .ZN(n6337) );
  INV_X1 U7448 ( .A(n6337), .ZN(n6339) );
  MUX2_X1 U7449 ( .A(n6313), .B(n6312), .S(n8516), .Z(n6335) );
  NAND2_X1 U7450 ( .A1(n6335), .A2(n6997), .ZN(n6334) );
  INV_X1 U7451 ( .A(n6334), .ZN(n6336) );
  MUX2_X1 U7452 ( .A(n7151), .B(n6314), .S(n6358), .Z(n6330) );
  NAND2_X1 U7453 ( .A1(n6330), .A2(n6329), .ZN(n6328) );
  INV_X1 U7454 ( .A(n6328), .ZN(n6333) );
  INV_X1 U7455 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10615) );
  MUX2_X1 U7456 ( .A(n5796), .B(n10615), .S(n6358), .Z(n6324) );
  MUX2_X1 U7457 ( .A(n6316), .B(n6315), .S(n8516), .Z(n6322) );
  MUX2_X1 U7458 ( .A(n5751), .B(n10575), .S(n6358), .Z(n6319) );
  XNOR2_X1 U7459 ( .A(n6319), .B(n6675), .ZN(n6674) );
  MUX2_X1 U7460 ( .A(n6318), .B(n6317), .S(n6358), .Z(n6495) );
  NAND2_X1 U7461 ( .A1(n6495), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6673) );
  INV_X1 U7462 ( .A(n6319), .ZN(n6320) );
  AOI22_X1 U7463 ( .A1(n6674), .A2(n6673), .B1(n6675), .B2(n6320), .ZN(n10443)
         );
  MUX2_X1 U7464 ( .A(n6271), .B(n6245), .S(n6358), .Z(n6321) );
  XNOR2_X1 U7465 ( .A(n6321), .B(n10433), .ZN(n10444) );
  OAI22_X1 U7466 ( .A1(n10443), .A2(n10444), .B1(n10433), .B2(n6321), .ZN(
        n10462) );
  XNOR2_X1 U7467 ( .A(n6322), .B(n6323), .ZN(n10463) );
  NOR2_X1 U7468 ( .A1(n10462), .A2(n10463), .ZN(n10461) );
  XNOR2_X1 U7469 ( .A(n6324), .B(n10471), .ZN(n10475) );
  NAND2_X1 U7470 ( .A1(n10476), .A2(n10475), .ZN(n10474) );
  OAI21_X1 U7471 ( .B1(n6325), .B2(n6324), .A(n10474), .ZN(n10501) );
  MUX2_X1 U7472 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8516), .Z(n6327) );
  XNOR2_X1 U7473 ( .A(n6327), .B(n6326), .ZN(n10502) );
  AOI22_X1 U7474 ( .A1(n10501), .A2(n10502), .B1(n6327), .B2(n10498), .ZN(
        n10517) );
  INV_X1 U7475 ( .A(n10517), .ZN(n6331) );
  OAI21_X1 U7476 ( .B1(n6330), .B2(n6329), .A(n6328), .ZN(n10518) );
  NOR2_X1 U7477 ( .A1(n6331), .A2(n10518), .ZN(n6332) );
  OAI21_X1 U7478 ( .B1(n6335), .B2(n6997), .A(n6334), .ZN(n6996) );
  NOR2_X1 U7479 ( .A1(n6995), .A2(n6996), .ZN(n6994) );
  NOR2_X1 U7480 ( .A1(n6336), .A2(n6994), .ZN(n7162) );
  OAI21_X1 U7481 ( .B1(n6338), .B2(n7165), .A(n6337), .ZN(n7163) );
  NOR2_X1 U7482 ( .A1(n7162), .A2(n7163), .ZN(n7161) );
  XNOR2_X1 U7483 ( .A(n6340), .B(n6464), .ZN(n7380) );
  NOR2_X1 U7484 ( .A1(n7379), .A2(n7380), .ZN(n7378) );
  MUX2_X1 U7485 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n6358), .Z(n6342) );
  OR2_X1 U7486 ( .A1(n6342), .A2(n6472), .ZN(n7665) );
  NAND2_X1 U7487 ( .A1(n6342), .A2(n6472), .ZN(n7666) );
  INV_X1 U7488 ( .A(n7666), .ZN(n6343) );
  AOI21_X1 U7489 ( .B1(n7669), .B2(n7665), .A(n6343), .ZN(n7582) );
  XNOR2_X1 U7490 ( .A(n6345), .B(n6344), .ZN(n7583) );
  NAND2_X1 U7491 ( .A1(n7582), .A2(n7583), .ZN(n7581) );
  NAND2_X1 U7492 ( .A1(n6346), .A2(n7581), .ZN(n8714) );
  NAND2_X1 U7493 ( .A1(n8715), .A2(n8714), .ZN(n8713) );
  NAND2_X1 U7494 ( .A1(n6347), .A2(n8713), .ZN(n8730) );
  NAND2_X1 U7495 ( .A1(n8731), .A2(n8730), .ZN(n8729) );
  OAI21_X1 U7496 ( .B1(n6348), .B2(n5050), .A(n8729), .ZN(n8747) );
  NAND2_X1 U7497 ( .A1(n8746), .A2(n8747), .ZN(n8745) );
  NAND2_X1 U7498 ( .A1(n6349), .A2(n8745), .ZN(n8770) );
  NAND2_X1 U7499 ( .A1(n8771), .A2(n8770), .ZN(n8769) );
  NAND2_X1 U7500 ( .A1(n6350), .A2(n8769), .ZN(n8780) );
  NAND2_X1 U7501 ( .A1(n8781), .A2(n8780), .ZN(n8779) );
  NAND2_X1 U7502 ( .A1(n6351), .A2(n8779), .ZN(n8797) );
  NAND2_X1 U7503 ( .A1(n8798), .A2(n8797), .ZN(n8796) );
  INV_X1 U7504 ( .A(n8796), .ZN(n6352) );
  MUX2_X1 U7505 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n6358), .Z(n6355) );
  NOR2_X1 U7506 ( .A1(n6356), .A2(n6355), .ZN(n8811) );
  NAND2_X1 U7507 ( .A1(n6356), .A2(n6355), .ZN(n8809) );
  OAI21_X1 U7508 ( .B1(n8811), .B2(n8821), .A(n8809), .ZN(n6362) );
  INV_X1 U7509 ( .A(n6357), .ZN(n6359) );
  MUX2_X1 U7510 ( .A(n6360), .B(n6359), .S(n8516), .Z(n6361) );
  XNOR2_X1 U7511 ( .A(n6362), .B(n6361), .ZN(n6364) );
  NAND2_X1 U7512 ( .A1(P2_U3893), .A2(n6363), .ZN(n10464) );
  INV_X1 U7513 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U7514 ( .A1(n6758), .A2(n6368), .ZN(n6369) );
  OR2_X1 U7515 ( .A1(n6370), .A2(n6369), .ZN(n7091) );
  OAI21_X1 U7516 ( .B1(n5487), .B2(n10643), .A(n6767), .ZN(n6374) );
  NOR2_X1 U7517 ( .A1(n6371), .A2(n8512), .ZN(n6372) );
  NAND2_X1 U7518 ( .A1(n7094), .A2(n6743), .ZN(n7092) );
  NAND2_X1 U7519 ( .A1(n6374), .A2(n7092), .ZN(n6376) );
  NAND2_X1 U7520 ( .A1(n7093), .A2(n7094), .ZN(n6375) );
  NAND3_X1 U7521 ( .A1(n6459), .A2(n6457), .A3(n6383), .ZN(n6565) );
  INV_X1 U7522 ( .A(n6565), .ZN(n6387) );
  NAND4_X1 U7523 ( .A1(n6387), .A2(n6386), .A3(n6385), .A4(n6384), .ZN(n6388)
         );
  NAND3_X1 U7524 ( .A1(n6404), .A2(n6406), .A3(n6408), .ZN(n6399) );
  NAND2_X1 U7525 ( .A1(n6396), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6397) );
  MUX2_X1 U7526 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6397), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n6398) );
  NAND2_X1 U7527 ( .A1(n6398), .A2(n4965), .ZN(n7744) );
  INV_X1 U7528 ( .A(n7744), .ZN(n6403) );
  NAND2_X1 U7529 ( .A1(n6399), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U7530 ( .A1(n6483), .A2(n6400), .ZN(n6401) );
  INV_X1 U7531 ( .A(n7700), .ZN(n6402) );
  NOR2_X1 U7532 ( .A1(n6969), .A2(P1_U3086), .ZN(n6410) );
  NAND2_X1 U7533 ( .A1(n6483), .A2(n6404), .ZN(n6405) );
  NAND2_X1 U7534 ( .A1(n6482), .A2(n6406), .ZN(n6407) );
  NAND2_X1 U7535 ( .A1(n6407), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6409) );
  NAND2_X2 U7536 ( .A1(n7890), .A2(P2_U3151), .ZN(n9162) );
  NOR2_X1 U7537 ( .A1(n7890), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9160) );
  AOI22_X1 U7538 ( .A1(n10433), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n9160), .ZN(n6411) );
  OAI21_X1 U7539 ( .B1(n6843), .B2(n9162), .A(n6411), .ZN(P2_U3293) );
  NAND2_X1 U7540 ( .A1(n5056), .A2(P1_U3086), .ZN(n10132) );
  INV_X1 U7541 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7031) );
  NAND2_X1 U7542 ( .A1(n6412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6413) );
  XNOR2_X1 U7543 ( .A(n6413), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10541) );
  INV_X1 U7544 ( .A(n10541), .ZN(n7034) );
  OAI222_X1 U7545 ( .A1(n10132), .A2(n7031), .B1(n10138), .B2(n7030), .C1(
        P1_U3086), .C2(n7034), .ZN(P1_U3351) );
  INV_X1 U7546 ( .A(n9160), .ZN(n9153) );
  INV_X1 U7547 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6414) );
  OAI222_X1 U7548 ( .A1(n9153), .A2(n6414), .B1(n9162), .B2(n6716), .C1(n6675), 
        .C2(P2_U3151), .ZN(P2_U3294) );
  INV_X1 U7549 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6415) );
  OAI222_X1 U7550 ( .A1(n10471), .A2(P2_U3151), .B1(n9162), .B2(n7030), .C1(
        n6415), .C2(n9153), .ZN(P2_U3291) );
  INV_X1 U7551 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6416) );
  OAI222_X1 U7552 ( .A1(n10498), .A2(P2_U3151), .B1(n9162), .B2(n7194), .C1(
        n6416), .C2(n9153), .ZN(P2_U3290) );
  INV_X1 U7553 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6417) );
  OAI222_X1 U7554 ( .A1(n9153), .A2(n6417), .B1(n9162), .B2(n6942), .C1(n10459), .C2(P2_U3151), .ZN(P2_U3292) );
  INV_X1 U7555 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6418) );
  OAI222_X1 U7556 ( .A1(n10512), .A2(P2_U3151), .B1(n9162), .B2(n7222), .C1(
        n6418), .C2(n9153), .ZN(P2_U3289) );
  INV_X1 U7557 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6844) );
  OR2_X1 U7558 ( .A1(n6419), .A2(n10124), .ZN(n6427) );
  INV_X1 U7559 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6426) );
  XNOR2_X1 U7560 ( .A(n6427), .B(n6426), .ZN(n6847) );
  OAI222_X1 U7561 ( .A1(n10132), .A2(n6844), .B1(n10138), .B2(n6843), .C1(
        P1_U3086), .C2(n6847), .ZN(P1_U3353) );
  INV_X1 U7562 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7195) );
  NAND2_X1 U7563 ( .A1(n6420), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6421) );
  MUX2_X1 U7564 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6421), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n6424) );
  INV_X1 U7565 ( .A(n6422), .ZN(n6423) );
  INV_X1 U7566 ( .A(n6528), .ZN(n7198) );
  OAI222_X1 U7567 ( .A1(n10132), .A2(n7195), .B1(n10138), .B2(n7194), .C1(
        P1_U3086), .C2(n7198), .ZN(P1_U3350) );
  INV_X1 U7568 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7223) );
  OR2_X1 U7569 ( .A1(n6422), .A2(n10124), .ZN(n6425) );
  XNOR2_X1 U7570 ( .A(n6425), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6544) );
  INV_X1 U7571 ( .A(n6544), .ZN(n7226) );
  OAI222_X1 U7572 ( .A1(n10132), .A2(n7223), .B1(n10138), .B2(n7222), .C1(
        P1_U3086), .C2(n7226), .ZN(P1_U3349) );
  INV_X1 U7573 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U7574 ( .A1(n6427), .A2(n6426), .ZN(n6428) );
  NAND2_X1 U7575 ( .A1(n6428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6430) );
  INV_X1 U7576 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6429) );
  XNOR2_X1 U7577 ( .A(n6430), .B(n6429), .ZN(n6947) );
  OAI222_X1 U7578 ( .A1(n10132), .A2(n6944), .B1(n10138), .B2(n6942), .C1(
        P1_U3086), .C2(n6947), .ZN(P1_U3352) );
  INV_X1 U7579 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U7580 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6431) );
  XNOR2_X1 U7581 ( .A(n6432), .B(n6431), .ZN(n6719) );
  OAI222_X1 U7582 ( .A1(P1_U3086), .A2(n6719), .B1(n10138), .B2(n6716), .C1(
        n5044), .C2(n10132), .ZN(P1_U3354) );
  INV_X1 U7583 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7347) );
  OR2_X1 U7584 ( .A1(n6433), .A2(n10124), .ZN(n6434) );
  XNOR2_X1 U7585 ( .A(n6434), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6555) );
  INV_X1 U7586 ( .A(n6555), .ZN(n7350) );
  OAI222_X1 U7587 ( .A1(n10132), .A2(n7347), .B1(n10138), .B2(n7346), .C1(
        P1_U3086), .C2(n7350), .ZN(P1_U3348) );
  OAI222_X1 U7588 ( .A1(n6436), .A2(P2_U3151), .B1(n9162), .B2(n7346), .C1(
        n6435), .C2(n9153), .ZN(P2_U3288) );
  INV_X1 U7589 ( .A(n7395), .ZN(n6441) );
  NAND2_X1 U7590 ( .A1(n6437), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6438) );
  XNOR2_X1 U7591 ( .A(n6438), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7393) );
  INV_X1 U7592 ( .A(n10132), .ZN(n10126) );
  AOI22_X1 U7593 ( .A1(n7393), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10126), .ZN(n6439) );
  OAI21_X1 U7594 ( .B1(n6441), .B2(n10138), .A(n6439), .ZN(P1_U3347) );
  OAI222_X1 U7595 ( .A1(n6442), .A2(P2_U3151), .B1(n9162), .B2(n6441), .C1(
        n6440), .C2(n9153), .ZN(P2_U3287) );
  INV_X1 U7596 ( .A(n6444), .ZN(n6445) );
  AOI22_X1 U7597 ( .A1(n6450), .A2(n5356), .B1(n6448), .B2(n6445), .ZN(
        P2_U3376) );
  INV_X1 U7598 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6449) );
  INV_X1 U7599 ( .A(n6446), .ZN(n6447) );
  AOI22_X1 U7600 ( .A1(n6450), .A2(n6449), .B1(n6448), .B2(n6447), .ZN(
        P2_U3377) );
  AND2_X1 U7601 ( .A1(n6450), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U7602 ( .A1(n6450), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U7603 ( .A1(n6450), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U7604 ( .A1(n6450), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U7605 ( .A1(n6450), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U7606 ( .A1(n6450), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U7607 ( .A1(n6450), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U7608 ( .A1(n6450), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U7609 ( .A1(n6450), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U7610 ( .A1(n6450), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U7611 ( .A1(n6450), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U7612 ( .A1(n6450), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U7613 ( .A1(n6450), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U7614 ( .A1(n6450), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U7615 ( .A1(n6450), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U7616 ( .A1(n6450), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U7617 ( .A1(n6450), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U7618 ( .A1(n6450), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U7619 ( .A1(n6450), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U7620 ( .A1(n6450), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U7621 ( .A1(n6450), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U7622 ( .A1(n6450), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U7623 ( .A1(n6450), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U7624 ( .A1(n6450), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U7625 ( .A1(n6450), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U7626 ( .A1(n6450), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U7627 ( .A1(n6450), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U7628 ( .A1(n6450), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U7629 ( .A1(n6450), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U7630 ( .A1(n6450), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U7631 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U7632 ( .A1(n7744), .A2(P1_B_REG_SCAN_IN), .ZN(n6451) );
  MUX2_X1 U7633 ( .A(P1_B_REG_SCAN_IN), .B(n6451), .S(n7700), .Z(n6452) );
  INV_X1 U7634 ( .A(n6453), .ZN(n7821) );
  AND2_X1 U7635 ( .A1(n7821), .A2(n7744), .ZN(n6454) );
  NAND2_X1 U7636 ( .A1(n6827), .A2(n6651), .ZN(n6455) );
  OAI21_X1 U7637 ( .B1(n6651), .B2(n6456), .A(n6455), .ZN(P1_U3440) );
  INV_X1 U7638 ( .A(n7511), .ZN(n6471) );
  OR2_X1 U7639 ( .A1(n6437), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6566) );
  NAND2_X1 U7640 ( .A1(n6566), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U7641 ( .A1(n6465), .A2(n6457), .ZN(n6458) );
  NAND2_X1 U7642 ( .A1(n6458), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U7643 ( .A1(n6460), .A2(n6459), .ZN(n6490) );
  OR2_X1 U7644 ( .A1(n6460), .A2(n6459), .ZN(n6461) );
  AOI22_X1 U7645 ( .A1(n7512), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10126), .ZN(n6462) );
  OAI21_X1 U7646 ( .B1(n6471), .B2(n10138), .A(n6462), .ZN(P1_U3345) );
  INV_X1 U7647 ( .A(n7483), .ZN(n6466) );
  OAI222_X1 U7648 ( .A1(P2_U3151), .A2(n6464), .B1(n9162), .B2(n6466), .C1(
        n6463), .C2(n9153), .ZN(P2_U3286) );
  XNOR2_X1 U7649 ( .A(n6465), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7484) );
  INV_X1 U7650 ( .A(n7484), .ZN(n6587) );
  OAI222_X1 U7651 ( .A1(n10132), .A2(n6467), .B1(n10138), .B2(n6466), .C1(
        n6587), .C2(P1_U3086), .ZN(P1_U3346) );
  AND2_X1 U7652 ( .A1(n7821), .A2(n7700), .ZN(n6628) );
  NAND2_X1 U7653 ( .A1(n10141), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6469) );
  OAI21_X1 U7654 ( .B1(n10141), .B2(n6628), .A(n6469), .ZN(P1_U3439) );
  OAI222_X1 U7655 ( .A1(P2_U3151), .A2(n6472), .B1(n9162), .B2(n6471), .C1(
        n6470), .C2(n9153), .ZN(P2_U3285) );
  INV_X1 U7656 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6477) );
  INV_X1 U7657 ( .A(n6594), .ZN(n6474) );
  NAND2_X1 U7658 ( .A1(n6474), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6475) );
  XNOR2_X1 U7659 ( .A(n6480), .B(P1_IR_REG_27__SCAN_IN), .ZN(n9684) );
  INV_X1 U7660 ( .A(n9684), .ZN(n10139) );
  OR2_X1 U7661 ( .A1(n10135), .A2(n10139), .ZN(n8295) );
  OR2_X1 U7662 ( .A1(n10135), .A2(n9684), .ZN(n9581) );
  INV_X1 U7663 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10568) );
  OAI22_X1 U7664 ( .A1(n6477), .A2(n8295), .B1(n9581), .B2(n10568), .ZN(n6478)
         );
  XNOR2_X1 U7665 ( .A(n6478), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6489) );
  INV_X1 U7666 ( .A(n7559), .ZN(n6479) );
  OAI21_X1 U7667 ( .B1(n6479), .B2(n6969), .A(P1_STATE_REG_SCAN_IN), .ZN(n6486) );
  NAND2_X1 U7668 ( .A1(n8223), .A2(n7559), .ZN(n6484) );
  NAND2_X1 U7669 ( .A1(n7392), .A2(n6484), .ZN(n6485) );
  OR2_X1 U7670 ( .A1(n6486), .A2(n6485), .ZN(n6516) );
  INV_X1 U7671 ( .A(n6485), .ZN(n6487) );
  INV_X1 U7672 ( .A(n9669), .ZN(n10532) );
  AOI22_X1 U7673 ( .A1(n10532), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6488) );
  OAI21_X1 U7674 ( .B1(n6489), .B2(n6516), .A(n6488), .ZN(P1_U3243) );
  INV_X1 U7675 ( .A(n7610), .ZN(n6494) );
  NAND2_X1 U7676 ( .A1(n6490), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6491) );
  XNOR2_X1 U7677 ( .A(n6491), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7611) );
  AOI22_X1 U7678 ( .A1(n7611), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10126), .ZN(n6492) );
  OAI21_X1 U7679 ( .B1(n6494), .B2(n10138), .A(n6492), .ZN(P1_U3344) );
  OAI222_X1 U7680 ( .A1(n7578), .A2(P2_U3151), .B1(n9162), .B2(n6494), .C1(
        n6493), .C2(n9153), .ZN(P2_U3284) );
  INV_X1 U7681 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6500) );
  AOI22_X1 U7682 ( .A1(n10516), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n6499) );
  OAI21_X1 U7683 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6495), .A(n6673), .ZN(n6496) );
  OAI21_X1 U7684 ( .B1(n6497), .B2(n10519), .A(n6496), .ZN(n6498) );
  OAI211_X1 U7685 ( .C1(n10511), .C2(n6500), .A(n6499), .B(n6498), .ZN(
        P2_U3182) );
  XNOR2_X1 U7686 ( .A(n6847), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9589) );
  XNOR2_X1 U7687 ( .A(n6719), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9570) );
  INV_X1 U7688 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6622) );
  NOR2_X1 U7689 ( .A1(n6622), .A2(n6477), .ZN(n9578) );
  NAND2_X1 U7690 ( .A1(n9570), .A2(n9578), .ZN(n9569) );
  INV_X1 U7691 ( .A(n6719), .ZN(n9568) );
  NAND2_X1 U7692 ( .A1(n9568), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6501) );
  NAND2_X1 U7693 ( .A1(n9569), .A2(n6501), .ZN(n9588) );
  NAND2_X1 U7694 ( .A1(n9589), .A2(n9588), .ZN(n9587) );
  INV_X1 U7695 ( .A(n6847), .ZN(n9586) );
  NAND2_X1 U7696 ( .A1(n9586), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U7697 ( .A1(n9587), .A2(n6502), .ZN(n9604) );
  XNOR2_X1 U7698 ( .A(n6947), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9605) );
  NAND2_X1 U7699 ( .A1(n9604), .A2(n9605), .ZN(n9603) );
  INV_X1 U7700 ( .A(n6947), .ZN(n9599) );
  NAND2_X1 U7701 ( .A1(n9599), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U7702 ( .A1(n9603), .A2(n6503), .ZN(n10539) );
  INV_X1 U7703 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6504) );
  MUX2_X1 U7704 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6504), .S(n10541), .Z(n10540) );
  AND2_X1 U7705 ( .A1(n10539), .A2(n10540), .ZN(n10536) );
  AOI21_X1 U7706 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n10541), .A(n10536), .ZN(
        n6507) );
  NAND2_X1 U7707 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6528), .ZN(n6505) );
  OAI21_X1 U7708 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6528), .A(n6505), .ZN(
        n6506) );
  NOR2_X1 U7709 ( .A1(n6507), .A2(n6506), .ZN(n6522) );
  INV_X1 U7710 ( .A(n10538), .ZN(n9623) );
  AOI211_X1 U7711 ( .C1(n6507), .C2(n6506), .A(n6522), .B(n9623), .ZN(n6521)
         );
  XNOR2_X1 U7712 ( .A(n6847), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9592) );
  XNOR2_X1 U7713 ( .A(n6719), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9567) );
  AND2_X1 U7714 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9566) );
  NAND2_X1 U7715 ( .A1(n9567), .A2(n9566), .ZN(n9565) );
  NAND2_X1 U7716 ( .A1(n9568), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U7717 ( .A1(n9565), .A2(n6508), .ZN(n9591) );
  NAND2_X1 U7718 ( .A1(n9592), .A2(n9591), .ZN(n9590) );
  NAND2_X1 U7719 ( .A1(n9586), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U7720 ( .A1(n9590), .A2(n6509), .ZN(n9601) );
  XNOR2_X1 U7721 ( .A(n6947), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9602) );
  NAND2_X1 U7722 ( .A1(n9601), .A2(n9602), .ZN(n9600) );
  NAND2_X1 U7723 ( .A1(n9599), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U7724 ( .A1(n9600), .A2(n6510), .ZN(n10534) );
  INV_X1 U7725 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10625) );
  MUX2_X1 U7726 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10625), .S(n10541), .Z(
        n10535) );
  NAND2_X1 U7727 ( .A1(n10534), .A2(n10535), .ZN(n10533) );
  INV_X1 U7728 ( .A(n10533), .ZN(n6511) );
  AOI21_X1 U7729 ( .B1(n10541), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6511), .ZN(
        n6515) );
  NAND2_X1 U7730 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6528), .ZN(n6512) );
  OAI21_X1 U7731 ( .B1(n6528), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6512), .ZN(
        n6514) );
  NOR2_X1 U7732 ( .A1(n6515), .A2(n6514), .ZN(n6527) );
  INV_X1 U7733 ( .A(n6516), .ZN(n6513) );
  AOI211_X1 U7734 ( .C1(n6515), .C2(n6514), .A(n6527), .B(n10546), .ZN(n6520)
         );
  INV_X1 U7735 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6518) );
  INV_X1 U7736 ( .A(n10135), .ZN(n9576) );
  NOR2_X2 U7737 ( .A1(n6516), .A2(n9576), .ZN(n10542) );
  NAND2_X1 U7738 ( .A1(n10542), .A2(n6528), .ZN(n6517) );
  NAND2_X1 U7739 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7205) );
  OAI211_X1 U7740 ( .C1(n6518), .C2(n9669), .A(n6517), .B(n7205), .ZN(n6519)
         );
  OR3_X1 U7741 ( .A1(n6521), .A2(n6520), .A3(n6519), .ZN(P1_U3248) );
  AOI21_X1 U7742 ( .B1(n6528), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6522), .ZN(
        n6540) );
  NAND2_X1 U7743 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n6544), .ZN(n6523) );
  OAI21_X1 U7744 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6544), .A(n6523), .ZN(
        n6539) );
  NOR2_X1 U7745 ( .A1(n6540), .A2(n6539), .ZN(n6538) );
  AOI21_X1 U7746 ( .B1(n6544), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6538), .ZN(
        n6526) );
  INV_X1 U7747 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6524) );
  AOI22_X1 U7748 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n7350), .B1(n6555), .B2(
        n6524), .ZN(n6525) );
  NOR2_X1 U7749 ( .A1(n6526), .A2(n6525), .ZN(n6550) );
  AOI211_X1 U7750 ( .C1(n6526), .C2(n6525), .A(n6550), .B(n9623), .ZN(n6537)
         );
  AOI21_X1 U7751 ( .B1(n6528), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6527), .ZN(
        n6543) );
  NAND2_X1 U7752 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(n6544), .ZN(n6529) );
  OAI21_X1 U7753 ( .B1(n6544), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6529), .ZN(
        n6542) );
  NOR2_X1 U7754 ( .A1(n6543), .A2(n6542), .ZN(n6541) );
  AOI21_X1 U7755 ( .B1(n6544), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6541), .ZN(
        n6532) );
  INV_X1 U7756 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6530) );
  MUX2_X1 U7757 ( .A(n6530), .B(P1_REG1_REG_7__SCAN_IN), .S(n6555), .Z(n6531)
         );
  NOR2_X1 U7758 ( .A1(n6532), .A2(n6531), .ZN(n6554) );
  AOI211_X1 U7759 ( .C1(n6532), .C2(n6531), .A(n6554), .B(n10546), .ZN(n6536)
         );
  INV_X1 U7760 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U7761 ( .A1(n10542), .A2(n6555), .ZN(n6533) );
  NAND2_X1 U7762 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n7443) );
  OAI211_X1 U7763 ( .C1(n6534), .C2(n9669), .A(n6533), .B(n7443), .ZN(n6535)
         );
  OR3_X1 U7764 ( .A1(n6537), .A2(n6536), .A3(n6535), .ZN(P1_U3250) );
  AOI211_X1 U7765 ( .C1(n6540), .C2(n6539), .A(n6538), .B(n9623), .ZN(n6549)
         );
  AOI211_X1 U7766 ( .C1(n6543), .C2(n6542), .A(n6541), .B(n10546), .ZN(n6548)
         );
  INV_X1 U7767 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U7768 ( .A1(n10542), .A2(n6544), .ZN(n6545) );
  NAND2_X1 U7769 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7232) );
  OAI211_X1 U7770 ( .C1(n6546), .C2(n9669), .A(n6545), .B(n7232), .ZN(n6547)
         );
  OR3_X1 U7771 ( .A1(n6549), .A2(n6548), .A3(n6547), .ZN(P1_U3249) );
  AOI21_X1 U7772 ( .B1(n6555), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6550), .ZN(
        n6553) );
  NAND2_X1 U7773 ( .A1(n7393), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6551) );
  OAI21_X1 U7774 ( .B1(n7393), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6551), .ZN(
        n6552) );
  NOR2_X1 U7775 ( .A1(n6553), .A2(n6552), .ZN(n6578) );
  AOI211_X1 U7776 ( .C1(n6553), .C2(n6552), .A(n6578), .B(n9623), .ZN(n6563)
         );
  AOI21_X1 U7777 ( .B1(n6555), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6554), .ZN(
        n6558) );
  NAND2_X1 U7778 ( .A1(n7393), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6556) );
  OAI21_X1 U7779 ( .B1(n7393), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6556), .ZN(
        n6557) );
  NOR2_X1 U7780 ( .A1(n6558), .A2(n6557), .ZN(n6581) );
  AOI211_X1 U7781 ( .C1(n6558), .C2(n6557), .A(n6581), .B(n10546), .ZN(n6562)
         );
  INV_X1 U7782 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6560) );
  NAND2_X1 U7783 ( .A1(n10542), .A2(n7393), .ZN(n6559) );
  NAND2_X1 U7784 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9393) );
  OAI211_X1 U7785 ( .C1(n6560), .C2(n9669), .A(n6559), .B(n9393), .ZN(n6561)
         );
  OR3_X1 U7786 ( .A1(n6563), .A2(n6562), .A3(n6561), .ZN(P1_U3251) );
  INV_X1 U7787 ( .A(n7703), .ZN(n6571) );
  INV_X1 U7788 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6564) );
  OAI222_X1 U7789 ( .A1(P2_U3151), .A2(n8718), .B1(n9162), .B2(n6571), .C1(
        n6564), .C2(n9153), .ZN(P2_U3283) );
  INV_X1 U7790 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6572) );
  NOR2_X1 U7791 ( .A1(n6566), .A2(n6565), .ZN(n6569) );
  OR2_X1 U7792 ( .A1(n6569), .A2(n10124), .ZN(n6567) );
  MUX2_X1 U7793 ( .A(n6567), .B(P1_IR_REG_31__SCAN_IN), .S(n6568), .Z(n6570)
         );
  NAND2_X1 U7794 ( .A1(n6569), .A2(n6568), .ZN(n6574) );
  INV_X1 U7795 ( .A(n7704), .ZN(n6878) );
  OAI222_X1 U7796 ( .A1(n10132), .A2(n6572), .B1(n10138), .B2(n6571), .C1(
        n6878), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U7797 ( .A(n7707), .ZN(n6592) );
  NAND2_X1 U7798 ( .A1(n6574), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6573) );
  MUX2_X1 U7799 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6573), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n6575) );
  AOI22_X1 U7800 ( .A1(n7708), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10126), .ZN(n6576) );
  OAI21_X1 U7801 ( .B1(n6592), .B2(n10138), .A(n6576), .ZN(P1_U3342) );
  NOR2_X1 U7802 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n7484), .ZN(n6577) );
  AOI21_X1 U7803 ( .B1(n7484), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6577), .ZN(
        n6580) );
  AOI21_X1 U7804 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7393), .A(n6578), .ZN(
        n6579) );
  NAND2_X1 U7805 ( .A1(n6580), .A2(n6579), .ZN(n6660) );
  OAI21_X1 U7806 ( .B1(n6580), .B2(n6579), .A(n6660), .ZN(n6589) );
  INV_X1 U7807 ( .A(n10542), .ZN(n9617) );
  INV_X1 U7808 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U7809 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n7484), .B1(n6587), .B2(
        n10716), .ZN(n6583) );
  AOI21_X1 U7810 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7393), .A(n6581), .ZN(
        n6582) );
  NAND2_X1 U7811 ( .A1(n6583), .A2(n6582), .ZN(n6664) );
  OAI21_X1 U7812 ( .B1(n6583), .B2(n6582), .A(n6664), .ZN(n6584) );
  INV_X1 U7813 ( .A(n10546), .ZN(n9644) );
  NAND2_X1 U7814 ( .A1(n6584), .A2(n9644), .ZN(n6586) );
  NOR2_X1 U7815 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7403), .ZN(n9460) );
  AOI21_X1 U7816 ( .B1(n10532), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9460), .ZN(
        n6585) );
  OAI211_X1 U7817 ( .C1(n9617), .C2(n6587), .A(n6586), .B(n6585), .ZN(n6588)
         );
  AOI21_X1 U7818 ( .B1(n6589), .B2(n10538), .A(n6588), .ZN(n6590) );
  INV_X1 U7819 ( .A(n6590), .ZN(P1_U3252) );
  INV_X1 U7820 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6591) );
  OAI222_X1 U7821 ( .A1(n5050), .A2(P2_U3151), .B1(n9162), .B2(n6592), .C1(
        n6591), .C2(n9153), .ZN(P2_U3282) );
  NOR2_X1 U7822 ( .A1(n10532), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U7823 ( .A(n6600), .ZN(n8302) );
  NAND2_X1 U7824 ( .A1(n6596), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U7825 ( .A1(n7206), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6604) );
  AND2_X2 U7826 ( .A1(n8302), .A2(n6599), .ZN(n7898) );
  NAND2_X1 U7827 ( .A1(n7898), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U7828 ( .A1(n5558), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U7829 ( .A1(n8054), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6601) );
  AND2_X1 U7830 ( .A1(n6831), .A2(n8227), .ZN(n6607) );
  AND2_X1 U7831 ( .A1(n6969), .A2(n6607), .ZN(n6608) );
  INV_X1 U7832 ( .A(SI_0_), .ZN(n6610) );
  INV_X1 U7833 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6609) );
  OAI21_X1 U7834 ( .B1(n7890), .B2(n6610), .A(n6609), .ZN(n6612) );
  AND2_X1 U7835 ( .A1(n6612), .A2(n6611), .ZN(n10140) );
  MUX2_X1 U7836 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10140), .S(n7392), .Z(n10567)
         );
  NAND2_X1 U7837 ( .A1(n6614), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7005) );
  NAND2_X1 U7838 ( .A1(n7005), .A2(n6615), .ZN(n7007) );
  NAND2_X1 U7839 ( .A1(n7007), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6617) );
  XNOR2_X2 U7840 ( .A(n6617), .B(n6616), .ZN(n9674) );
  NAND2_X1 U7841 ( .A1(n7546), .A2(n8227), .ZN(n6618) );
  NAND2_X1 U7842 ( .A1(n6969), .A2(n6618), .ZN(n9370) );
  AND2_X1 U7843 ( .A1(n10567), .A2(n6725), .ZN(n6619) );
  AOI21_X1 U7844 ( .B1(n6799), .B2(n4948), .A(n6619), .ZN(n6722) );
  INV_X1 U7845 ( .A(n6969), .ZN(n6620) );
  NAND2_X1 U7846 ( .A1(n6620), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U7847 ( .A1(n6722), .A2(n6621), .ZN(n6627) );
  NAND2_X1 U7848 ( .A1(n6799), .A2(n9307), .ZN(n6625) );
  NOR2_X1 U7849 ( .A1(n6969), .A2(n6622), .ZN(n6623) );
  AOI21_X1 U7850 ( .B1(n10567), .B2(n4948), .A(n6623), .ZN(n6624) );
  NAND2_X1 U7851 ( .A1(n6625), .A2(n6624), .ZN(n6626) );
  NAND2_X1 U7852 ( .A1(n6627), .A2(n6626), .ZN(n6724) );
  OAI21_X1 U7853 ( .B1(n6627), .B2(n6626), .A(n6724), .ZN(n9575) );
  INV_X1 U7854 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6629) );
  NOR4_X1 U7855 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6638) );
  NOR4_X1 U7856 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6637) );
  NOR4_X1 U7857 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6633) );
  NOR4_X1 U7858 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6632) );
  NOR4_X1 U7859 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6631) );
  NOR4_X1 U7860 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6630) );
  NAND4_X1 U7861 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .ZN(n6634)
         );
  NOR4_X1 U7862 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n6635), .A4(n6634), .ZN(n6636) );
  NAND3_X1 U7863 ( .A1(n6638), .A2(n6637), .A3(n6636), .ZN(n6639) );
  NAND2_X1 U7864 ( .A1(n6640), .A2(n6639), .ZN(n6815) );
  NAND3_X1 U7865 ( .A1(n6821), .A2(n6827), .A3(n6815), .ZN(n6652) );
  INV_X1 U7866 ( .A(n6652), .ZN(n6644) );
  INV_X1 U7867 ( .A(n6651), .ZN(n6641) );
  INV_X1 U7868 ( .A(n8223), .ZN(n6805) );
  NAND2_X1 U7869 ( .A1(n10765), .A2(n6805), .ZN(n6648) );
  NOR2_X1 U7870 ( .A1(n6641), .A2(n6648), .ZN(n6642) );
  NAND2_X1 U7871 ( .A1(n6651), .A2(n10566), .ZN(n6645) );
  NOR2_X1 U7872 ( .A1(n6645), .A2(n8227), .ZN(n6643) );
  NAND2_X1 U7873 ( .A1(n6644), .A2(n6643), .ZN(n6647) );
  INV_X1 U7874 ( .A(n6645), .ZN(n6646) );
  NAND2_X1 U7875 ( .A1(n6651), .A2(n10555), .ZN(n8296) );
  NAND2_X1 U7876 ( .A1(n6836), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7247) );
  NAND3_X1 U7877 ( .A1(n8296), .A2(n6648), .A3(n7247), .ZN(n6649) );
  AND2_X1 U7878 ( .A1(n6652), .A2(n6649), .ZN(n6972) );
  INV_X1 U7879 ( .A(n6650), .ZN(n8293) );
  NAND2_X1 U7880 ( .A1(n8223), .A2(n8293), .ZN(n6970) );
  NAND2_X1 U7881 ( .A1(n6651), .A2(n6970), .ZN(n6814) );
  OR2_X1 U7882 ( .A1(n6972), .A2(n6814), .ZN(n6860) );
  AOI22_X1 U7883 ( .A1(n9473), .A2(n10567), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n6860), .ZN(n6659) );
  OR2_X1 U7884 ( .A1(n6652), .A2(n8296), .ZN(n6738) );
  INV_X1 U7885 ( .A(n6738), .ZN(n6653) );
  NAND2_X1 U7886 ( .A1(n7898), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U7887 ( .A1(n7206), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U7888 ( .A1(n5558), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U7889 ( .A1(n8054), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6654) );
  NAND4_X1 U7890 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n6798)
         );
  NAND2_X1 U7891 ( .A1(n9496), .A2(n9564), .ZN(n6658) );
  OAI211_X1 U7892 ( .C1(n9575), .C2(n9548), .A(n6659), .B(n6658), .ZN(P1_U3232) );
  OAI21_X1 U7893 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7484), .A(n6660), .ZN(
        n6663) );
  NAND2_X1 U7894 ( .A1(n7512), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6661) );
  OAI21_X1 U7895 ( .B1(n7512), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6661), .ZN(
        n6662) );
  NOR2_X1 U7896 ( .A1(n6663), .A2(n6662), .ZN(n6703) );
  AOI211_X1 U7897 ( .C1(n6663), .C2(n6662), .A(n6703), .B(n9623), .ZN(n6672)
         );
  OAI21_X1 U7898 ( .B1(n7484), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6664), .ZN(
        n6667) );
  INV_X1 U7899 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6665) );
  MUX2_X1 U7900 ( .A(n6665), .B(P1_REG1_REG_10__SCAN_IN), .S(n7512), .Z(n6666)
         );
  NOR2_X1 U7901 ( .A1(n6667), .A2(n6666), .ZN(n6707) );
  AOI211_X1 U7902 ( .C1(n6667), .C2(n6666), .A(n6707), .B(n10546), .ZN(n6671)
         );
  INV_X1 U7903 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U7904 ( .A1(n10542), .A2(n7512), .ZN(n6668) );
  NAND2_X1 U7905 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9353) );
  OAI211_X1 U7906 ( .C1(n6669), .C2(n9669), .A(n6668), .B(n9353), .ZN(n6670)
         );
  OR3_X1 U7907 ( .A1(n6672), .A2(n6671), .A3(n6670), .ZN(P1_U3253) );
  XNOR2_X1 U7908 ( .A(n6674), .B(n6673), .ZN(n6688) );
  NOR2_X1 U7909 ( .A1(n10511), .A2(n6675), .ZN(n6686) );
  INV_X1 U7910 ( .A(n10496), .ZN(n10525) );
  NAND2_X1 U7911 ( .A1(n6677), .A2(n6676), .ZN(n6678) );
  NAND2_X1 U7912 ( .A1(n10525), .A2(n6678), .ZN(n6684) );
  NAND2_X1 U7913 ( .A1(n6679), .A2(n10575), .ZN(n6680) );
  NAND2_X1 U7914 ( .A1(n6681), .A2(n6680), .ZN(n6682) );
  NAND2_X1 U7915 ( .A1(n10492), .A2(n6682), .ZN(n6683) );
  OAI211_X1 U7916 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6795), .A(n6684), .B(n6683), .ZN(n6685) );
  AOI211_X1 U7917 ( .C1(n10516), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6686), .B(
        n6685), .ZN(n6687) );
  OAI21_X1 U7918 ( .B1(n6688), .B2(n10464), .A(n6687), .ZN(P2_U3183) );
  INV_X1 U7919 ( .A(n7780), .ZN(n6695) );
  NAND2_X1 U7920 ( .A1(n6697), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6689) );
  XNOR2_X1 U7921 ( .A(n6689), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7781) );
  AOI22_X1 U7922 ( .A1(n7781), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10126), .ZN(n6690) );
  OAI21_X1 U7923 ( .B1(n6695), .B2(n10138), .A(n6690), .ZN(P1_U3341) );
  INV_X1 U7924 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U7925 ( .A1(n8709), .A2(n6773), .ZN(n8368) );
  NAND2_X1 U7926 ( .A1(n8363), .A2(n8368), .ZN(n9025) );
  OAI21_X1 U7927 ( .B1(n10641), .B2(n10720), .A(n9025), .ZN(n6691) );
  NAND2_X1 U7928 ( .A1(n10591), .A2(n6190), .ZN(n9020) );
  OAI211_X1 U7929 ( .C1(n10799), .C2(n6773), .A(n6691), .B(n9020), .ZN(n6785)
         );
  NAND2_X1 U7930 ( .A1(n6785), .A2(n10810), .ZN(n6692) );
  OAI21_X1 U7931 ( .B1(n10810), .B2(n6693), .A(n6692), .ZN(P2_U3390) );
  OAI222_X1 U7932 ( .A1(n8750), .A2(P2_U3151), .B1(n9162), .B2(n6695), .C1(
        n6694), .C2(n9153), .ZN(P2_U3281) );
  INV_X1 U7933 ( .A(n8022), .ZN(n6701) );
  INV_X1 U7934 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6696) );
  OAI222_X1 U7935 ( .A1(P2_U3151), .A2(n8766), .B1(n9162), .B2(n6701), .C1(
        n6696), .C2(n9153), .ZN(P2_U3280) );
  INV_X1 U7936 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U7937 ( .A1(n6698), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6700) );
  INV_X1 U7938 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U7939 ( .A1(n6700), .A2(n6699), .ZN(n6896) );
  OAI21_X1 U7940 ( .B1(n6700), .B2(n6699), .A(n6896), .ZN(n9618) );
  OAI222_X1 U7941 ( .A1(n10132), .A2(n6702), .B1(n10138), .B2(n6701), .C1(
        n9618), .C2(P1_U3086), .ZN(P1_U3340) );
  AOI21_X1 U7942 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7512), .A(n6703), .ZN(
        n6706) );
  NAND2_X1 U7943 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7611), .ZN(n6704) );
  OAI21_X1 U7944 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7611), .A(n6704), .ZN(
        n6705) );
  NOR2_X1 U7945 ( .A1(n6706), .A2(n6705), .ZN(n6869) );
  AOI211_X1 U7946 ( .C1(n6706), .C2(n6705), .A(n6869), .B(n9623), .ZN(n6715)
         );
  AOI21_X1 U7947 ( .B1(n7512), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6707), .ZN(
        n6710) );
  INV_X1 U7948 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6708) );
  MUX2_X1 U7949 ( .A(n6708), .B(P1_REG1_REG_11__SCAN_IN), .S(n7611), .Z(n6709)
         );
  NOR2_X1 U7950 ( .A1(n6710), .A2(n6709), .ZN(n6872) );
  AOI211_X1 U7951 ( .C1(n6710), .C2(n6709), .A(n6872), .B(n10546), .ZN(n6714)
         );
  INV_X1 U7952 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U7953 ( .A1(n10542), .A2(n7611), .ZN(n6711) );
  NAND2_X1 U7954 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9508) );
  OAI211_X1 U7955 ( .C1(n6712), .C2(n9669), .A(n6711), .B(n9508), .ZN(n6713)
         );
  OR3_X1 U7956 ( .A1(n6715), .A2(n6714), .A3(n6713), .ZN(P1_U3254) );
  NAND2_X1 U7957 ( .A1(n9564), .A2(n9307), .ZN(n6721) );
  OR2_X1 U7958 ( .A1(n6943), .A2(n5044), .ZN(n6718) );
  OAI211_X1 U7959 ( .C1(n7392), .C2(n6719), .A(n6718), .B(n6717), .ZN(n6797)
         );
  NAND2_X1 U7960 ( .A1(n6726), .A2(n4948), .ZN(n6720) );
  NAND2_X1 U7961 ( .A1(n6721), .A2(n6720), .ZN(n6852) );
  INV_X2 U7962 ( .A(n9314), .ZN(n9373) );
  NAND2_X1 U7963 ( .A1(n6722), .A2(n9373), .ZN(n6723) );
  NAND2_X1 U7964 ( .A1(n6724), .A2(n6723), .ZN(n6733) );
  INV_X1 U7965 ( .A(n6733), .ZN(n6731) );
  NAND2_X1 U7966 ( .A1(n6798), .A2(n4948), .ZN(n6728) );
  NAND2_X1 U7967 ( .A1(n6726), .A2(n6725), .ZN(n6727) );
  NAND2_X1 U7968 ( .A1(n6728), .A2(n6727), .ZN(n6729) );
  XNOR2_X1 U7969 ( .A(n6729), .B(n9314), .ZN(n6732) );
  INV_X1 U7970 ( .A(n6732), .ZN(n6730) );
  NAND2_X1 U7971 ( .A1(n6731), .A2(n6730), .ZN(n6853) );
  NAND2_X1 U7972 ( .A1(n6733), .A2(n6732), .ZN(n6854) );
  NAND2_X1 U7973 ( .A1(n6853), .A2(n6854), .ZN(n6734) );
  XOR2_X1 U7974 ( .A(n6852), .B(n6734), .Z(n6741) );
  AOI22_X1 U7975 ( .A1(n9473), .A2(n6726), .B1(n6860), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U7976 ( .A1(n7898), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U7977 ( .A1(n7206), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6735) );
  NAND3_X1 U7978 ( .A1(n6737), .A2(n6736), .A3(n6735), .ZN(n6941) );
  INV_X1 U7979 ( .A(n6983), .ZN(n9563) );
  NOR2_X2 U7980 ( .A1(n6738), .A2(n10135), .ZN(n9539) );
  AOI22_X1 U7981 ( .A1(n9496), .A2(n9563), .B1(n9539), .B2(n6799), .ZN(n6739)
         );
  OAI211_X1 U7982 ( .C1(n6741), .C2(n9548), .A(n6740), .B(n6739), .ZN(P1_U3222) );
  NAND2_X1 U7983 ( .A1(n6759), .A2(n6742), .ZN(n6747) );
  NAND3_X1 U7984 ( .A1(n6744), .A2(n7561), .A3(n6743), .ZN(n6745) );
  AOI21_X1 U7985 ( .B1(n6756), .B2(n6751), .A(n6745), .ZN(n6746) );
  NAND2_X1 U7986 ( .A1(n6747), .A2(n6746), .ZN(n6748) );
  NAND2_X1 U7987 ( .A1(n6748), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6750) );
  NAND2_X1 U7988 ( .A1(n6758), .A2(n9022), .ZN(n6755) );
  INV_X1 U7989 ( .A(n6755), .ZN(n8518) );
  NAND2_X1 U7990 ( .A1(n6756), .A2(n8518), .ZN(n6749) );
  AND2_X2 U7991 ( .A1(n6750), .A2(n6749), .ZN(n8683) );
  INV_X1 U7992 ( .A(n8683), .ZN(n8615) );
  NOR2_X1 U7993 ( .A1(n8615), .A2(P2_U3151), .ZN(n6796) );
  INV_X1 U7994 ( .A(n6751), .ZN(n6752) );
  OAI22_X1 U7995 ( .A1(n6759), .A2(n6753), .B1(n6756), .B2(n6752), .ZN(n6754)
         );
  INV_X1 U7996 ( .A(n10591), .ZN(n6781) );
  NOR2_X1 U7997 ( .A1(n6756), .A2(n6755), .ZN(n6780) );
  INV_X1 U7998 ( .A(n6779), .ZN(n6757) );
  NAND2_X1 U7999 ( .A1(n6758), .A2(n10747), .ZN(n6760) );
  OR2_X1 U8000 ( .A1(n6759), .A2(n6760), .ZN(n6762) );
  OAI22_X1 U8001 ( .A1(n6781), .A2(n8660), .B1(n8689), .B2(n6773), .ZN(n6763)
         );
  AOI21_X1 U8002 ( .B1(n8624), .B2(n9025), .A(n6763), .ZN(n6764) );
  OAI21_X1 U8003 ( .B1(n6796), .B2(n6765), .A(n6764), .ZN(P2_U3172) );
  AND2_X1 U8004 ( .A1(n8362), .A2(n7098), .ZN(n6766) );
  NAND2_X1 U8005 ( .A1(n5487), .A2(n8512), .ZN(n6768) );
  AND2_X4 U8006 ( .A1(n6769), .A2(n6768), .ZN(n7870) );
  XNOR2_X1 U8007 ( .A(n7138), .B(n7870), .ZN(n6771) );
  NAND2_X1 U8008 ( .A1(n6771), .A2(n10591), .ZN(n6772) );
  NAND2_X1 U8009 ( .A1(n6773), .A2(n7874), .ZN(n6774) );
  NAND2_X1 U8010 ( .A1(n6788), .A2(n6789), .ZN(n6787) );
  NAND2_X1 U8011 ( .A1(n6787), .A2(n6775), .ZN(n6776) );
  OAI21_X1 U8012 ( .B1(n6777), .B2(n6776), .A(n6885), .ZN(n6778) );
  NAND2_X1 U8013 ( .A1(n6778), .A2(n8624), .ZN(n6784) );
  NAND2_X1 U8014 ( .A1(n6780), .A2(n6779), .ZN(n8680) );
  OAI22_X1 U8015 ( .A1(n6781), .A2(n8680), .B1(n8689), .B2(n10599), .ZN(n6782)
         );
  AOI21_X1 U8016 ( .B1(n8686), .B2(n10592), .A(n6782), .ZN(n6783) );
  OAI211_X1 U8017 ( .C1(n6796), .C2(n10597), .A(n6784), .B(n6783), .ZN(
        P2_U3177) );
  NAND2_X1 U8018 ( .A1(n6785), .A2(n10806), .ZN(n6786) );
  OAI21_X1 U8019 ( .B1(n10806), .B2(n6317), .A(n6786), .ZN(P2_U3459) );
  OAI21_X1 U8020 ( .B1(n6789), .B2(n6788), .A(n6787), .ZN(n6790) );
  NAND2_X1 U8021 ( .A1(n6790), .A2(n8624), .ZN(n6794) );
  INV_X1 U8022 ( .A(n8709), .ZN(n6791) );
  OAI22_X1 U8023 ( .A1(n6791), .A2(n8680), .B1(n8689), .B2(n10571), .ZN(n6792)
         );
  AOI21_X1 U8024 ( .B1(n8686), .B2(n8708), .A(n6792), .ZN(n6793) );
  OAI211_X1 U8025 ( .C1(n6796), .C2(n6795), .A(n6794), .B(n6793), .ZN(P2_U3162) );
  INV_X1 U8026 ( .A(n10553), .ZN(n6812) );
  INV_X1 U8027 ( .A(n7316), .ZN(n10693) );
  NAND2_X1 U8028 ( .A1(n6799), .A2(n10567), .ZN(n6801) );
  NAND2_X1 U8029 ( .A1(n6800), .A2(n6801), .ZN(n6940) );
  OAI21_X1 U8030 ( .B1(n6800), .B2(n6801), .A(n6940), .ZN(n6811) );
  AOI211_X1 U8031 ( .C1(n10567), .C2(n6726), .A(n9915), .B(n7085), .ZN(n6839)
         );
  INV_X1 U8032 ( .A(n6811), .ZN(n6842) );
  NAND2_X1 U8033 ( .A1(n6613), .A2(n9674), .ZN(n6802) );
  NAND2_X1 U8034 ( .A1(n6802), .A2(n8293), .ZN(n6803) );
  NAND2_X1 U8035 ( .A1(n6803), .A2(n10556), .ZN(n6804) );
  OR2_X1 U8036 ( .A1(n10555), .A2(n6804), .ZN(n7629) );
  AOI22_X1 U8037 ( .A1(n10759), .A2(n6799), .B1(n9563), .B2(n10756), .ZN(n6810) );
  INV_X1 U8038 ( .A(n10567), .ZN(n10554) );
  NOR2_X1 U8039 ( .A1(n6799), .A2(n10554), .ZN(n6806) );
  NAND2_X1 U8040 ( .A1(n8029), .A2(n6806), .ZN(n6956) );
  OAI21_X1 U8041 ( .B1(n8029), .B2(n6806), .A(n6956), .ZN(n6808) );
  NAND2_X1 U8042 ( .A1(n6613), .A2(n9671), .ZN(n8186) );
  NAND2_X1 U8043 ( .A1(n6808), .A2(n10752), .ZN(n6809) );
  OAI211_X1 U8044 ( .C1(n6842), .C2(n7629), .A(n6810), .B(n6809), .ZN(n6833)
         );
  AOI211_X1 U8045 ( .C1(n10693), .C2(n6811), .A(n6839), .B(n6833), .ZN(n6826)
         );
  NOR2_X1 U8046 ( .A1(n10556), .A2(n6812), .ZN(n6813) );
  NOR2_X1 U8047 ( .A1(n6827), .A2(n6813), .ZN(n6817) );
  INV_X1 U8048 ( .A(n6814), .ZN(n6816) );
  INV_X1 U8049 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6818) );
  OAI22_X1 U8050 ( .A1(n10069), .A2(n6938), .B1(n10770), .B2(n6818), .ZN(n6819) );
  INV_X1 U8051 ( .A(n6819), .ZN(n6820) );
  OAI21_X1 U8052 ( .B1(n6826), .B2(n10768), .A(n6820), .ZN(P1_U3523) );
  INV_X1 U8053 ( .A(n6821), .ZN(n6828) );
  INV_X1 U8054 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6823) );
  OAI22_X1 U8055 ( .A1(n10122), .A2(n6938), .B1(n10774), .B2(n6823), .ZN(n6824) );
  INV_X1 U8056 ( .A(n6824), .ZN(n6825) );
  OAI21_X1 U8057 ( .B1(n6826), .B2(n10771), .A(n6825), .ZN(P1_U3456) );
  NAND3_X1 U8058 ( .A1(n6829), .A2(n6828), .A3(n6827), .ZN(n6830) );
  AND2_X1 U8059 ( .A1(n10553), .A2(n6831), .ZN(n6832) );
  NAND2_X1 U8060 ( .A1(n10560), .A2(n6832), .ZN(n7635) );
  NAND2_X1 U8061 ( .A1(n6833), .A2(n10560), .ZN(n6841) );
  AND2_X2 U8062 ( .A1(n10560), .A2(n9674), .ZN(n9972) );
  INV_X1 U8063 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6835) );
  INV_X1 U8064 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6834) );
  OAI22_X1 U8065 ( .A1(n10560), .A2(n6835), .B1(n6834), .B2(n7126), .ZN(n6838)
         );
  NAND3_X2 U8066 ( .A1(n10560), .A2(n10566), .A3(n6836), .ZN(n9976) );
  NOR2_X1 U8067 ( .A1(n9976), .A2(n6938), .ZN(n6837) );
  AOI211_X1 U8068 ( .C1(n6839), .C2(n9972), .A(n6838), .B(n6837), .ZN(n6840)
         );
  OAI211_X1 U8069 ( .C1(n6842), .C2(n7635), .A(n6841), .B(n6840), .ZN(P1_U3292) );
  NAND2_X1 U8070 ( .A1(n6941), .A2(n4948), .ZN(n6849) );
  OR2_X1 U8071 ( .A1(n7394), .A2(n6843), .ZN(n6846) );
  OR2_X1 U8072 ( .A1(n6943), .A2(n6844), .ZN(n6845) );
  NAND2_X1 U8073 ( .A1(n8079), .A2(n6725), .ZN(n6848) );
  NAND2_X1 U8074 ( .A1(n6849), .A2(n6848), .ZN(n6850) );
  XNOR2_X1 U8075 ( .A(n6850), .B(n9373), .ZN(n6975) );
  AND2_X1 U8076 ( .A1(n8079), .A2(n4948), .ZN(n6851) );
  AOI21_X1 U8077 ( .B1(n9563), .B2(n9307), .A(n6851), .ZN(n6974) );
  XNOR2_X1 U8078 ( .A(n6975), .B(n6974), .ZN(n6859) );
  NAND2_X1 U8079 ( .A1(n6853), .A2(n6852), .ZN(n6855) );
  NAND2_X1 U8080 ( .A1(n6855), .A2(n6854), .ZN(n6858) );
  INV_X1 U8081 ( .A(n6859), .ZN(n6856) );
  INV_X1 U8082 ( .A(n6977), .ZN(n6857) );
  AOI21_X1 U8083 ( .B1(n6859), .B2(n6858), .A(n6857), .ZN(n6867) );
  AOI22_X1 U8084 ( .A1(n9473), .A2(n8079), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6860), .ZN(n6866) );
  NAND2_X1 U8085 ( .A1(n5558), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6863) );
  INV_X1 U8086 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U8087 ( .A1(n8054), .A2(n6949), .ZN(n6861) );
  AOI22_X1 U8088 ( .A1(n9496), .A2(n9562), .B1(n9539), .B2(n9564), .ZN(n6865)
         );
  OAI211_X1 U8089 ( .C1(n6867), .C2(n9548), .A(n6866), .B(n6865), .ZN(P1_U3237) );
  NOR2_X1 U8090 ( .A1(n7704), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6868) );
  AOI21_X1 U8091 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7704), .A(n6868), .ZN(
        n6871) );
  AOI21_X1 U8092 ( .B1(n7611), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6869), .ZN(
        n6870) );
  NAND2_X1 U8093 ( .A1(n6871), .A2(n6870), .ZN(n7053) );
  OAI21_X1 U8094 ( .B1(n6871), .B2(n6870), .A(n7053), .ZN(n6880) );
  INV_X1 U8095 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U8096 ( .A1(n7704), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n10769), .B2(
        n6878), .ZN(n6874) );
  AOI21_X1 U8097 ( .B1(n7611), .B2(P1_REG1_REG_11__SCAN_IN), .A(n6872), .ZN(
        n6873) );
  NAND2_X1 U8098 ( .A1(n6874), .A2(n6873), .ZN(n7057) );
  OAI21_X1 U8099 ( .B1(n6874), .B2(n6873), .A(n7057), .ZN(n6875) );
  NAND2_X1 U8100 ( .A1(n6875), .A2(n9644), .ZN(n6877) );
  AND2_X1 U8101 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9412) );
  AOI21_X1 U8102 ( .B1(n10532), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9412), .ZN(
        n6876) );
  OAI211_X1 U8103 ( .C1(n9617), .C2(n6878), .A(n6877), .B(n6876), .ZN(n6879)
         );
  AOI21_X1 U8104 ( .B1(n6880), .B2(n10538), .A(n6879), .ZN(n6881) );
  INV_X1 U8105 ( .A(n6881), .ZN(P1_U3255) );
  INV_X1 U8106 ( .A(n8708), .ZN(n6883) );
  NAND2_X1 U8107 ( .A1(n6883), .A2(n6882), .ZN(n6884) );
  NAND2_X1 U8108 ( .A1(n6885), .A2(n6884), .ZN(n6887) );
  XNOR2_X1 U8109 ( .A(n6886), .B(n7870), .ZN(n6901) );
  XNOR2_X1 U8110 ( .A(n6901), .B(n10592), .ZN(n6888) );
  AOI21_X1 U8111 ( .B1(n6887), .B2(n6888), .A(n8676), .ZN(n6891) );
  INV_X1 U8112 ( .A(n6887), .ZN(n6890) );
  NAND2_X1 U8113 ( .A1(n6891), .A2(n6903), .ZN(n6895) );
  INV_X1 U8114 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10244) );
  NOR2_X1 U8115 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10244), .ZN(n10450) );
  INV_X1 U8116 ( .A(n10636), .ZN(n6892) );
  OAI22_X1 U8117 ( .A1(n6892), .A2(n8660), .B1(n8689), .B2(n10605), .ZN(n6893)
         );
  AOI211_X1 U8118 ( .C1(n8663), .C2(n8708), .A(n10450), .B(n6893), .ZN(n6894)
         );
  OAI211_X1 U8119 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8683), .A(n6895), .B(
        n6894), .ZN(P2_U3158) );
  INV_X1 U8120 ( .A(n8011), .ZN(n6900) );
  NAND2_X1 U8121 ( .A1(n6896), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6897) );
  XNOR2_X1 U8122 ( .A(n6897), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9636) );
  INV_X1 U8123 ( .A(n9636), .ZN(n9616) );
  OAI222_X1 U8124 ( .A1(n10132), .A2(n6898), .B1(n10138), .B2(n6900), .C1(
        P1_U3086), .C2(n9616), .ZN(P1_U3339) );
  OAI222_X1 U8125 ( .A1(n8784), .A2(P2_U3151), .B1(n9162), .B2(n6900), .C1(
        n6899), .C2(n9153), .ZN(P2_U3279) );
  NAND2_X1 U8126 ( .A1(n6901), .A2(n10592), .ZN(n6902) );
  XNOR2_X1 U8127 ( .A(n6904), .B(n7870), .ZN(n6905) );
  OR2_X1 U8128 ( .A1(n6905), .A2(n10636), .ZN(n7015) );
  NAND2_X1 U8129 ( .A1(n6905), .A2(n10636), .ZN(n6906) );
  AND2_X1 U8130 ( .A1(n7015), .A2(n6906), .ZN(n6907) );
  OAI21_X1 U8131 ( .B1(n5036), .B2(n6907), .A(n7016), .ZN(n6908) );
  NAND2_X1 U8132 ( .A1(n6908), .A2(n8624), .ZN(n6912) );
  NAND2_X1 U8133 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10483) );
  INV_X1 U8134 ( .A(n10483), .ZN(n6910) );
  INV_X1 U8135 ( .A(n8707), .ZN(n7253) );
  OAI22_X1 U8136 ( .A1(n7253), .A2(n8660), .B1(n8689), .B2(n10612), .ZN(n6909)
         );
  AOI211_X1 U8137 ( .C1(n8663), .C2(n10592), .A(n6910), .B(n6909), .ZN(n6911)
         );
  OAI211_X1 U8138 ( .C1(n7103), .C2(n8683), .A(n6912), .B(n6911), .ZN(P2_U3170) );
  INV_X1 U8139 ( .A(n8001), .ZN(n6917) );
  OAI222_X1 U8140 ( .A1(P2_U3151), .A2(n8799), .B1(n9162), .B2(n6917), .C1(
        n6913), .C2(n9153), .ZN(P2_U3278) );
  NAND2_X1 U8141 ( .A1(n6914), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6915) );
  XNOR2_X1 U8142 ( .A(n6915), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9634) );
  INV_X1 U8143 ( .A(n9634), .ZN(n9654) );
  OAI222_X1 U8144 ( .A1(P1_U3086), .A2(n9654), .B1(n10138), .B2(n6917), .C1(
        n6916), .C2(n10132), .ZN(P1_U3338) );
  NOR2_X1 U8145 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n6918) );
  AOI21_X1 U8146 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n6918), .ZN(n10428) );
  INV_X1 U8147 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9632) );
  INV_X1 U8148 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n6919) );
  AOI22_X1 U8149 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n9632), .B2(n6919), .ZN(n10425) );
  NOR2_X1 U8150 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6920) );
  AOI21_X1 U8151 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6920), .ZN(n10422) );
  NOR2_X1 U8152 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6921) );
  AOI21_X1 U8153 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6921), .ZN(n10419) );
  NOR2_X1 U8154 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6922) );
  AOI21_X1 U8155 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6922), .ZN(n10416) );
  NOR2_X1 U8156 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6923) );
  AOI21_X1 U8157 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6923), .ZN(n10413) );
  NOR2_X1 U8158 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6924) );
  AOI21_X1 U8159 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6924), .ZN(n10410) );
  NOR2_X1 U8160 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n6925) );
  AOI21_X1 U8161 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6925), .ZN(n10407) );
  NOR2_X1 U8162 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n6926) );
  AOI21_X1 U8163 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6926), .ZN(n10404) );
  NOR2_X1 U8164 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n6927) );
  AOI21_X1 U8165 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n6927), .ZN(n10401) );
  NOR2_X1 U8166 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n6928) );
  AOI21_X1 U8167 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n6928), .ZN(n10398) );
  NOR2_X1 U8168 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n6929) );
  AOI21_X1 U8169 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n6929), .ZN(n10395) );
  NOR2_X1 U8170 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n6930) );
  AOI21_X1 U8171 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n6930), .ZN(n10392) );
  NOR2_X1 U8172 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n6931) );
  AOI21_X1 U8173 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n6931), .ZN(n10389) );
  AND2_X1 U8174 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n6932) );
  NOR2_X1 U8175 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n6932), .ZN(n10374) );
  INV_X1 U8176 ( .A(n10374), .ZN(n10375) );
  INV_X1 U8177 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10377) );
  NAND3_X1 U8178 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10376) );
  NAND2_X1 U8179 ( .A1(n10377), .A2(n10376), .ZN(n10373) );
  NAND2_X1 U8180 ( .A1(n10375), .A2(n10373), .ZN(n10380) );
  NAND2_X1 U8181 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n6933) );
  OAI21_X1 U8182 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n6933), .ZN(n10379) );
  NOR2_X1 U8183 ( .A1(n10380), .A2(n10379), .ZN(n10378) );
  AOI21_X1 U8184 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10378), .ZN(n10383) );
  NAND2_X1 U8185 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n6934) );
  OAI21_X1 U8186 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n6934), .ZN(n10382) );
  NOR2_X1 U8187 ( .A1(n10383), .A2(n10382), .ZN(n10381) );
  AOI21_X1 U8188 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10381), .ZN(n10386) );
  NOR2_X1 U8189 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6935) );
  AOI21_X1 U8190 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n6935), .ZN(n10385) );
  NAND2_X1 U8191 ( .A1(n10386), .A2(n10385), .ZN(n10384) );
  OAI21_X1 U8192 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10384), .ZN(n10388) );
  NAND2_X1 U8193 ( .A1(n10389), .A2(n10388), .ZN(n10387) );
  OAI21_X1 U8194 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10387), .ZN(n10391) );
  NAND2_X1 U8195 ( .A1(n10392), .A2(n10391), .ZN(n10390) );
  OAI21_X1 U8196 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10390), .ZN(n10394) );
  NAND2_X1 U8197 ( .A1(n10395), .A2(n10394), .ZN(n10393) );
  OAI21_X1 U8198 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10393), .ZN(n10397) );
  NAND2_X1 U8199 ( .A1(n10398), .A2(n10397), .ZN(n10396) );
  OAI21_X1 U8200 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10396), .ZN(n10400) );
  NAND2_X1 U8201 ( .A1(n10401), .A2(n10400), .ZN(n10399) );
  OAI21_X1 U8202 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10399), .ZN(n10403) );
  NAND2_X1 U8203 ( .A1(n10404), .A2(n10403), .ZN(n10402) );
  OAI21_X1 U8204 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10402), .ZN(n10406) );
  NAND2_X1 U8205 ( .A1(n10407), .A2(n10406), .ZN(n10405) );
  OAI21_X1 U8206 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10405), .ZN(n10409) );
  NAND2_X1 U8207 ( .A1(n10410), .A2(n10409), .ZN(n10408) );
  OAI21_X1 U8208 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10408), .ZN(n10412) );
  NAND2_X1 U8209 ( .A1(n10413), .A2(n10412), .ZN(n10411) );
  OAI21_X1 U8210 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10411), .ZN(n10415) );
  NAND2_X1 U8211 ( .A1(n10416), .A2(n10415), .ZN(n10414) );
  OAI21_X1 U8212 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10414), .ZN(n10418) );
  NAND2_X1 U8213 ( .A1(n10419), .A2(n10418), .ZN(n10417) );
  OAI21_X1 U8214 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10417), .ZN(n10421) );
  NAND2_X1 U8215 ( .A1(n10422), .A2(n10421), .ZN(n10420) );
  OAI21_X1 U8216 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10420), .ZN(n10424) );
  NAND2_X1 U8217 ( .A1(n10425), .A2(n10424), .ZN(n10423) );
  OAI21_X1 U8218 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10423), .ZN(n10427) );
  NAND2_X1 U8219 ( .A1(n10428), .A2(n10427), .ZN(n10426) );
  OAI21_X1 U8220 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10426), .ZN(n6937) );
  XNOR2_X1 U8221 ( .A(n5245), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n6936) );
  XNOR2_X1 U8222 ( .A(n6937), .B(n6936), .ZN(ADD_1068_U4) );
  NAND2_X1 U8223 ( .A1(n10552), .A2(n6938), .ZN(n6939) );
  NAND2_X1 U8224 ( .A1(n6940), .A2(n6939), .ZN(n7082) );
  NAND2_X1 U8225 ( .A1(n6941), .A2(n10578), .ZN(n8085) );
  NAND2_X1 U8226 ( .A1(n8232), .A2(n8085), .ZN(n6957) );
  NAND2_X1 U8227 ( .A1(n7082), .A2(n6957), .ZN(n7081) );
  NAND2_X1 U8228 ( .A1(n6983), .A2(n10578), .ZN(n8081) );
  NAND2_X1 U8229 ( .A1(n7081), .A2(n8081), .ZN(n6948) );
  OR2_X1 U8230 ( .A1(n7394), .A2(n6942), .ZN(n6946) );
  OR2_X1 U8231 ( .A1(n6943), .A2(n6944), .ZN(n6945) );
  OAI211_X1 U8232 ( .C1(n7392), .C2(n6947), .A(n6946), .B(n6945), .ZN(n6986)
         );
  NAND2_X1 U8233 ( .A1(n7119), .A2(n6986), .ZN(n8088) );
  INV_X1 U8234 ( .A(n6986), .ZN(n7118) );
  NAND2_X1 U8235 ( .A1(n9562), .A2(n7118), .ZN(n8083) );
  NAND2_X1 U8236 ( .A1(n8088), .A2(n8083), .ZN(n6959) );
  NAND2_X1 U8237 ( .A1(n6948), .A2(n6959), .ZN(n7121) );
  OAI21_X1 U8238 ( .B1(n6948), .B2(n6959), .A(n7121), .ZN(n7066) );
  NAND2_X1 U8239 ( .A1(n7206), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U8240 ( .A1(n7898), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6953) );
  INV_X1 U8241 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7041) );
  NAND2_X1 U8242 ( .A1(n6949), .A2(n7041), .ZN(n6950) );
  AND2_X1 U8243 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7042) );
  INV_X1 U8244 ( .A(n7042), .ZN(n7044) );
  AND2_X1 U8245 ( .A1(n6950), .A2(n7044), .ZN(n7024) );
  NAND2_X1 U8246 ( .A1(n8054), .A2(n7024), .ZN(n6952) );
  NAND2_X1 U8247 ( .A1(n5558), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6951) );
  NAND4_X1 U8248 ( .A1(n6954), .A2(n6953), .A3(n6952), .A4(n6951), .ZN(n9561)
         );
  OAI22_X1 U8249 ( .A1(n6983), .A2(n9949), .B1(n7272), .B2(n10551), .ZN(n6962)
         );
  NAND2_X1 U8250 ( .A1(n10552), .A2(n6726), .ZN(n6955) );
  INV_X1 U8251 ( .A(n6957), .ZN(n8030) );
  NAND2_X1 U8252 ( .A1(n7077), .A2(n8232), .ZN(n6958) );
  INV_X1 U8253 ( .A(n6959), .ZN(n8031) );
  NAND3_X1 U8254 ( .A1(n7077), .A2(n6959), .A3(n8232), .ZN(n6960) );
  AOI21_X1 U8255 ( .B1(n7123), .B2(n6960), .A(n10563), .ZN(n6961) );
  AOI211_X1 U8256 ( .C1(n7400), .C2(n7066), .A(n6962), .B(n6961), .ZN(n7068)
         );
  INV_X2 U8257 ( .A(n10560), .ZN(n10786) );
  INV_X1 U8258 ( .A(n7635), .ZN(n7421) );
  INV_X1 U8259 ( .A(n9972), .ZN(n10658) );
  NAND2_X1 U8260 ( .A1(n7085), .A2(n10578), .ZN(n7084) );
  INV_X1 U8261 ( .A(n7084), .ZN(n6963) );
  OR2_X1 U8262 ( .A1(n7084), .A2(n6986), .ZN(n7125) );
  OAI211_X1 U8263 ( .C1(n6963), .C2(n7118), .A(n10762), .B(n7125), .ZN(n7067)
         );
  INV_X1 U8264 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6964) );
  OAI22_X1 U8265 ( .A1(n10560), .A2(n6964), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n7126), .ZN(n6965) );
  AOI21_X1 U8266 ( .B1(n10777), .B2(n6986), .A(n6965), .ZN(n6966) );
  OAI21_X1 U8267 ( .B1(n10658), .B2(n7067), .A(n6966), .ZN(n6967) );
  AOI21_X1 U8268 ( .B1(n7066), .B2(n7421), .A(n6967), .ZN(n6968) );
  OAI21_X1 U8269 ( .B1(n7068), .B2(n10786), .A(n6968), .ZN(P1_U3290) );
  NAND3_X1 U8270 ( .A1(n6970), .A2(n7559), .A3(n6969), .ZN(n6971) );
  OR2_X1 U8271 ( .A1(n6972), .A2(n6971), .ZN(n6973) );
  NAND2_X1 U8272 ( .A1(n6973), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7446) );
  NAND2_X1 U8273 ( .A1(n6975), .A2(n6974), .ZN(n6976) );
  NAND2_X1 U8274 ( .A1(n9562), .A2(n4948), .ZN(n6979) );
  NAND2_X1 U8275 ( .A1(n6986), .A2(n6725), .ZN(n6978) );
  NAND2_X1 U8276 ( .A1(n6979), .A2(n6978), .ZN(n6980) );
  XNOR2_X1 U8277 ( .A(n6980), .B(n9314), .ZN(n7025) );
  AND2_X1 U8278 ( .A1(n6986), .A2(n4948), .ZN(n6981) );
  AOI21_X1 U8279 ( .B1(n9562), .B2(n9307), .A(n6981), .ZN(n7026) );
  XNOR2_X1 U8280 ( .A(n7025), .B(n7026), .ZN(n7028) );
  XNOR2_X1 U8281 ( .A(n7029), .B(n7028), .ZN(n6982) );
  NAND2_X1 U8282 ( .A1(n6982), .A2(n9529), .ZN(n6988) );
  NAND2_X1 U8283 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9596) );
  INV_X1 U8284 ( .A(n9596), .ZN(n6985) );
  OAI22_X1 U8285 ( .A1(n9498), .A2(n6983), .B1(n7272), .B2(n9542), .ZN(n6984)
         );
  AOI211_X1 U8286 ( .C1(n6986), .C2(n9473), .A(n6985), .B(n6984), .ZN(n6987)
         );
  OAI211_X1 U8287 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n7446), .A(n6988), .B(
        n6987), .ZN(P1_U3218) );
  AOI21_X1 U8288 ( .B1(n6312), .B2(n6990), .A(n6989), .ZN(n7004) );
  AOI21_X1 U8289 ( .B1(n6313), .B2(n6992), .A(n6991), .ZN(n6993) );
  NOR2_X1 U8290 ( .A1(n6993), .A2(n10496), .ZN(n7002) );
  AOI21_X1 U8291 ( .B1(n6996), .B2(n6995), .A(n6994), .ZN(n7000) );
  INV_X1 U8292 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10317) );
  NOR2_X1 U8293 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10317), .ZN(n7296) );
  AOI21_X1 U8294 ( .B1(n10516), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7296), .ZN(
        n6999) );
  INV_X1 U8295 ( .A(n10511), .ZN(n10434) );
  NAND2_X1 U8296 ( .A1(n10434), .A2(n6997), .ZN(n6998) );
  OAI211_X1 U8297 ( .C1(n7000), .C2(n10464), .A(n6999), .B(n6998), .ZN(n7001)
         );
  NOR2_X1 U8298 ( .A1(n7002), .A2(n7001), .ZN(n7003) );
  OAI21_X1 U8299 ( .B1(n7004), .B2(n10514), .A(n7003), .ZN(P2_U3189) );
  INV_X1 U8300 ( .A(n7005), .ZN(n7006) );
  NAND2_X1 U8301 ( .A1(n7006), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n7008) );
  AND2_X1 U8302 ( .A1(n7008), .A2(n7007), .ZN(n9650) );
  INV_X1 U8303 ( .A(n9650), .ZN(n9643) );
  INV_X1 U8304 ( .A(n8044), .ZN(n7011) );
  INV_X1 U8305 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7009) );
  OAI222_X1 U8306 ( .A1(P1_U3086), .A2(n9643), .B1(n10138), .B2(n7011), .C1(
        n7009), .C2(n10132), .ZN(P1_U3337) );
  INV_X1 U8307 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7012) );
  OAI222_X1 U8308 ( .A1(n9153), .A2(n7012), .B1(n9162), .B2(n7011), .C1(
        P2_U3151), .C2(n7010), .ZN(P2_U3277) );
  INV_X1 U8309 ( .A(n7016), .ZN(n7014) );
  XNOR2_X1 U8310 ( .A(n7013), .B(n7874), .ZN(n7252) );
  XNOR2_X1 U8311 ( .A(n7252), .B(n8707), .ZN(n7017) );
  NOR3_X1 U8312 ( .A1(n7014), .A2(n5332), .A3(n7017), .ZN(n7020) );
  NAND2_X1 U8313 ( .A1(n7018), .A2(n7017), .ZN(n7255) );
  INV_X1 U8314 ( .A(n7255), .ZN(n7019) );
  OAI21_X1 U8315 ( .B1(n7020), .B2(n7019), .A(n8624), .ZN(n7023) );
  NOR2_X1 U8316 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5814), .ZN(n10493) );
  INV_X1 U8317 ( .A(n10635), .ZN(n7307) );
  OAI22_X1 U8318 ( .A1(n7307), .A2(n8660), .B1(n8689), .B2(n10652), .ZN(n7021)
         );
  AOI211_X1 U8319 ( .C1(n8663), .C2(n10636), .A(n10493), .B(n7021), .ZN(n7022)
         );
  OAI211_X1 U8320 ( .C1(n10651), .C2(n8683), .A(n7023), .B(n7022), .ZN(
        P2_U3167) );
  INV_X1 U8321 ( .A(n7024), .ZN(n7127) );
  INV_X1 U8322 ( .A(n7025), .ZN(n7027) );
  NAND2_X1 U8323 ( .A1(n9561), .A2(n4948), .ZN(n7036) );
  OR2_X1 U8324 ( .A1(n7394), .A2(n7030), .ZN(n7033) );
  OR2_X1 U8325 ( .A1(n6943), .A2(n7031), .ZN(n7032) );
  OAI211_X1 U8326 ( .C1(n7392), .C2(n7034), .A(n7033), .B(n7032), .ZN(n10618)
         );
  NAND2_X1 U8327 ( .A1(n10618), .A2(n6725), .ZN(n7035) );
  NAND2_X1 U8328 ( .A1(n7036), .A2(n7035), .ZN(n7037) );
  XNOR2_X1 U8329 ( .A(n7037), .B(n9314), .ZN(n7191) );
  AND2_X1 U8330 ( .A1(n10618), .A2(n4948), .ZN(n7038) );
  AOI21_X1 U8331 ( .B1(n9561), .B2(n9307), .A(n7038), .ZN(n7189) );
  XNOR2_X1 U8332 ( .A(n7191), .B(n7189), .ZN(n7039) );
  NAND2_X1 U8333 ( .A1(n7040), .A2(n7039), .ZN(n7193) );
  OAI211_X1 U8334 ( .C1(n7040), .C2(n7039), .A(n7193), .B(n9529), .ZN(n7052)
         );
  NOR2_X1 U8335 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7041), .ZN(n10531) );
  NAND2_X1 U8336 ( .A1(n7206), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7049) );
  NAND2_X1 U8337 ( .A1(n7898), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7048) );
  NAND2_X1 U8338 ( .A1(n7042), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7208) );
  INV_X1 U8339 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7043) );
  NAND2_X1 U8340 ( .A1(n7044), .A2(n7043), .ZN(n7045) );
  AND2_X1 U8341 ( .A1(n7208), .A2(n7045), .ZN(n10660) );
  NAND2_X1 U8342 ( .A1(n8054), .A2(n10660), .ZN(n7047) );
  NAND2_X1 U8343 ( .A1(n5558), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7046) );
  INV_X1 U8344 ( .A(n9560), .ZN(n7270) );
  OAI22_X1 U8345 ( .A1(n9498), .A2(n7119), .B1(n7270), .B2(n9542), .ZN(n7050)
         );
  AOI211_X1 U8346 ( .C1(n10618), .C2(n9473), .A(n10531), .B(n7050), .ZN(n7051)
         );
  OAI211_X1 U8347 ( .C1(n7446), .C2(n7127), .A(n7052), .B(n7051), .ZN(P1_U3230) );
  OAI21_X1 U8348 ( .B1(n7704), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7053), .ZN(
        n7056) );
  NAND2_X1 U8349 ( .A1(n7708), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7054) );
  OAI21_X1 U8350 ( .B1(n7708), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7054), .ZN(
        n7055) );
  NOR2_X1 U8351 ( .A1(n7055), .A2(n7056), .ZN(n7177) );
  AOI211_X1 U8352 ( .C1(n7056), .C2(n7055), .A(n7177), .B(n9623), .ZN(n7065)
         );
  OAI21_X1 U8353 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n7704), .A(n7057), .ZN(
        n7060) );
  INV_X1 U8354 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7058) );
  MUX2_X1 U8355 ( .A(n7058), .B(P1_REG1_REG_13__SCAN_IN), .S(n7708), .Z(n7059)
         );
  NOR2_X1 U8356 ( .A1(n7059), .A2(n7060), .ZN(n7181) );
  AOI211_X1 U8357 ( .C1(n7060), .C2(n7059), .A(n7181), .B(n10546), .ZN(n7064)
         );
  INV_X1 U8358 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7062) );
  NAND2_X1 U8359 ( .A1(n10542), .A2(n7708), .ZN(n7061) );
  NAND2_X1 U8360 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9481) );
  OAI211_X1 U8361 ( .C1(n7062), .C2(n9669), .A(n7061), .B(n9481), .ZN(n7063)
         );
  OR3_X1 U8362 ( .A1(n7065), .A2(n7064), .A3(n7063), .ZN(P1_U3256) );
  INV_X1 U8363 ( .A(n7066), .ZN(n7069) );
  OAI211_X1 U8364 ( .C1(n7069), .C2(n7316), .A(n7068), .B(n7067), .ZN(n7075)
         );
  INV_X1 U8365 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7070) );
  OAI22_X1 U8366 ( .A1(n10122), .A2(n7118), .B1(n10774), .B2(n7070), .ZN(n7071) );
  AOI21_X1 U8367 ( .B1(n7075), .B2(n10774), .A(n7071), .ZN(n7072) );
  INV_X1 U8368 ( .A(n7072), .ZN(P1_U3462) );
  INV_X1 U8369 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7073) );
  OAI22_X1 U8370 ( .A1(n10069), .A2(n7118), .B1(n10770), .B2(n7073), .ZN(n7074) );
  AOI21_X1 U8371 ( .B1(n7075), .B2(n10770), .A(n7074), .ZN(n7076) );
  INV_X1 U8372 ( .A(n7076), .ZN(P1_U3525) );
  INV_X2 U8373 ( .A(n7126), .ZN(n10775) );
  INV_X1 U8374 ( .A(n8092), .ZN(n7079) );
  INV_X1 U8375 ( .A(n7077), .ZN(n7078) );
  AOI21_X1 U8376 ( .B1(n7079), .B2(n6957), .A(n7078), .ZN(n7080) );
  OAI222_X1 U8377 ( .A1(n10551), .A2(n7119), .B1(n9949), .B2(n10552), .C1(
        n10563), .C2(n7080), .ZN(n10579) );
  AOI21_X1 U8378 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n10775), .A(n10579), .ZN(
        n7089) );
  OAI21_X1 U8379 ( .B1(n7082), .B2(n6957), .A(n7081), .ZN(n10581) );
  NAND2_X1 U8380 ( .A1(n10560), .A2(n7400), .ZN(n7083) );
  OAI211_X1 U8381 ( .C1(n7085), .C2(n10578), .A(n7084), .B(n10762), .ZN(n10577) );
  AOI22_X1 U8382 ( .A1(n10777), .A2(n8079), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n10786), .ZN(n7086) );
  OAI21_X1 U8383 ( .B1(n10658), .B2(n10577), .A(n7086), .ZN(n7087) );
  AOI21_X1 U8384 ( .B1(n10581), .B2(n10781), .A(n7087), .ZN(n7088) );
  OAI21_X1 U8385 ( .B1(n7089), .B2(n10786), .A(n7088), .ZN(P1_U3291) );
  XNOR2_X1 U8386 ( .A(n7090), .B(n8377), .ZN(n10614) );
  INV_X1 U8387 ( .A(n10614), .ZN(n7108) );
  INV_X1 U8388 ( .A(n7091), .ZN(n7097) );
  AOI22_X1 U8389 ( .A1(n7095), .A2(n7094), .B1(n7093), .B2(n7092), .ZN(n7096)
         );
  OR2_X1 U8390 ( .A1(n8362), .A2(n7098), .ZN(n10648) );
  INV_X1 U8391 ( .A(n10648), .ZN(n8832) );
  OR2_X1 U8392 ( .A1(n10634), .A2(n8832), .ZN(n10700) );
  AOI21_X1 U8393 ( .B1(n7099), .B2(n8377), .A(n9000), .ZN(n7102) );
  INV_X1 U8394 ( .A(n10592), .ZN(n7100) );
  OAI22_X1 U8395 ( .A1(n7253), .A2(n9005), .B1(n7100), .B2(n9003), .ZN(n7101)
         );
  AOI21_X1 U8396 ( .B1(n7102), .B2(n10629), .A(n7101), .ZN(n10611) );
  INV_X1 U8397 ( .A(n10611), .ZN(n7106) );
  NOR2_X1 U8398 ( .A1(n10709), .A2(n5796), .ZN(n7105) );
  OAI22_X1 U8399 ( .A1(n10653), .A2(n10612), .B1(n7103), .B2(n10650), .ZN(
        n7104) );
  AOI211_X1 U8400 ( .C1(n7106), .C2(n10709), .A(n7105), .B(n7104), .ZN(n7107)
         );
  OAI21_X1 U8401 ( .B1(n7108), .B2(n8968), .A(n7107), .ZN(P2_U3229) );
  XNOR2_X1 U8402 ( .A(n7109), .B(n8329), .ZN(n10608) );
  OAI22_X1 U8403 ( .A1(n10653), .A2(n10605), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10650), .ZN(n7116) );
  INV_X1 U8404 ( .A(n8329), .ZN(n7110) );
  XNOR2_X1 U8405 ( .A(n7111), .B(n7110), .ZN(n7112) );
  NAND2_X1 U8406 ( .A1(n7112), .A2(n10641), .ZN(n7114) );
  AOI22_X1 U8407 ( .A1(n10637), .A2(n8708), .B1(n10636), .B2(n6190), .ZN(n7113) );
  NAND2_X1 U8408 ( .A1(n7114), .A2(n7113), .ZN(n10606) );
  MUX2_X1 U8409 ( .A(n10606), .B(P2_REG2_REG_3__SCAN_IN), .S(n9017), .Z(n7115)
         );
  AOI211_X1 U8410 ( .C1(n9015), .C2(n10608), .A(n7116), .B(n7115), .ZN(n7117)
         );
  INV_X1 U8411 ( .A(n7117), .ZN(P2_U3230) );
  NAND2_X1 U8412 ( .A1(n7119), .A2(n7118), .ZN(n7120) );
  NAND2_X1 U8413 ( .A1(n7121), .A2(n7120), .ZN(n7268) );
  NAND2_X1 U8414 ( .A1(n9561), .A2(n7271), .ZN(n8087) );
  NAND2_X1 U8415 ( .A1(n8096), .A2(n8087), .ZN(n7266) );
  NAND2_X1 U8416 ( .A1(n7268), .A2(n7266), .ZN(n7317) );
  OAI21_X1 U8417 ( .B1(n7268), .B2(n7266), .A(n7317), .ZN(n7122) );
  INV_X1 U8418 ( .A(n7122), .ZN(n10622) );
  NAND2_X1 U8419 ( .A1(n7123), .A2(n8088), .ZN(n7264) );
  INV_X1 U8420 ( .A(n7266), .ZN(n8027) );
  XNOR2_X1 U8421 ( .A(n7264), .B(n8027), .ZN(n7124) );
  AOI222_X1 U8422 ( .A1(n10752), .A2(n7124), .B1(n9560), .B2(n10756), .C1(
        n9562), .C2(n10759), .ZN(n10621) );
  MUX2_X1 U8423 ( .A(n6504), .B(n10621), .S(n10560), .Z(n7130) );
  AOI211_X1 U8424 ( .C1(n10618), .C2(n7125), .A(n9915), .B(n7327), .ZN(n10617)
         );
  OAI22_X1 U8425 ( .A1(n9976), .A2(n7271), .B1(n7127), .B2(n7126), .ZN(n7128)
         );
  AOI21_X1 U8426 ( .B1(n10617), .B2(n9972), .A(n7128), .ZN(n7129) );
  OAI211_X1 U8427 ( .C1(n9979), .C2(n10622), .A(n7130), .B(n7129), .ZN(
        P1_U3289) );
  OAI21_X1 U8428 ( .B1(n7131), .B2(n6138), .A(n10588), .ZN(n7132) );
  NAND2_X1 U8429 ( .A1(n7132), .A2(n10641), .ZN(n7134) );
  AOI22_X1 U8430 ( .A1(n10637), .A2(n8709), .B1(n8708), .B2(n6190), .ZN(n7133)
         );
  NAND2_X1 U8431 ( .A1(n7134), .A2(n7133), .ZN(n10572) );
  INV_X1 U8432 ( .A(n10572), .ZN(n7142) );
  OAI21_X1 U8433 ( .B1(n7137), .B2(n7136), .A(n7135), .ZN(n10574) );
  INV_X1 U8434 ( .A(n10653), .ZN(n10704) );
  AOI22_X1 U8435 ( .A1(n10704), .A2(n7138), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10706), .ZN(n7139) );
  OAI21_X1 U8436 ( .B1(n5751), .B2(n10709), .A(n7139), .ZN(n7140) );
  AOI21_X1 U8437 ( .B1(n10574), .B2(n9015), .A(n7140), .ZN(n7141) );
  OAI21_X1 U8438 ( .B1(n7142), .B2(n9017), .A(n7141), .ZN(P2_U3232) );
  INV_X1 U8439 ( .A(n7143), .ZN(n7144) );
  NOR2_X1 U8440 ( .A1(n7144), .A2(n8380), .ZN(n10633) );
  NAND2_X1 U8441 ( .A1(n7145), .A2(n8384), .ZN(n10632) );
  NOR2_X1 U8442 ( .A1(n10633), .A2(n10632), .ZN(n10631) );
  INV_X1 U8443 ( .A(n7145), .ZN(n8381) );
  NOR2_X1 U8444 ( .A1(n10631), .A2(n8381), .ZN(n7146) );
  XNOR2_X1 U8445 ( .A(n7146), .B(n8331), .ZN(n10669) );
  INV_X1 U8446 ( .A(n7251), .ZN(n7147) );
  AOI22_X1 U8447 ( .A1(n10704), .A2(n7260), .B1(n10706), .B2(n7147), .ZN(n7153) );
  XNOR2_X1 U8448 ( .A(n7469), .B(n8331), .ZN(n7150) );
  NAND2_X1 U8449 ( .A1(n8707), .A2(n10637), .ZN(n7148) );
  OAI21_X1 U8450 ( .B1(n7290), .B2(n9005), .A(n7148), .ZN(n7149) );
  AOI21_X1 U8451 ( .B1(n7150), .B2(n10641), .A(n7149), .ZN(n10670) );
  MUX2_X1 U8452 ( .A(n7151), .B(n10670), .S(n10709), .Z(n7152) );
  OAI211_X1 U8453 ( .C1(n10669), .C2(n8968), .A(n7153), .B(n7152), .ZN(
        P2_U3227) );
  AOI21_X1 U8454 ( .B1(n7156), .B2(n7155), .A(n7154), .ZN(n7172) );
  AOI21_X1 U8455 ( .B1(n7159), .B2(n7158), .A(n7157), .ZN(n7160) );
  NOR2_X1 U8456 ( .A1(n7160), .A2(n10496), .ZN(n7170) );
  AOI21_X1 U8457 ( .B1(n7163), .B2(n7162), .A(n7161), .ZN(n7168) );
  NOR2_X1 U8458 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7164), .ZN(n7459) );
  AOI21_X1 U8459 ( .B1(n10516), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7459), .ZN(
        n7167) );
  NAND2_X1 U8460 ( .A1(n10434), .A2(n7165), .ZN(n7166) );
  OAI211_X1 U8461 ( .C1(n7168), .C2(n10464), .A(n7167), .B(n7166), .ZN(n7169)
         );
  NOR2_X1 U8462 ( .A1(n7170), .A2(n7169), .ZN(n7171) );
  OAI21_X1 U8463 ( .B1(n7172), .B2(n10514), .A(n7171), .ZN(P2_U3190) );
  INV_X1 U8464 ( .A(n7990), .ZN(n7175) );
  OAI222_X1 U8465 ( .A1(n10132), .A2(n7173), .B1(n10138), .B2(n7175), .C1(
        n9674), .C2(P1_U3086), .ZN(P1_U3336) );
  OAI222_X1 U8466 ( .A1(n7176), .A2(P2_U3151), .B1(n9162), .B2(n7175), .C1(
        n7174), .C2(n9153), .ZN(P2_U3276) );
  AOI21_X1 U8467 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7708), .A(n7177), .ZN(
        n7180) );
  NAND2_X1 U8468 ( .A1(n7781), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7178) );
  OAI21_X1 U8469 ( .B1(n7781), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7178), .ZN(
        n7179) );
  NOR2_X1 U8470 ( .A1(n7180), .A2(n7179), .ZN(n7640) );
  AOI211_X1 U8471 ( .C1(n7180), .C2(n7179), .A(n7640), .B(n9623), .ZN(n7188)
         );
  AOI21_X1 U8472 ( .B1(n7708), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7181), .ZN(
        n7183) );
  XNOR2_X1 U8473 ( .A(n7781), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7182) );
  NOR2_X1 U8474 ( .A1(n7183), .A2(n7182), .ZN(n7636) );
  AOI211_X1 U8475 ( .C1(n7183), .C2(n7182), .A(n7636), .B(n10546), .ZN(n7187)
         );
  INV_X1 U8476 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7185) );
  NAND2_X1 U8477 ( .A1(n10542), .A2(n7781), .ZN(n7184) );
  NAND2_X1 U8478 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9335) );
  OAI211_X1 U8479 ( .C1(n7185), .C2(n9669), .A(n7184), .B(n9335), .ZN(n7186)
         );
  OR3_X1 U8480 ( .A1(n7188), .A2(n7187), .A3(n7186), .ZN(P1_U3257) );
  INV_X1 U8481 ( .A(n7189), .ZN(n7190) );
  NAND2_X1 U8482 ( .A1(n7191), .A2(n7190), .ZN(n7192) );
  NAND2_X1 U8483 ( .A1(n9560), .A2(n9309), .ZN(n7200) );
  OR2_X1 U8484 ( .A1(n7394), .A2(n7194), .ZN(n7197) );
  OR2_X1 U8485 ( .A1(n6943), .A2(n7195), .ZN(n7196) );
  OAI211_X1 U8486 ( .C1(n7392), .C2(n7198), .A(n7197), .B(n7196), .ZN(n7269)
         );
  NAND2_X1 U8487 ( .A1(n7269), .A2(n6725), .ZN(n7199) );
  NAND2_X1 U8488 ( .A1(n7200), .A2(n7199), .ZN(n7201) );
  XNOR2_X1 U8489 ( .A(n7201), .B(n9314), .ZN(n7202) );
  NAND2_X1 U8490 ( .A1(n7221), .A2(n7220), .ZN(n7204) );
  AND2_X1 U8491 ( .A1(n7269), .A2(n4948), .ZN(n7203) );
  AOI21_X1 U8492 ( .B1(n9560), .B2(n9307), .A(n7203), .ZN(n7219) );
  XNOR2_X1 U8493 ( .A(n7204), .B(n7219), .ZN(n7218) );
  INV_X1 U8494 ( .A(n7205), .ZN(n7215) );
  NAND2_X1 U8495 ( .A1(n7898), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7213) );
  NAND2_X1 U8496 ( .A1(n8072), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7212) );
  INV_X1 U8497 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7207) );
  NOR2_X1 U8498 ( .A1(n7208), .A2(n7207), .ZN(n7233) );
  INV_X1 U8499 ( .A(n7233), .ZN(n7235) );
  NAND2_X1 U8500 ( .A1(n7208), .A2(n7207), .ZN(n7209) );
  AND2_X1 U8501 ( .A1(n7235), .A2(n7209), .ZN(n7281) );
  NAND2_X1 U8502 ( .A1(n7948), .A2(n7281), .ZN(n7211) );
  NAND2_X1 U8503 ( .A1(n8071), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7210) );
  NAND4_X1 U8504 ( .A1(n7213), .A2(n7212), .A3(n7211), .A4(n7210), .ZN(n9559)
         );
  INV_X1 U8505 ( .A(n9559), .ZN(n7343) );
  OAI22_X1 U8506 ( .A1(n9498), .A2(n7272), .B1(n7343), .B2(n9542), .ZN(n7214)
         );
  AOI211_X1 U8507 ( .C1(n7269), .C2(n9473), .A(n7215), .B(n7214), .ZN(n7217)
         );
  NAND2_X1 U8508 ( .A1(n9546), .A2(n10660), .ZN(n7216) );
  OAI211_X1 U8509 ( .C1(n7218), .C2(n9548), .A(n7217), .B(n7216), .ZN(P1_U3227) );
  NAND2_X1 U8510 ( .A1(n9559), .A2(n4948), .ZN(n7228) );
  OR2_X1 U8511 ( .A1(n7394), .A2(n7222), .ZN(n7225) );
  OR2_X1 U8512 ( .A1(n6943), .A2(n7223), .ZN(n7224) );
  OAI211_X1 U8513 ( .C1(n7392), .C2(n7226), .A(n7225), .B(n7224), .ZN(n7262)
         );
  NAND2_X1 U8514 ( .A1(n7262), .A2(n6725), .ZN(n7227) );
  NAND2_X1 U8515 ( .A1(n7228), .A2(n7227), .ZN(n7229) );
  XNOR2_X1 U8516 ( .A(n7229), .B(n9373), .ZN(n7424) );
  AND2_X1 U8517 ( .A1(n7262), .A2(n4948), .ZN(n7230) );
  AOI21_X1 U8518 ( .B1(n9559), .B2(n9307), .A(n7230), .ZN(n7425) );
  XNOR2_X1 U8519 ( .A(n7424), .B(n7425), .ZN(n7231) );
  XNOR2_X1 U8520 ( .A(n7423), .B(n7231), .ZN(n7245) );
  INV_X1 U8521 ( .A(n7232), .ZN(n7242) );
  NAND2_X1 U8522 ( .A1(n8072), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7240) );
  NAND2_X1 U8523 ( .A1(n7898), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7239) );
  NAND2_X1 U8524 ( .A1(n7233), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7353) );
  INV_X1 U8525 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7234) );
  NAND2_X1 U8526 ( .A1(n7235), .A2(n7234), .ZN(n7236) );
  AND2_X1 U8527 ( .A1(n7353), .A2(n7236), .ZN(n7444) );
  NAND2_X1 U8528 ( .A1(n7948), .A2(n7444), .ZN(n7238) );
  NAND2_X1 U8529 ( .A1(n8071), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7237) );
  NAND4_X1 U8530 ( .A1(n7240), .A2(n7239), .A3(n7238), .A4(n7237), .ZN(n9558)
         );
  INV_X1 U8531 ( .A(n9558), .ZN(n7390) );
  OAI22_X1 U8532 ( .A1(n9498), .A2(n7270), .B1(n7390), .B2(n9542), .ZN(n7241)
         );
  AOI211_X1 U8533 ( .C1(n7262), .C2(n9473), .A(n7242), .B(n7241), .ZN(n7244)
         );
  NAND2_X1 U8534 ( .A1(n9546), .A2(n7281), .ZN(n7243) );
  OAI211_X1 U8535 ( .C1(n7245), .C2(n9548), .A(n7244), .B(n7243), .ZN(P1_U3239) );
  INV_X1 U8536 ( .A(n7981), .ZN(n7315) );
  NAND2_X1 U8537 ( .A1(n10126), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7246) );
  OAI211_X1 U8538 ( .C1(n7315), .C2(n10138), .A(n7247), .B(n7246), .ZN(
        P1_U3335) );
  NAND2_X1 U8539 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10528) );
  INV_X1 U8540 ( .A(n10528), .ZN(n7248) );
  AOI21_X1 U8541 ( .B1(n8663), .B2(n8707), .A(n7248), .ZN(n7250) );
  OR2_X1 U8542 ( .A1(n7290), .A2(n8660), .ZN(n7249) );
  OAI211_X1 U8543 ( .C1(n8683), .C2(n7251), .A(n7250), .B(n7249), .ZN(n7259)
         );
  XNOR2_X1 U8544 ( .A(n7260), .B(n7870), .ZN(n7287) );
  XNOR2_X1 U8545 ( .A(n7287), .B(n10635), .ZN(n7257) );
  NAND2_X1 U8546 ( .A1(n7253), .A2(n7252), .ZN(n7254) );
  AOI211_X1 U8547 ( .C1(n7257), .C2(n7256), .A(n8676), .B(n7288), .ZN(n7258)
         );
  AOI211_X1 U8548 ( .C1(n7260), .C2(n8673), .A(n7259), .B(n7258), .ZN(n7261)
         );
  INV_X1 U8549 ( .A(n7261), .ZN(P2_U3179) );
  NAND2_X1 U8550 ( .A1(n7343), .A2(n7262), .ZN(n8238) );
  INV_X1 U8551 ( .A(n7262), .ZN(n10676) );
  NAND2_X1 U8552 ( .A1(n9559), .A2(n10676), .ZN(n8104) );
  NAND2_X1 U8553 ( .A1(n8238), .A2(n8104), .ZN(n8099) );
  NAND2_X1 U8554 ( .A1(n7270), .A2(n7269), .ZN(n8239) );
  INV_X1 U8555 ( .A(n8096), .ZN(n7263) );
  INV_X1 U8556 ( .A(n7269), .ZN(n10662) );
  NAND2_X1 U8557 ( .A1(n9560), .A2(n10662), .ZN(n8242) );
  INV_X1 U8558 ( .A(n8242), .ZN(n8098) );
  XOR2_X1 U8559 ( .A(n8099), .B(n5029), .Z(n7280) );
  AOI22_X1 U8560 ( .A1(n10759), .A2(n9560), .B1(n9558), .B2(n10756), .ZN(n7279) );
  NAND2_X1 U8561 ( .A1(n8239), .A2(n8242), .ZN(n8102) );
  AND2_X1 U8562 ( .A1(n7266), .A2(n8102), .ZN(n7267) );
  NAND2_X1 U8563 ( .A1(n7268), .A2(n7267), .ZN(n7318) );
  AND2_X1 U8564 ( .A1(n8239), .A2(n7269), .ZN(n7275) );
  NAND2_X1 U8565 ( .A1(n7270), .A2(n10662), .ZN(n7273) );
  NAND2_X1 U8566 ( .A1(n7272), .A2(n7271), .ZN(n7319) );
  AND2_X1 U8567 ( .A1(n7273), .A2(n7319), .ZN(n7274) );
  OR2_X1 U8568 ( .A1(n7275), .A2(n7274), .ZN(n7276) );
  NAND2_X1 U8569 ( .A1(n7318), .A2(n7276), .ZN(n7277) );
  NAND2_X1 U8570 ( .A1(n7277), .A2(n8099), .ZN(n7345) );
  OAI21_X1 U8571 ( .B1(n7277), .B2(n8099), .A(n7345), .ZN(n10679) );
  NAND2_X1 U8572 ( .A1(n10679), .A2(n7400), .ZN(n7278) );
  OAI211_X1 U8573 ( .C1(n7280), .C2(n10563), .A(n7279), .B(n7278), .ZN(n10677)
         );
  INV_X1 U8574 ( .A(n10677), .ZN(n7286) );
  NAND2_X1 U8575 ( .A1(n7325), .A2(n10676), .ZN(n7367) );
  OAI211_X1 U8576 ( .C1(n7325), .C2(n10676), .A(n10762), .B(n7367), .ZN(n10675) );
  NOR2_X1 U8577 ( .A1(n10675), .A2(n10658), .ZN(n7284) );
  AOI22_X1 U8578 ( .A1(n10786), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7281), .B2(
        n10775), .ZN(n7282) );
  OAI21_X1 U8579 ( .B1(n10676), .B2(n9976), .A(n7282), .ZN(n7283) );
  AOI211_X1 U8580 ( .C1(n10679), .C2(n7421), .A(n7284), .B(n7283), .ZN(n7285)
         );
  OAI21_X1 U8581 ( .B1(n7286), .B2(n10786), .A(n7285), .ZN(P1_U3287) );
  XNOR2_X1 U8582 ( .A(n10687), .B(n7874), .ZN(n7289) );
  NAND2_X1 U8583 ( .A1(n7290), .A2(n7289), .ZN(n7453) );
  INV_X1 U8584 ( .A(n7289), .ZN(n7291) );
  INV_X1 U8585 ( .A(n7290), .ZN(n8706) );
  NAND2_X1 U8586 ( .A1(n7291), .A2(n8706), .ZN(n7292) );
  AND2_X1 U8587 ( .A1(n7453), .A2(n7292), .ZN(n7293) );
  OAI21_X1 U8588 ( .B1(n7294), .B2(n7293), .A(n7454), .ZN(n7295) );
  NAND2_X1 U8589 ( .A1(n7295), .A2(n8624), .ZN(n7301) );
  AOI21_X1 U8590 ( .B1(n8663), .B2(n10635), .A(n7296), .ZN(n7298) );
  NAND2_X1 U8591 ( .A1(n8705), .A2(n8686), .ZN(n7297) );
  OAI211_X1 U8592 ( .C1(n8683), .C2(n7308), .A(n7298), .B(n7297), .ZN(n7299)
         );
  INV_X1 U8593 ( .A(n7299), .ZN(n7300) );
  OAI211_X1 U8594 ( .C1(n7302), .C2(n8689), .A(n7301), .B(n7300), .ZN(P2_U3153) );
  INV_X1 U8595 ( .A(n7469), .ZN(n7303) );
  OAI21_X1 U8596 ( .B1(n7303), .B2(n7307), .A(n10668), .ZN(n7304) );
  OAI21_X1 U8597 ( .B1(n7469), .B2(n10635), .A(n7304), .ZN(n7305) );
  XNOR2_X1 U8598 ( .A(n7305), .B(n8403), .ZN(n7306) );
  OAI222_X1 U8599 ( .A1(n9005), .A2(n5437), .B1(n9003), .B2(n7307), .C1(n9000), 
        .C2(n7306), .ZN(n10685) );
  INV_X1 U8600 ( .A(n10685), .ZN(n7313) );
  OAI22_X1 U8601 ( .A1(n10709), .A2(n6313), .B1(n7308), .B2(n10650), .ZN(n7311) );
  NOR2_X1 U8602 ( .A1(n7309), .A2(n8403), .ZN(n10684) );
  INV_X1 U8603 ( .A(n7466), .ZN(n10683) );
  NOR3_X1 U8604 ( .A1(n10684), .A2(n10683), .A3(n8968), .ZN(n7310) );
  AOI211_X1 U8605 ( .C1(n10704), .C2(n10687), .A(n7311), .B(n7310), .ZN(n7312)
         );
  OAI21_X1 U8606 ( .B1(n7313), .B2(n9017), .A(n7312), .ZN(P2_U3226) );
  OAI222_X1 U8607 ( .A1(P2_U3151), .A2(n8512), .B1(n9162), .B2(n7315), .C1(
        n7314), .C2(n9153), .ZN(P2_U3275) );
  NAND2_X1 U8608 ( .A1(n7317), .A2(n7319), .ZN(n7322) );
  INV_X1 U8609 ( .A(n8102), .ZN(n8028) );
  OR2_X1 U8610 ( .A1(n8028), .A2(n7319), .ZN(n7320) );
  AND2_X1 U8611 ( .A1(n7318), .A2(n7320), .ZN(n7321) );
  OAI21_X1 U8612 ( .B1(n7322), .B2(n8102), .A(n7321), .ZN(n10665) );
  INV_X1 U8613 ( .A(n10665), .ZN(n7328) );
  XNOR2_X1 U8614 ( .A(n8102), .B(n7323), .ZN(n7324) );
  AOI222_X1 U8615 ( .A1(n10752), .A2(n7324), .B1(n9559), .B2(n10756), .C1(
        n9561), .C2(n10759), .ZN(n10667) );
  INV_X1 U8616 ( .A(n7325), .ZN(n7326) );
  OAI211_X1 U8617 ( .C1(n10662), .C2(n7327), .A(n7326), .B(n10762), .ZN(n10659) );
  OAI211_X1 U8618 ( .C1(n10623), .C2(n7328), .A(n10667), .B(n10659), .ZN(n7334) );
  INV_X1 U8619 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7329) );
  OAI22_X1 U8620 ( .A1(n10069), .A2(n10662), .B1(n10770), .B2(n7329), .ZN(
        n7330) );
  AOI21_X1 U8621 ( .B1(n7334), .B2(n10770), .A(n7330), .ZN(n7331) );
  INV_X1 U8622 ( .A(n7331), .ZN(P1_U3527) );
  INV_X1 U8623 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7332) );
  OAI22_X1 U8624 ( .A1(n10122), .A2(n10662), .B1(n10774), .B2(n7332), .ZN(
        n7333) );
  AOI21_X1 U8625 ( .B1(n7334), .B2(n10774), .A(n7333), .ZN(n7335) );
  INV_X1 U8626 ( .A(n7335), .ZN(P1_U3468) );
  XOR2_X1 U8627 ( .A(n8334), .B(n7336), .Z(n7337) );
  OAI222_X1 U8628 ( .A1(n9005), .A2(n8641), .B1(n9003), .B2(n5437), .C1(n9000), 
        .C2(n7337), .ZN(n10722) );
  INV_X1 U8629 ( .A(n10722), .ZN(n7342) );
  OAI22_X1 U8630 ( .A1(n10709), .A2(n5879), .B1(n7650), .B2(n10650), .ZN(n7338) );
  AOI21_X1 U8631 ( .B1(n10704), .B2(n10724), .A(n7338), .ZN(n7341) );
  NAND2_X1 U8632 ( .A1(n7339), .A2(n8334), .ZN(n10719) );
  NAND3_X1 U8633 ( .A1(n10721), .A2(n10719), .A3(n9015), .ZN(n7340) );
  OAI211_X1 U8634 ( .C1(n7342), .C2(n9017), .A(n7341), .B(n7340), .ZN(P2_U3224) );
  NAND2_X1 U8635 ( .A1(n7343), .A2(n10676), .ZN(n7344) );
  OR2_X1 U8636 ( .A1(n7394), .A2(n7346), .ZN(n7349) );
  OR2_X1 U8637 ( .A1(n6943), .A2(n7347), .ZN(n7348) );
  OAI211_X1 U8638 ( .C1(n7392), .C2(n7350), .A(n7349), .B(n7348), .ZN(n7601)
         );
  NAND2_X1 U8639 ( .A1(n7390), .A2(n7601), .ZN(n8112) );
  NAND2_X1 U8640 ( .A1(n9558), .A2(n7605), .ZN(n8113) );
  NAND2_X1 U8641 ( .A1(n8112), .A2(n8113), .ZN(n7361) );
  OAI21_X1 U8642 ( .B1(n7351), .B2(n7361), .A(n7391), .ZN(n7600) );
  INV_X1 U8643 ( .A(n7600), .ZN(n7372) );
  NAND2_X1 U8644 ( .A1(n8070), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7358) );
  NAND2_X1 U8645 ( .A1(n8072), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7357) );
  NAND2_X1 U8646 ( .A1(n7353), .A2(n7352), .ZN(n7354) );
  AND2_X1 U8647 ( .A1(n7404), .A2(n7354), .ZN(n9395) );
  NAND2_X1 U8648 ( .A1(n7948), .A2(n9395), .ZN(n7356) );
  NAND2_X1 U8649 ( .A1(n8071), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7355) );
  NAND4_X1 U8650 ( .A1(n7358), .A2(n7357), .A3(n7356), .A4(n7355), .ZN(n9557)
         );
  AOI22_X1 U8651 ( .A1(n10759), .A2(n9559), .B1(n9557), .B2(n10756), .ZN(n7365) );
  INV_X1 U8652 ( .A(n8104), .ZN(n7359) );
  NOR2_X1 U8653 ( .A1(n7361), .A2(n7359), .ZN(n7360) );
  NAND2_X1 U8654 ( .A1(n7519), .A2(n7360), .ZN(n7488) );
  INV_X1 U8655 ( .A(n7488), .ZN(n7363) );
  AOI21_X1 U8656 ( .B1(n7519), .B2(n8104), .A(n5497), .ZN(n7362) );
  OAI21_X1 U8657 ( .B1(n7363), .B2(n7362), .A(n10752), .ZN(n7364) );
  OAI211_X1 U8658 ( .C1(n7372), .C2(n7629), .A(n7365), .B(n7364), .ZN(n7598)
         );
  NAND2_X1 U8659 ( .A1(n7598), .A2(n10560), .ZN(n7371) );
  INV_X1 U8660 ( .A(n7416), .ZN(n7366) );
  AOI211_X1 U8661 ( .C1(n7601), .C2(n7367), .A(n9915), .B(n7366), .ZN(n7599)
         );
  AOI22_X1 U8662 ( .A1(n10786), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7444), .B2(
        n10775), .ZN(n7368) );
  OAI21_X1 U8663 ( .B1(n7605), .B2(n9976), .A(n7368), .ZN(n7369) );
  AOI21_X1 U8664 ( .B1(n7599), .B2(n9972), .A(n7369), .ZN(n7370) );
  OAI211_X1 U8665 ( .C1(n7372), .C2(n7635), .A(n7371), .B(n7370), .ZN(P1_U3286) );
  AOI21_X1 U8666 ( .B1(n10725), .B2(n7374), .A(n7373), .ZN(n7388) );
  AOI21_X1 U8667 ( .B1(n5879), .B2(n7376), .A(n7375), .ZN(n7377) );
  NOR2_X1 U8668 ( .A1(n7377), .A2(n10496), .ZN(n7386) );
  AOI21_X1 U8669 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n7384) );
  AND2_X1 U8670 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7647) );
  AOI21_X1 U8671 ( .B1(n10516), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7647), .ZN(
        n7383) );
  NAND2_X1 U8672 ( .A1(n10434), .A2(n7381), .ZN(n7382) );
  OAI211_X1 U8673 ( .C1(n7384), .C2(n10464), .A(n7383), .B(n7382), .ZN(n7385)
         );
  NOR2_X1 U8674 ( .A1(n7386), .A2(n7385), .ZN(n7387) );
  OAI21_X1 U8675 ( .B1(n7388), .B2(n10514), .A(n7387), .ZN(P2_U3191) );
  INV_X1 U8676 ( .A(n7972), .ZN(n7481) );
  INV_X1 U8677 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7389) );
  OAI222_X1 U8678 ( .A1(P2_U3151), .A2(n8362), .B1(n9162), .B2(n7481), .C1(
        n7389), .C2(n9153), .ZN(P2_U3274) );
  INV_X1 U8679 ( .A(n9557), .ZN(n9463) );
  AOI22_X1 U8680 ( .A1(n8046), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8045), .B2(
        n7393), .ZN(n7397) );
  NAND2_X1 U8681 ( .A1(n7395), .A2(n8043), .ZN(n7396) );
  NAND2_X1 U8682 ( .A1(n7397), .A2(n7396), .ZN(n9179) );
  NAND2_X1 U8683 ( .A1(n9463), .A2(n9179), .ZN(n8106) );
  INV_X1 U8684 ( .A(n9179), .ZN(n10691) );
  NAND2_X1 U8685 ( .A1(n9557), .A2(n10691), .ZN(n7517) );
  NAND2_X1 U8686 ( .A1(n8106), .A2(n7517), .ZN(n7401) );
  OR2_X1 U8687 ( .A1(n7398), .A2(n7401), .ZN(n7399) );
  NAND2_X1 U8688 ( .A1(n7504), .A2(n7399), .ZN(n10694) );
  NAND2_X1 U8689 ( .A1(n10694), .A2(n7400), .ZN(n7415) );
  NAND2_X1 U8690 ( .A1(n7488), .A2(n8112), .ZN(n7402) );
  INV_X1 U8691 ( .A(n7401), .ZN(n8118) );
  XNOR2_X1 U8692 ( .A(n7402), .B(n8118), .ZN(n7413) );
  NAND2_X1 U8693 ( .A1(n9558), .A2(n10759), .ZN(n7411) );
  NAND2_X1 U8694 ( .A1(n8070), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U8695 ( .A1(n8071), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7408) );
  NOR2_X1 U8696 ( .A1(n7404), .A2(n7403), .ZN(n7491) );
  INV_X1 U8697 ( .A(n7491), .ZN(n7493) );
  NAND2_X1 U8698 ( .A1(n7404), .A2(n7403), .ZN(n7405) );
  AND2_X1 U8699 ( .A1(n7493), .A2(n7405), .ZN(n9459) );
  NAND2_X1 U8700 ( .A1(n7948), .A2(n9459), .ZN(n7407) );
  NAND2_X1 U8701 ( .A1(n8072), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7406) );
  NAND4_X1 U8702 ( .A1(n7409), .A2(n7408), .A3(n7407), .A4(n7406), .ZN(n9556)
         );
  NAND2_X1 U8703 ( .A1(n9556), .A2(n10756), .ZN(n7410) );
  NAND2_X1 U8704 ( .A1(n7411), .A2(n7410), .ZN(n7412) );
  AOI21_X1 U8705 ( .B1(n7413), .B2(n10752), .A(n7412), .ZN(n7414) );
  AOI21_X1 U8706 ( .B1(n7416), .B2(n9179), .A(n9915), .ZN(n7417) );
  NAND2_X1 U8707 ( .A1(n7417), .A2(n7537), .ZN(n10690) );
  NOR2_X1 U8708 ( .A1(n10690), .A2(n10658), .ZN(n7420) );
  AOI22_X1 U8709 ( .A1(n10786), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9395), .B2(
        n10775), .ZN(n7418) );
  OAI21_X1 U8710 ( .B1(n10691), .B2(n9976), .A(n7418), .ZN(n7419) );
  AOI211_X1 U8711 ( .C1(n10694), .C2(n7421), .A(n7420), .B(n7419), .ZN(n7422)
         );
  OAI21_X1 U8712 ( .B1(n10696), .B2(n10786), .A(n7422), .ZN(P1_U3285) );
  INV_X1 U8713 ( .A(n7424), .ZN(n7427) );
  INV_X1 U8714 ( .A(n7425), .ZN(n7426) );
  NAND2_X1 U8715 ( .A1(n7427), .A2(n7426), .ZN(n7428) );
  NAND2_X1 U8716 ( .A1(n7429), .A2(n7428), .ZN(n9167) );
  NAND2_X1 U8717 ( .A1(n9558), .A2(n9309), .ZN(n7431) );
  NAND2_X1 U8718 ( .A1(n7601), .A2(n6725), .ZN(n7430) );
  NAND2_X1 U8719 ( .A1(n7431), .A2(n7430), .ZN(n7432) );
  XNOR2_X1 U8720 ( .A(n7432), .B(n9314), .ZN(n7435) );
  NAND2_X1 U8721 ( .A1(n9558), .A2(n9307), .ZN(n7434) );
  NAND2_X1 U8722 ( .A1(n7601), .A2(n9309), .ZN(n7433) );
  NAND2_X1 U8723 ( .A1(n7434), .A2(n7433), .ZN(n7436) );
  AND2_X1 U8724 ( .A1(n7435), .A2(n7436), .ZN(n9165) );
  INV_X1 U8725 ( .A(n9165), .ZN(n7439) );
  INV_X1 U8726 ( .A(n7435), .ZN(n7438) );
  INV_X1 U8727 ( .A(n7436), .ZN(n7437) );
  NAND2_X1 U8728 ( .A1(n7438), .A2(n7437), .ZN(n9166) );
  NAND2_X1 U8729 ( .A1(n7439), .A2(n9166), .ZN(n7440) );
  XNOR2_X1 U8730 ( .A(n9167), .B(n7440), .ZN(n7441) );
  NAND2_X1 U8731 ( .A1(n7441), .A2(n9529), .ZN(n7450) );
  NAND2_X1 U8732 ( .A1(n9539), .A2(n9559), .ZN(n7442) );
  OAI211_X1 U8733 ( .C1(n9463), .C2(n9542), .A(n7443), .B(n7442), .ZN(n7448)
         );
  INV_X1 U8734 ( .A(n7444), .ZN(n7445) );
  NOR2_X1 U8735 ( .A1(n7446), .A2(n7445), .ZN(n7447) );
  NOR2_X1 U8736 ( .A1(n7448), .A2(n7447), .ZN(n7449) );
  OAI211_X1 U8737 ( .C1(n7605), .C2(n9543), .A(n7450), .B(n7449), .ZN(P1_U3213) );
  INV_X1 U8738 ( .A(n7454), .ZN(n7452) );
  INV_X1 U8739 ( .A(n7453), .ZN(n7451) );
  XNOR2_X1 U8740 ( .A(n10705), .B(n7874), .ZN(n7651) );
  XNOR2_X1 U8741 ( .A(n7651), .B(n8705), .ZN(n7455) );
  NOR3_X1 U8742 ( .A1(n7452), .A2(n7451), .A3(n7455), .ZN(n7458) );
  NAND2_X1 U8743 ( .A1(n7454), .A2(n7453), .ZN(n7456) );
  NAND2_X1 U8744 ( .A1(n7456), .A2(n7455), .ZN(n7653) );
  INV_X1 U8745 ( .A(n7653), .ZN(n7457) );
  OAI21_X1 U8746 ( .B1(n7458), .B2(n7457), .A(n8624), .ZN(n7464) );
  AOI21_X1 U8747 ( .B1(n8706), .B2(n8663), .A(n7459), .ZN(n7460) );
  OAI21_X1 U8748 ( .B1(n7461), .B2(n8660), .A(n7460), .ZN(n7462) );
  AOI21_X1 U8749 ( .B1(n10707), .B2(n8615), .A(n7462), .ZN(n7463) );
  OAI211_X1 U8750 ( .C1(n7477), .C2(n8689), .A(n7464), .B(n7463), .ZN(P2_U3161) );
  NAND2_X1 U8751 ( .A1(n7466), .A2(n7465), .ZN(n7467) );
  XOR2_X1 U8752 ( .A(n8333), .B(n7467), .Z(n10702) );
  OR2_X1 U8753 ( .A1(n7469), .A2(n7468), .ZN(n7471) );
  NAND2_X1 U8754 ( .A1(n7471), .A2(n7470), .ZN(n7472) );
  XNOR2_X1 U8755 ( .A(n7472), .B(n8333), .ZN(n7473) );
  AOI222_X1 U8756 ( .A1(n10641), .A2(n7473), .B1(n8704), .B2(n6190), .C1(n8706), .C2(n10637), .ZN(n10701) );
  OAI21_X1 U8757 ( .B1(n10801), .B2(n10702), .A(n10701), .ZN(n7479) );
  INV_X1 U8758 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7474) );
  OAI22_X1 U8759 ( .A1(n9143), .A2(n7477), .B1(n10810), .B2(n7474), .ZN(n7475)
         );
  AOI21_X1 U8760 ( .B1(n7479), .B2(n10810), .A(n7475), .ZN(n7476) );
  INV_X1 U8761 ( .A(n7476), .ZN(P2_U3414) );
  OAI22_X1 U8762 ( .A1(n9089), .A2(n7477), .B1(n10806), .B2(n6310), .ZN(n7478)
         );
  AOI21_X1 U8763 ( .B1(n7479), .B2(n10806), .A(n7478), .ZN(n7480) );
  INV_X1 U8764 ( .A(n7480), .ZN(P2_U3467) );
  INV_X1 U8765 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7482) );
  OAI222_X1 U8766 ( .A1(n10132), .A2(n7482), .B1(P1_U3086), .B2(n8231), .C1(
        n10138), .C2(n7481), .ZN(P1_U3334) );
  INV_X1 U8767 ( .A(n9556), .ZN(n7487) );
  NAND2_X1 U8768 ( .A1(n7483), .A2(n8043), .ZN(n7486) );
  AOI22_X1 U8769 ( .A1(n8046), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8045), .B2(
        n7484), .ZN(n7485) );
  NAND2_X1 U8770 ( .A1(n7486), .A2(n7485), .ZN(n9465) );
  NAND2_X1 U8771 ( .A1(n7487), .A2(n9465), .ZN(n8107) );
  INV_X1 U8772 ( .A(n9465), .ZN(n10713) );
  NAND2_X1 U8773 ( .A1(n9556), .A2(n10713), .ZN(n8105) );
  NAND2_X1 U8774 ( .A1(n8107), .A2(n8105), .ZN(n7505) );
  NAND2_X1 U8775 ( .A1(n8112), .A2(n8106), .ZN(n7522) );
  INV_X1 U8776 ( .A(n7522), .ZN(n8034) );
  INV_X1 U8777 ( .A(n7517), .ZN(n8132) );
  AOI21_X1 U8778 ( .B1(n7488), .B2(n8034), .A(n8132), .ZN(n7489) );
  XOR2_X1 U8779 ( .A(n7505), .B(n7489), .Z(n7490) );
  AOI22_X1 U8780 ( .A1(n7490), .A2(n10752), .B1(n10759), .B2(n9557), .ZN(
        n10712) );
  XNOR2_X1 U8781 ( .A(n7537), .B(n10713), .ZN(n7499) );
  NAND2_X1 U8782 ( .A1(n8070), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7498) );
  NAND2_X1 U8783 ( .A1(n8071), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7497) );
  INV_X1 U8784 ( .A(n7527), .ZN(n7529) );
  INV_X1 U8785 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U8786 ( .A1(n7493), .A2(n7492), .ZN(n7494) );
  AND2_X1 U8787 ( .A1(n7529), .A2(n7494), .ZN(n9355) );
  NAND2_X1 U8788 ( .A1(n7948), .A2(n9355), .ZN(n7496) );
  NAND2_X1 U8789 ( .A1(n8072), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7495) );
  NAND4_X1 U8790 ( .A1(n7498), .A2(n7497), .A3(n7496), .A4(n7495), .ZN(n9555)
         );
  AOI22_X1 U8791 ( .A1(n7499), .A2(n10762), .B1(n10756), .B2(n9555), .ZN(
        n10711) );
  INV_X1 U8792 ( .A(n10711), .ZN(n7502) );
  AOI22_X1 U8793 ( .A1(n10786), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9459), .B2(
        n10775), .ZN(n7500) );
  OAI21_X1 U8794 ( .B1(n10713), .B2(n9976), .A(n7500), .ZN(n7501) );
  AOI21_X1 U8795 ( .B1(n7502), .B2(n9972), .A(n7501), .ZN(n7508) );
  OR2_X1 U8796 ( .A1(n9557), .A2(n9179), .ZN(n7503) );
  NAND2_X1 U8797 ( .A1(n7504), .A2(n7503), .ZN(n7506) );
  NAND2_X1 U8798 ( .A1(n7506), .A2(n7505), .ZN(n7510) );
  OAI21_X1 U8799 ( .B1(n7506), .B2(n7505), .A(n7510), .ZN(n10715) );
  NAND2_X1 U8800 ( .A1(n10715), .A2(n10781), .ZN(n7507) );
  OAI211_X1 U8801 ( .C1(n10712), .C2(n10786), .A(n7508), .B(n7507), .ZN(
        P1_U3284) );
  NAND2_X1 U8802 ( .A1(n7487), .A2(n10713), .ZN(n7509) );
  NAND2_X1 U8803 ( .A1(n7510), .A2(n7509), .ZN(n7516) );
  INV_X1 U8804 ( .A(n9555), .ZN(n7515) );
  NAND2_X1 U8805 ( .A1(n7511), .A2(n8043), .ZN(n7514) );
  AOI22_X1 U8806 ( .A1(n8046), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8045), .B2(
        n7512), .ZN(n7513) );
  NAND2_X1 U8807 ( .A1(n7514), .A2(n7513), .ZN(n9188) );
  NAND2_X1 U8808 ( .A1(n7515), .A2(n9188), .ZN(n8119) );
  NAND2_X1 U8809 ( .A1(n8119), .A2(n8250), .ZN(n8036) );
  NAND2_X1 U8810 ( .A1(n7516), .A2(n8036), .ZN(n7609) );
  OAI21_X1 U8811 ( .B1(n7516), .B2(n8036), .A(n7609), .ZN(n10732) );
  INV_X1 U8812 ( .A(n10732), .ZN(n7543) );
  INV_X1 U8813 ( .A(n8036), .ZN(n7525) );
  NAND2_X1 U8814 ( .A1(n7517), .A2(n8105), .ZN(n7520) );
  NAND2_X1 U8815 ( .A1(n8104), .A2(n8113), .ZN(n7518) );
  NOR2_X1 U8816 ( .A1(n7520), .A2(n7518), .ZN(n8244) );
  INV_X1 U8817 ( .A(n7520), .ZN(n7521) );
  INV_X1 U8818 ( .A(n8107), .ZN(n8125) );
  AOI21_X1 U8819 ( .B1(n7522), .B2(n7521), .A(n8125), .ZN(n8245) );
  NAND2_X1 U8820 ( .A1(n7523), .A2(n8245), .ZN(n7524) );
  OAI21_X1 U8821 ( .B1(n7525), .B2(n7524), .A(n7621), .ZN(n7526) );
  NAND2_X1 U8822 ( .A1(n7526), .A2(n10752), .ZN(n7536) );
  NAND2_X1 U8823 ( .A1(n8072), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7534) );
  NAND2_X1 U8824 ( .A1(n8070), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U8825 ( .A1(n7527), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7615) );
  INV_X1 U8826 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U8827 ( .A1(n7529), .A2(n7528), .ZN(n7530) );
  AND2_X1 U8828 ( .A1(n7615), .A2(n7530), .ZN(n9513) );
  NAND2_X1 U8829 ( .A1(n7948), .A2(n9513), .ZN(n7532) );
  NAND2_X1 U8830 ( .A1(n8071), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7531) );
  NAND4_X1 U8831 ( .A1(n7534), .A2(n7533), .A3(n7532), .A4(n7531), .ZN(n10758)
         );
  AOI22_X1 U8832 ( .A1(n10759), .A2(n9556), .B1(n10758), .B2(n10756), .ZN(
        n7535) );
  NAND2_X1 U8833 ( .A1(n7536), .A2(n7535), .ZN(n10731) );
  OAI211_X1 U8834 ( .C1(n7538), .C2(n10729), .A(n7630), .B(n10762), .ZN(n10728) );
  NOR2_X1 U8835 ( .A1(n10728), .A2(n10658), .ZN(n7541) );
  AOI22_X1 U8836 ( .A1(n10786), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n9355), .B2(
        n10775), .ZN(n7539) );
  OAI21_X1 U8837 ( .B1(n10729), .B2(n9976), .A(n7539), .ZN(n7540) );
  AOI211_X1 U8838 ( .C1(n10731), .C2(n10560), .A(n7541), .B(n7540), .ZN(n7542)
         );
  OAI21_X1 U8839 ( .B1(n7543), .B2(n9979), .A(n7542), .ZN(P1_U3283) );
  INV_X1 U8840 ( .A(n7962), .ZN(n7547) );
  INV_X1 U8841 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7544) );
  OAI222_X1 U8842 ( .A1(n7545), .A2(P2_U3151), .B1(n9162), .B2(n7547), .C1(
        n7544), .C2(n9153), .ZN(P2_U3273) );
  INV_X1 U8843 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7548) );
  OAI222_X1 U8844 ( .A1(n10132), .A2(n7548), .B1(n10138), .B2(n7547), .C1(
        n7546), .C2(P1_U3086), .ZN(P1_U3333) );
  XNOR2_X1 U8845 ( .A(n7551), .B(n8335), .ZN(n10740) );
  XOR2_X1 U8846 ( .A(n7552), .B(n8335), .Z(n7555) );
  AOI22_X1 U8847 ( .A1(n10637), .A2(n8704), .B1(n8702), .B2(n6190), .ZN(n7554)
         );
  NAND2_X1 U8848 ( .A1(n10740), .A2(n10634), .ZN(n7553) );
  OAI211_X1 U8849 ( .C1(n7555), .C2(n9000), .A(n7554), .B(n7553), .ZN(n10737)
         );
  AOI21_X1 U8850 ( .B1(n8832), .B2(n10740), .A(n10737), .ZN(n7558) );
  OAI22_X1 U8851 ( .A1(n10709), .A2(n6283), .B1(n7774), .B2(n10650), .ZN(n7556) );
  AOI21_X1 U8852 ( .B1(n10704), .B2(n10735), .A(n7556), .ZN(n7557) );
  OAI21_X1 U8853 ( .B1(n7558), .B2(n9017), .A(n7557), .ZN(P2_U3223) );
  INV_X1 U8854 ( .A(n7953), .ZN(n7563) );
  OR2_X1 U8855 ( .A1(n7559), .A2(P1_U3086), .ZN(n8297) );
  INV_X1 U8856 ( .A(n8297), .ZN(n8291) );
  AOI21_X1 U8857 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10126), .A(n8291), .ZN(
        n7560) );
  OAI21_X1 U8858 ( .B1(n7563), .B2(n10138), .A(n7560), .ZN(P1_U3332) );
  NAND2_X1 U8859 ( .A1(n9160), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7562) );
  OR2_X1 U8860 ( .A1(n7561), .A2(P2_U3151), .ZN(n8522) );
  OAI211_X1 U8861 ( .C1(n7563), .C2(n9162), .A(n7562), .B(n8522), .ZN(P2_U3272) );
  XOR2_X1 U8862 ( .A(n7564), .B(n8339), .Z(n10743) );
  XNOR2_X1 U8863 ( .A(n7565), .B(n8339), .ZN(n7566) );
  OAI222_X1 U8864 ( .A1(n9005), .A2(n8627), .B1(n9003), .B2(n8641), .C1(n9000), 
        .C2(n7566), .ZN(n10745) );
  NAND2_X1 U8865 ( .A1(n10745), .A2(n10709), .ZN(n7570) );
  OAI22_X1 U8866 ( .A1(n10709), .A2(n7567), .B1(n8645), .B2(n10650), .ZN(n7568) );
  AOI21_X1 U8867 ( .B1(n10746), .B2(n10704), .A(n7568), .ZN(n7569) );
  OAI211_X1 U8868 ( .C1(n8968), .C2(n10743), .A(n7570), .B(n7569), .ZN(
        P2_U3222) );
  AOI21_X1 U8869 ( .B1(n5916), .B2(n7572), .A(n7571), .ZN(n7587) );
  AOI21_X1 U8870 ( .B1(n7574), .B2(n7567), .A(n7573), .ZN(n7577) );
  NAND2_X1 U8871 ( .A1(n10516), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7576) );
  AND2_X1 U8872 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8643) );
  INV_X1 U8873 ( .A(n8643), .ZN(n7575) );
  OAI211_X1 U8874 ( .C1(n7577), .C2(n10496), .A(n7576), .B(n7575), .ZN(n7580)
         );
  NOR2_X1 U8875 ( .A1(n10511), .A2(n7578), .ZN(n7579) );
  NOR2_X1 U8876 ( .A1(n7580), .A2(n7579), .ZN(n7586) );
  OAI21_X1 U8877 ( .B1(n7583), .B2(n7582), .A(n7581), .ZN(n7584) );
  NAND2_X1 U8878 ( .A1(n7584), .A2(n10519), .ZN(n7585) );
  OAI211_X1 U8879 ( .C1(n7587), .C2(n10514), .A(n7586), .B(n7585), .ZN(
        P2_U3193) );
  AND2_X1 U8880 ( .A1(n7589), .A2(n7588), .ZN(n8433) );
  XNOR2_X1 U8881 ( .A(n7590), .B(n8433), .ZN(n7593) );
  NAND2_X1 U8882 ( .A1(n8702), .A2(n10637), .ZN(n7591) );
  OAI21_X1 U8883 ( .B1(n8566), .B2(n9005), .A(n7591), .ZN(n7592) );
  AOI21_X1 U8884 ( .B1(n7593), .B2(n10641), .A(n7592), .ZN(n7691) );
  OAI22_X1 U8885 ( .A1(n10709), .A2(n6285), .B1(n8569), .B2(n10650), .ZN(n7594) );
  AOI21_X1 U8886 ( .B1(n8575), .B2(n10704), .A(n7594), .ZN(n7597) );
  INV_X1 U8887 ( .A(n8433), .ZN(n8337) );
  XNOR2_X1 U8888 ( .A(n7595), .B(n8337), .ZN(n7690) );
  NAND2_X1 U8889 ( .A1(n7690), .A2(n9015), .ZN(n7596) );
  OAI211_X1 U8890 ( .C1(n7691), .C2(n9017), .A(n7597), .B(n7596), .ZN(P2_U3221) );
  AOI211_X1 U8891 ( .C1(n10693), .C2(n7600), .A(n7599), .B(n7598), .ZN(n7608)
         );
  INV_X1 U8892 ( .A(n10069), .ZN(n7602) );
  AOI22_X1 U8893 ( .A1(n7602), .A2(n7601), .B1(n10768), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7603) );
  OAI21_X1 U8894 ( .B1(n7608), .B2(n10768), .A(n7603), .ZN(P1_U3529) );
  INV_X1 U8895 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7604) );
  OAI22_X1 U8896 ( .A1(n10122), .A2(n7605), .B1(n10774), .B2(n7604), .ZN(n7606) );
  INV_X1 U8897 ( .A(n7606), .ZN(n7607) );
  OAI21_X1 U8898 ( .B1(n7608), .B2(n10771), .A(n7607), .ZN(P1_U3474) );
  OAI21_X1 U8899 ( .B1(n9555), .B2(n9188), .A(n7609), .ZN(n7702) );
  INV_X1 U8900 ( .A(n10758), .ZN(n9415) );
  NAND2_X1 U8901 ( .A1(n7610), .A2(n8043), .ZN(n7613) );
  AOI22_X1 U8902 ( .A1(n8046), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8045), .B2(
        n7611), .ZN(n7612) );
  OR2_X1 U8903 ( .A1(n9415), .A2(n9197), .ZN(n8130) );
  NAND2_X1 U8904 ( .A1(n9197), .A2(n9415), .ZN(n8128) );
  XNOR2_X1 U8905 ( .A(n7702), .B(n8038), .ZN(n7754) );
  NAND2_X1 U8906 ( .A1(n8070), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7620) );
  NAND2_X1 U8907 ( .A1(n8071), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7619) );
  INV_X1 U8908 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7614) );
  NAND2_X1 U8909 ( .A1(n7615), .A2(n7614), .ZN(n7616) );
  AND2_X1 U8910 ( .A1(n7712), .A2(n7616), .ZN(n10776) );
  NAND2_X1 U8911 ( .A1(n7948), .A2(n10776), .ZN(n7618) );
  NAND2_X1 U8912 ( .A1(n8072), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7617) );
  NAND4_X1 U8913 ( .A1(n7620), .A2(n7619), .A3(n7618), .A4(n7617), .ZN(n9554)
         );
  AOI22_X1 U8914 ( .A1(n10759), .A2(n9555), .B1(n9554), .B2(n10756), .ZN(n7628) );
  INV_X1 U8915 ( .A(n8130), .ZN(n7626) );
  AND2_X1 U8916 ( .A1(n8128), .A2(n8119), .ZN(n8248) );
  NAND2_X1 U8917 ( .A1(n7621), .A2(n8248), .ZN(n7718) );
  INV_X1 U8918 ( .A(n7621), .ZN(n7624) );
  INV_X1 U8919 ( .A(n8119), .ZN(n7623) );
  INV_X1 U8920 ( .A(n8038), .ZN(n7622) );
  OAI21_X1 U8921 ( .B1(n7624), .B2(n7623), .A(n7622), .ZN(n7625) );
  OAI211_X1 U8922 ( .C1(n7626), .C2(n7718), .A(n7625), .B(n10752), .ZN(n7627)
         );
  OAI211_X1 U8923 ( .C1(n7754), .C2(n7629), .A(n7628), .B(n7627), .ZN(n7755)
         );
  NAND2_X1 U8924 ( .A1(n7755), .A2(n10560), .ZN(n7634) );
  INV_X1 U8925 ( .A(n7733), .ZN(n10764) );
  AOI211_X1 U8926 ( .C1(n9197), .C2(n7630), .A(n10764), .B(n9915), .ZN(n7756)
         );
  INV_X1 U8927 ( .A(n9197), .ZN(n9510) );
  AOI22_X1 U8928 ( .A1(n10786), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9513), .B2(
        n10775), .ZN(n7631) );
  OAI21_X1 U8929 ( .B1(n9510), .B2(n9976), .A(n7631), .ZN(n7632) );
  AOI21_X1 U8930 ( .B1(n7756), .B2(n9972), .A(n7632), .ZN(n7633) );
  OAI211_X1 U8931 ( .C1(n7754), .C2(n7635), .A(n7634), .B(n7633), .ZN(P1_U3282) );
  AOI21_X1 U8932 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n7781), .A(n7636), .ZN(
        n9609) );
  XNOR2_X1 U8933 ( .A(n9618), .B(n9609), .ZN(n7637) );
  INV_X1 U8934 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U8935 ( .A1(n10062), .A2(n7637), .ZN(n9610) );
  AOI21_X1 U8936 ( .B1(n7637), .B2(n10062), .A(n9610), .ZN(n7645) );
  INV_X1 U8937 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7639) );
  INV_X1 U8938 ( .A(n9618), .ZN(n8023) );
  NAND2_X1 U8939 ( .A1(n10542), .A2(n8023), .ZN(n7638) );
  NAND2_X1 U8940 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9540) );
  OAI211_X1 U8941 ( .C1(n7639), .C2(n9669), .A(n7638), .B(n9540), .ZN(n7644)
         );
  AOI21_X1 U8942 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7781), .A(n7640), .ZN(
        n9619) );
  XNOR2_X1 U8943 ( .A(n9618), .B(n9619), .ZN(n7642) );
  INV_X1 U8944 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7641) );
  NOR2_X1 U8945 ( .A1(n7641), .A2(n7642), .ZN(n9620) );
  AOI211_X1 U8946 ( .C1(n7642), .C2(n7641), .A(n9620), .B(n9623), .ZN(n7643)
         );
  AOI211_X1 U8947 ( .C1(n9644), .C2(n7645), .A(n7644), .B(n7643), .ZN(n7646)
         );
  INV_X1 U8948 ( .A(n7646), .ZN(P1_U3258) );
  AOI21_X1 U8949 ( .B1(n8663), .B2(n8705), .A(n7647), .ZN(n7649) );
  OR2_X1 U8950 ( .A1(n8641), .A2(n8660), .ZN(n7648) );
  OAI211_X1 U8951 ( .C1(n8683), .C2(n7650), .A(n7649), .B(n7648), .ZN(n7660)
         );
  XNOR2_X1 U8952 ( .A(n10724), .B(n7870), .ZN(n7762) );
  XNOR2_X1 U8953 ( .A(n7762), .B(n8704), .ZN(n7658) );
  NAND2_X1 U8954 ( .A1(n7651), .A2(n5437), .ZN(n7652) );
  NAND2_X1 U8955 ( .A1(n7653), .A2(n7652), .ZN(n7657) );
  INV_X1 U8956 ( .A(n7657), .ZN(n7655) );
  INV_X1 U8957 ( .A(n7764), .ZN(n7656) );
  AOI211_X1 U8958 ( .C1(n7658), .C2(n7657), .A(n8676), .B(n7656), .ZN(n7659)
         );
  AOI211_X1 U8959 ( .C1(n10724), .C2(n8673), .A(n7660), .B(n7659), .ZN(n7661)
         );
  INV_X1 U8960 ( .A(n7661), .ZN(P2_U3171) );
  AOI21_X1 U8961 ( .B1(n7664), .B2(n7663), .A(n7662), .ZN(n7680) );
  INV_X1 U8962 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7672) );
  AND2_X1 U8963 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3151), .ZN(n7771) );
  AND2_X1 U8964 ( .A1(n7666), .A2(n7665), .ZN(n7668) );
  OAI21_X1 U8965 ( .B1(n7669), .B2(n7668), .A(n10519), .ZN(n7667) );
  AOI21_X1 U8966 ( .B1(n7669), .B2(n7668), .A(n7667), .ZN(n7670) );
  NOR2_X1 U8967 ( .A1(n7771), .A2(n7670), .ZN(n7671) );
  OAI21_X1 U8968 ( .B1(n10506), .B2(n7672), .A(n7671), .ZN(n7677) );
  AOI21_X1 U8969 ( .B1(n5034), .B2(n7674), .A(n7673), .ZN(n7675) );
  NOR2_X1 U8970 ( .A1(n7675), .A2(n10496), .ZN(n7676) );
  AOI211_X1 U8971 ( .C1(n10434), .C2(n7678), .A(n7677), .B(n7676), .ZN(n7679)
         );
  OAI21_X1 U8972 ( .B1(n7680), .B2(n10514), .A(n7679), .ZN(P2_U3192) );
  INV_X1 U8973 ( .A(n8432), .ZN(n8342) );
  XNOR2_X1 U8974 ( .A(n7681), .B(n8342), .ZN(n10788) );
  XNOR2_X1 U8975 ( .A(n7682), .B(n8342), .ZN(n7683) );
  NAND2_X1 U8976 ( .A1(n7683), .A2(n10641), .ZN(n7685) );
  AOI22_X1 U8977 ( .A1(n6190), .A2(n8699), .B1(n8701), .B2(n10637), .ZN(n7684)
         );
  NAND2_X1 U8978 ( .A1(n7685), .A2(n7684), .ZN(n10789) );
  INV_X1 U8979 ( .A(n8361), .ZN(n10787) );
  OAI22_X1 U8980 ( .A1(n10787), .A2(n10598), .B1(n8628), .B2(n10650), .ZN(
        n7686) );
  OAI21_X1 U8981 ( .B1(n10789), .B2(n7686), .A(n10709), .ZN(n7688) );
  NAND2_X1 U8982 ( .A1(n9017), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7687) );
  OAI211_X1 U8983 ( .C1(n10788), .C2(n8968), .A(n7688), .B(n7687), .ZN(
        P2_U3220) );
  INV_X1 U8984 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7693) );
  AND2_X1 U8985 ( .A1(n8575), .A2(n10747), .ZN(n7689) );
  AOI21_X1 U8986 ( .B1(n7690), .B2(n10720), .A(n7689), .ZN(n7692) );
  AND2_X1 U8987 ( .A1(n7692), .A2(n7691), .ZN(n7695) );
  MUX2_X1 U8988 ( .A(n7693), .B(n7695), .S(n10810), .Z(n7694) );
  INV_X1 U8989 ( .A(n7694), .ZN(P2_U3426) );
  MUX2_X1 U8990 ( .A(n5932), .B(n7695), .S(n10806), .Z(n7696) );
  INV_X1 U8991 ( .A(n7696), .ZN(P2_U3471) );
  INV_X1 U8992 ( .A(n7943), .ZN(n7699) );
  OAI222_X1 U8993 ( .A1(n7698), .A2(P2_U3151), .B1(n9162), .B2(n7699), .C1(
        n7697), .C2(n9153), .ZN(P2_U3271) );
  OAI222_X1 U8994 ( .A1(n10132), .A2(n7701), .B1(P1_U3086), .B2(n7700), .C1(
        n7699), .C2(n10138), .ZN(P1_U3331) );
  NAND2_X1 U8995 ( .A1(n7703), .A2(n8043), .ZN(n7706) );
  AOI22_X1 U8996 ( .A1(n8046), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8045), .B2(
        n7704), .ZN(n7705) );
  INV_X1 U8997 ( .A(n9554), .ZN(n9509) );
  NAND2_X1 U8998 ( .A1(n10778), .A2(n9509), .ZN(n8136) );
  NAND2_X1 U8999 ( .A1(n7707), .A2(n8043), .ZN(n7710) );
  AOI22_X1 U9000 ( .A1(n8046), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8045), .B2(
        n7708), .ZN(n7709) );
  NAND2_X1 U9001 ( .A1(n8070), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U9002 ( .A1(n8071), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7716) );
  INV_X1 U9003 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7711) );
  NAND2_X1 U9004 ( .A1(n7712), .A2(n7711), .ZN(n7713) );
  AND2_X1 U9005 ( .A1(n7725), .A2(n7713), .ZN(n9485) );
  NAND2_X1 U9006 ( .A1(n7948), .A2(n9485), .ZN(n7715) );
  NAND2_X1 U9007 ( .A1(n8072), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7714) );
  NAND4_X1 U9008 ( .A1(n7717), .A2(n7716), .A3(n7715), .A4(n7714), .ZN(n10757)
         );
  INV_X1 U9009 ( .A(n10757), .ZN(n7778) );
  OR2_X1 U9010 ( .A1(n9212), .A2(n7778), .ZN(n8138) );
  NAND2_X1 U9011 ( .A1(n9212), .A2(n7778), .ZN(n8142) );
  NAND2_X1 U9012 ( .A1(n8138), .A2(n8142), .ZN(n8026) );
  XNOR2_X1 U9013 ( .A(n7779), .B(n8026), .ZN(n7806) );
  INV_X1 U9014 ( .A(n7806), .ZN(n7739) );
  NAND2_X1 U9015 ( .A1(n7718), .A2(n8130), .ZN(n10754) );
  NAND2_X1 U9016 ( .A1(n10754), .A2(n10755), .ZN(n10753) );
  NAND2_X1 U9017 ( .A1(n10753), .A2(n8139), .ZN(n7719) );
  NAND2_X1 U9018 ( .A1(n7719), .A2(n8026), .ZN(n7722) );
  INV_X1 U9019 ( .A(n8139), .ZN(n7720) );
  NOR2_X1 U9020 ( .A1(n8026), .A2(n7720), .ZN(n7721) );
  NAND2_X1 U9021 ( .A1(n7722), .A2(n7784), .ZN(n7723) );
  NAND2_X1 U9022 ( .A1(n7723), .A2(n10752), .ZN(n7732) );
  NAND2_X1 U9023 ( .A1(n8070), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7730) );
  NAND2_X1 U9024 ( .A1(n8072), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7729) );
  INV_X1 U9025 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7724) );
  INV_X1 U9026 ( .A(n7786), .ZN(n7788) );
  NAND2_X1 U9027 ( .A1(n7725), .A2(n7724), .ZN(n7726) );
  AND2_X1 U9028 ( .A1(n7788), .A2(n7726), .ZN(n9334) );
  NAND2_X1 U9029 ( .A1(n7948), .A2(n9334), .ZN(n7728) );
  NAND2_X1 U9030 ( .A1(n8071), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7727) );
  NAND4_X1 U9031 ( .A1(n7730), .A2(n7729), .A3(n7728), .A4(n7727), .ZN(n9965)
         );
  AOI22_X1 U9032 ( .A1(n10756), .A2(n9965), .B1(n9554), .B2(n10759), .ZN(n7731) );
  NAND2_X1 U9033 ( .A1(n7732), .A2(n7731), .ZN(n7804) );
  INV_X1 U9034 ( .A(n7734), .ZN(n10763) );
  AOI211_X1 U9035 ( .C1(n9212), .C2(n10763), .A(n9915), .B(n7796), .ZN(n7805)
         );
  NAND2_X1 U9036 ( .A1(n7805), .A2(n9972), .ZN(n7736) );
  AOI22_X1 U9037 ( .A1(n10786), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9485), .B2(
        n10775), .ZN(n7735) );
  OAI211_X1 U9038 ( .C1(n9488), .C2(n9976), .A(n7736), .B(n7735), .ZN(n7737)
         );
  AOI21_X1 U9039 ( .B1(n7804), .B2(n10560), .A(n7737), .ZN(n7738) );
  OAI21_X1 U9040 ( .B1(n7739), .B2(n9979), .A(n7738), .ZN(P1_U3280) );
  INV_X1 U9041 ( .A(n7934), .ZN(n7743) );
  OAI222_X1 U9042 ( .A1(n7741), .A2(P2_U3151), .B1(n9162), .B2(n7743), .C1(
        n7740), .C2(n9153), .ZN(P2_U3270) );
  OAI222_X1 U9043 ( .A1(P1_U3086), .A2(n7744), .B1(n10138), .B2(n7743), .C1(
        n7742), .C2(n10132), .ZN(P1_U3330) );
  INV_X1 U9044 ( .A(n8438), .ZN(n8340) );
  OAI21_X1 U9045 ( .B1(n5026), .B2(n8340), .A(n7745), .ZN(n10794) );
  XNOR2_X1 U9046 ( .A(n7746), .B(n8438), .ZN(n7747) );
  NAND2_X1 U9047 ( .A1(n7747), .A2(n10641), .ZN(n7749) );
  AOI22_X1 U9048 ( .A1(n8700), .A2(n10637), .B1(n6190), .B2(n8698), .ZN(n7748)
         );
  NAND2_X1 U9049 ( .A1(n7749), .A2(n7748), .ZN(n10795) );
  INV_X1 U9050 ( .A(n8357), .ZN(n10793) );
  NOR2_X1 U9051 ( .A1(n10793), .A2(n10598), .ZN(n7750) );
  OAI21_X1 U9052 ( .B1(n10795), .B2(n7750), .A(n10709), .ZN(n7753) );
  INV_X1 U9053 ( .A(n8538), .ZN(n7751) );
  AOI22_X1 U9054 ( .A1(n9017), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n10706), .B2(
        n7751), .ZN(n7752) );
  OAI211_X1 U9055 ( .C1(n8968), .C2(n10794), .A(n7753), .B(n7752), .ZN(
        P2_U3219) );
  INV_X1 U9056 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7758) );
  INV_X1 U9057 ( .A(n7754), .ZN(n7757) );
  AOI211_X1 U9058 ( .C1(n10693), .C2(n7757), .A(n7756), .B(n7755), .ZN(n7760)
         );
  MUX2_X1 U9059 ( .A(n7758), .B(n7760), .S(n10774), .Z(n7759) );
  OAI21_X1 U9060 ( .B1(n9510), .B2(n10122), .A(n7759), .ZN(P1_U3486) );
  MUX2_X1 U9061 ( .A(n6708), .B(n7760), .S(n10770), .Z(n7761) );
  OAI21_X1 U9062 ( .B1(n9510), .B2(n10069), .A(n7761), .ZN(P1_U3533) );
  NAND2_X1 U9063 ( .A1(n7762), .A2(n8704), .ZN(n7763) );
  XNOR2_X1 U9064 ( .A(n10735), .B(n7874), .ZN(n7765) );
  INV_X1 U9065 ( .A(n7765), .ZN(n7766) );
  INV_X1 U9066 ( .A(n7768), .ZN(n7770) );
  INV_X1 U9067 ( .A(n8649), .ZN(n7769) );
  AOI21_X1 U9068 ( .B1(n8703), .B2(n7770), .A(n7769), .ZN(n7777) );
  AOI21_X1 U9069 ( .B1(n8663), .B2(n8704), .A(n7771), .ZN(n7773) );
  NAND2_X1 U9070 ( .A1(n8702), .A2(n8686), .ZN(n7772) );
  OAI211_X1 U9071 ( .C1(n8683), .C2(n7774), .A(n7773), .B(n7772), .ZN(n7775)
         );
  AOI21_X1 U9072 ( .B1(n10735), .B2(n8673), .A(n7775), .ZN(n7776) );
  OAI21_X1 U9073 ( .B1(n7777), .B2(n8676), .A(n7776), .ZN(P2_U3157) );
  NAND2_X1 U9074 ( .A1(n7780), .A2(n8043), .ZN(n7783) );
  AOI22_X1 U9075 ( .A1(n8046), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8045), .B2(
        n7781), .ZN(n7782) );
  XNOR2_X1 U9076 ( .A(n9708), .B(n9707), .ZN(n8141) );
  XOR2_X1 U9077 ( .A(n9711), .B(n8141), .Z(n10066) );
  INV_X1 U9078 ( .A(n10066), .ZN(n7803) );
  INV_X1 U9079 ( .A(n8141), .ZN(n7785) );
  OAI211_X1 U9080 ( .C1(n5028), .C2(n7785), .A(n10752), .B(n9961), .ZN(n7795)
         );
  NAND2_X1 U9081 ( .A1(n8070), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7793) );
  NAND2_X1 U9082 ( .A1(n8071), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U9083 ( .A1(n7786), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8015) );
  INV_X1 U9084 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U9085 ( .A1(n7788), .A2(n7787), .ZN(n7789) );
  AND2_X1 U9086 ( .A1(n8015), .A2(n7789), .ZN(n9973) );
  NAND2_X1 U9087 ( .A1(n7948), .A2(n9973), .ZN(n7791) );
  NAND2_X1 U9088 ( .A1(n8072), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7790) );
  NAND4_X1 U9089 ( .A1(n7793), .A2(n7792), .A3(n7791), .A4(n7790), .ZN(n9553)
         );
  AOI22_X1 U9090 ( .A1(n10759), .A2(n10757), .B1(n9553), .B2(n10756), .ZN(
        n7794) );
  NAND2_X1 U9091 ( .A1(n7795), .A2(n7794), .ZN(n10064) );
  INV_X1 U9092 ( .A(n7796), .ZN(n7798) );
  NAND2_X1 U9093 ( .A1(n7796), .A2(n10123), .ZN(n9970) );
  INV_X1 U9094 ( .A(n9970), .ZN(n7797) );
  AOI211_X1 U9095 ( .C1(n9708), .C2(n7798), .A(n9915), .B(n7797), .ZN(n10065)
         );
  NAND2_X1 U9096 ( .A1(n10065), .A2(n9972), .ZN(n7800) );
  AOI22_X1 U9097 ( .A1(n10786), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9334), .B2(
        n10775), .ZN(n7799) );
  OAI211_X1 U9098 ( .C1(n10123), .C2(n9976), .A(n7800), .B(n7799), .ZN(n7801)
         );
  AOI21_X1 U9099 ( .B1(n10064), .B2(n10560), .A(n7801), .ZN(n7802) );
  OAI21_X1 U9100 ( .B1(n7803), .B2(n9979), .A(n7802), .ZN(P1_U3279) );
  INV_X1 U9101 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7807) );
  AOI211_X1 U9102 ( .C1(n7806), .C2(n10767), .A(n7805), .B(n7804), .ZN(n7809)
         );
  MUX2_X1 U9103 ( .A(n7807), .B(n7809), .S(n10774), .Z(n7808) );
  OAI21_X1 U9104 ( .B1(n9488), .B2(n10122), .A(n7808), .ZN(P1_U3492) );
  MUX2_X1 U9105 ( .A(n7058), .B(n7809), .S(n10770), .Z(n7810) );
  OAI21_X1 U9106 ( .B1(n9488), .B2(n10069), .A(n7810), .ZN(P1_U3535) );
  INV_X1 U9107 ( .A(n9007), .ZN(n7811) );
  AOI21_X1 U9108 ( .B1(n8341), .B2(n7812), .A(n7811), .ZN(n10802) );
  OAI22_X1 U9109 ( .A1(n10709), .A2(n7813), .B1(n8682), .B2(n10650), .ZN(n7814) );
  AOI21_X1 U9110 ( .B1(n8356), .B2(n10704), .A(n7814), .ZN(n7820) );
  INV_X1 U9111 ( .A(n8341), .ZN(n8445) );
  XNOR2_X1 U9112 ( .A(n7815), .B(n8445), .ZN(n7816) );
  NAND2_X1 U9113 ( .A1(n7816), .A2(n10641), .ZN(n7818) );
  AOI22_X1 U9114 ( .A1(n8697), .A2(n6190), .B1(n10637), .B2(n8699), .ZN(n7817)
         );
  NAND2_X1 U9115 ( .A1(n7818), .A2(n7817), .ZN(n10803) );
  NAND2_X1 U9116 ( .A1(n10803), .A2(n10709), .ZN(n7819) );
  OAI211_X1 U9117 ( .C1(n10802), .C2(n8968), .A(n7820), .B(n7819), .ZN(
        P2_U3218) );
  INV_X1 U9118 ( .A(n7925), .ZN(n7824) );
  OAI222_X1 U9119 ( .A1(n10132), .A2(n7822), .B1(n10138), .B2(n7824), .C1(
        P1_U3086), .C2(n7821), .ZN(P1_U3329) );
  OAI222_X1 U9120 ( .A1(P2_U3151), .A2(n7825), .B1(n9162), .B2(n7824), .C1(
        n7823), .C2(n9153), .ZN(P2_U3269) );
  NAND2_X1 U9121 ( .A1(n7826), .A2(n8647), .ZN(n7827) );
  XNOR2_X1 U9122 ( .A(n10746), .B(n7874), .ZN(n7829) );
  XNOR2_X1 U9123 ( .A(n7829), .B(n8702), .ZN(n8646) );
  NAND2_X1 U9124 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  XNOR2_X1 U9125 ( .A(n8575), .B(n7870), .ZN(n7835) );
  XNOR2_X1 U9126 ( .A(n7835), .B(n8701), .ZN(n8572) );
  XNOR2_X1 U9127 ( .A(n8361), .B(n7874), .ZN(n7832) );
  NAND2_X1 U9128 ( .A1(n7832), .A2(n8566), .ZN(n8532) );
  INV_X1 U9129 ( .A(n7832), .ZN(n7833) );
  NAND2_X1 U9130 ( .A1(n7833), .A2(n8700), .ZN(n7834) );
  NAND2_X1 U9131 ( .A1(n8532), .A2(n7834), .ZN(n8620) );
  AND2_X1 U9132 ( .A1(n7835), .A2(n8701), .ZN(n8619) );
  NOR2_X1 U9133 ( .A1(n8620), .A2(n8619), .ZN(n7836) );
  NAND2_X1 U9134 ( .A1(n8623), .A2(n7836), .ZN(n8531) );
  NAND2_X1 U9135 ( .A1(n8531), .A2(n8532), .ZN(n7837) );
  XNOR2_X1 U9136 ( .A(n8357), .B(n7874), .ZN(n7838) );
  XNOR2_X1 U9137 ( .A(n7838), .B(n8699), .ZN(n8533) );
  NAND2_X1 U9138 ( .A1(n7838), .A2(n8681), .ZN(n7839) );
  XNOR2_X1 U9139 ( .A(n8356), .B(n7870), .ZN(n7841) );
  XNOR2_X1 U9140 ( .A(n7841), .B(n8698), .ZN(n8677) );
  XNOR2_X1 U9141 ( .A(n9010), .B(n7870), .ZN(n8590) );
  INV_X1 U9142 ( .A(n8590), .ZN(n7840) );
  AND2_X1 U9143 ( .A1(n7840), .A2(n8988), .ZN(n7846) );
  XNOR2_X1 U9144 ( .A(n8599), .B(n7870), .ZN(n8593) );
  NAND2_X1 U9145 ( .A1(n7841), .A2(n8698), .ZN(n8584) );
  NAND2_X1 U9146 ( .A1(n8584), .A2(n8988), .ZN(n7842) );
  NAND2_X1 U9147 ( .A1(n8590), .A2(n7842), .ZN(n7843) );
  OAI21_X1 U9148 ( .B1(n8988), .B2(n8584), .A(n7843), .ZN(n7844) );
  AOI21_X1 U9149 ( .B1(n8593), .B2(n8696), .A(n7844), .ZN(n7845) );
  INV_X1 U9150 ( .A(n8593), .ZN(n7847) );
  NAND2_X1 U9151 ( .A1(n7847), .A2(n9004), .ZN(n7848) );
  NAND2_X1 U9152 ( .A1(n7849), .A2(n7848), .ZN(n8657) );
  XNOR2_X1 U9153 ( .A(n8655), .B(n7870), .ZN(n7853) );
  XNOR2_X1 U9154 ( .A(n7853), .B(n8958), .ZN(n8656) );
  XNOR2_X1 U9155 ( .A(n8956), .B(n7870), .ZN(n8551) );
  INV_X1 U9156 ( .A(n8551), .ZN(n7850) );
  NAND2_X1 U9157 ( .A1(n7850), .A2(n8944), .ZN(n7854) );
  INV_X1 U9158 ( .A(n7854), .ZN(n7851) );
  OR2_X1 U9159 ( .A1(n8656), .A2(n5566), .ZN(n7852) );
  NOR2_X1 U9160 ( .A1(n8657), .A2(n7852), .ZN(n7857) );
  NAND2_X1 U9161 ( .A1(n7853), .A2(n8958), .ZN(n8549) );
  AND2_X1 U9162 ( .A1(n8549), .A2(n7854), .ZN(n7855) );
  NOR2_X1 U9163 ( .A1(n5566), .A2(n7855), .ZN(n7856) );
  NOR2_X1 U9164 ( .A1(n7857), .A2(n7856), .ZN(n8611) );
  XNOR2_X1 U9165 ( .A(n8950), .B(n7874), .ZN(n7858) );
  XNOR2_X1 U9166 ( .A(n7858), .B(n8959), .ZN(n8610) );
  NAND2_X1 U9167 ( .A1(n7858), .A2(n8554), .ZN(n7859) );
  XNOR2_X1 U9168 ( .A(n9062), .B(n7874), .ZN(n7860) );
  XNOR2_X1 U9169 ( .A(n7860), .B(n8943), .ZN(n8559) );
  NAND2_X1 U9170 ( .A1(n8560), .A2(n8559), .ZN(n7862) );
  NAND2_X1 U9171 ( .A1(n7860), .A2(n8913), .ZN(n7861) );
  XNOR2_X1 U9172 ( .A(n8347), .B(n7870), .ZN(n7863) );
  XNOR2_X1 U9173 ( .A(n7863), .B(n8927), .ZN(n8633) );
  NAND2_X1 U9174 ( .A1(n7863), .A2(n8927), .ZN(n7864) );
  XOR2_X1 U9175 ( .A(n7874), .B(n8904), .Z(n7866) );
  XNOR2_X1 U9176 ( .A(n8891), .B(n7874), .ZN(n7867) );
  XNOR2_X1 U9177 ( .A(n7867), .B(n8694), .ZN(n8603) );
  XNOR2_X1 U9178 ( .A(n9045), .B(n7874), .ZN(n7868) );
  XOR2_X1 U9179 ( .A(n8693), .B(n7868), .Z(n8578) );
  INV_X1 U9180 ( .A(n7868), .ZN(n7869) );
  OAI22_X2 U9181 ( .A1(n8577), .A2(n8578), .B1(n7869), .B2(n8693), .ZN(n8666)
         );
  XNOR2_X1 U9182 ( .A(n8871), .B(n7870), .ZN(n7871) );
  NAND2_X1 U9183 ( .A1(n7871), .A2(n8692), .ZN(n8668) );
  NOR2_X1 U9184 ( .A1(n7871), .A2(n8692), .ZN(n8667) );
  XNOR2_X1 U9185 ( .A(n8859), .B(n7874), .ZN(n7872) );
  XNOR2_X1 U9186 ( .A(n7872), .B(n8843), .ZN(n8524) );
  INV_X1 U9187 ( .A(n7872), .ZN(n7873) );
  XNOR2_X1 U9188 ( .A(n8840), .B(n7874), .ZN(n7875) );
  OAI22_X1 U9189 ( .A1(n8868), .A2(n8680), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10325), .ZN(n7876) );
  AOI21_X1 U9190 ( .B1(n8686), .B2(n8844), .A(n7876), .ZN(n7877) );
  OAI21_X1 U9191 ( .B1(n7878), .B2(n8683), .A(n7877), .ZN(n7879) );
  AOI21_X1 U9192 ( .B1(n8839), .B2(n8673), .A(n7879), .ZN(n7880) );
  INV_X1 U9193 ( .A(SI_29_), .ZN(n10266) );
  INV_X1 U9194 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8303) );
  INV_X1 U9195 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7885) );
  MUX2_X1 U9196 ( .A(n8303), .B(n7885), .S(n5056), .Z(n7886) );
  INV_X1 U9197 ( .A(SI_30_), .ZN(n10262) );
  NAND2_X1 U9198 ( .A1(n7886), .A2(n10262), .ZN(n7889) );
  INV_X1 U9199 ( .A(n7886), .ZN(n7887) );
  NAND2_X1 U9200 ( .A1(n7887), .A2(SI_30_), .ZN(n7888) );
  NAND2_X1 U9201 ( .A1(n7889), .A2(n7888), .ZN(n8066) );
  MUX2_X1 U9202 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n5056), .Z(n7892) );
  INV_X1 U9203 ( .A(SI_31_), .ZN(n7891) );
  XNOR2_X1 U9204 ( .A(n7892), .B(n7891), .ZN(n7893) );
  NAND2_X1 U9205 ( .A1(n9145), .A2(n8043), .ZN(n7897) );
  INV_X1 U9206 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7895) );
  OR2_X1 U9207 ( .A1(n6943), .A2(n7895), .ZN(n7896) );
  NAND2_X1 U9208 ( .A1(n7898), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7901) );
  NAND2_X1 U9209 ( .A1(n8071), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U9210 ( .A1(n8072), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7899) );
  OR2_X1 U9211 ( .A1(n9682), .A2(n9686), .ZN(n8218) );
  INV_X1 U9212 ( .A(n8218), .ZN(n8285) );
  NAND2_X1 U9213 ( .A1(n9682), .A2(n9686), .ZN(n8222) );
  INV_X1 U9214 ( .A(n8222), .ZN(n8289) );
  OR2_X1 U9215 ( .A1(n6943), .A2(n10131), .ZN(n7902) );
  NAND2_X1 U9216 ( .A1(n8072), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7907) );
  NAND2_X1 U9217 ( .A1(n8070), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7906) );
  INV_X1 U9218 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8014) );
  INV_X1 U9219 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8005) );
  NAND2_X1 U9220 ( .A1(n8049), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7995) );
  INV_X1 U9221 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U9222 ( .A1(n7984), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7975) );
  NAND2_X1 U9223 ( .A1(n7947), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7937) );
  INV_X1 U9224 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7929) );
  NAND3_X1 U9225 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .A3(n7928), .ZN(n7913) );
  INV_X1 U9226 ( .A(n7913), .ZN(n9732) );
  NAND2_X1 U9227 ( .A1(n7948), .A2(n9732), .ZN(n7905) );
  NAND2_X1 U9228 ( .A1(n5558), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U9229 ( .A1(n9155), .A2(n8043), .ZN(n7909) );
  INV_X1 U9230 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10133) );
  OR2_X1 U9231 ( .A1(n6943), .A2(n10133), .ZN(n7908) );
  NAND2_X1 U9232 ( .A1(n8070), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7917) );
  NAND2_X1 U9233 ( .A1(n8072), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7916) );
  INV_X1 U9234 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U9235 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n7928), .ZN(n7910) );
  NAND2_X1 U9236 ( .A1(n7911), .A2(n7910), .ZN(n7912) );
  NAND2_X1 U9237 ( .A1(n7948), .A2(n9749), .ZN(n7915) );
  NAND2_X1 U9238 ( .A1(n8071), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7914) );
  NAND2_X1 U9239 ( .A1(n9995), .A2(n9728), .ZN(n9703) );
  NAND2_X1 U9240 ( .A1(n9158), .A2(n8043), .ZN(n7919) );
  NAND2_X1 U9241 ( .A1(n8046), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7918) );
  NAND2_X1 U9242 ( .A1(n8072), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7924) );
  NAND2_X1 U9243 ( .A1(n8070), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7923) );
  INV_X1 U9244 ( .A(n7928), .ZN(n7920) );
  XNOR2_X1 U9245 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n7920), .ZN(n9766) );
  NAND2_X1 U9246 ( .A1(n8054), .A2(n9766), .ZN(n7922) );
  NAND2_X1 U9247 ( .A1(n8071), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7921) );
  NAND4_X1 U9248 ( .A1(n7924), .A2(n7923), .A3(n7922), .A4(n7921), .ZN(n9552)
         );
  NAND2_X1 U9249 ( .A1(n9765), .A2(n9780), .ZN(n8189) );
  NAND2_X1 U9250 ( .A1(n7925), .A2(n8043), .ZN(n7927) );
  NAND2_X1 U9251 ( .A1(n8046), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7926) );
  NAND2_X1 U9252 ( .A1(n8070), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n7933) );
  NAND2_X1 U9253 ( .A1(n8072), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7932) );
  AOI21_X1 U9254 ( .B1(n7929), .B2(n7937), .A(n7928), .ZN(n9784) );
  NAND2_X1 U9255 ( .A1(n7948), .A2(n9784), .ZN(n7931) );
  NAND2_X1 U9256 ( .A1(n8071), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7930) );
  NAND4_X1 U9257 ( .A1(n7933), .A2(n7932), .A3(n7931), .A4(n7930), .ZN(n9761)
         );
  INV_X1 U9258 ( .A(n9761), .ZN(n9795) );
  OR2_X1 U9259 ( .A1(n10005), .A2(n9795), .ZN(n8209) );
  NAND2_X1 U9260 ( .A1(n10005), .A2(n9795), .ZN(n9756) );
  NAND2_X1 U9261 ( .A1(n7934), .A2(n8043), .ZN(n7936) );
  NAND2_X1 U9262 ( .A1(n8046), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U9263 ( .A1(n8072), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U9264 ( .A1(n8070), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n7941) );
  OAI21_X1 U9265 ( .B1(n7947), .B2(P1_REG3_REG_25__SCAN_IN), .A(n7937), .ZN(
        n7938) );
  INV_X1 U9266 ( .A(n7938), .ZN(n9798) );
  NAND2_X1 U9267 ( .A1(n7948), .A2(n9798), .ZN(n7940) );
  NAND2_X1 U9268 ( .A1(n8071), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7939) );
  NAND4_X1 U9269 ( .A1(n7942), .A2(n7941), .A3(n7940), .A4(n7939), .ZN(n9723)
         );
  NAND2_X1 U9270 ( .A1(n9797), .A2(n9809), .ZN(n8172) );
  NAND2_X1 U9271 ( .A1(n7943), .A2(n8043), .ZN(n7945) );
  NAND2_X1 U9272 ( .A1(n8046), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7944) );
  NAND2_X1 U9273 ( .A1(n8070), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U9274 ( .A1(n8072), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7951) );
  NOR2_X1 U9275 ( .A1(n7957), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n7946) );
  NOR2_X1 U9276 ( .A1(n7947), .A2(n7946), .ZN(n9812) );
  NAND2_X1 U9277 ( .A1(n7948), .A2(n9812), .ZN(n7950) );
  NAND2_X1 U9278 ( .A1(n8071), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7949) );
  NAND4_X1 U9279 ( .A1(n7952), .A2(n7951), .A3(n7950), .A4(n7949), .ZN(n9825)
         );
  NAND2_X1 U9280 ( .A1(n10015), .A2(n9794), .ZN(n8206) );
  NAND2_X1 U9281 ( .A1(n9699), .A2(n8206), .ZN(n9806) );
  INV_X1 U9282 ( .A(n9806), .ZN(n8167) );
  NAND2_X1 U9283 ( .A1(n7953), .A2(n8043), .ZN(n7955) );
  NAND2_X1 U9284 ( .A1(n8046), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7954) );
  NAND2_X1 U9285 ( .A1(n8070), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U9286 ( .A1(n8072), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7960) );
  NOR2_X1 U9287 ( .A1(n7967), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7956) );
  NOR2_X1 U9288 ( .A1(n7957), .A2(n7956), .ZN(n9832) );
  NAND2_X1 U9289 ( .A1(n7948), .A2(n9832), .ZN(n7959) );
  NAND2_X1 U9290 ( .A1(n8071), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7958) );
  NAND4_X1 U9291 ( .A1(n7961), .A2(n7960), .A3(n7959), .A4(n7958), .ZN(n9722)
         );
  OR2_X1 U9292 ( .A1(n9831), .A2(n9847), .ZN(n8164) );
  NAND2_X1 U9293 ( .A1(n9831), .A2(n9847), .ZN(n9805) );
  NAND2_X1 U9294 ( .A1(n8164), .A2(n9805), .ZN(n9820) );
  NAND2_X1 U9295 ( .A1(n7962), .A2(n8043), .ZN(n7964) );
  NAND2_X1 U9296 ( .A1(n8046), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U9297 ( .A1(n8072), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U9298 ( .A1(n8070), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7970) );
  NOR2_X1 U9299 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n7965), .ZN(n7966) );
  NOR2_X1 U9300 ( .A1(n7967), .A2(n7966), .ZN(n9842) );
  NAND2_X1 U9301 ( .A1(n7948), .A2(n9842), .ZN(n7969) );
  NAND2_X1 U9302 ( .A1(n8071), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7968) );
  NAND4_X1 U9303 ( .A1(n7971), .A2(n7970), .A3(n7969), .A4(n7968), .ZN(n9826)
         );
  XNOR2_X1 U9304 ( .A(n10024), .B(n9862), .ZN(n9845) );
  NAND2_X1 U9305 ( .A1(n7972), .A2(n8043), .ZN(n7974) );
  NAND2_X1 U9306 ( .A1(n8046), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U9307 ( .A1(n8072), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7980) );
  NAND2_X1 U9308 ( .A1(n8070), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7979) );
  OAI21_X1 U9309 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n7984), .A(n7975), .ZN(
        n7976) );
  INV_X1 U9310 ( .A(n7976), .ZN(n9865) );
  NAND2_X1 U9311 ( .A1(n8054), .A2(n9865), .ZN(n7978) );
  NAND2_X1 U9312 ( .A1(n8071), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7977) );
  NAND4_X1 U9313 ( .A1(n7980), .A2(n7979), .A3(n7978), .A4(n7977), .ZN(n9876)
         );
  INV_X1 U9314 ( .A(n9876), .ZN(n9848) );
  NAND2_X1 U9315 ( .A1(n10030), .A2(n9848), .ZN(n8197) );
  NAND2_X1 U9316 ( .A1(n8198), .A2(n8197), .ZN(n9858) );
  INV_X1 U9317 ( .A(n9858), .ZN(n9855) );
  NAND2_X1 U9318 ( .A1(n7981), .A2(n8043), .ZN(n7983) );
  NAND2_X1 U9319 ( .A1(n8046), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U9320 ( .A1(n8072), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U9321 ( .A1(n8070), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n7988) );
  AOI21_X1 U9322 ( .B1(n7995), .B2(n7985), .A(n7984), .ZN(n9882) );
  NAND2_X1 U9323 ( .A1(n7948), .A2(n9882), .ZN(n7987) );
  NAND2_X1 U9324 ( .A1(n8071), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7986) );
  NAND4_X1 U9325 ( .A1(n7989), .A2(n7988), .A3(n7987), .A4(n7986), .ZN(n9893)
         );
  INV_X1 U9326 ( .A(n9893), .ZN(n9861) );
  NAND2_X1 U9327 ( .A1(n9881), .A2(n9861), .ZN(n8196) );
  NAND2_X1 U9328 ( .A1(n9857), .A2(n8196), .ZN(n9873) );
  INV_X1 U9329 ( .A(n9873), .ZN(n8061) );
  NAND2_X1 U9330 ( .A1(n7990), .A2(n8043), .ZN(n7992) );
  AOI22_X1 U9331 ( .A1(n8046), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8045), .B2(
        n9671), .ZN(n7991) );
  NAND2_X1 U9332 ( .A1(n8072), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U9333 ( .A1(n8070), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n7998) );
  OR2_X1 U9334 ( .A1(n8049), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7994) );
  AND2_X1 U9335 ( .A1(n7995), .A2(n7994), .ZN(n9898) );
  NAND2_X1 U9336 ( .A1(n7948), .A2(n9898), .ZN(n7997) );
  NAND2_X1 U9337 ( .A1(n8071), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7996) );
  NAND4_X1 U9338 ( .A1(n7999), .A2(n7998), .A3(n7997), .A4(n7996), .ZN(n9910)
         );
  AND2_X1 U9339 ( .A1(n9897), .A2(n9910), .ZN(n9717) );
  INV_X1 U9340 ( .A(n9717), .ZN(n8000) );
  OR2_X1 U9341 ( .A1(n9897), .A2(n9910), .ZN(n9716) );
  NAND2_X1 U9342 ( .A1(n8000), .A2(n9716), .ZN(n9889) );
  NAND2_X1 U9343 ( .A1(n8001), .A2(n8043), .ZN(n8003) );
  AOI22_X1 U9344 ( .A1(n8046), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8045), .B2(
        n9634), .ZN(n8002) );
  NAND2_X1 U9345 ( .A1(n8072), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8010) );
  NAND2_X1 U9346 ( .A1(n8070), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8009) );
  INV_X1 U9347 ( .A(n8004), .ZN(n8051) );
  NAND2_X1 U9348 ( .A1(n8017), .A2(n8005), .ZN(n8006) );
  AND2_X1 U9349 ( .A1(n8051), .A2(n8006), .ZN(n9933) );
  NAND2_X1 U9350 ( .A1(n7948), .A2(n9933), .ZN(n8008) );
  NAND2_X1 U9351 ( .A1(n8071), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8007) );
  NAND4_X1 U9352 ( .A1(n8010), .A2(n8009), .A3(n8008), .A4(n8007), .ZN(n9911)
         );
  NAND2_X1 U9353 ( .A1(n9932), .A2(n9950), .ZN(n8153) );
  NAND2_X1 U9354 ( .A1(n8011), .A2(n8043), .ZN(n8013) );
  AOI22_X1 U9355 ( .A1(n8046), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8045), .B2(
        n9636), .ZN(n8012) );
  NAND2_X1 U9356 ( .A1(n8070), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U9357 ( .A1(n8072), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U9358 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  AND2_X1 U9359 ( .A1(n8017), .A2(n8016), .ZN(n9953) );
  NAND2_X1 U9360 ( .A1(n7948), .A2(n9953), .ZN(n8019) );
  NAND2_X1 U9361 ( .A1(n8071), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8018) );
  NAND4_X1 U9362 ( .A1(n8021), .A2(n8020), .A3(n8019), .A4(n8018), .ZN(n9964)
         );
  OR2_X1 U9363 ( .A1(n9952), .A2(n9712), .ZN(n8264) );
  NAND2_X1 U9364 ( .A1(n9952), .A2(n9712), .ZN(n8259) );
  NAND2_X1 U9365 ( .A1(n8264), .A2(n8259), .ZN(n9940) );
  INV_X1 U9366 ( .A(n9940), .ZN(n9943) );
  NAND2_X1 U9367 ( .A1(n8022), .A2(n8043), .ZN(n8025) );
  AOI22_X1 U9368 ( .A1(n8046), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8045), .B2(
        n8023), .ZN(n8024) );
  NAND2_X1 U9369 ( .A1(n9971), .A2(n9948), .ZN(n8150) );
  NAND2_X1 U9370 ( .A1(n9944), .A2(n8150), .ZN(n9960) );
  INV_X1 U9371 ( .A(n8026), .ZN(n8040) );
  XNOR2_X1 U9372 ( .A(n6799), .B(n10567), .ZN(n10562) );
  NAND4_X1 U9373 ( .A1(n8028), .A2(n8027), .A3(n10562), .A4(n8231), .ZN(n8033)
         );
  NAND4_X1 U9374 ( .A1(n8031), .A2(n8030), .A3(n8238), .A4(n8029), .ZN(n8032)
         );
  NOR2_X1 U9375 ( .A1(n8033), .A2(n8032), .ZN(n8035) );
  NAND4_X1 U9376 ( .A1(n8035), .A2(n8244), .A3(n8034), .A4(n8107), .ZN(n8037)
         );
  NOR2_X1 U9377 ( .A1(n8037), .A2(n8036), .ZN(n8039) );
  NAND4_X1 U9378 ( .A1(n8040), .A2(n8039), .A3(n10755), .A4(n8038), .ZN(n8041)
         );
  NOR3_X1 U9379 ( .A1(n9960), .A2(n8141), .A3(n8041), .ZN(n8042) );
  AND4_X1 U9380 ( .A1(n9889), .A2(n5309), .A3(n9943), .A4(n8042), .ZN(n8060)
         );
  NAND2_X1 U9381 ( .A1(n8044), .A2(n8043), .ZN(n8048) );
  AOI22_X1 U9382 ( .A1(n8046), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8045), .B2(
        n9650), .ZN(n8047) );
  NAND2_X1 U9383 ( .A1(n8070), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U9384 ( .A1(n8071), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8057) );
  INV_X1 U9385 ( .A(n8049), .ZN(n8053) );
  INV_X1 U9386 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8050) );
  NAND2_X1 U9387 ( .A1(n8051), .A2(n8050), .ZN(n8052) );
  AND2_X1 U9388 ( .A1(n8053), .A2(n8052), .ZN(n9918) );
  NAND2_X1 U9389 ( .A1(n8054), .A2(n9918), .ZN(n8056) );
  NAND2_X1 U9390 ( .A1(n8072), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8055) );
  NAND4_X1 U9391 ( .A1(n8058), .A2(n8057), .A3(n8056), .A4(n8055), .ZN(n9927)
         );
  XNOR2_X1 U9392 ( .A(n9917), .B(n9714), .ZN(n9905) );
  INV_X1 U9393 ( .A(n9905), .ZN(n8059) );
  NAND4_X1 U9394 ( .A1(n9855), .A2(n8061), .A3(n8060), .A4(n8059), .ZN(n8062)
         );
  NOR3_X1 U9395 ( .A1(n9820), .A2(n9845), .A3(n8062), .ZN(n8063) );
  NAND3_X1 U9396 ( .A1(n9791), .A2(n8167), .A3(n8063), .ZN(n8064) );
  NOR2_X1 U9397 ( .A1(n9778), .A2(n8064), .ZN(n8065) );
  NAND4_X1 U9398 ( .A1(n9729), .A2(n9744), .A3(n9754), .A4(n8065), .ZN(n8078)
         );
  NAND2_X1 U9399 ( .A1(n8306), .A2(n8043), .ZN(n8069) );
  OR2_X1 U9400 ( .A1(n6943), .A2(n8303), .ZN(n8068) );
  NAND2_X1 U9401 ( .A1(n8070), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8075) );
  NAND2_X1 U9402 ( .A1(n8071), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U9403 ( .A1(n8072), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8073) );
  AND3_X1 U9404 ( .A1(n8075), .A2(n8074), .A3(n8073), .ZN(n9705) );
  NAND2_X1 U9405 ( .A1(n8076), .A2(n9705), .ZN(n8284) );
  NAND2_X1 U9406 ( .A1(n8288), .A2(n8284), .ZN(n8077) );
  NOR4_X1 U9407 ( .A1(n8285), .A2(n8289), .A3(n8078), .A4(n8077), .ZN(n8188)
         );
  OR2_X1 U9408 ( .A1(n6613), .A2(n9674), .ZN(n8174) );
  INV_X1 U9409 ( .A(n8174), .ZN(n8181) );
  MUX2_X1 U9410 ( .A(n8281), .B(n8213), .S(n8174), .Z(n8178) );
  MUX2_X1 U9411 ( .A(n9703), .B(n8212), .S(n8181), .Z(n8177) );
  NAND2_X1 U9412 ( .A1(n9563), .A2(n8079), .ZN(n8080) );
  NAND2_X1 U9413 ( .A1(n8081), .A2(n8080), .ZN(n8093) );
  NAND2_X1 U9414 ( .A1(n8092), .A2(n8093), .ZN(n8082) );
  NAND3_X1 U9415 ( .A1(n8082), .A2(n8088), .A3(n8232), .ZN(n8084) );
  AND2_X1 U9416 ( .A1(n8087), .A2(n8083), .ZN(n8086) );
  NAND2_X1 U9417 ( .A1(n8084), .A2(n8086), .ZN(n8095) );
  INV_X1 U9418 ( .A(n8091), .ZN(n8236) );
  INV_X1 U9419 ( .A(n8087), .ZN(n8089) );
  OAI21_X1 U9420 ( .B1(n8089), .B2(n8088), .A(n8096), .ZN(n8090) );
  AOI21_X1 U9421 ( .B1(n8092), .B2(n8091), .A(n8090), .ZN(n8235) );
  OAI21_X1 U9422 ( .B1(n8093), .B2(n8236), .A(n8235), .ZN(n8094) );
  OAI21_X1 U9423 ( .B1(n8098), .B2(n8096), .A(n8239), .ZN(n8097) );
  MUX2_X1 U9424 ( .A(n8098), .B(n8097), .S(n8174), .Z(n8100) );
  NOR2_X1 U9425 ( .A1(n8100), .A2(n8099), .ZN(n8101) );
  MUX2_X1 U9426 ( .A(n8238), .B(n8104), .S(n8174), .Z(n8109) );
  NAND3_X1 U9427 ( .A1(n8119), .A2(n8107), .A3(n8106), .ZN(n8108) );
  NAND2_X1 U9428 ( .A1(n8108), .A2(n8181), .ZN(n8123) );
  AND4_X1 U9429 ( .A1(n8109), .A2(n5497), .A3(n8116), .A4(n8123), .ZN(n8110)
         );
  NAND2_X1 U9430 ( .A1(n8111), .A2(n8110), .ZN(n8127) );
  NAND2_X1 U9431 ( .A1(n8112), .A2(n8174), .ZN(n8115) );
  NAND2_X1 U9432 ( .A1(n8113), .A2(n8181), .ZN(n8114) );
  NAND2_X1 U9433 ( .A1(n8115), .A2(n8114), .ZN(n8117) );
  AOI21_X1 U9434 ( .B1(n8118), .B2(n8117), .A(n8120), .ZN(n8124) );
  NAND3_X1 U9435 ( .A1(n8120), .A2(n8181), .A3(n8119), .ZN(n8121) );
  NAND2_X1 U9436 ( .A1(n8121), .A2(n8130), .ZN(n8122) );
  NAND2_X1 U9437 ( .A1(n8125), .A2(n8250), .ZN(n8126) );
  NAND2_X1 U9438 ( .A1(n8248), .A2(n8126), .ZN(n8129) );
  AND2_X1 U9439 ( .A1(n8136), .A2(n8128), .ZN(n8134) );
  INV_X1 U9440 ( .A(n8129), .ZN(n8131) );
  NAND2_X1 U9441 ( .A1(n8139), .A2(n8130), .ZN(n8253) );
  AOI21_X1 U9442 ( .B1(n8132), .B2(n8131), .A(n8253), .ZN(n8133) );
  MUX2_X1 U9443 ( .A(n8134), .B(n8133), .S(n8174), .Z(n8135) );
  AND2_X1 U9444 ( .A1(n8142), .A2(n8136), .ZN(n8252) );
  OR2_X1 U9445 ( .A1(n9708), .A2(n9707), .ZN(n9959) );
  NAND2_X1 U9446 ( .A1(n9959), .A2(n8138), .ZN(n8255) );
  AOI21_X1 U9447 ( .B1(n8140), .B2(n8252), .A(n8255), .ZN(n8137) );
  AND2_X1 U9448 ( .A1(n9708), .A2(n9707), .ZN(n8144) );
  OAI211_X1 U9449 ( .C1(n8137), .C2(n8144), .A(n9944), .B(n8174), .ZN(n8148)
         );
  AOI21_X1 U9450 ( .B1(n8143), .B2(n8142), .A(n8141), .ZN(n8146) );
  INV_X1 U9451 ( .A(n8144), .ZN(n8145) );
  NAND2_X1 U9452 ( .A1(n8150), .A2(n8145), .ZN(n8256) );
  NAND2_X1 U9453 ( .A1(n8264), .A2(n9944), .ZN(n8149) );
  NAND2_X1 U9454 ( .A1(n8259), .A2(n8150), .ZN(n8151) );
  NAND2_X1 U9455 ( .A1(n8152), .A2(n5309), .ZN(n8155) );
  INV_X1 U9456 ( .A(n8155), .ZN(n8154) );
  NAND2_X1 U9457 ( .A1(n9917), .A2(n9714), .ZN(n8156) );
  NAND2_X1 U9458 ( .A1(n8156), .A2(n8153), .ZN(n8193) );
  OR2_X1 U9459 ( .A1(n9917), .A2(n9714), .ZN(n8262) );
  INV_X1 U9460 ( .A(n9910), .ZN(n9521) );
  NAND2_X1 U9461 ( .A1(n9897), .A2(n9521), .ZN(n8267) );
  NAND3_X1 U9462 ( .A1(n8155), .A2(n8263), .A3(n8262), .ZN(n8157) );
  NAND3_X1 U9463 ( .A1(n8157), .A2(n8267), .A3(n8156), .ZN(n8158) );
  OR2_X1 U9464 ( .A1(n9897), .A2(n9521), .ZN(n9872) );
  AND2_X1 U9465 ( .A1(n9857), .A2(n9872), .ZN(n8194) );
  AOI21_X1 U9466 ( .B1(n8158), .B2(n8194), .A(n5202), .ZN(n8159) );
  OAI21_X1 U9467 ( .B1(n8174), .B2(n8198), .A(n8160), .ZN(n8163) );
  NAND2_X1 U9468 ( .A1(n10024), .A2(n9862), .ZN(n8161) );
  AND2_X1 U9469 ( .A1(n9805), .A2(n8161), .ZN(n8195) );
  OAI21_X1 U9470 ( .B1(n9845), .B2(n8197), .A(n8195), .ZN(n8162) );
  AOI22_X1 U9471 ( .A1(n8163), .A2(n5506), .B1(n8174), .B2(n8162), .ZN(n8166)
         );
  INV_X1 U9472 ( .A(n8164), .ZN(n8165) );
  NOR2_X1 U9473 ( .A1(n10024), .A2(n9862), .ZN(n9695) );
  INV_X1 U9474 ( .A(n9695), .ZN(n9819) );
  AND2_X1 U9475 ( .A1(n9819), .A2(n8164), .ZN(n8203) );
  OAI22_X1 U9476 ( .A1(n8166), .A2(n8165), .B1(n8203), .B2(n8174), .ZN(n8168)
         );
  OAI211_X1 U9477 ( .C1(n9805), .C2(n8174), .A(n8168), .B(n8167), .ZN(n8170)
         );
  NAND2_X1 U9478 ( .A1(n8172), .A2(n8206), .ZN(n8169) );
  INV_X1 U9479 ( .A(n9773), .ZN(n9700) );
  AOI21_X1 U9480 ( .B1(n9791), .B2(n9699), .A(n8174), .ZN(n8171) );
  NAND2_X1 U9481 ( .A1(n9756), .A2(n8172), .ZN(n8273) );
  OAI211_X1 U9482 ( .C1(n8209), .C2(n8174), .A(n8173), .B(n9754), .ZN(n8176)
         );
  MUX2_X1 U9483 ( .A(n8189), .B(n9745), .S(n8174), .Z(n8175) );
  INV_X1 U9484 ( .A(n9705), .ZN(n9551) );
  INV_X1 U9485 ( .A(n9686), .ZN(n9550) );
  NAND2_X1 U9486 ( .A1(n9551), .A2(n9550), .ZN(n8179) );
  NAND2_X1 U9487 ( .A1(n8076), .A2(n8179), .ZN(n8219) );
  NAND2_X1 U9488 ( .A1(n8180), .A2(n8222), .ZN(n8184) );
  NAND2_X1 U9489 ( .A1(n8222), .A2(n8217), .ZN(n8182) );
  NAND2_X1 U9490 ( .A1(n8182), .A2(n8181), .ZN(n8183) );
  AOI211_X1 U9491 ( .C1(n8186), .C2(n8185), .A(n8188), .B(n8187), .ZN(n8229)
         );
  INV_X1 U9492 ( .A(n8188), .ZN(n8226) );
  AND2_X1 U9493 ( .A1(n9703), .A2(n8189), .ZN(n8277) );
  INV_X1 U9494 ( .A(n9960), .ZN(n8190) );
  NAND2_X1 U9495 ( .A1(n8191), .A2(n8190), .ZN(n9963) );
  INV_X1 U9496 ( .A(n9944), .ZN(n8260) );
  NOR2_X1 U9497 ( .A1(n9940), .A2(n8260), .ZN(n8192) );
  NAND2_X1 U9498 ( .A1(n9963), .A2(n8192), .ZN(n9942) );
  NAND2_X1 U9499 ( .A1(n9942), .A2(n8259), .ZN(n9925) );
  NAND2_X1 U9500 ( .A1(n8193), .A2(n8262), .ZN(n8266) );
  NAND2_X1 U9501 ( .A1(n9891), .A2(n8267), .ZN(n9874) );
  AND2_X1 U9502 ( .A1(n8194), .A2(n8198), .ZN(n8272) );
  NAND2_X1 U9503 ( .A1(n9874), .A2(n8272), .ZN(n9694) );
  INV_X1 U9504 ( .A(n8195), .ZN(n8201) );
  NAND2_X1 U9505 ( .A1(n8197), .A2(n8196), .ZN(n8199) );
  NAND2_X1 U9506 ( .A1(n8199), .A2(n8198), .ZN(n9693) );
  INV_X1 U9507 ( .A(n9693), .ZN(n8200) );
  NOR2_X1 U9508 ( .A1(n8201), .A2(n8200), .ZN(n8202) );
  AND2_X1 U9509 ( .A1(n8206), .A2(n8202), .ZN(n8269) );
  INV_X1 U9510 ( .A(n8203), .ZN(n8204) );
  NAND2_X1 U9511 ( .A1(n8204), .A2(n9805), .ZN(n8205) );
  NAND2_X1 U9512 ( .A1(n9699), .A2(n8205), .ZN(n8207) );
  NAND2_X1 U9513 ( .A1(n8207), .A2(n8206), .ZN(n8208) );
  NAND2_X1 U9514 ( .A1(n9773), .A2(n8208), .ZN(n8275) );
  AOI21_X1 U9515 ( .B1(n9694), .B2(n8269), .A(n8275), .ZN(n8211) );
  INV_X1 U9516 ( .A(n9745), .ZN(n8210) );
  NOR2_X1 U9517 ( .A1(n8210), .A2(n5179), .ZN(n8280) );
  OAI21_X1 U9518 ( .B1(n8211), .B2(n8273), .A(n8280), .ZN(n8214) );
  NAND2_X1 U9519 ( .A1(n8213), .A2(n8212), .ZN(n8283) );
  AOI21_X1 U9520 ( .B1(n8277), .B2(n8214), .A(n8283), .ZN(n8216) );
  INV_X1 U9521 ( .A(n8281), .ZN(n8215) );
  NOR2_X1 U9522 ( .A1(n8216), .A2(n8215), .ZN(n8221) );
  INV_X1 U9523 ( .A(n8217), .ZN(n8220) );
  OAI211_X1 U9524 ( .C1(n8221), .C2(n8220), .A(n8219), .B(n8218), .ZN(n8224)
         );
  NAND3_X1 U9525 ( .A1(n8224), .A2(n8223), .A3(n8222), .ZN(n8225) );
  AOI21_X1 U9526 ( .B1(n8226), .B2(n8225), .A(n9671), .ZN(n8228) );
  NOR2_X1 U9527 ( .A1(n10552), .A2(n6726), .ZN(n8230) );
  AOI211_X1 U9528 ( .C1(n10554), .C2(n6799), .A(n8231), .B(n8230), .ZN(n8234)
         );
  INV_X1 U9529 ( .A(n8232), .ZN(n8233) );
  NOR2_X1 U9530 ( .A1(n8234), .A2(n8233), .ZN(n8237) );
  OAI21_X1 U9531 ( .B1(n8237), .B2(n8236), .A(n8235), .ZN(n8243) );
  INV_X1 U9532 ( .A(n8238), .ZN(n8241) );
  INV_X1 U9533 ( .A(n8239), .ZN(n8240) );
  AOI211_X1 U9534 ( .C1(n8243), .C2(n8242), .A(n8241), .B(n8240), .ZN(n8247)
         );
  INV_X1 U9535 ( .A(n8244), .ZN(n8246) );
  OAI21_X1 U9536 ( .B1(n8247), .B2(n8246), .A(n8245), .ZN(n8251) );
  INV_X1 U9537 ( .A(n8248), .ZN(n8249) );
  AOI21_X1 U9538 ( .B1(n8251), .B2(n8250), .A(n8249), .ZN(n8254) );
  OAI21_X1 U9539 ( .B1(n8254), .B2(n8253), .A(n8252), .ZN(n8258) );
  INV_X1 U9540 ( .A(n8255), .ZN(n8257) );
  AOI21_X1 U9541 ( .B1(n8258), .B2(n8257), .A(n8256), .ZN(n8261) );
  OAI21_X1 U9542 ( .B1(n8261), .B2(n8260), .A(n8259), .ZN(n8265) );
  NAND4_X1 U9543 ( .A1(n8265), .A2(n8264), .A3(n8263), .A4(n8262), .ZN(n8268)
         );
  NAND3_X1 U9544 ( .A1(n8268), .A2(n8267), .A3(n8266), .ZN(n8271) );
  INV_X1 U9545 ( .A(n8269), .ZN(n8270) );
  AOI21_X1 U9546 ( .B1(n8272), .B2(n8271), .A(n8270), .ZN(n8276) );
  INV_X1 U9547 ( .A(n8273), .ZN(n8274) );
  OAI21_X1 U9548 ( .B1(n8276), .B2(n8275), .A(n8274), .ZN(n8279) );
  INV_X1 U9549 ( .A(n8277), .ZN(n8278) );
  AOI21_X1 U9550 ( .B1(n8280), .B2(n8279), .A(n8278), .ZN(n8282) );
  OAI21_X1 U9551 ( .B1(n8283), .B2(n8282), .A(n8281), .ZN(n8287) );
  INV_X1 U9552 ( .A(n8284), .ZN(n8286) );
  AOI211_X1 U9553 ( .C1(n8288), .C2(n8287), .A(n8286), .B(n8285), .ZN(n8290)
         );
  NOR2_X1 U9554 ( .A1(n8290), .A2(n8289), .ZN(n8294) );
  NAND2_X1 U9555 ( .A1(n8294), .A2(n10553), .ZN(n8292) );
  OAI211_X1 U9556 ( .C1(n8294), .C2(n8293), .A(n8292), .B(n8291), .ZN(n8300)
         );
  NOR2_X1 U9557 ( .A1(n8296), .A2(n8295), .ZN(n8299) );
  OAI21_X1 U9558 ( .B1(n8297), .B2(n6613), .A(P1_B_REG_SCAN_IN), .ZN(n8298) );
  OAI22_X1 U9559 ( .A1(n8301), .A2(n8300), .B1(n8299), .B2(n8298), .ZN(
        P1_U3242) );
  INV_X1 U9560 ( .A(n8306), .ZN(n9151) );
  OAI222_X1 U9561 ( .A1(n10132), .A2(n8303), .B1(n10138), .B2(n9151), .C1(
        n8302), .C2(P1_U3086), .ZN(P1_U3325) );
  NAND2_X1 U9562 ( .A1(n9145), .A2(n6113), .ZN(n8305) );
  NAND2_X1 U9563 ( .A1(n8307), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8304) );
  INV_X1 U9564 ( .A(n9094), .ZN(n8327) );
  NAND2_X1 U9565 ( .A1(n8306), .A2(n6113), .ZN(n8309) );
  NAND2_X1 U9566 ( .A1(n8307), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8308) );
  INV_X1 U9567 ( .A(n8690), .ZN(n8324) );
  NOR2_X1 U9568 ( .A1(n8828), .A2(n8324), .ZN(n8502) );
  INV_X1 U9569 ( .A(n8502), .ZN(n8353) );
  NAND2_X1 U9570 ( .A1(n8310), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8317) );
  INV_X1 U9571 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8311) );
  OR2_X1 U9572 ( .A1(n8312), .A2(n8311), .ZN(n8316) );
  INV_X1 U9573 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8313) );
  OR2_X1 U9574 ( .A1(n8314), .A2(n8313), .ZN(n8315) );
  NAND4_X1 U9575 ( .A1(n8318), .A2(n8317), .A3(n8316), .A4(n8315), .ZN(n8826)
         );
  NAND2_X1 U9576 ( .A1(n8353), .A2(n8826), .ZN(n8326) );
  INV_X1 U9577 ( .A(n8826), .ZN(n8319) );
  NOR2_X1 U9578 ( .A1(n8327), .A2(n8319), .ZN(n8510) );
  INV_X1 U9579 ( .A(n8320), .ZN(n8321) );
  NAND2_X1 U9580 ( .A1(n8828), .A2(n8324), .ZN(n8508) );
  NOR2_X1 U9581 ( .A1(n9094), .A2(n8826), .ZN(n8507) );
  AND2_X2 U9582 ( .A1(n8491), .A2(n8490), .ZN(n8857) );
  INV_X1 U9583 ( .A(n8857), .ZN(n8351) );
  INV_X1 U9584 ( .A(n8869), .ZN(n8350) );
  NAND2_X1 U9585 ( .A1(n8477), .A2(n8476), .ZN(n8903) );
  NAND3_X1 U9586 ( .A1(n10587), .A2(n8329), .A3(n8377), .ZN(n8330) );
  NOR4_X1 U9587 ( .A1(n8330), .A2(n10632), .A3(n9025), .A4(n6138), .ZN(n8332)
         );
  NAND3_X1 U9588 ( .A1(n8332), .A2(n8403), .A3(n8331), .ZN(n8336) );
  NOR4_X1 U9589 ( .A1(n8336), .A2(n8335), .A3(n8334), .A4(n8333), .ZN(n8338)
         );
  NAND4_X1 U9590 ( .A1(n8340), .A2(n8339), .A3(n8338), .A4(n8337), .ZN(n8343)
         );
  NOR4_X1 U9591 ( .A1(n8998), .A2(n8343), .A3(n8342), .A4(n8341), .ZN(n8345)
         );
  NAND4_X1 U9592 ( .A1(n8966), .A2(n8978), .A3(n8345), .A4(n8344), .ZN(n8346)
         );
  NOR4_X1 U9593 ( .A1(n8903), .A2(n5476), .A3(n8924), .A4(n8346), .ZN(n8348)
         );
  XNOR2_X1 U9594 ( .A(n8347), .B(n8927), .ZN(n8914) );
  NAND2_X1 U9595 ( .A1(n8483), .A2(n8479), .ZN(n8894) );
  NAND4_X1 U9596 ( .A1(n5005), .A2(n8348), .A3(n8914), .A4(n8894), .ZN(n8349)
         );
  NAND4_X1 U9597 ( .A1(n6128), .A2(n8353), .A3(n8352), .A4(n8508), .ZN(n8354)
         );
  NOR3_X1 U9598 ( .A1(n8507), .A2(n8510), .A3(n8354), .ZN(n8355) );
  INV_X1 U9599 ( .A(n8512), .ZN(n8513) );
  MUX2_X1 U9600 ( .A(n8691), .B(n8839), .S(n8506), .Z(n8497) );
  MUX2_X1 U9601 ( .A(n8694), .B(n8891), .S(n8500), .Z(n8478) );
  INV_X1 U9602 ( .A(n8478), .ZN(n8484) );
  INV_X1 U9603 ( .A(n8356), .ZN(n10800) );
  AOI21_X1 U9604 ( .B1(n9002), .B2(n8681), .A(n8506), .ZN(n8443) );
  OAI211_X1 U9605 ( .C1(n9002), .C2(n8357), .A(n8356), .B(n8506), .ZN(n8360)
         );
  NAND3_X1 U9606 ( .A1(n8698), .A2(n8699), .A3(n8500), .ZN(n8359) );
  NAND3_X1 U9607 ( .A1(n8357), .A2(n9002), .A3(n8506), .ZN(n8358) );
  NAND3_X1 U9608 ( .A1(n8360), .A2(n8359), .A3(n8358), .ZN(n8442) );
  NAND2_X1 U9609 ( .A1(n10800), .A2(n9002), .ZN(n8439) );
  MUX2_X1 U9610 ( .A(n8506), .B(n8361), .S(n8700), .Z(n8437) );
  NOR2_X1 U9611 ( .A1(n8361), .A2(n8506), .ZN(n8436) );
  NAND3_X1 U9612 ( .A1(n8363), .A2(n8365), .A3(n8362), .ZN(n8364) );
  NAND2_X1 U9613 ( .A1(n8364), .A2(n8506), .ZN(n8370) );
  INV_X1 U9614 ( .A(n8365), .ZN(n8366) );
  AOI21_X1 U9615 ( .B1(n8368), .B2(n8367), .A(n8366), .ZN(n8369) );
  MUX2_X1 U9616 ( .A(n8370), .B(n8506), .S(n8369), .Z(n8372) );
  NOR2_X1 U9617 ( .A1(n8372), .A2(n8371), .ZN(n8379) );
  NAND2_X1 U9618 ( .A1(n8388), .A2(n8373), .ZN(n8376) );
  NAND2_X1 U9619 ( .A1(n8382), .A2(n8374), .ZN(n8375) );
  MUX2_X1 U9620 ( .A(n8376), .B(n8375), .S(n8500), .Z(n8378) );
  INV_X1 U9621 ( .A(n8390), .ZN(n8383) );
  AOI211_X1 U9622 ( .C1(n8383), .C2(n8382), .A(n8381), .B(n8380), .ZN(n8387)
         );
  NAND2_X1 U9623 ( .A1(n8393), .A2(n8384), .ZN(n8386) );
  OAI21_X1 U9624 ( .B1(n8387), .B2(n8386), .A(n8385), .ZN(n8397) );
  INV_X1 U9625 ( .A(n8388), .ZN(n8389) );
  NOR2_X1 U9626 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  AOI211_X1 U9627 ( .C1(n10612), .C2(n10636), .A(n8392), .B(n8391), .ZN(n8395)
         );
  OAI21_X1 U9628 ( .B1(n8395), .B2(n8394), .A(n8393), .ZN(n8396) );
  MUX2_X1 U9629 ( .A(n8397), .B(n8396), .S(n8500), .Z(n8412) );
  NAND2_X1 U9630 ( .A1(n8406), .A2(n8404), .ZN(n8400) );
  INV_X1 U9631 ( .A(n8398), .ZN(n8399) );
  MUX2_X1 U9632 ( .A(n8400), .B(n8399), .S(n8500), .Z(n8402) );
  INV_X1 U9633 ( .A(n8417), .ZN(n8401) );
  NOR2_X1 U9634 ( .A1(n8402), .A2(n8401), .ZN(n8415) );
  NAND2_X1 U9635 ( .A1(n8415), .A2(n8403), .ZN(n8411) );
  NAND2_X1 U9636 ( .A1(n8405), .A2(n8404), .ZN(n8409) );
  INV_X1 U9637 ( .A(n8420), .ZN(n8408) );
  INV_X1 U9638 ( .A(n8406), .ZN(n8407) );
  INV_X1 U9639 ( .A(n8413), .ZN(n8416) );
  NAND3_X1 U9640 ( .A1(n8422), .A2(n8425), .A3(n8416), .ZN(n8414) );
  NAND2_X1 U9641 ( .A1(n8414), .A2(n8423), .ZN(n8428) );
  INV_X1 U9642 ( .A(n8415), .ZN(n8419) );
  OAI211_X1 U9643 ( .C1(n8419), .C2(n8418), .A(n8417), .B(n8416), .ZN(n8421)
         );
  OAI21_X1 U9644 ( .B1(n8422), .B2(n8421), .A(n8420), .ZN(n8426) );
  INV_X1 U9645 ( .A(n8423), .ZN(n8424) );
  AOI21_X1 U9646 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8427) );
  MUX2_X1 U9647 ( .A(n8430), .B(n8429), .S(n8500), .Z(n8431) );
  OAI21_X1 U9648 ( .B1(n8437), .B2(n8436), .A(n8435), .ZN(n8446) );
  AOI211_X1 U9649 ( .C1(n8440), .C2(n8439), .A(n8438), .B(n8446), .ZN(n8441)
         );
  NAND3_X1 U9650 ( .A1(n8446), .A2(n5428), .A3(n8445), .ZN(n8447) );
  INV_X1 U9651 ( .A(n8998), .ZN(n9008) );
  NAND2_X1 U9652 ( .A1(n8447), .A2(n9008), .ZN(n8451) );
  MUX2_X1 U9653 ( .A(n8449), .B(n8448), .S(n8500), .Z(n8450) );
  MUX2_X1 U9654 ( .A(n8696), .B(n8599), .S(n8506), .Z(n8455) );
  INV_X1 U9655 ( .A(n8599), .ZN(n9139) );
  NAND2_X1 U9656 ( .A1(n8456), .A2(n9139), .ZN(n8454) );
  NAND2_X1 U9657 ( .A1(n8964), .A2(n9004), .ZN(n8453) );
  MUX2_X1 U9658 ( .A(n8456), .B(n8964), .S(n8500), .Z(n8457) );
  INV_X1 U9659 ( .A(n8459), .ZN(n8461) );
  MUX2_X1 U9660 ( .A(n8461), .B(n8460), .S(n8500), .Z(n8462) );
  INV_X1 U9661 ( .A(n8924), .ZN(n8922) );
  NAND2_X1 U9662 ( .A1(n8950), .A2(n8554), .ZN(n8463) );
  MUX2_X1 U9663 ( .A(n8464), .B(n8463), .S(n8506), .Z(n8465) );
  OAI211_X1 U9664 ( .C1(n8466), .C2(n5476), .A(n8922), .B(n8465), .ZN(n8470)
         );
  MUX2_X1 U9665 ( .A(n8468), .B(n8467), .S(n8506), .Z(n8469) );
  NAND3_X1 U9666 ( .A1(n8470), .A2(n8914), .A3(n8469), .ZN(n8474) );
  MUX2_X1 U9667 ( .A(n8472), .B(n8471), .S(n8500), .Z(n8473) );
  AOI21_X1 U9668 ( .B1(n8474), .B2(n8473), .A(n8903), .ZN(n8475) );
  INV_X1 U9669 ( .A(n8475), .ZN(n8481) );
  MUX2_X1 U9670 ( .A(n8477), .B(n8476), .S(n8506), .Z(n8480) );
  AOI22_X1 U9671 ( .A1(n8481), .A2(n8480), .B1(n8479), .B2(n8478), .ZN(n8482)
         );
  MUX2_X1 U9672 ( .A(n8486), .B(n8485), .S(n8506), .Z(n8487) );
  MUX2_X1 U9673 ( .A(n8488), .B(n8855), .S(n8500), .Z(n8489) );
  MUX2_X1 U9674 ( .A(n8491), .B(n8490), .S(n8506), .Z(n8492) );
  INV_X1 U9675 ( .A(n8497), .ZN(n8494) );
  MUX2_X1 U9676 ( .A(n8691), .B(n8839), .S(n8500), .Z(n8493) );
  INV_X1 U9677 ( .A(n8498), .ZN(n8501) );
  OAI21_X1 U9678 ( .B1(n8501), .B2(n8500), .A(n8499), .ZN(n8503) );
  OAI21_X1 U9679 ( .B1(n8506), .B2(n8505), .A(n8504), .ZN(n8509) );
  AOI21_X1 U9680 ( .B1(n8509), .B2(n8508), .A(n8507), .ZN(n8511) );
  NAND3_X1 U9681 ( .A1(n8518), .A2(n8517), .A3(n8516), .ZN(n8519) );
  OAI211_X1 U9682 ( .C1(n8520), .C2(n8522), .A(n8519), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8521) );
  OAI21_X1 U9683 ( .B1(n8523), .B2(n8522), .A(n8521), .ZN(P2_U3296) );
  XNOR2_X1 U9684 ( .A(n8525), .B(n8524), .ZN(n8530) );
  AOI22_X1 U9685 ( .A1(n8691), .A2(n8686), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8527) );
  NAND2_X1 U9686 ( .A1(n8663), .A2(n8692), .ZN(n8526) );
  OAI211_X1 U9687 ( .C1(n8860), .C2(n8683), .A(n8527), .B(n8526), .ZN(n8528)
         );
  AOI21_X1 U9688 ( .B1(n8859), .B2(n8673), .A(n8528), .ZN(n8529) );
  OAI21_X1 U9689 ( .B1(n8530), .B2(n8676), .A(n8529), .ZN(P2_U3154) );
  INV_X1 U9690 ( .A(n8531), .ZN(n8626) );
  INV_X1 U9691 ( .A(n8532), .ZN(n8534) );
  NOR3_X1 U9692 ( .A1(n8626), .A2(n8534), .A3(n8533), .ZN(n8537) );
  INV_X1 U9693 ( .A(n8535), .ZN(n8536) );
  OAI21_X1 U9694 ( .B1(n8537), .B2(n8536), .A(n8624), .ZN(n8542) );
  NAND2_X1 U9695 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n8748) );
  OAI21_X1 U9696 ( .B1(n8566), .B2(n8680), .A(n8748), .ZN(n8540) );
  NOR2_X1 U9697 ( .A1(n8683), .A2(n8538), .ZN(n8539) );
  AOI211_X1 U9698 ( .C1(n8686), .C2(n8698), .A(n8540), .B(n8539), .ZN(n8541)
         );
  OAI211_X1 U9699 ( .C1(n10793), .C2(n8689), .A(n8542), .B(n8541), .ZN(
        P2_U3155) );
  XNOR2_X1 U9700 ( .A(n8543), .B(n8912), .ZN(n8548) );
  AOI22_X1 U9701 ( .A1(n8694), .A2(n8686), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8545) );
  NAND2_X1 U9702 ( .A1(n8663), .A2(n8927), .ZN(n8544) );
  OAI211_X1 U9703 ( .C1(n8683), .C2(n8905), .A(n8545), .B(n8544), .ZN(n8546)
         );
  AOI21_X1 U9704 ( .B1(n8904), .B2(n8673), .A(n8546), .ZN(n8547) );
  OAI21_X1 U9705 ( .B1(n8548), .B2(n8676), .A(n8547), .ZN(P2_U3156) );
  INV_X1 U9706 ( .A(n8972), .ZN(n9131) );
  NAND2_X1 U9707 ( .A1(n8658), .A2(n8549), .ZN(n8552) );
  NAND2_X1 U9708 ( .A1(n8552), .A2(n8551), .ZN(n8550) );
  OAI211_X1 U9709 ( .C1(n8552), .C2(n8551), .A(n8550), .B(n8624), .ZN(n8558)
         );
  OAI21_X1 U9710 ( .B1(n8554), .B2(n8660), .A(n8553), .ZN(n8556) );
  NOR2_X1 U9711 ( .A1(n8683), .A2(n8962), .ZN(n8555) );
  AOI211_X1 U9712 ( .C1(n8663), .C2(n8958), .A(n8556), .B(n8555), .ZN(n8557)
         );
  OAI211_X1 U9713 ( .C1(n9131), .C2(n8689), .A(n8558), .B(n8557), .ZN(P2_U3159) );
  XOR2_X1 U9714 ( .A(n8560), .B(n8559), .Z(n8565) );
  AOI22_X1 U9715 ( .A1(n8927), .A2(n8686), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8562) );
  NAND2_X1 U9716 ( .A1(n8663), .A2(n8959), .ZN(n8561) );
  OAI211_X1 U9717 ( .C1(n8683), .C2(n8930), .A(n8562), .B(n8561), .ZN(n8563)
         );
  AOI21_X1 U9718 ( .B1(n9062), .B2(n8673), .A(n8563), .ZN(n8564) );
  OAI21_X1 U9719 ( .B1(n8565), .B2(n8676), .A(n8564), .ZN(P2_U3163) );
  INV_X1 U9720 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10341) );
  NOR2_X1 U9721 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10341), .ZN(n8716) );
  NOR2_X1 U9722 ( .A1(n8566), .A2(n8660), .ZN(n8567) );
  AOI211_X1 U9723 ( .C1(n8663), .C2(n8702), .A(n8716), .B(n8567), .ZN(n8568)
         );
  OAI21_X1 U9724 ( .B1(n8569), .B2(n8683), .A(n8568), .ZN(n8574) );
  INV_X1 U9725 ( .A(n8623), .ZN(n8570) );
  AOI211_X1 U9726 ( .C1(n8572), .C2(n8571), .A(n8676), .B(n8570), .ZN(n8573)
         );
  AOI211_X1 U9727 ( .C1(n8575), .C2(n8673), .A(n8574), .B(n8573), .ZN(n8576)
         );
  INV_X1 U9728 ( .A(n8576), .ZN(P2_U3164) );
  XOR2_X1 U9729 ( .A(n8578), .B(n8577), .Z(n8583) );
  AOI22_X1 U9730 ( .A1(n8692), .A2(n8686), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8580) );
  NAND2_X1 U9731 ( .A1(n8663), .A2(n8694), .ZN(n8579) );
  OAI211_X1 U9732 ( .C1(n8683), .C2(n8883), .A(n8580), .B(n8579), .ZN(n8581)
         );
  AOI21_X1 U9733 ( .B1(n9045), .B2(n8673), .A(n8581), .ZN(n8582) );
  OAI21_X1 U9734 ( .B1(n8583), .B2(n8676), .A(n8582), .ZN(P2_U3165) );
  NAND2_X1 U9735 ( .A1(n5556), .A2(n8584), .ZN(n8592) );
  XNOR2_X1 U9736 ( .A(n8590), .B(n8988), .ZN(n8591) );
  XNOR2_X1 U9737 ( .A(n8592), .B(n8591), .ZN(n8589) );
  OR2_X1 U9738 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10340), .ZN(n8782) );
  OAI21_X1 U9739 ( .B1(n9004), .B2(n8660), .A(n8782), .ZN(n8585) );
  AOI21_X1 U9740 ( .B1(n8663), .B2(n8698), .A(n8585), .ZN(n8586) );
  OAI21_X1 U9741 ( .B1(n9011), .B2(n8683), .A(n8586), .ZN(n8587) );
  AOI21_X1 U9742 ( .B1(n9010), .B2(n8673), .A(n8587), .ZN(n8588) );
  OAI21_X1 U9743 ( .B1(n8589), .B2(n8676), .A(n8588), .ZN(P2_U3166) );
  AOI22_X1 U9744 ( .A1(n8592), .A2(n8591), .B1(n8590), .B2(n8697), .ZN(n8595)
         );
  XNOR2_X1 U9745 ( .A(n8593), .B(n8696), .ZN(n8594) );
  XNOR2_X1 U9746 ( .A(n8595), .B(n8594), .ZN(n8601) );
  INV_X1 U9747 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10229) );
  OR2_X1 U9748 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10229), .ZN(n8801) );
  OAI21_X1 U9749 ( .B1(n8988), .B2(n8680), .A(n8801), .ZN(n8596) );
  AOI21_X1 U9750 ( .B1(n8686), .B2(n8958), .A(n8596), .ZN(n8597) );
  OAI21_X1 U9751 ( .B1(n8992), .B2(n8683), .A(n8597), .ZN(n8598) );
  AOI21_X1 U9752 ( .B1(n8599), .B2(n8673), .A(n8598), .ZN(n8600) );
  OAI21_X1 U9753 ( .B1(n8601), .B2(n8676), .A(n8600), .ZN(P2_U3168) );
  XOR2_X1 U9754 ( .A(n8603), .B(n8602), .Z(n8608) );
  AOI22_X1 U9755 ( .A1(n8693), .A2(n8686), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8605) );
  NAND2_X1 U9756 ( .A1(n8663), .A2(n8695), .ZN(n8604) );
  OAI211_X1 U9757 ( .C1(n8683), .C2(n8892), .A(n8605), .B(n8604), .ZN(n8606)
         );
  AOI21_X1 U9758 ( .B1(n8891), .B2(n8673), .A(n8606), .ZN(n8607) );
  OAI21_X1 U9759 ( .B1(n8608), .B2(n8676), .A(n8607), .ZN(P2_U3169) );
  INV_X1 U9760 ( .A(n8950), .ZN(n9067) );
  OAI21_X1 U9761 ( .B1(n8611), .B2(n8610), .A(n8609), .ZN(n8612) );
  NAND2_X1 U9762 ( .A1(n8612), .A2(n8624), .ZN(n8618) );
  INV_X1 U9763 ( .A(n8947), .ZN(n8616) );
  AOI22_X1 U9764 ( .A1(n8943), .A2(n8686), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8613) );
  OAI21_X1 U9765 ( .B1(n8977), .B2(n8680), .A(n8613), .ZN(n8614) );
  AOI21_X1 U9766 ( .B1(n8616), .B2(n8615), .A(n8614), .ZN(n8617) );
  OAI211_X1 U9767 ( .C1(n9067), .C2(n8689), .A(n8618), .B(n8617), .ZN(P2_U3173) );
  INV_X1 U9768 ( .A(n8619), .ZN(n8622) );
  INV_X1 U9769 ( .A(n8620), .ZN(n8621) );
  AOI21_X1 U9770 ( .B1(n8623), .B2(n8622), .A(n8621), .ZN(n8625) );
  OAI21_X1 U9771 ( .B1(n8626), .B2(n8625), .A(n8624), .ZN(n8632) );
  OR2_X1 U9772 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5947), .ZN(n8734) );
  OAI21_X1 U9773 ( .B1(n8627), .B2(n8680), .A(n8734), .ZN(n8630) );
  NOR2_X1 U9774 ( .A1(n8683), .A2(n8628), .ZN(n8629) );
  AOI211_X1 U9775 ( .C1(n8686), .C2(n8699), .A(n8630), .B(n8629), .ZN(n8631)
         );
  OAI211_X1 U9776 ( .C1(n10787), .C2(n8689), .A(n8632), .B(n8631), .ZN(
        P2_U3174) );
  AOI21_X1 U9777 ( .B1(n8634), .B2(n8633), .A(n8676), .ZN(n8636) );
  NAND2_X1 U9778 ( .A1(n8636), .A2(n8635), .ZN(n8640) );
  OAI22_X1 U9779 ( .A1(n8913), .A2(n8680), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10235), .ZN(n8638) );
  NOR2_X1 U9780 ( .A1(n8683), .A2(n8916), .ZN(n8637) );
  AOI211_X1 U9781 ( .C1(n8686), .C2(n8695), .A(n8638), .B(n8637), .ZN(n8639)
         );
  OAI211_X1 U9782 ( .C1(n9125), .C2(n8689), .A(n8640), .B(n8639), .ZN(P2_U3175) );
  NOR2_X1 U9783 ( .A1(n8641), .A2(n8680), .ZN(n8642) );
  AOI211_X1 U9784 ( .C1(n8686), .C2(n8701), .A(n8643), .B(n8642), .ZN(n8644)
         );
  OAI21_X1 U9785 ( .B1(n8645), .B2(n8683), .A(n8644), .ZN(n8653) );
  INV_X1 U9786 ( .A(n8646), .ZN(n8648) );
  NAND3_X1 U9787 ( .A1(n8649), .A2(n8648), .A3(n8647), .ZN(n8650) );
  AOI21_X1 U9788 ( .B1(n8651), .B2(n8650), .A(n8676), .ZN(n8652) );
  AOI211_X1 U9789 ( .C1(n10746), .C2(n8673), .A(n8653), .B(n8652), .ZN(n8654)
         );
  INV_X1 U9790 ( .A(n8654), .ZN(P2_U3176) );
  AOI21_X1 U9791 ( .B1(n8657), .B2(n8656), .A(n8676), .ZN(n8659) );
  NAND2_X1 U9792 ( .A1(n8659), .A2(n8658), .ZN(n8665) );
  NAND2_X1 U9793 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8817) );
  OAI21_X1 U9794 ( .B1(n8977), .B2(n8660), .A(n8817), .ZN(n8662) );
  NOR2_X1 U9795 ( .A1(n8683), .A2(n8980), .ZN(n8661) );
  AOI211_X1 U9796 ( .C1(n8663), .C2(n8696), .A(n8662), .B(n8661), .ZN(n8664)
         );
  OAI211_X1 U9797 ( .C1(n9135), .C2(n8689), .A(n8665), .B(n8664), .ZN(P2_U3178) );
  NAND2_X1 U9798 ( .A1(n5353), .A2(n8668), .ZN(n8669) );
  XNOR2_X1 U9799 ( .A(n8666), .B(n8669), .ZN(n8675) );
  OAI22_X1 U9800 ( .A1(n8890), .A2(n8680), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10364), .ZN(n8670) );
  AOI21_X1 U9801 ( .B1(n8686), .B2(n8843), .A(n8670), .ZN(n8671) );
  OAI21_X1 U9802 ( .B1(n8872), .B2(n8683), .A(n8671), .ZN(n8672) );
  AOI21_X1 U9803 ( .B1(n8871), .B2(n8673), .A(n8672), .ZN(n8674) );
  OAI21_X1 U9804 ( .B1(n8675), .B2(n8676), .A(n8674), .ZN(P2_U3180) );
  AOI21_X1 U9805 ( .B1(n8678), .B2(n8677), .A(n8676), .ZN(n8679) );
  NAND2_X1 U9806 ( .A1(n8679), .A2(n5556), .ZN(n8688) );
  INV_X1 U9807 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10363) );
  OR2_X1 U9808 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10363), .ZN(n8763) );
  OAI21_X1 U9809 ( .B1(n8681), .B2(n8680), .A(n8763), .ZN(n8685) );
  NOR2_X1 U9810 ( .A1(n8683), .A2(n8682), .ZN(n8684) );
  AOI211_X1 U9811 ( .C1(n8686), .C2(n8697), .A(n8685), .B(n8684), .ZN(n8687)
         );
  OAI211_X1 U9812 ( .C1(n10800), .C2(n8689), .A(n8688), .B(n8687), .ZN(
        P2_U3181) );
  MUX2_X1 U9813 ( .A(n8826), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8812), .Z(
        P2_U3522) );
  MUX2_X1 U9814 ( .A(n8690), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8812), .Z(
        P2_U3521) );
  MUX2_X1 U9815 ( .A(n8844), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8812), .Z(
        P2_U3520) );
  MUX2_X1 U9816 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8691), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9817 ( .A(n8843), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8812), .Z(
        P2_U3518) );
  MUX2_X1 U9818 ( .A(n8692), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8812), .Z(
        P2_U3517) );
  MUX2_X1 U9819 ( .A(n8693), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8812), .Z(
        P2_U3516) );
  MUX2_X1 U9820 ( .A(n8694), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8812), .Z(
        P2_U3515) );
  MUX2_X1 U9821 ( .A(n8695), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8812), .Z(
        P2_U3514) );
  MUX2_X1 U9822 ( .A(n8927), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8812), .Z(
        P2_U3513) );
  MUX2_X1 U9823 ( .A(n8943), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8812), .Z(
        P2_U3512) );
  MUX2_X1 U9824 ( .A(n8959), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8812), .Z(
        P2_U3511) );
  MUX2_X1 U9825 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8944), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9826 ( .A(n8958), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8812), .Z(
        P2_U3509) );
  MUX2_X1 U9827 ( .A(n8696), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8812), .Z(
        P2_U3508) );
  MUX2_X1 U9828 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8697), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9829 ( .A(n8698), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8812), .Z(
        P2_U3506) );
  MUX2_X1 U9830 ( .A(n8699), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8812), .Z(
        P2_U3505) );
  MUX2_X1 U9831 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8700), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9832 ( .A(n8701), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8812), .Z(
        P2_U3503) );
  MUX2_X1 U9833 ( .A(n8702), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8812), .Z(
        P2_U3502) );
  MUX2_X1 U9834 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8703), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9835 ( .A(n8704), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8812), .Z(
        P2_U3500) );
  MUX2_X1 U9836 ( .A(n8705), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8812), .Z(
        P2_U3499) );
  MUX2_X1 U9837 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8706), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9838 ( .A(n10635), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8812), .Z(
        P2_U3497) );
  MUX2_X1 U9839 ( .A(n8707), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8812), .Z(
        P2_U3496) );
  MUX2_X1 U9840 ( .A(n10636), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8812), .Z(
        P2_U3495) );
  MUX2_X1 U9841 ( .A(n10592), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8812), .Z(
        P2_U3494) );
  MUX2_X1 U9842 ( .A(n8708), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8812), .Z(
        P2_U3493) );
  MUX2_X1 U9843 ( .A(n10591), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8812), .Z(
        P2_U3492) );
  MUX2_X1 U9844 ( .A(n8709), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8812), .Z(
        P2_U3491) );
  AOI21_X1 U9845 ( .B1(n8712), .B2(n8711), .A(n8710), .ZN(n8726) );
  OAI21_X1 U9846 ( .B1(n8715), .B2(n8714), .A(n8713), .ZN(n8724) );
  AOI21_X1 U9847 ( .B1(n10516), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8716), .ZN(
        n8717) );
  OAI21_X1 U9848 ( .B1(n8718), .B2(n10511), .A(n8717), .ZN(n8723) );
  AOI21_X1 U9849 ( .B1(n5031), .B2(n8720), .A(n8719), .ZN(n8721) );
  NOR2_X1 U9850 ( .A1(n8721), .A2(n10514), .ZN(n8722) );
  AOI211_X1 U9851 ( .C1(n10519), .C2(n8724), .A(n8723), .B(n8722), .ZN(n8725)
         );
  OAI21_X1 U9852 ( .B1(n8726), .B2(n10496), .A(n8725), .ZN(P2_U3194) );
  AOI21_X1 U9853 ( .B1(n5946), .B2(n8728), .A(n8727), .ZN(n8741) );
  OAI21_X1 U9854 ( .B1(n8731), .B2(n8730), .A(n8729), .ZN(n8739) );
  NOR2_X1 U9855 ( .A1(n10511), .A2(n5050), .ZN(n8738) );
  AOI21_X1 U9856 ( .B1(n8733), .B2(n5950), .A(n8732), .ZN(n8736) );
  NAND2_X1 U9857 ( .A1(n10516), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8735) );
  OAI211_X1 U9858 ( .C1(n8736), .C2(n10496), .A(n8735), .B(n8734), .ZN(n8737)
         );
  AOI211_X1 U9859 ( .C1(n10519), .C2(n8739), .A(n8738), .B(n8737), .ZN(n8740)
         );
  OAI21_X1 U9860 ( .B1(n8741), .B2(n10514), .A(n8740), .ZN(P2_U3195) );
  AOI21_X1 U9861 ( .B1(n8744), .B2(n8743), .A(n8742), .ZN(n8758) );
  OAI21_X1 U9862 ( .B1(n8747), .B2(n8746), .A(n8745), .ZN(n8756) );
  NAND2_X1 U9863 ( .A1(n10516), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8749) );
  OAI211_X1 U9864 ( .C1(n10511), .C2(n8750), .A(n8749), .B(n8748), .ZN(n8755)
         );
  AOI21_X1 U9865 ( .B1(n4985), .B2(n8752), .A(n8751), .ZN(n8753) );
  NOR2_X1 U9866 ( .A1(n8753), .A2(n10514), .ZN(n8754) );
  AOI211_X1 U9867 ( .C1(n10519), .C2(n8756), .A(n8755), .B(n8754), .ZN(n8757)
         );
  OAI21_X1 U9868 ( .B1(n8758), .B2(n10496), .A(n8757), .ZN(P2_U3196) );
  AOI21_X1 U9869 ( .B1(n5977), .B2(n8760), .A(n8759), .ZN(n8775) );
  AOI21_X1 U9870 ( .B1(n8762), .B2(n7813), .A(n8761), .ZN(n8765) );
  NAND2_X1 U9871 ( .A1(n10516), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8764) );
  OAI211_X1 U9872 ( .C1(n8765), .C2(n10496), .A(n8764), .B(n8763), .ZN(n8768)
         );
  NOR2_X1 U9873 ( .A1(n10511), .A2(n8766), .ZN(n8767) );
  NOR2_X1 U9874 ( .A1(n8768), .A2(n8767), .ZN(n8774) );
  OAI21_X1 U9875 ( .B1(n8771), .B2(n8770), .A(n8769), .ZN(n8772) );
  NAND2_X1 U9876 ( .A1(n8772), .A2(n10519), .ZN(n8773) );
  OAI211_X1 U9877 ( .C1(n8775), .C2(n10514), .A(n8774), .B(n8773), .ZN(
        P2_U3197) );
  AOI21_X1 U9878 ( .B1(n8778), .B2(n8777), .A(n8776), .ZN(n8793) );
  OAI21_X1 U9879 ( .B1(n8781), .B2(n8780), .A(n8779), .ZN(n8791) );
  NAND2_X1 U9880 ( .A1(n10516), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8783) );
  OAI211_X1 U9881 ( .C1(n10511), .C2(n8784), .A(n8783), .B(n8782), .ZN(n8790)
         );
  AOI21_X1 U9882 ( .B1(n8787), .B2(n8786), .A(n8785), .ZN(n8788) );
  NOR2_X1 U9883 ( .A1(n8788), .A2(n10496), .ZN(n8789) );
  AOI211_X1 U9884 ( .C1(n10519), .C2(n8791), .A(n8790), .B(n8789), .ZN(n8792)
         );
  OAI21_X1 U9885 ( .B1(n8793), .B2(n10514), .A(n8792), .ZN(P2_U3198) );
  AOI21_X1 U9886 ( .B1(n9083), .B2(n8795), .A(n8794), .ZN(n8805) );
  OAI21_X1 U9887 ( .B1(n8798), .B2(n8797), .A(n8796), .ZN(n8803) );
  NOR2_X1 U9888 ( .A1(n10511), .A2(n8799), .ZN(n8802) );
  OAI21_X1 U9889 ( .B1(n8805), .B2(n10514), .A(n8804), .ZN(P2_U3199) );
  AOI21_X1 U9890 ( .B1(n8808), .B2(n8807), .A(n8806), .ZN(n8823) );
  INV_X1 U9891 ( .A(n8809), .ZN(n8810) );
  NOR2_X1 U9892 ( .A1(n8811), .A2(n8810), .ZN(n8819) );
  INV_X1 U9893 ( .A(n8819), .ZN(n8813) );
  OAI21_X1 U9894 ( .B1(n8813), .B2(n8812), .A(n10511), .ZN(n8820) );
  NAND2_X1 U9895 ( .A1(n10516), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8818) );
  OAI21_X1 U9896 ( .B1(n8823), .B2(n10514), .A(n8822), .ZN(P2_U3200) );
  NOR2_X1 U9897 ( .A1(n10650), .A2(n8824), .ZN(n8836) );
  NOR2_X1 U9898 ( .A1(n9017), .A2(n8836), .ZN(n8847) );
  NAND2_X1 U9899 ( .A1(n8826), .A2(n8825), .ZN(n9092) );
  NAND2_X1 U9900 ( .A1(n8847), .A2(n9092), .ZN(n8829) );
  OAI21_X1 U9901 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(n10709), .A(n8829), .ZN(
        n8827) );
  OAI21_X1 U9902 ( .B1(n9094), .B2(n10653), .A(n8827), .ZN(P2_U3202) );
  OAI21_X1 U9903 ( .B1(P2_REG2_REG_30__SCAN_IN), .B2(n10709), .A(n8829), .ZN(
        n8830) );
  OAI21_X1 U9904 ( .B1(n9098), .B2(n10653), .A(n8830), .ZN(P2_U3203) );
  AOI21_X1 U9905 ( .B1(n8833), .B2(n8832), .A(n8831), .ZN(n8838) );
  NOR2_X1 U9906 ( .A1(n8834), .A2(n10653), .ZN(n8835) );
  AOI211_X1 U9907 ( .C1(n9017), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8836), .B(
        n8835), .ZN(n8837) );
  OAI21_X1 U9908 ( .B1(n8838), .B2(n9017), .A(n8837), .ZN(P2_U3204) );
  XNOR2_X1 U9909 ( .A(n8841), .B(n6127), .ZN(n8842) );
  NAND2_X1 U9910 ( .A1(n8842), .A2(n10641), .ZN(n8846) );
  AOI22_X1 U9911 ( .A1(n6190), .A2(n8844), .B1(n8843), .B2(n10637), .ZN(n8845)
         );
  NAND2_X1 U9912 ( .A1(n8846), .A2(n8845), .ZN(n9034) );
  OAI21_X1 U9913 ( .B1(n8848), .B2(n10650), .A(n8847), .ZN(n8849) );
  OAI22_X1 U9914 ( .A1(n9034), .A2(n8849), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10709), .ZN(n8852) );
  XNOR2_X1 U9915 ( .A(n8850), .B(n6127), .ZN(n9032) );
  NAND2_X1 U9916 ( .A1(n9032), .A2(n9015), .ZN(n8851) );
  OAI211_X1 U9917 ( .C1(n9102), .C2(n10653), .A(n8852), .B(n8851), .ZN(
        P2_U3205) );
  INV_X1 U9918 ( .A(n9037), .ZN(n8865) );
  NAND2_X1 U9919 ( .A1(n8856), .A2(n8855), .ZN(n8858) );
  XNOR2_X1 U9920 ( .A(n8858), .B(n8857), .ZN(n9038) );
  NOR2_X1 U9921 ( .A1(n9105), .A2(n10653), .ZN(n8863) );
  OAI22_X1 U9922 ( .A1(n10709), .A2(n8861), .B1(n8860), .B2(n10650), .ZN(n8862) );
  AOI211_X1 U9923 ( .C1(n9038), .C2(n9015), .A(n8863), .B(n8862), .ZN(n8864)
         );
  OAI21_X1 U9924 ( .B1(n8865), .B2(n9017), .A(n8864), .ZN(P2_U3206) );
  XNOR2_X1 U9925 ( .A(n8866), .B(n8869), .ZN(n8867) );
  OAI222_X1 U9926 ( .A1(n9003), .A2(n8890), .B1(n9005), .B2(n8868), .C1(n9000), 
        .C2(n8867), .ZN(n9041) );
  INV_X1 U9927 ( .A(n9041), .ZN(n8877) );
  XNOR2_X1 U9928 ( .A(n8870), .B(n8869), .ZN(n9042) );
  INV_X1 U9929 ( .A(n8871), .ZN(n9109) );
  NOR2_X1 U9930 ( .A1(n9109), .A2(n10653), .ZN(n8875) );
  OAI22_X1 U9931 ( .A1(n10709), .A2(n8873), .B1(n8872), .B2(n10650), .ZN(n8874) );
  AOI211_X1 U9932 ( .C1(n9042), .C2(n9015), .A(n8875), .B(n8874), .ZN(n8876)
         );
  OAI21_X1 U9933 ( .B1(n8877), .B2(n9017), .A(n8876), .ZN(P2_U3207) );
  INV_X1 U9934 ( .A(n10598), .ZN(n8881) );
  XNOR2_X1 U9935 ( .A(n8878), .B(n5005), .ZN(n8879) );
  OAI222_X1 U9936 ( .A1(n9005), .A2(n8880), .B1(n9003), .B2(n8901), .C1(n9000), 
        .C2(n8879), .ZN(n9046) );
  AOI21_X1 U9937 ( .B1(n8881), .B2(n9045), .A(n9046), .ZN(n8887) );
  XNOR2_X1 U9938 ( .A(n8882), .B(n5005), .ZN(n9047) );
  OAI22_X1 U9939 ( .A1(n10709), .A2(n8884), .B1(n8883), .B2(n10650), .ZN(n8885) );
  AOI21_X1 U9940 ( .B1(n9047), .B2(n9015), .A(n8885), .ZN(n8886) );
  OAI21_X1 U9941 ( .B1(n8887), .B2(n9017), .A(n8886), .ZN(P2_U3208) );
  XNOR2_X1 U9942 ( .A(n8888), .B(n8894), .ZN(n8889) );
  OAI222_X1 U9943 ( .A1(n9003), .A2(n8912), .B1(n9005), .B2(n8890), .C1(n8889), 
        .C2(n9000), .ZN(n9050) );
  INV_X1 U9944 ( .A(n8891), .ZN(n9117) );
  OAI22_X1 U9945 ( .A1(n9117), .A2(n10598), .B1(n8892), .B2(n10650), .ZN(n8893) );
  OAI21_X1 U9946 ( .B1(n9050), .B2(n8893), .A(n10709), .ZN(n8897) );
  XNOR2_X1 U9947 ( .A(n8895), .B(n8894), .ZN(n9051) );
  AOI22_X1 U9948 ( .A1(n9051), .A2(n9015), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9017), .ZN(n8896) );
  NAND2_X1 U9949 ( .A1(n8897), .A2(n8896), .ZN(P2_U3209) );
  XNOR2_X1 U9950 ( .A(n8898), .B(n8903), .ZN(n8899) );
  OAI222_X1 U9951 ( .A1(n9005), .A2(n8901), .B1(n9003), .B2(n8900), .C1(n8899), 
        .C2(n9000), .ZN(n9054) );
  INV_X1 U9952 ( .A(n9054), .ZN(n8910) );
  XOR2_X1 U9953 ( .A(n8903), .B(n8902), .Z(n9055) );
  INV_X1 U9954 ( .A(n8904), .ZN(n9121) );
  NOR2_X1 U9955 ( .A1(n9121), .A2(n10653), .ZN(n8908) );
  OAI22_X1 U9956 ( .A1(n10709), .A2(n8906), .B1(n8905), .B2(n10650), .ZN(n8907) );
  AOI211_X1 U9957 ( .C1(n9055), .C2(n9015), .A(n8908), .B(n8907), .ZN(n8909)
         );
  OAI21_X1 U9958 ( .B1(n8910), .B2(n9017), .A(n8909), .ZN(P2_U3210) );
  OAI222_X1 U9959 ( .A1(n9003), .A2(n8913), .B1(n9005), .B2(n8912), .C1(n8911), 
        .C2(n9000), .ZN(n9058) );
  INV_X1 U9960 ( .A(n9058), .ZN(n8921) );
  XNOR2_X1 U9961 ( .A(n8915), .B(n8914), .ZN(n9059) );
  NOR2_X1 U9962 ( .A1(n9125), .A2(n10653), .ZN(n8919) );
  OAI22_X1 U9963 ( .A1(n10709), .A2(n8917), .B1(n8916), .B2(n10650), .ZN(n8918) );
  AOI211_X1 U9964 ( .C1(n9059), .C2(n9015), .A(n8919), .B(n8918), .ZN(n8920)
         );
  OAI21_X1 U9965 ( .B1(n8921), .B2(n9017), .A(n8920), .ZN(P2_U3211) );
  XNOR2_X1 U9966 ( .A(n8923), .B(n8922), .ZN(n9064) );
  XNOR2_X1 U9967 ( .A(n8925), .B(n8924), .ZN(n8926) );
  NAND2_X1 U9968 ( .A1(n8926), .A2(n10641), .ZN(n8929) );
  AOI22_X1 U9969 ( .A1(n6190), .A2(n8927), .B1(n8959), .B2(n10637), .ZN(n8928)
         );
  NAND2_X1 U9970 ( .A1(n8929), .A2(n8928), .ZN(n9066) );
  NAND2_X1 U9971 ( .A1(n9066), .A2(n10709), .ZN(n8934) );
  OAI22_X1 U9972 ( .A1(n10709), .A2(n8931), .B1(n8930), .B2(n10650), .ZN(n8932) );
  AOI21_X1 U9973 ( .B1(n9062), .B2(n10704), .A(n8932), .ZN(n8933) );
  OAI211_X1 U9974 ( .C1(n9064), .C2(n8968), .A(n8934), .B(n8933), .ZN(P2_U3212) );
  OR2_X1 U9975 ( .A1(n8935), .A2(n8938), .ZN(n8936) );
  NAND2_X1 U9976 ( .A1(n8937), .A2(n8936), .ZN(n9068) );
  NAND2_X1 U9977 ( .A1(n8939), .A2(n8938), .ZN(n8940) );
  NAND2_X1 U9978 ( .A1(n8941), .A2(n8940), .ZN(n8942) );
  NAND2_X1 U9979 ( .A1(n8942), .A2(n10641), .ZN(n8946) );
  AOI22_X1 U9980 ( .A1(n8944), .A2(n10637), .B1(n6190), .B2(n8943), .ZN(n8945)
         );
  NAND2_X1 U9981 ( .A1(n8946), .A2(n8945), .ZN(n9070) );
  NAND2_X1 U9982 ( .A1(n9070), .A2(n10709), .ZN(n8952) );
  OAI22_X1 U9983 ( .A1(n10709), .A2(n8948), .B1(n8947), .B2(n10650), .ZN(n8949) );
  AOI21_X1 U9984 ( .B1(n8950), .B2(n10704), .A(n8949), .ZN(n8951) );
  OAI211_X1 U9985 ( .C1(n9068), .C2(n8968), .A(n8952), .B(n8951), .ZN(P2_U3213) );
  AND2_X1 U9986 ( .A1(n8954), .A2(n8953), .ZN(n8957) );
  OAI211_X1 U9987 ( .C1(n8957), .C2(n8956), .A(n10641), .B(n8955), .ZN(n8961)
         );
  AOI22_X1 U9988 ( .A1(n6190), .A2(n8959), .B1(n8958), .B2(n10637), .ZN(n8960)
         );
  NAND2_X1 U9989 ( .A1(n8961), .A2(n8960), .ZN(n9072) );
  INV_X1 U9990 ( .A(n9072), .ZN(n8974) );
  OAI22_X1 U9991 ( .A1(n10709), .A2(n8963), .B1(n8962), .B2(n10650), .ZN(n8971) );
  NAND2_X1 U9992 ( .A1(n8965), .A2(n8964), .ZN(n8967) );
  NOR2_X1 U9993 ( .A1(n8967), .A2(n8966), .ZN(n9071) );
  NAND2_X1 U9994 ( .A1(n8967), .A2(n8966), .ZN(n9073) );
  INV_X1 U9995 ( .A(n9073), .ZN(n8969) );
  NOR3_X1 U9996 ( .A1(n9071), .A2(n8969), .A3(n8968), .ZN(n8970) );
  AOI211_X1 U9997 ( .C1(n10704), .C2(n8972), .A(n8971), .B(n8970), .ZN(n8973)
         );
  OAI21_X1 U9998 ( .B1(n9017), .B2(n8974), .A(n8973), .ZN(P2_U3214) );
  XOR2_X1 U9999 ( .A(n8978), .B(n8975), .Z(n8976) );
  OAI222_X1 U10000 ( .A1(n9005), .A2(n8977), .B1(n9003), .B2(n9004), .C1(n8976), .C2(n9000), .ZN(n9077) );
  INV_X1 U10001 ( .A(n9077), .ZN(n8985) );
  XOR2_X1 U10002 ( .A(n8979), .B(n8978), .Z(n9078) );
  NOR2_X1 U10003 ( .A1(n9135), .A2(n10653), .ZN(n8983) );
  OAI22_X1 U10004 ( .A1(n10709), .A2(n8981), .B1(n8980), .B2(n10650), .ZN(
        n8982) );
  AOI211_X1 U10005 ( .C1(n9078), .C2(n9015), .A(n8983), .B(n8982), .ZN(n8984)
         );
  OAI21_X1 U10006 ( .B1(n8985), .B2(n9017), .A(n8984), .ZN(P2_U3215) );
  XNOR2_X1 U10007 ( .A(n8986), .B(n8990), .ZN(n8987) );
  OAI222_X1 U10008 ( .A1(n9005), .A2(n8989), .B1(n9003), .B2(n8988), .C1(n9000), .C2(n8987), .ZN(n9081) );
  INV_X1 U10009 ( .A(n9081), .ZN(n8997) );
  XNOR2_X1 U10010 ( .A(n8991), .B(n8990), .ZN(n9082) );
  NOR2_X1 U10011 ( .A1(n9139), .A2(n10653), .ZN(n8995) );
  OAI22_X1 U10012 ( .A1(n10709), .A2(n8993), .B1(n8992), .B2(n10650), .ZN(
        n8994) );
  AOI211_X1 U10013 ( .C1(n9082), .C2(n9015), .A(n8995), .B(n8994), .ZN(n8996)
         );
  OAI21_X1 U10014 ( .B1(n8997), .B2(n9017), .A(n8996), .ZN(P2_U3216) );
  XNOR2_X1 U10015 ( .A(n8999), .B(n8998), .ZN(n9001) );
  OAI222_X1 U10016 ( .A1(n9005), .A2(n9004), .B1(n9003), .B2(n9002), .C1(n9001), .C2(n9000), .ZN(n9085) );
  INV_X1 U10017 ( .A(n9085), .ZN(n9018) );
  NAND2_X1 U10018 ( .A1(n9007), .A2(n9006), .ZN(n9009) );
  XNOR2_X1 U10019 ( .A(n9009), .B(n9008), .ZN(n9086) );
  INV_X1 U10020 ( .A(n9010), .ZN(n9144) );
  NOR2_X1 U10021 ( .A1(n9144), .A2(n10653), .ZN(n9014) );
  OAI22_X1 U10022 ( .A1(n10709), .A2(n9012), .B1(n9011), .B2(n10650), .ZN(
        n9013) );
  AOI211_X1 U10023 ( .C1(n9086), .C2(n9015), .A(n9014), .B(n9013), .ZN(n9016)
         );
  OAI21_X1 U10024 ( .B1(n9018), .B2(n9017), .A(n9016), .ZN(P2_U3217) );
  AOI22_X1 U10025 ( .A1(n10704), .A2(n9019), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10706), .ZN(n9028) );
  MUX2_X1 U10026 ( .A(n6318), .B(n9020), .S(n10709), .Z(n9027) );
  INV_X1 U10027 ( .A(n9021), .ZN(n9024) );
  INV_X1 U10028 ( .A(n9022), .ZN(n9023) );
  NAND4_X1 U10029 ( .A1(n9025), .A2(n9024), .A3(n9023), .A4(n10799), .ZN(n9026) );
  NAND3_X1 U10030 ( .A1(n9028), .A2(n9027), .A3(n9026), .ZN(P2_U3233) );
  NOR2_X1 U10031 ( .A1(n10805), .A2(n9092), .ZN(n9030) );
  AOI21_X1 U10032 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10805), .A(n9030), .ZN(
        n9029) );
  OAI21_X1 U10033 ( .B1(n9094), .B2(n9089), .A(n9029), .ZN(P2_U3490) );
  AOI21_X1 U10034 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10805), .A(n9030), .ZN(
        n9031) );
  OAI21_X1 U10035 ( .B1(n9098), .B2(n9089), .A(n9031), .ZN(P2_U3489) );
  INV_X1 U10036 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9035) );
  AND2_X1 U10037 ( .A1(n9032), .A2(n10720), .ZN(n9033) );
  NOR2_X1 U10038 ( .A1(n9034), .A2(n9033), .ZN(n9099) );
  MUX2_X1 U10039 ( .A(n9035), .B(n9099), .S(n10748), .Z(n9036) );
  OAI21_X1 U10040 ( .B1(n9102), .B2(n9089), .A(n9036), .ZN(P2_U3487) );
  MUX2_X1 U10041 ( .A(n9039), .B(n9103), .S(n10806), .Z(n9040) );
  OAI21_X1 U10042 ( .B1(n9105), .B2(n9089), .A(n9040), .ZN(P2_U3486) );
  AOI21_X1 U10043 ( .B1(n9042), .B2(n10720), .A(n9041), .ZN(n9106) );
  MUX2_X1 U10044 ( .A(n9043), .B(n9106), .S(n10748), .Z(n9044) );
  OAI21_X1 U10045 ( .B1(n9109), .B2(n9089), .A(n9044), .ZN(P2_U3485) );
  INV_X1 U10046 ( .A(n9045), .ZN(n9113) );
  AOI21_X1 U10047 ( .B1(n9047), .B2(n10720), .A(n9046), .ZN(n9110) );
  MUX2_X1 U10048 ( .A(n9048), .B(n9110), .S(n10806), .Z(n9049) );
  OAI21_X1 U10049 ( .B1(n9113), .B2(n9089), .A(n9049), .ZN(P2_U3484) );
  AOI21_X1 U10050 ( .B1(n10720), .B2(n9051), .A(n9050), .ZN(n9114) );
  MUX2_X1 U10051 ( .A(n9052), .B(n9114), .S(n10806), .Z(n9053) );
  OAI21_X1 U10052 ( .B1(n9117), .B2(n9089), .A(n9053), .ZN(P2_U3483) );
  AOI21_X1 U10053 ( .B1(n9055), .B2(n10720), .A(n9054), .ZN(n9118) );
  MUX2_X1 U10054 ( .A(n9056), .B(n9118), .S(n10806), .Z(n9057) );
  OAI21_X1 U10055 ( .B1(n9121), .B2(n9089), .A(n9057), .ZN(P2_U3482) );
  INV_X1 U10056 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9060) );
  AOI21_X1 U10057 ( .B1(n10720), .B2(n9059), .A(n9058), .ZN(n9122) );
  MUX2_X1 U10058 ( .A(n9060), .B(n9122), .S(n10806), .Z(n9061) );
  OAI21_X1 U10059 ( .B1(n9125), .B2(n9089), .A(n9061), .ZN(P2_U3481) );
  INV_X1 U10060 ( .A(n9062), .ZN(n9063) );
  OAI22_X1 U10061 ( .A1(n9064), .A2(n10801), .B1(n9063), .B2(n10799), .ZN(
        n9065) );
  MUX2_X1 U10062 ( .A(n9126), .B(P2_REG1_REG_21__SCAN_IN), .S(n10805), .Z(
        P2_U3480) );
  OAI22_X1 U10063 ( .A1(n9068), .A2(n10801), .B1(n9067), .B2(n10799), .ZN(
        n9069) );
  MUX2_X1 U10064 ( .A(n9127), .B(P2_REG1_REG_20__SCAN_IN), .S(n10805), .Z(
        P2_U3479) );
  NOR2_X1 U10065 ( .A1(n9071), .A2(n10801), .ZN(n9074) );
  AOI21_X1 U10066 ( .B1(n9074), .B2(n9073), .A(n9072), .ZN(n9128) );
  MUX2_X1 U10067 ( .A(n9075), .B(n9128), .S(n10806), .Z(n9076) );
  OAI21_X1 U10068 ( .B1(n9131), .B2(n9089), .A(n9076), .ZN(P2_U3478) );
  INV_X1 U10069 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9079) );
  AOI21_X1 U10070 ( .B1(n10720), .B2(n9078), .A(n9077), .ZN(n9132) );
  MUX2_X1 U10071 ( .A(n9079), .B(n9132), .S(n10806), .Z(n9080) );
  OAI21_X1 U10072 ( .B1(n9135), .B2(n9089), .A(n9080), .ZN(P2_U3477) );
  AOI21_X1 U10073 ( .B1(n9082), .B2(n10720), .A(n9081), .ZN(n9136) );
  MUX2_X1 U10074 ( .A(n9083), .B(n9136), .S(n10806), .Z(n9084) );
  OAI21_X1 U10075 ( .B1(n9139), .B2(n9089), .A(n9084), .ZN(P2_U3476) );
  AOI21_X1 U10076 ( .B1(n9086), .B2(n10720), .A(n9085), .ZN(n9140) );
  MUX2_X1 U10077 ( .A(n9087), .B(n9140), .S(n10806), .Z(n9088) );
  OAI21_X1 U10078 ( .B1(n9144), .B2(n9089), .A(n9088), .ZN(P2_U3475) );
  NAND2_X1 U10079 ( .A1(n9091), .A2(n9090), .ZN(n9097) );
  NOR2_X1 U10080 ( .A1(n10807), .A2(n9092), .ZN(n9095) );
  AOI21_X1 U10081 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(n10807), .A(n9095), .ZN(
        n9093) );
  OAI21_X1 U10082 ( .B1(n9094), .B2(n9097), .A(n9093), .ZN(P2_U3458) );
  AOI21_X1 U10083 ( .B1(P2_REG0_REG_30__SCAN_IN), .B2(n10807), .A(n9095), .ZN(
        n9096) );
  OAI21_X1 U10084 ( .B1(n9098), .B2(n9097), .A(n9096), .ZN(P2_U3457) );
  MUX2_X1 U10085 ( .A(n9100), .B(n9099), .S(n10810), .Z(n9101) );
  OAI21_X1 U10086 ( .B1(n9102), .B2(n9143), .A(n9101), .ZN(P2_U3455) );
  INV_X1 U10087 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9104) );
  INV_X1 U10088 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9107) );
  MUX2_X1 U10089 ( .A(n9107), .B(n9106), .S(n10810), .Z(n9108) );
  OAI21_X1 U10090 ( .B1(n9109), .B2(n9143), .A(n9108), .ZN(P2_U3453) );
  INV_X1 U10091 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9111) );
  MUX2_X1 U10092 ( .A(n9111), .B(n9110), .S(n10810), .Z(n9112) );
  OAI21_X1 U10093 ( .B1(n9113), .B2(n9143), .A(n9112), .ZN(P2_U3452) );
  INV_X1 U10094 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9115) );
  MUX2_X1 U10095 ( .A(n9115), .B(n9114), .S(n10810), .Z(n9116) );
  OAI21_X1 U10096 ( .B1(n9117), .B2(n9143), .A(n9116), .ZN(P2_U3451) );
  INV_X1 U10097 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9119) );
  MUX2_X1 U10098 ( .A(n9119), .B(n9118), .S(n10810), .Z(n9120) );
  OAI21_X1 U10099 ( .B1(n9121), .B2(n9143), .A(n9120), .ZN(P2_U3450) );
  MUX2_X1 U10100 ( .A(n9123), .B(n9122), .S(n10810), .Z(n9124) );
  OAI21_X1 U10101 ( .B1(n9125), .B2(n9143), .A(n9124), .ZN(P2_U3449) );
  MUX2_X1 U10102 ( .A(n9126), .B(P2_REG0_REG_21__SCAN_IN), .S(n10807), .Z(
        P2_U3448) );
  MUX2_X1 U10103 ( .A(n9127), .B(P2_REG0_REG_20__SCAN_IN), .S(n10807), .Z(
        P2_U3447) );
  INV_X1 U10104 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9129) );
  MUX2_X1 U10105 ( .A(n9129), .B(n9128), .S(n10810), .Z(n9130) );
  OAI21_X1 U10106 ( .B1(n9131), .B2(n9143), .A(n9130), .ZN(P2_U3446) );
  MUX2_X1 U10107 ( .A(n9133), .B(n9132), .S(n10810), .Z(n9134) );
  OAI21_X1 U10108 ( .B1(n9135), .B2(n9143), .A(n9134), .ZN(P2_U3444) );
  INV_X1 U10109 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9137) );
  MUX2_X1 U10110 ( .A(n9137), .B(n9136), .S(n10810), .Z(n9138) );
  OAI21_X1 U10111 ( .B1(n9139), .B2(n9143), .A(n9138), .ZN(P2_U3441) );
  INV_X1 U10112 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9141) );
  MUX2_X1 U10113 ( .A(n9141), .B(n9140), .S(n10810), .Z(n9142) );
  OAI21_X1 U10114 ( .B1(n9144), .B2(n9143), .A(n9142), .ZN(P2_U3438) );
  INV_X1 U10115 ( .A(n9145), .ZN(n10128) );
  NOR4_X1 U10116 ( .A1(n9146), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5807), .ZN(n9147) );
  AOI21_X1 U10117 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9160), .A(n9147), .ZN(
        n9148) );
  OAI21_X1 U10118 ( .B1(n10128), .B2(n9162), .A(n9148), .ZN(P2_U3264) );
  AOI22_X1 U10119 ( .A1(n9149), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9160), .ZN(n9150) );
  OAI21_X1 U10120 ( .B1(n9151), .B2(n9162), .A(n9150), .ZN(P2_U3265) );
  INV_X1 U10121 ( .A(n9152), .ZN(n10129) );
  OAI222_X1 U10122 ( .A1(P2_U3151), .A2(n9154), .B1(n9162), .B2(n10129), .C1(
        n10370), .C2(n9153), .ZN(P2_U3266) );
  INV_X1 U10123 ( .A(n9155), .ZN(n10134) );
  AOI21_X1 U10124 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9160), .A(n9156), .ZN(
        n9157) );
  OAI21_X1 U10125 ( .B1(n10134), .B2(n9162), .A(n9157), .ZN(P2_U3267) );
  INV_X1 U10126 ( .A(n9158), .ZN(n10137) );
  AOI21_X1 U10127 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9160), .A(n9159), .ZN(
        n9161) );
  OAI21_X1 U10128 ( .B1(n10137), .B2(n9162), .A(n9161), .ZN(P2_U3268) );
  MUX2_X1 U10129 ( .A(n9163), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI22_X1 U10130 ( .A1(n9831), .A2(n4948), .B1(n9307), .B2(n9722), .ZN(n9294)
         );
  AOI22_X1 U10131 ( .A1(n9831), .A2(n6725), .B1(n4948), .B2(n9722), .ZN(n9164)
         );
  XNOR2_X1 U10132 ( .A(n9164), .B(n9314), .ZN(n9293) );
  AOI21_X1 U10133 ( .B1(n9167), .B2(n9166), .A(n9165), .ZN(n9178) );
  INV_X1 U10134 ( .A(n9178), .ZN(n9172) );
  NAND2_X1 U10135 ( .A1(n9557), .A2(n9309), .ZN(n9169) );
  NAND2_X1 U10136 ( .A1(n9179), .A2(n6725), .ZN(n9168) );
  NAND2_X1 U10137 ( .A1(n9169), .A2(n9168), .ZN(n9170) );
  XNOR2_X1 U10138 ( .A(n9170), .B(n9373), .ZN(n9177) );
  INV_X1 U10139 ( .A(n9177), .ZN(n9171) );
  NAND2_X1 U10140 ( .A1(n9172), .A2(n9171), .ZN(n9389) );
  NAND2_X1 U10141 ( .A1(n9556), .A2(n9309), .ZN(n9174) );
  NAND2_X1 U10142 ( .A1(n9465), .A2(n6725), .ZN(n9173) );
  NAND2_X1 U10143 ( .A1(n9174), .A2(n9173), .ZN(n9175) );
  XNOR2_X1 U10144 ( .A(n9175), .B(n9373), .ZN(n9183) );
  AOI22_X1 U10145 ( .A1(n9556), .A2(n9307), .B1(n4948), .B2(n9465), .ZN(n9182)
         );
  XNOR2_X1 U10146 ( .A(n9183), .B(n9182), .ZN(n9458) );
  INV_X1 U10147 ( .A(n9458), .ZN(n9176) );
  NAND2_X1 U10148 ( .A1(n9178), .A2(n9177), .ZN(n9390) );
  NAND2_X1 U10149 ( .A1(n9557), .A2(n9307), .ZN(n9181) );
  NAND2_X1 U10150 ( .A1(n9179), .A2(n9309), .ZN(n9180) );
  NAND2_X1 U10151 ( .A1(n9181), .A2(n9180), .ZN(n9391) );
  NAND2_X1 U10152 ( .A1(n9390), .A2(n9391), .ZN(n9455) );
  NAND2_X1 U10153 ( .A1(n9183), .A2(n9182), .ZN(n9184) );
  NAND2_X1 U10154 ( .A1(n9555), .A2(n9309), .ZN(n9186) );
  NAND2_X1 U10155 ( .A1(n9188), .A2(n6725), .ZN(n9185) );
  NAND2_X1 U10156 ( .A1(n9186), .A2(n9185), .ZN(n9187) );
  XNOR2_X1 U10157 ( .A(n9187), .B(n9373), .ZN(n9191) );
  NAND2_X1 U10158 ( .A1(n9555), .A2(n9307), .ZN(n9190) );
  NAND2_X1 U10159 ( .A1(n9188), .A2(n4948), .ZN(n9189) );
  AND2_X1 U10160 ( .A1(n9190), .A2(n9189), .ZN(n9352) );
  NAND2_X1 U10161 ( .A1(n9350), .A2(n9352), .ZN(n9193) );
  NAND2_X1 U10162 ( .A1(n9192), .A2(n9191), .ZN(n9349) );
  NAND2_X1 U10163 ( .A1(n9193), .A2(n9349), .ZN(n9503) );
  NAND2_X1 U10164 ( .A1(n9197), .A2(n6725), .ZN(n9195) );
  NAND2_X1 U10165 ( .A1(n10758), .A2(n9309), .ZN(n9194) );
  NAND2_X1 U10166 ( .A1(n9195), .A2(n9194), .ZN(n9196) );
  XNOR2_X1 U10167 ( .A(n9196), .B(n9373), .ZN(n9505) );
  NAND2_X1 U10168 ( .A1(n9197), .A2(n9309), .ZN(n9199) );
  NAND2_X1 U10169 ( .A1(n10758), .A2(n9307), .ZN(n9198) );
  NAND2_X1 U10170 ( .A1(n10778), .A2(n6725), .ZN(n9201) );
  NAND2_X1 U10171 ( .A1(n9554), .A2(n9309), .ZN(n9200) );
  NAND2_X1 U10172 ( .A1(n9201), .A2(n9200), .ZN(n9202) );
  XNOR2_X1 U10173 ( .A(n9202), .B(n9373), .ZN(n9223) );
  AND2_X1 U10174 ( .A1(n9554), .A2(n9307), .ZN(n9203) );
  AOI21_X1 U10175 ( .B1(n10778), .B2(n4948), .A(n9203), .ZN(n9222) );
  XNOR2_X1 U10176 ( .A(n9223), .B(n9222), .ZN(n9411) );
  NAND2_X1 U10177 ( .A1(n9708), .A2(n6725), .ZN(n9205) );
  NAND2_X1 U10178 ( .A1(n9965), .A2(n9309), .ZN(n9204) );
  NAND2_X1 U10179 ( .A1(n9205), .A2(n9204), .ZN(n9206) );
  XNOR2_X1 U10180 ( .A(n9206), .B(n9373), .ZN(n9331) );
  AND2_X1 U10181 ( .A1(n9965), .A2(n9307), .ZN(n9207) );
  AOI21_X1 U10182 ( .B1(n9708), .B2(n9309), .A(n9207), .ZN(n9214) );
  NAND2_X1 U10183 ( .A1(n9331), .A2(n9214), .ZN(n9224) );
  INV_X1 U10184 ( .A(n9224), .ZN(n9218) );
  NAND2_X1 U10185 ( .A1(n9212), .A2(n6725), .ZN(n9209) );
  NAND2_X1 U10186 ( .A1(n10757), .A2(n9309), .ZN(n9208) );
  NAND2_X1 U10187 ( .A1(n9209), .A2(n9208), .ZN(n9210) );
  XNOR2_X1 U10188 ( .A(n9210), .B(n9314), .ZN(n9221) );
  AND2_X1 U10189 ( .A1(n10757), .A2(n9307), .ZN(n9211) );
  AOI21_X1 U10190 ( .B1(n9212), .B2(n9309), .A(n9211), .ZN(n9220) );
  INV_X1 U10191 ( .A(n9220), .ZN(n9213) );
  NAND2_X1 U10192 ( .A1(n9221), .A2(n9213), .ZN(n9329) );
  INV_X1 U10193 ( .A(n9331), .ZN(n9215) );
  INV_X1 U10194 ( .A(n9214), .ZN(n9330) );
  NAND2_X1 U10195 ( .A1(n9215), .A2(n9330), .ZN(n9216) );
  AND2_X1 U10196 ( .A1(n9329), .A2(n9216), .ZN(n9217) );
  NOR2_X1 U10197 ( .A1(n9218), .A2(n9217), .ZN(n9226) );
  OR2_X1 U10198 ( .A1(n9411), .A2(n9226), .ZN(n9219) );
  XNOR2_X1 U10199 ( .A(n9221), .B(n9220), .ZN(n9479) );
  NAND2_X1 U10200 ( .A1(n9223), .A2(n9222), .ZN(n9476) );
  AND2_X1 U10201 ( .A1(n9479), .A2(n9476), .ZN(n9328) );
  AND2_X1 U10202 ( .A1(n9328), .A2(n9224), .ZN(n9225) );
  NAND2_X1 U10203 ( .A1(n9971), .A2(n6725), .ZN(n9229) );
  NAND2_X1 U10204 ( .A1(n9553), .A2(n9309), .ZN(n9228) );
  NAND2_X1 U10205 ( .A1(n9229), .A2(n9228), .ZN(n9230) );
  XNOR2_X1 U10206 ( .A(n9230), .B(n9314), .ZN(n9536) );
  NAND2_X1 U10207 ( .A1(n9971), .A2(n9309), .ZN(n9232) );
  NAND2_X1 U10208 ( .A1(n9553), .A2(n9307), .ZN(n9231) );
  NAND2_X1 U10209 ( .A1(n9232), .A2(n9231), .ZN(n9537) );
  NAND2_X1 U10210 ( .A1(n9952), .A2(n6725), .ZN(n9234) );
  NAND2_X1 U10211 ( .A1(n9964), .A2(n4948), .ZN(n9233) );
  NAND2_X1 U10212 ( .A1(n9234), .A2(n9233), .ZN(n9235) );
  XNOR2_X1 U10213 ( .A(n9235), .B(n9373), .ZN(n9237) );
  AND2_X1 U10214 ( .A1(n9964), .A2(n9307), .ZN(n9236) );
  AOI21_X1 U10215 ( .B1(n9952), .B2(n9309), .A(n9236), .ZN(n9238) );
  NAND2_X1 U10216 ( .A1(n9237), .A2(n9238), .ZN(n9434) );
  INV_X1 U10217 ( .A(n9237), .ZN(n9240) );
  INV_X1 U10218 ( .A(n9238), .ZN(n9239) );
  NAND2_X1 U10219 ( .A1(n9240), .A2(n9239), .ZN(n9241) );
  NAND2_X1 U10220 ( .A1(n9434), .A2(n9241), .ZN(n9428) );
  NAND2_X1 U10221 ( .A1(n9932), .A2(n6725), .ZN(n9243) );
  NAND2_X1 U10222 ( .A1(n9911), .A2(n9309), .ZN(n9242) );
  NAND2_X1 U10223 ( .A1(n9243), .A2(n9242), .ZN(n9244) );
  XNOR2_X1 U10224 ( .A(n9244), .B(n9314), .ZN(n9251) );
  NAND2_X1 U10225 ( .A1(n9932), .A2(n4948), .ZN(n9246) );
  NAND2_X1 U10226 ( .A1(n9911), .A2(n9307), .ZN(n9245) );
  NAND2_X1 U10227 ( .A1(n9246), .A2(n9245), .ZN(n9252) );
  NAND2_X1 U10228 ( .A1(n9251), .A2(n9252), .ZN(n9437) );
  INV_X1 U10229 ( .A(n9437), .ZN(n9256) );
  OR2_X1 U10230 ( .A1(n9428), .A2(n9256), .ZN(n9261) );
  NAND2_X1 U10231 ( .A1(n9917), .A2(n6725), .ZN(n9248) );
  NAND2_X1 U10232 ( .A1(n9927), .A2(n4948), .ZN(n9247) );
  NAND2_X1 U10233 ( .A1(n9248), .A2(n9247), .ZN(n9249) );
  OR2_X1 U10234 ( .A1(n9261), .A2(n5562), .ZN(n9250) );
  INV_X1 U10235 ( .A(n9251), .ZN(n9254) );
  INV_X1 U10236 ( .A(n9252), .ZN(n9253) );
  NAND2_X1 U10237 ( .A1(n9254), .A2(n9253), .ZN(n9436) );
  AND2_X1 U10238 ( .A1(n9434), .A2(n9436), .ZN(n9255) );
  OR2_X1 U10239 ( .A1(n9256), .A2(n9255), .ZN(n9259) );
  OR2_X1 U10240 ( .A1(n5562), .A2(n9259), .ZN(n9257) );
  AND2_X1 U10241 ( .A1(n9259), .A2(n5562), .ZN(n9260) );
  OAI21_X1 U10242 ( .B1(n9426), .B2(n9261), .A(n9260), .ZN(n9516) );
  AND2_X1 U10243 ( .A1(n9927), .A2(n9307), .ZN(n9262) );
  AOI21_X1 U10244 ( .B1(n9917), .B2(n9309), .A(n9262), .ZN(n9518) );
  NAND2_X1 U10245 ( .A1(n9516), .A2(n9518), .ZN(n9263) );
  NAND2_X1 U10246 ( .A1(n9517), .A2(n9263), .ZN(n9363) );
  NAND2_X1 U10247 ( .A1(n9897), .A2(n6725), .ZN(n9265) );
  NAND2_X1 U10248 ( .A1(n9910), .A2(n6608), .ZN(n9264) );
  NAND2_X1 U10249 ( .A1(n9265), .A2(n9264), .ZN(n9266) );
  XNOR2_X1 U10250 ( .A(n9266), .B(n9314), .ZN(n9268) );
  AND2_X1 U10251 ( .A1(n9910), .A2(n9307), .ZN(n9267) );
  AOI21_X1 U10252 ( .B1(n9897), .B2(n9309), .A(n9267), .ZN(n9269) );
  XNOR2_X1 U10253 ( .A(n9268), .B(n9269), .ZN(n9364) );
  INV_X1 U10254 ( .A(n9268), .ZN(n9270) );
  NAND2_X1 U10255 ( .A1(n9270), .A2(n9269), .ZN(n9271) );
  NAND2_X1 U10256 ( .A1(n9881), .A2(n6725), .ZN(n9273) );
  NAND2_X1 U10257 ( .A1(n9893), .A2(n4948), .ZN(n9272) );
  NAND2_X1 U10258 ( .A1(n9273), .A2(n9272), .ZN(n9274) );
  XNOR2_X1 U10259 ( .A(n9274), .B(n9314), .ZN(n9276) );
  AND2_X1 U10260 ( .A1(n9893), .A2(n9307), .ZN(n9275) );
  AOI21_X1 U10261 ( .B1(n9881), .B2(n9309), .A(n9275), .ZN(n9277) );
  XNOR2_X1 U10262 ( .A(n9276), .B(n9277), .ZN(n9469) );
  INV_X1 U10263 ( .A(n9276), .ZN(n9278) );
  NAND2_X1 U10264 ( .A1(n9278), .A2(n9277), .ZN(n9279) );
  NAND2_X1 U10265 ( .A1(n10030), .A2(n6725), .ZN(n9281) );
  NAND2_X1 U10266 ( .A1(n9876), .A2(n6608), .ZN(n9280) );
  NAND2_X1 U10267 ( .A1(n9281), .A2(n9280), .ZN(n9282) );
  XNOR2_X1 U10268 ( .A(n9282), .B(n9314), .ZN(n9284) );
  AND2_X1 U10269 ( .A1(n9876), .A2(n9307), .ZN(n9283) );
  AOI21_X1 U10270 ( .B1(n10030), .B2(n9309), .A(n9283), .ZN(n9285) );
  XNOR2_X1 U10271 ( .A(n9284), .B(n9285), .ZN(n9403) );
  INV_X1 U10272 ( .A(n9284), .ZN(n9286) );
  NAND2_X1 U10273 ( .A1(n9286), .A2(n9285), .ZN(n9287) );
  NAND2_X1 U10274 ( .A1(n10024), .A2(n6725), .ZN(n9289) );
  NAND2_X1 U10275 ( .A1(n9826), .A2(n6608), .ZN(n9288) );
  NAND2_X1 U10276 ( .A1(n9289), .A2(n9288), .ZN(n9290) );
  XNOR2_X1 U10277 ( .A(n9290), .B(n9373), .ZN(n9291) );
  NAND2_X1 U10278 ( .A1(n9292), .A2(n9291), .ZN(n9494) );
  OAI22_X1 U10279 ( .A1(n9844), .A2(n9376), .B1(n9862), .B2(n9370), .ZN(n9492)
         );
  NAND2_X1 U10280 ( .A1(n9494), .A2(n9492), .ZN(n9490) );
  XNOR2_X1 U10281 ( .A(n9293), .B(n9294), .ZN(n9343) );
  NAND2_X1 U10282 ( .A1(n10015), .A2(n6725), .ZN(n9296) );
  NAND2_X1 U10283 ( .A1(n9825), .A2(n6608), .ZN(n9295) );
  NAND2_X1 U10284 ( .A1(n9296), .A2(n9295), .ZN(n9297) );
  XNOR2_X1 U10285 ( .A(n9297), .B(n9373), .ZN(n9300) );
  AND2_X1 U10286 ( .A1(n9825), .A2(n9307), .ZN(n9298) );
  AOI21_X1 U10287 ( .B1(n10015), .B2(n9309), .A(n9298), .ZN(n9299) );
  NOR2_X1 U10288 ( .A1(n9300), .A2(n9299), .ZN(n9447) );
  NAND2_X1 U10289 ( .A1(n9300), .A2(n9299), .ZN(n9445) );
  NAND2_X1 U10290 ( .A1(n9797), .A2(n6725), .ZN(n9302) );
  NAND2_X1 U10291 ( .A1(n9723), .A2(n6608), .ZN(n9301) );
  NAND2_X1 U10292 ( .A1(n9302), .A2(n9301), .ZN(n9303) );
  XNOR2_X1 U10293 ( .A(n9303), .B(n9314), .ZN(n9310) );
  AOI22_X1 U10294 ( .A1(n9797), .A2(n4948), .B1(n9307), .B2(n9723), .ZN(n9311)
         );
  XNOR2_X1 U10295 ( .A(n9310), .B(n9311), .ZN(n9420) );
  NAND2_X1 U10296 ( .A1(n9419), .A2(n9420), .ZN(n9527) );
  NAND2_X1 U10297 ( .A1(n10005), .A2(n6725), .ZN(n9305) );
  NAND2_X1 U10298 ( .A1(n9761), .A2(n6608), .ZN(n9304) );
  NAND2_X1 U10299 ( .A1(n9305), .A2(n9304), .ZN(n9306) );
  XNOR2_X1 U10300 ( .A(n9306), .B(n9314), .ZN(n9319) );
  AND2_X1 U10301 ( .A1(n9761), .A2(n9307), .ZN(n9308) );
  AOI21_X1 U10302 ( .B1(n10005), .B2(n9309), .A(n9308), .ZN(n9317) );
  XNOR2_X1 U10303 ( .A(n9319), .B(n9317), .ZN(n9530) );
  INV_X1 U10304 ( .A(n9310), .ZN(n9312) );
  NAND2_X1 U10305 ( .A1(n9312), .A2(n9311), .ZN(n9526) );
  AOI22_X1 U10306 ( .A1(n9765), .A2(n6725), .B1(n4948), .B2(n9552), .ZN(n9313)
         );
  XOR2_X1 U10307 ( .A(n9314), .B(n9313), .Z(n9316) );
  OAI22_X1 U10308 ( .A1(n10083), .A2(n9376), .B1(n9780), .B2(n9370), .ZN(n9315) );
  NOR2_X1 U10309 ( .A1(n9316), .A2(n9315), .ZN(n9384) );
  AOI21_X1 U10310 ( .B1(n9316), .B2(n9315), .A(n9384), .ZN(n9320) );
  INV_X1 U10311 ( .A(n9317), .ZN(n9318) );
  NAND2_X1 U10312 ( .A1(n9319), .A2(n9318), .ZN(n9321) );
  AOI21_X1 U10313 ( .B1(n9528), .B2(n9321), .A(n9320), .ZN(n9322) );
  OAI21_X1 U10314 ( .B1(n9379), .B2(n9322), .A(n9529), .ZN(n9326) );
  AOI22_X1 U10315 ( .A1(n9539), .A2(n9761), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n9323) );
  OAI21_X1 U10316 ( .B1(n9728), .B2(n9542), .A(n9323), .ZN(n9324) );
  AOI21_X1 U10317 ( .B1(n9766), .B2(n9546), .A(n9324), .ZN(n9325) );
  OAI211_X1 U10318 ( .C1(n10083), .C2(n9543), .A(n9326), .B(n9325), .ZN(
        P1_U3214) );
  OR2_X1 U10319 ( .A1(n9327), .A2(n9411), .ZN(n9477) );
  NAND2_X1 U10320 ( .A1(n9477), .A2(n9328), .ZN(n9478) );
  NAND2_X1 U10321 ( .A1(n9478), .A2(n9329), .ZN(n9333) );
  XNOR2_X1 U10322 ( .A(n9331), .B(n9330), .ZN(n9332) );
  XNOR2_X1 U10323 ( .A(n9333), .B(n9332), .ZN(n9341) );
  NAND2_X1 U10324 ( .A1(n9546), .A2(n9334), .ZN(n9338) );
  INV_X1 U10325 ( .A(n9335), .ZN(n9336) );
  AOI21_X1 U10326 ( .B1(n9539), .B2(n10757), .A(n9336), .ZN(n9337) );
  OAI211_X1 U10327 ( .C1(n9948), .C2(n9542), .A(n9338), .B(n9337), .ZN(n9339)
         );
  AOI21_X1 U10328 ( .B1(n9708), .B2(n9473), .A(n9339), .ZN(n9340) );
  OAI21_X1 U10329 ( .B1(n9341), .B2(n9548), .A(n9340), .ZN(P1_U3215) );
  AOI21_X1 U10330 ( .B1(n9343), .B2(n9489), .A(n9342), .ZN(n9348) );
  AOI22_X1 U10331 ( .A1(n9496), .A2(n9825), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9344) );
  OAI21_X1 U10332 ( .B1(n9862), .B2(n9498), .A(n9344), .ZN(n9346) );
  NOR2_X1 U10333 ( .A1(n10093), .A2(n9543), .ZN(n9345) );
  AOI211_X1 U10334 ( .C1(n9546), .C2(n9832), .A(n9346), .B(n9345), .ZN(n9347)
         );
  OAI21_X1 U10335 ( .B1(n9348), .B2(n9548), .A(n9347), .ZN(P1_U3216) );
  NAND2_X1 U10336 ( .A1(n9350), .A2(n9349), .ZN(n9351) );
  XOR2_X1 U10337 ( .A(n9352), .B(n9351), .Z(n9361) );
  NOR2_X1 U10338 ( .A1(n10729), .A2(n9543), .ZN(n9360) );
  INV_X1 U10339 ( .A(n9353), .ZN(n9354) );
  AOI21_X1 U10340 ( .B1(n9496), .B2(n10758), .A(n9354), .ZN(n9358) );
  NAND2_X1 U10341 ( .A1(n9546), .A2(n9355), .ZN(n9357) );
  NAND2_X1 U10342 ( .A1(n9539), .A2(n9556), .ZN(n9356) );
  NAND3_X1 U10343 ( .A1(n9358), .A2(n9357), .A3(n9356), .ZN(n9359) );
  AOI211_X1 U10344 ( .C1(n9361), .C2(n9529), .A(n9360), .B(n9359), .ZN(n9362)
         );
  INV_X1 U10345 ( .A(n9362), .ZN(P1_U3217) );
  XOR2_X1 U10346 ( .A(n9364), .B(n9363), .Z(n9369) );
  NAND2_X1 U10347 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9668) );
  NAND2_X1 U10348 ( .A1(n9539), .A2(n9927), .ZN(n9365) );
  OAI211_X1 U10349 ( .C1(n9861), .C2(n9542), .A(n9668), .B(n9365), .ZN(n9366)
         );
  AOI21_X1 U10350 ( .B1(n9898), .B2(n9546), .A(n9366), .ZN(n9368) );
  NAND2_X1 U10351 ( .A1(n9897), .A2(n9473), .ZN(n9367) );
  OAI211_X1 U10352 ( .C1(n9369), .C2(n9548), .A(n9368), .B(n9367), .ZN(
        P1_U3219) );
  NAND2_X1 U10353 ( .A1(n9995), .A2(n6608), .ZN(n9372) );
  OR2_X1 U10354 ( .A1(n9728), .A2(n9370), .ZN(n9371) );
  NAND2_X1 U10355 ( .A1(n9372), .A2(n9371), .ZN(n9374) );
  XNOR2_X1 U10356 ( .A(n9374), .B(n9373), .ZN(n9378) );
  NAND2_X1 U10357 ( .A1(n9995), .A2(n6725), .ZN(n9375) );
  OAI21_X1 U10358 ( .B1(n9728), .B2(n9376), .A(n9375), .ZN(n9377) );
  XNOR2_X1 U10359 ( .A(n9378), .B(n9377), .ZN(n9383) );
  OR4_X2 U10360 ( .A1(n9379), .A2(n9384), .A3(n9383), .A4(n9548), .ZN(n9388)
         );
  NAND3_X1 U10361 ( .A1(n9379), .A2(n9529), .A3(n9383), .ZN(n9387) );
  AOI22_X1 U10362 ( .A1(n9539), .A2(n9552), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9380) );
  OAI21_X1 U10363 ( .B1(n10369), .B2(n9542), .A(n9380), .ZN(n9382) );
  NOR2_X1 U10364 ( .A1(n9742), .A2(n9543), .ZN(n9381) );
  AOI211_X1 U10365 ( .C1(n9546), .C2(n9749), .A(n9382), .B(n9381), .ZN(n9386)
         );
  NAND3_X1 U10366 ( .A1(n9384), .A2(n9529), .A3(n9383), .ZN(n9385) );
  NAND4_X1 U10367 ( .A1(n9388), .A2(n9387), .A3(n9386), .A4(n9385), .ZN(
        P1_U3220) );
  NAND2_X1 U10368 ( .A1(n9390), .A2(n9389), .ZN(n9392) );
  XNOR2_X1 U10369 ( .A(n9392), .B(n9391), .ZN(n9401) );
  NOR2_X1 U10370 ( .A1(n9543), .A2(n10691), .ZN(n9400) );
  INV_X1 U10371 ( .A(n9393), .ZN(n9394) );
  AOI21_X1 U10372 ( .B1(n9496), .B2(n9556), .A(n9394), .ZN(n9398) );
  NAND2_X1 U10373 ( .A1(n9546), .A2(n9395), .ZN(n9397) );
  NAND2_X1 U10374 ( .A1(n9539), .A2(n9558), .ZN(n9396) );
  NAND3_X1 U10375 ( .A1(n9398), .A2(n9397), .A3(n9396), .ZN(n9399) );
  AOI211_X1 U10376 ( .C1(n9401), .C2(n9529), .A(n9400), .B(n9399), .ZN(n9402)
         );
  INV_X1 U10377 ( .A(n9402), .ZN(P1_U3221) );
  XOR2_X1 U10378 ( .A(n9404), .B(n9403), .Z(n9409) );
  AOI22_X1 U10379 ( .A1(n9496), .A2(n9826), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9405) );
  OAI21_X1 U10380 ( .B1(n9861), .B2(n9498), .A(n9405), .ZN(n9407) );
  INV_X1 U10381 ( .A(n10030), .ZN(n9868) );
  NOR2_X1 U10382 ( .A1(n9868), .A2(n9543), .ZN(n9406) );
  AOI211_X1 U10383 ( .C1(n9546), .C2(n9865), .A(n9407), .B(n9406), .ZN(n9408)
         );
  OAI21_X1 U10384 ( .B1(n9409), .B2(n9548), .A(n9408), .ZN(P1_U3223) );
  INV_X1 U10385 ( .A(n9477), .ZN(n9410) );
  AOI21_X1 U10386 ( .B1(n9411), .B2(n9327), .A(n9410), .ZN(n9418) );
  AOI21_X1 U10387 ( .B1(n9496), .B2(n10757), .A(n9412), .ZN(n9414) );
  NAND2_X1 U10388 ( .A1(n9546), .A2(n10776), .ZN(n9413) );
  OAI211_X1 U10389 ( .C1(n9415), .C2(n9498), .A(n9414), .B(n9413), .ZN(n9416)
         );
  AOI21_X1 U10390 ( .B1(n10778), .B2(n9473), .A(n9416), .ZN(n9417) );
  OAI21_X1 U10391 ( .B1(n9418), .B2(n9548), .A(n9417), .ZN(P1_U3224) );
  OAI21_X1 U10392 ( .B1(n9420), .B2(n9419), .A(n9527), .ZN(n9421) );
  NAND2_X1 U10393 ( .A1(n9421), .A2(n9529), .ZN(n9425) );
  AOI22_X1 U10394 ( .A1(n9496), .A2(n9761), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9422) );
  OAI21_X1 U10395 ( .B1(n9794), .B2(n9498), .A(n9422), .ZN(n9423) );
  AOI21_X1 U10396 ( .B1(n9798), .B2(n9546), .A(n9423), .ZN(n9424) );
  OAI211_X1 U10397 ( .C1(n10088), .C2(n9543), .A(n9425), .B(n9424), .ZN(
        P1_U3225) );
  OR2_X1 U10398 ( .A1(n9426), .A2(n9428), .ZN(n9435) );
  INV_X1 U10399 ( .A(n9435), .ZN(n9427) );
  AOI21_X1 U10400 ( .B1(n9428), .B2(n9426), .A(n9427), .ZN(n9433) );
  AND2_X1 U10401 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9614) );
  AOI21_X1 U10402 ( .B1(n9496), .B2(n9911), .A(n9614), .ZN(n9430) );
  NAND2_X1 U10403 ( .A1(n9546), .A2(n9953), .ZN(n9429) );
  OAI211_X1 U10404 ( .C1(n9948), .C2(n9498), .A(n9430), .B(n9429), .ZN(n9431)
         );
  AOI21_X1 U10405 ( .B1(n9952), .B2(n9473), .A(n9431), .ZN(n9432) );
  OAI21_X1 U10406 ( .B1(n9433), .B2(n9548), .A(n9432), .ZN(P1_U3226) );
  NAND2_X1 U10407 ( .A1(n9435), .A2(n9434), .ZN(n9439) );
  NAND2_X1 U10408 ( .A1(n9437), .A2(n9436), .ZN(n9438) );
  XNOR2_X1 U10409 ( .A(n9439), .B(n9438), .ZN(n9444) );
  NAND2_X1 U10410 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9631) );
  NAND2_X1 U10411 ( .A1(n9539), .A2(n9964), .ZN(n9440) );
  OAI211_X1 U10412 ( .C1(n9714), .C2(n9542), .A(n9631), .B(n9440), .ZN(n9442)
         );
  NOR2_X1 U10413 ( .A1(n10110), .A2(n9543), .ZN(n9441) );
  AOI211_X1 U10414 ( .C1(n9546), .C2(n9933), .A(n9442), .B(n9441), .ZN(n9443)
         );
  OAI21_X1 U10415 ( .B1(n9444), .B2(n9548), .A(n9443), .ZN(P1_U3228) );
  INV_X1 U10416 ( .A(n9445), .ZN(n9446) );
  NOR2_X1 U10417 ( .A1(n9447), .A2(n9446), .ZN(n9448) );
  XNOR2_X1 U10418 ( .A(n9449), .B(n9448), .ZN(n9454) );
  AOI22_X1 U10419 ( .A1(n9496), .A2(n9723), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9450) );
  OAI21_X1 U10420 ( .B1(n9847), .B2(n9498), .A(n9450), .ZN(n9452) );
  NOR2_X1 U10421 ( .A1(n9815), .A2(n9543), .ZN(n9451) );
  AOI211_X1 U10422 ( .C1(n9546), .C2(n9812), .A(n9452), .B(n9451), .ZN(n9453)
         );
  OAI21_X1 U10423 ( .B1(n9454), .B2(n9548), .A(n9453), .ZN(P1_U3229) );
  NAND2_X1 U10424 ( .A1(n9455), .A2(n9389), .ZN(n9457) );
  AOI21_X1 U10425 ( .B1(n9458), .B2(n9457), .A(n9456), .ZN(n9467) );
  NAND2_X1 U10426 ( .A1(n9546), .A2(n9459), .ZN(n9462) );
  AOI21_X1 U10427 ( .B1(n9496), .B2(n9555), .A(n9460), .ZN(n9461) );
  OAI211_X1 U10428 ( .C1(n9463), .C2(n9498), .A(n9462), .B(n9461), .ZN(n9464)
         );
  AOI21_X1 U10429 ( .B1(n9465), .B2(n9473), .A(n9464), .ZN(n9466) );
  OAI21_X1 U10430 ( .B1(n9467), .B2(n9548), .A(n9466), .ZN(P1_U3231) );
  XOR2_X1 U10431 ( .A(n9468), .B(n9469), .Z(n9475) );
  AOI22_X1 U10432 ( .A1(n9496), .A2(n9876), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9471) );
  NAND2_X1 U10433 ( .A1(n9546), .A2(n9882), .ZN(n9470) );
  OAI211_X1 U10434 ( .C1(n9521), .C2(n9498), .A(n9471), .B(n9470), .ZN(n9472)
         );
  AOI21_X1 U10435 ( .B1(n9881), .B2(n9473), .A(n9472), .ZN(n9474) );
  OAI21_X1 U10436 ( .B1(n9475), .B2(n9548), .A(n9474), .ZN(P1_U3233) );
  AND2_X1 U10437 ( .A1(n9477), .A2(n9476), .ZN(n9480) );
  OAI211_X1 U10438 ( .C1(n9480), .C2(n9479), .A(n9529), .B(n9478), .ZN(n9487)
         );
  INV_X1 U10439 ( .A(n9481), .ZN(n9482) );
  AOI21_X1 U10440 ( .B1(n9539), .B2(n9554), .A(n9482), .ZN(n9483) );
  OAI21_X1 U10441 ( .B1(n9707), .B2(n9542), .A(n9483), .ZN(n9484) );
  AOI21_X1 U10442 ( .B1(n9485), .B2(n9546), .A(n9484), .ZN(n9486) );
  OAI211_X1 U10443 ( .C1(n9488), .C2(n9543), .A(n9487), .B(n9486), .ZN(
        P1_U3234) );
  INV_X1 U10444 ( .A(n9489), .ZN(n9495) );
  INV_X1 U10445 ( .A(n9490), .ZN(n9491) );
  NAND2_X1 U10446 ( .A1(n9491), .A2(n5563), .ZN(n9493) );
  AOI22_X1 U10447 ( .A1(n9495), .A2(n9494), .B1(n9493), .B2(n9492), .ZN(n9502)
         );
  AOI22_X1 U10448 ( .A1(n9496), .A2(n9722), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9497) );
  OAI21_X1 U10449 ( .B1(n9848), .B2(n9498), .A(n9497), .ZN(n9500) );
  NOR2_X1 U10450 ( .A1(n9844), .A2(n9543), .ZN(n9499) );
  AOI211_X1 U10451 ( .C1(n9546), .C2(n9842), .A(n9500), .B(n9499), .ZN(n9501)
         );
  OAI21_X1 U10452 ( .B1(n9502), .B2(n9548), .A(n9501), .ZN(P1_U3235) );
  XNOR2_X1 U10453 ( .A(n9505), .B(n9504), .ZN(n9506) );
  XNOR2_X1 U10454 ( .A(n9503), .B(n9506), .ZN(n9515) );
  NAND2_X1 U10455 ( .A1(n9539), .A2(n9555), .ZN(n9507) );
  OAI211_X1 U10456 ( .C1(n9509), .C2(n9542), .A(n9508), .B(n9507), .ZN(n9512)
         );
  NOR2_X1 U10457 ( .A1(n9510), .A2(n9543), .ZN(n9511) );
  AOI211_X1 U10458 ( .C1(n9546), .C2(n9513), .A(n9512), .B(n9511), .ZN(n9514)
         );
  OAI21_X1 U10459 ( .B1(n9515), .B2(n9548), .A(n9514), .ZN(P1_U3236) );
  NAND2_X1 U10460 ( .A1(n9516), .A2(n9517), .ZN(n9519) );
  XNOR2_X1 U10461 ( .A(n9519), .B(n9518), .ZN(n9525) );
  NAND2_X1 U10462 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9647) );
  NAND2_X1 U10463 ( .A1(n9539), .A2(n9911), .ZN(n9520) );
  OAI211_X1 U10464 ( .C1(n9521), .C2(n9542), .A(n9647), .B(n9520), .ZN(n9523)
         );
  NOR2_X1 U10465 ( .A1(n10106), .A2(n9543), .ZN(n9522) );
  AOI211_X1 U10466 ( .C1(n9546), .C2(n9918), .A(n9523), .B(n9522), .ZN(n9524)
         );
  OAI21_X1 U10467 ( .B1(n9525), .B2(n9548), .A(n9524), .ZN(P1_U3238) );
  AND2_X1 U10468 ( .A1(n9527), .A2(n9526), .ZN(n9531) );
  OAI211_X1 U10469 ( .C1(n9531), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9535)
         );
  AOI22_X1 U10470 ( .A1(n9539), .A2(n9723), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9532) );
  OAI21_X1 U10471 ( .B1(n9780), .B2(n9542), .A(n9532), .ZN(n9533) );
  AOI21_X1 U10472 ( .B1(n9784), .B2(n9546), .A(n9533), .ZN(n9534) );
  OAI211_X1 U10473 ( .C1(n9787), .C2(n9543), .A(n9535), .B(n9534), .ZN(
        P1_U3240) );
  XOR2_X1 U10474 ( .A(n9537), .B(n9536), .Z(n9538) );
  XNOR2_X1 U10475 ( .A(n5030), .B(n9538), .ZN(n9549) );
  NAND2_X1 U10476 ( .A1(n9539), .A2(n9965), .ZN(n9541) );
  OAI211_X1 U10477 ( .C1(n9712), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9545)
         );
  NOR2_X1 U10478 ( .A1(n10118), .A2(n9543), .ZN(n9544) );
  AOI211_X1 U10479 ( .C1(n9546), .C2(n9973), .A(n9545), .B(n9544), .ZN(n9547)
         );
  OAI21_X1 U10480 ( .B1(n9549), .B2(n9548), .A(n9547), .ZN(P1_U3241) );
  MUX2_X1 U10481 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9550), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10482 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9551), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10483 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n5550), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10484 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9552), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10485 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9761), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10486 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9723), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10487 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9825), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10488 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9722), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10489 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9826), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10490 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9876), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10491 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9893), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10492 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9910), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10493 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9927), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10494 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9911), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10495 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9964), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10496 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9553), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10497 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9965), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10498 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n10757), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10499 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9554), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10500 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n10758), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10501 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9555), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10502 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9556), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10503 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9557), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10504 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9558), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10505 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9559), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10506 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9560), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10507 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9561), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10508 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9562), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10509 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9563), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10510 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9564), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10511 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6799), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U10512 ( .C1(n9567), .C2(n9566), .A(n9644), .B(n9565), .ZN(n9574)
         );
  AOI22_X1 U10513 ( .A1(n10532), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9573) );
  NAND2_X1 U10514 ( .A1(n10542), .A2(n9568), .ZN(n9572) );
  OAI211_X1 U10515 ( .C1(n9570), .C2(n9578), .A(n10538), .B(n9569), .ZN(n9571)
         );
  NAND4_X1 U10516 ( .A1(n9574), .A2(n9573), .A3(n9572), .A4(n9571), .ZN(
        P1_U3244) );
  INV_X1 U10517 ( .A(n9575), .ZN(n9582) );
  AOI21_X1 U10518 ( .B1(n9576), .B2(P1_REG2_REG_0__SCAN_IN), .A(
        P1_IR_REG_0__SCAN_IN), .ZN(n9579) );
  NAND2_X1 U10519 ( .A1(n10135), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9577) );
  OAI211_X1 U10520 ( .C1(n9579), .C2(n9578), .A(n9581), .B(n9577), .ZN(n9580)
         );
  OAI211_X1 U10521 ( .C1(n9582), .C2(n9581), .A(P1_U3973), .B(n9580), .ZN(
        n10548) );
  INV_X1 U10522 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9584) );
  INV_X1 U10523 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9583) );
  OAI22_X1 U10524 ( .A1(n9669), .A2(n9584), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9583), .ZN(n9585) );
  AOI21_X1 U10525 ( .B1(n10542), .B2(n9586), .A(n9585), .ZN(n9595) );
  OAI211_X1 U10526 ( .C1(n9589), .C2(n9588), .A(n10538), .B(n9587), .ZN(n9594)
         );
  OAI211_X1 U10527 ( .C1(n9592), .C2(n9591), .A(n9644), .B(n9590), .ZN(n9593)
         );
  NAND4_X1 U10528 ( .A1(n10548), .A2(n9595), .A3(n9594), .A4(n9593), .ZN(
        P1_U3245) );
  INV_X1 U10529 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9597) );
  OAI21_X1 U10530 ( .B1(n9669), .B2(n9597), .A(n9596), .ZN(n9598) );
  AOI21_X1 U10531 ( .B1(n10542), .B2(n9599), .A(n9598), .ZN(n9608) );
  OAI211_X1 U10532 ( .C1(n9602), .C2(n9601), .A(n9644), .B(n9600), .ZN(n9607)
         );
  OAI211_X1 U10533 ( .C1(n9605), .C2(n9604), .A(n10538), .B(n9603), .ZN(n9606)
         );
  NAND3_X1 U10534 ( .A1(n9608), .A2(n9607), .A3(n9606), .ZN(P1_U3246) );
  NOR2_X1 U10535 ( .A1(n9609), .A2(n9618), .ZN(n9611) );
  NOR2_X1 U10536 ( .A1(n9611), .A2(n9610), .ZN(n9613) );
  INV_X1 U10537 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10057) );
  AOI22_X1 U10538 ( .A1(n9636), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n10057), 
        .B2(n9616), .ZN(n9612) );
  NAND2_X1 U10539 ( .A1(n9612), .A2(n9613), .ZN(n9630) );
  OAI21_X1 U10540 ( .B1(n9613), .B2(n9612), .A(n9630), .ZN(n9628) );
  AOI21_X1 U10541 ( .B1(n10532), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9614), .ZN(
        n9615) );
  OAI21_X1 U10542 ( .B1(n9617), .B2(n9616), .A(n9615), .ZN(n9627) );
  NOR2_X1 U10543 ( .A1(n9619), .A2(n9618), .ZN(n9621) );
  NOR2_X1 U10544 ( .A1(n9621), .A2(n9620), .ZN(n9625) );
  NAND2_X1 U10545 ( .A1(n9636), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9622) );
  OAI21_X1 U10546 ( .B1(n9636), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9622), .ZN(
        n9624) );
  NOR2_X1 U10547 ( .A1(n9625), .A2(n9624), .ZN(n9635) );
  AOI211_X1 U10548 ( .C1(n9625), .C2(n9624), .A(n9635), .B(n9623), .ZN(n9626)
         );
  AOI211_X1 U10549 ( .C1(n9644), .C2(n9628), .A(n9627), .B(n9626), .ZN(n9629)
         );
  INV_X1 U10550 ( .A(n9629), .ZN(P1_U3259) );
  INV_X1 U10551 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10051) );
  XNOR2_X1 U10552 ( .A(n9634), .B(n10051), .ZN(n9641) );
  OAI21_X1 U10553 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9636), .A(n9630), .ZN(
        n9642) );
  XOR2_X1 U10554 ( .A(n9641), .B(n9642), .Z(n9640) );
  OAI21_X1 U10555 ( .B1(n9669), .B2(n9632), .A(n9631), .ZN(n9633) );
  AOI21_X1 U10556 ( .B1(n10542), .B2(n9634), .A(n9633), .ZN(n9639) );
  INV_X1 U10557 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9653) );
  XNOR2_X1 U10558 ( .A(n9634), .B(n9653), .ZN(n9652) );
  AOI21_X1 U10559 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9636), .A(n9635), .ZN(
        n9651) );
  XNOR2_X1 U10560 ( .A(n9652), .B(n9651), .ZN(n9637) );
  NAND2_X1 U10561 ( .A1(n10538), .A2(n9637), .ZN(n9638) );
  OAI211_X1 U10562 ( .C1(n9640), .C2(n10546), .A(n9639), .B(n9638), .ZN(
        P1_U3260) );
  AOI22_X1 U10563 ( .A1(n9642), .A2(n9641), .B1(n10051), .B2(n9654), .ZN(n9646) );
  INV_X1 U10564 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10046) );
  AND2_X1 U10565 ( .A1(n9650), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9663) );
  AOI21_X1 U10566 ( .B1(n10046), .B2(n9643), .A(n9663), .ZN(n9645) );
  NAND2_X1 U10567 ( .A1(n9646), .A2(n9645), .ZN(n9665) );
  OAI211_X1 U10568 ( .C1(n9646), .C2(n9645), .A(n9665), .B(n9644), .ZN(n9662)
         );
  INV_X1 U10569 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9648) );
  OAI21_X1 U10570 ( .B1(n9669), .B2(n9648), .A(n9647), .ZN(n9649) );
  AOI21_X1 U10571 ( .B1(n10542), .B2(n9650), .A(n9649), .ZN(n9661) );
  NAND2_X1 U10572 ( .A1(n9650), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9672) );
  OAI21_X1 U10573 ( .B1(n9650), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9672), .ZN(
        n9658) );
  NAND2_X1 U10574 ( .A1(n9652), .A2(n9651), .ZN(n9656) );
  NAND2_X1 U10575 ( .A1(n9654), .A2(n9653), .ZN(n9655) );
  NAND2_X1 U10576 ( .A1(n9656), .A2(n9655), .ZN(n9657) );
  NAND2_X1 U10577 ( .A1(n9658), .A2(n9657), .ZN(n9659) );
  NAND3_X1 U10578 ( .A1(n10538), .A2(n9673), .A3(n9659), .ZN(n9660) );
  NAND3_X1 U10579 ( .A1(n9662), .A2(n9661), .A3(n9660), .ZN(P1_U3261) );
  INV_X1 U10580 ( .A(n9663), .ZN(n9664) );
  NAND2_X1 U10581 ( .A1(n9665), .A2(n9664), .ZN(n9667) );
  XNOR2_X1 U10582 ( .A(n9674), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9666) );
  XNOR2_X1 U10583 ( .A(n9667), .B(n9666), .ZN(n9681) );
  OAI21_X1 U10584 ( .B1(n9669), .B2(n5246), .A(n9668), .ZN(n9670) );
  AOI21_X1 U10585 ( .B1(n10542), .B2(n9671), .A(n9670), .ZN(n9680) );
  NAND2_X1 U10586 ( .A1(n9673), .A2(n9672), .ZN(n9677) );
  INV_X1 U10587 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9675) );
  MUX2_X1 U10588 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9675), .S(n9674), .Z(n9676) );
  XNOR2_X1 U10589 ( .A(n9677), .B(n9676), .ZN(n9678) );
  NAND2_X1 U10590 ( .A1(n10538), .A2(n9678), .ZN(n9679) );
  OAI211_X1 U10591 ( .C1(n9681), .C2(n10546), .A(n9680), .B(n9679), .ZN(
        P1_U3262) );
  OR2_X2 U10592 ( .A1(n9970), .A2(n9971), .ZN(n9968) );
  NAND2_X1 U10593 ( .A1(n9863), .A2(n9844), .ZN(n9839) );
  NAND2_X1 U10594 ( .A1(n10077), .A2(n9731), .ZN(n9689) );
  XNOR2_X1 U10595 ( .A(n9689), .B(n9682), .ZN(n9683) );
  NAND2_X1 U10596 ( .A1(n9982), .A2(n9972), .ZN(n9688) );
  AND2_X1 U10597 ( .A1(n9684), .A2(P1_B_REG_SCAN_IN), .ZN(n9685) );
  OR2_X1 U10598 ( .A1(n10551), .A2(n9685), .ZN(n9706) );
  NOR2_X1 U10599 ( .A1(n9686), .A2(n9706), .ZN(n9981) );
  INV_X1 U10600 ( .A(n9981), .ZN(n9985) );
  NOR2_X1 U10601 ( .A1(n9985), .A2(n10786), .ZN(n9691) );
  AOI21_X1 U10602 ( .B1(n10786), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9691), .ZN(
        n9687) );
  OAI211_X1 U10603 ( .C1(n10073), .C2(n9976), .A(n9688), .B(n9687), .ZN(
        P1_U3263) );
  OAI211_X1 U10604 ( .C1(n10077), .C2(n9731), .A(n10762), .B(n9689), .ZN(n9986) );
  NOR2_X1 U10605 ( .A1(n10077), .A2(n9976), .ZN(n9690) );
  AOI211_X1 U10606 ( .C1(n10786), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9691), .B(
        n9690), .ZN(n9692) );
  OAI21_X1 U10607 ( .B1(n10658), .B2(n9986), .A(n9692), .ZN(P1_U3264) );
  NAND2_X1 U10608 ( .A1(n9694), .A2(n9693), .ZN(n9846) );
  NOR2_X1 U10609 ( .A1(n9820), .A2(n9695), .ZN(n9696) );
  INV_X1 U10610 ( .A(n9805), .ZN(n9697) );
  NOR2_X1 U10611 ( .A1(n9806), .A2(n9697), .ZN(n9698) );
  NAND2_X1 U10612 ( .A1(n9792), .A2(n9791), .ZN(n9774) );
  NOR2_X1 U10613 ( .A1(n9778), .A2(n9700), .ZN(n9701) );
  INV_X1 U10614 ( .A(n9754), .ZN(n9757) );
  NOR2_X1 U10615 ( .A1(n9757), .A2(n5175), .ZN(n9702) );
  NAND2_X1 U10616 ( .A1(n9743), .A2(n9703), .ZN(n9704) );
  NAND2_X1 U10617 ( .A1(n10123), .A2(n9707), .ZN(n9710) );
  AOI21_X1 U10618 ( .B1(n9711), .B2(n9710), .A(n9709), .ZN(n9958) );
  AOI22_X1 U10619 ( .A1(n9958), .A2(n9960), .B1(n9948), .B2(n10118), .ZN(n9941) );
  NAND2_X1 U10620 ( .A1(n9941), .A2(n9940), .ZN(n9939) );
  NOR2_X1 U10621 ( .A1(n10110), .A2(n9950), .ZN(n9713) );
  NOR2_X1 U10622 ( .A1(n9917), .A2(n9927), .ZN(n9715) );
  NAND2_X1 U10623 ( .A1(n9871), .A2(n9873), .ZN(n9719) );
  NAND2_X1 U10624 ( .A1(n9719), .A2(n9718), .ZN(n9856) );
  NAND2_X1 U10625 ( .A1(n9856), .A2(n9858), .ZN(n9720) );
  NAND2_X1 U10626 ( .A1(n10093), .A2(n9847), .ZN(n9721) );
  NOR2_X1 U10627 ( .A1(n9797), .A2(n9723), .ZN(n9724) );
  OAI22_X1 U10628 ( .A1(n9790), .A2(n9724), .B1(n9809), .B2(n10088), .ZN(n9772) );
  NAND2_X1 U10629 ( .A1(n9772), .A2(n9778), .ZN(n9726) );
  NAND2_X1 U10630 ( .A1(n10005), .A2(n9761), .ZN(n9725) );
  NAND2_X1 U10631 ( .A1(n10083), .A2(n9780), .ZN(n9727) );
  XNOR2_X1 U10632 ( .A(n9730), .B(n9729), .ZN(n9989) );
  NAND2_X1 U10633 ( .A1(n9989), .A2(n10781), .ZN(n9736) );
  AOI211_X1 U10634 ( .C1(n9991), .C2(n9738), .A(n9915), .B(n9731), .ZN(n9990)
         );
  AOI22_X1 U10635 ( .A1(n10786), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9732), 
        .B2(n10775), .ZN(n9733) );
  OAI21_X1 U10636 ( .B1(n5123), .B2(n9976), .A(n9733), .ZN(n9734) );
  AOI21_X1 U10637 ( .B1(n9990), .B2(n9972), .A(n9734), .ZN(n9735) );
  OAI211_X1 U10638 ( .C1(n5002), .C2(n10786), .A(n9736), .B(n9735), .ZN(
        P1_U3356) );
  OAI21_X1 U10639 ( .B1(n4977), .B2(n5551), .A(n9737), .ZN(n9997) );
  INV_X1 U10640 ( .A(n9738), .ZN(n9739) );
  AOI211_X1 U10641 ( .C1(n9995), .C2(n9740), .A(n9915), .B(n9739), .ZN(n9994)
         );
  INV_X1 U10642 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9741) );
  OAI22_X1 U10643 ( .A1(n9742), .A2(n9976), .B1(n10560), .B2(n9741), .ZN(n9752) );
  INV_X1 U10644 ( .A(n9743), .ZN(n9747) );
  AOI21_X1 U10645 ( .B1(n9759), .B2(n9745), .A(n9744), .ZN(n9746) );
  OAI222_X1 U10646 ( .A1(n10551), .A2(n10369), .B1(n9949), .B2(n9780), .C1(
        n10563), .C2(n9748), .ZN(n9993) );
  AOI21_X1 U10647 ( .B1(n9749), .B2(n10775), .A(n9993), .ZN(n9750) );
  NOR2_X1 U10648 ( .A1(n9750), .A2(n10786), .ZN(n9751) );
  OAI21_X1 U10649 ( .B1(n9997), .B2(n9979), .A(n9753), .ZN(P1_U3265) );
  XNOR2_X1 U10650 ( .A(n9755), .B(n9754), .ZN(n10000) );
  INV_X1 U10651 ( .A(n10000), .ZN(n9771) );
  NAND2_X1 U10652 ( .A1(n9775), .A2(n9756), .ZN(n9758) );
  NAND2_X1 U10653 ( .A1(n9758), .A2(n9757), .ZN(n9760) );
  NAND3_X1 U10654 ( .A1(n9760), .A2(n10752), .A3(n9759), .ZN(n9763) );
  AOI22_X1 U10655 ( .A1(n5550), .A2(n10756), .B1(n10759), .B2(n9761), .ZN(
        n9762) );
  NAND2_X1 U10656 ( .A1(n9763), .A2(n9762), .ZN(n9998) );
  AOI211_X1 U10657 ( .C1(n9765), .C2(n9781), .A(n9915), .B(n9764), .ZN(n9999)
         );
  NAND2_X1 U10658 ( .A1(n9999), .A2(n9972), .ZN(n9768) );
  AOI22_X1 U10659 ( .A1(n10786), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9766), 
        .B2(n10775), .ZN(n9767) );
  OAI211_X1 U10660 ( .C1(n10083), .C2(n9976), .A(n9768), .B(n9767), .ZN(n9769)
         );
  AOI21_X1 U10661 ( .B1(n9998), .B2(n10560), .A(n9769), .ZN(n9770) );
  OAI21_X1 U10662 ( .B1(n9771), .B2(n9979), .A(n9770), .ZN(P1_U3266) );
  XNOR2_X1 U10663 ( .A(n9772), .B(n9778), .ZN(n10007) );
  NAND2_X1 U10664 ( .A1(n9774), .A2(n9773), .ZN(n9777) );
  INV_X1 U10665 ( .A(n9775), .ZN(n9776) );
  AOI21_X1 U10666 ( .B1(n9778), .B2(n9777), .A(n9776), .ZN(n9779) );
  OAI222_X1 U10667 ( .A1(n10551), .A2(n9780), .B1(n9949), .B2(n9809), .C1(
        n10563), .C2(n9779), .ZN(n10003) );
  INV_X1 U10668 ( .A(n9796), .ZN(n9783) );
  INV_X1 U10669 ( .A(n9781), .ZN(n9782) );
  AOI211_X1 U10670 ( .C1(n10005), .C2(n9783), .A(n9915), .B(n9782), .ZN(n10004) );
  NAND2_X1 U10671 ( .A1(n10004), .A2(n9972), .ZN(n9786) );
  AOI22_X1 U10672 ( .A1(n10786), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9784), 
        .B2(n10775), .ZN(n9785) );
  OAI211_X1 U10673 ( .C1(n9787), .C2(n9976), .A(n9786), .B(n9785), .ZN(n9788)
         );
  AOI21_X1 U10674 ( .B1(n10003), .B2(n10560), .A(n9788), .ZN(n9789) );
  OAI21_X1 U10675 ( .B1(n10007), .B2(n9979), .A(n9789), .ZN(P1_U3267) );
  XOR2_X1 U10676 ( .A(n9791), .B(n9790), .Z(n10010) );
  INV_X1 U10677 ( .A(n10010), .ZN(n9803) );
  XNOR2_X1 U10678 ( .A(n9792), .B(n9791), .ZN(n9793) );
  OAI222_X1 U10679 ( .A1(n10551), .A2(n9795), .B1(n9949), .B2(n9794), .C1(
        n10563), .C2(n9793), .ZN(n10008) );
  AOI211_X1 U10680 ( .C1(n9797), .C2(n9810), .A(n9915), .B(n9796), .ZN(n10009)
         );
  NAND2_X1 U10681 ( .A1(n10009), .A2(n9972), .ZN(n9800) );
  AOI22_X1 U10682 ( .A1(n10786), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9798), 
        .B2(n10775), .ZN(n9799) );
  OAI211_X1 U10683 ( .C1(n10088), .C2(n9976), .A(n9800), .B(n9799), .ZN(n9801)
         );
  AOI21_X1 U10684 ( .B1(n10008), .B2(n10560), .A(n9801), .ZN(n9802) );
  OAI21_X1 U10685 ( .B1(n9803), .B2(n9979), .A(n9802), .ZN(P1_U3268) );
  XNOR2_X1 U10686 ( .A(n9804), .B(n9806), .ZN(n10017) );
  NAND2_X1 U10687 ( .A1(n9822), .A2(n9805), .ZN(n9807) );
  XNOR2_X1 U10688 ( .A(n9807), .B(n9806), .ZN(n9808) );
  OAI222_X1 U10689 ( .A1(n10551), .A2(n9809), .B1(n9949), .B2(n9847), .C1(
        n9808), .C2(n10563), .ZN(n10013) );
  INV_X1 U10690 ( .A(n9810), .ZN(n9811) );
  AOI211_X1 U10691 ( .C1(n10015), .C2(n9829), .A(n9915), .B(n9811), .ZN(n10014) );
  NAND2_X1 U10692 ( .A1(n10014), .A2(n9972), .ZN(n9814) );
  AOI22_X1 U10693 ( .A1(n10786), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9812), 
        .B2(n10775), .ZN(n9813) );
  OAI211_X1 U10694 ( .C1(n9815), .C2(n9976), .A(n9814), .B(n9813), .ZN(n9816)
         );
  AOI21_X1 U10695 ( .B1(n10013), .B2(n10560), .A(n9816), .ZN(n9817) );
  OAI21_X1 U10696 ( .B1(n10017), .B2(n9979), .A(n9817), .ZN(P1_U3269) );
  XOR2_X1 U10697 ( .A(n9820), .B(n9818), .Z(n10020) );
  INV_X1 U10698 ( .A(n10020), .ZN(n9837) );
  NAND2_X1 U10699 ( .A1(n9850), .A2(n9819), .ZN(n9821) );
  NAND2_X1 U10700 ( .A1(n9821), .A2(n9820), .ZN(n9823) );
  NAND2_X1 U10701 ( .A1(n9823), .A2(n9822), .ZN(n9824) );
  NAND2_X1 U10702 ( .A1(n9824), .A2(n10752), .ZN(n9828) );
  AOI22_X1 U10703 ( .A1(n10759), .A2(n9826), .B1(n9825), .B2(n10756), .ZN(
        n9827) );
  NAND2_X1 U10704 ( .A1(n9828), .A2(n9827), .ZN(n10018) );
  INV_X1 U10705 ( .A(n9829), .ZN(n9830) );
  AOI211_X1 U10706 ( .C1(n9831), .C2(n9839), .A(n9915), .B(n9830), .ZN(n10019)
         );
  NAND2_X1 U10707 ( .A1(n10019), .A2(n9972), .ZN(n9834) );
  AOI22_X1 U10708 ( .A1(n10786), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9832), 
        .B2(n10775), .ZN(n9833) );
  OAI211_X1 U10709 ( .C1(n10093), .C2(n9976), .A(n9834), .B(n9833), .ZN(n9835)
         );
  AOI21_X1 U10710 ( .B1(n10018), .B2(n10560), .A(n9835), .ZN(n9836) );
  OAI21_X1 U10711 ( .B1(n9837), .B2(n9979), .A(n9836), .ZN(P1_U3270) );
  XNOR2_X1 U10712 ( .A(n9838), .B(n5506), .ZN(n10027) );
  INV_X1 U10713 ( .A(n9863), .ZN(n9841) );
  INV_X1 U10714 ( .A(n9839), .ZN(n9840) );
  AOI211_X1 U10715 ( .C1(n10024), .C2(n9841), .A(n9915), .B(n9840), .ZN(n10023) );
  AOI22_X1 U10716 ( .A1(n10786), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9842), 
        .B2(n10775), .ZN(n9843) );
  OAI21_X1 U10717 ( .B1(n9844), .B2(n9976), .A(n9843), .ZN(n9853) );
  AOI21_X1 U10718 ( .B1(n9846), .B2(n9845), .A(n10563), .ZN(n9851) );
  OAI22_X1 U10719 ( .A1(n9848), .A2(n9949), .B1(n9847), .B2(n10551), .ZN(n9849) );
  AOI21_X1 U10720 ( .B1(n9851), .B2(n9850), .A(n9849), .ZN(n10026) );
  NOR2_X1 U10721 ( .A1(n10026), .A2(n10786), .ZN(n9852) );
  AOI211_X1 U10722 ( .C1(n10023), .C2(n9972), .A(n9853), .B(n9852), .ZN(n9854)
         );
  OAI21_X1 U10723 ( .B1(n10027), .B2(n9979), .A(n9854), .ZN(P1_U3271) );
  XNOR2_X1 U10724 ( .A(n9856), .B(n9855), .ZN(n10032) );
  AOI21_X1 U10725 ( .B1(n9874), .B2(n9872), .A(n9873), .ZN(n9879) );
  NOR2_X1 U10726 ( .A1(n9879), .A2(n5199), .ZN(n9859) );
  XNOR2_X1 U10727 ( .A(n9859), .B(n9858), .ZN(n9860) );
  OAI222_X1 U10728 ( .A1(n10551), .A2(n9862), .B1(n9949), .B2(n9861), .C1(
        n10563), .C2(n9860), .ZN(n10028) );
  INV_X1 U10729 ( .A(n9880), .ZN(n9864) );
  AOI211_X1 U10730 ( .C1(n10030), .C2(n9864), .A(n9915), .B(n9863), .ZN(n10029) );
  NAND2_X1 U10731 ( .A1(n10029), .A2(n9972), .ZN(n9867) );
  AOI22_X1 U10732 ( .A1(n10786), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9865), 
        .B2(n10775), .ZN(n9866) );
  OAI211_X1 U10733 ( .C1(n9868), .C2(n9976), .A(n9867), .B(n9866), .ZN(n9869)
         );
  AOI21_X1 U10734 ( .B1(n10028), .B2(n10560), .A(n9869), .ZN(n9870) );
  OAI21_X1 U10735 ( .B1(n10032), .B2(n9979), .A(n9870), .ZN(P1_U3272) );
  XNOR2_X1 U10736 ( .A(n9871), .B(n9873), .ZN(n10035) );
  INV_X1 U10737 ( .A(n10035), .ZN(n9887) );
  NAND3_X1 U10738 ( .A1(n9874), .A2(n9873), .A3(n9872), .ZN(n9875) );
  NAND2_X1 U10739 ( .A1(n9875), .A2(n10752), .ZN(n9878) );
  AOI22_X1 U10740 ( .A1(n10759), .A2(n9910), .B1(n9876), .B2(n10756), .ZN(
        n9877) );
  OAI21_X1 U10741 ( .B1(n9879), .B2(n9878), .A(n9877), .ZN(n10033) );
  INV_X1 U10742 ( .A(n9881), .ZN(n10099) );
  AOI211_X1 U10743 ( .C1(n9881), .C2(n9896), .A(n9915), .B(n9880), .ZN(n10034)
         );
  NAND2_X1 U10744 ( .A1(n10034), .A2(n9972), .ZN(n9884) );
  AOI22_X1 U10745 ( .A1(n10786), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9882), 
        .B2(n10775), .ZN(n9883) );
  OAI211_X1 U10746 ( .C1(n10099), .C2(n9976), .A(n9884), .B(n9883), .ZN(n9885)
         );
  AOI21_X1 U10747 ( .B1(n10033), .B2(n10560), .A(n9885), .ZN(n9886) );
  OAI21_X1 U10748 ( .B1(n9887), .B2(n9979), .A(n9886), .ZN(P1_U3273) );
  XNOR2_X1 U10749 ( .A(n9888), .B(n9889), .ZN(n10040) );
  INV_X1 U10750 ( .A(n10040), .ZN(n9903) );
  INV_X1 U10751 ( .A(n9889), .ZN(n9890) );
  XNOR2_X1 U10752 ( .A(n9891), .B(n9890), .ZN(n9892) );
  NAND2_X1 U10753 ( .A1(n9892), .A2(n10752), .ZN(n9895) );
  AOI22_X1 U10754 ( .A1(n10759), .A2(n9927), .B1(n9893), .B2(n10756), .ZN(
        n9894) );
  NAND2_X1 U10755 ( .A1(n9895), .A2(n9894), .ZN(n10038) );
  AOI211_X1 U10756 ( .C1(n9897), .C2(n9914), .A(n9915), .B(n5114), .ZN(n10039)
         );
  NAND2_X1 U10757 ( .A1(n10039), .A2(n9972), .ZN(n9900) );
  AOI22_X1 U10758 ( .A1(n10786), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9898), 
        .B2(n10775), .ZN(n9899) );
  OAI211_X1 U10759 ( .C1(n5120), .C2(n9976), .A(n9900), .B(n9899), .ZN(n9901)
         );
  AOI21_X1 U10760 ( .B1(n10038), .B2(n10560), .A(n9901), .ZN(n9902) );
  OAI21_X1 U10761 ( .B1(n9903), .B2(n9979), .A(n9902), .ZN(P1_U3274) );
  XNOR2_X1 U10762 ( .A(n9904), .B(n9905), .ZN(n10045) );
  INV_X1 U10763 ( .A(n10045), .ZN(n9923) );
  NAND2_X1 U10764 ( .A1(n9906), .A2(n9905), .ZN(n9907) );
  NAND2_X1 U10765 ( .A1(n9908), .A2(n9907), .ZN(n9909) );
  NAND2_X1 U10766 ( .A1(n9909), .A2(n10752), .ZN(n9913) );
  AOI22_X1 U10767 ( .A1(n10759), .A2(n9911), .B1(n9910), .B2(n10756), .ZN(
        n9912) );
  NAND2_X1 U10768 ( .A1(n9913), .A2(n9912), .ZN(n10043) );
  INV_X1 U10769 ( .A(n9930), .ZN(n9916) );
  AOI211_X1 U10770 ( .C1(n9917), .C2(n9916), .A(n9915), .B(n5121), .ZN(n10044)
         );
  NAND2_X1 U10771 ( .A1(n10044), .A2(n9972), .ZN(n9920) );
  AOI22_X1 U10772 ( .A1(n10786), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9918), 
        .B2(n10775), .ZN(n9919) );
  OAI211_X1 U10773 ( .C1(n10106), .C2(n9976), .A(n9920), .B(n9919), .ZN(n9921)
         );
  AOI21_X1 U10774 ( .B1(n10043), .B2(n10560), .A(n9921), .ZN(n9922) );
  OAI21_X1 U10775 ( .B1(n9923), .B2(n9979), .A(n9922), .ZN(P1_U3275) );
  XNOR2_X1 U10776 ( .A(n9924), .B(n5309), .ZN(n10050) );
  INV_X1 U10777 ( .A(n10050), .ZN(n9938) );
  XNOR2_X1 U10778 ( .A(n9925), .B(n5309), .ZN(n9926) );
  NAND2_X1 U10779 ( .A1(n9926), .A2(n10752), .ZN(n9929) );
  AOI22_X1 U10780 ( .A1(n10759), .A2(n9964), .B1(n9927), .B2(n10756), .ZN(
        n9928) );
  NAND2_X1 U10781 ( .A1(n9929), .A2(n9928), .ZN(n10048) );
  INV_X1 U10782 ( .A(n9951), .ZN(n9931) );
  AOI211_X1 U10783 ( .C1(n9932), .C2(n9931), .A(n9915), .B(n9930), .ZN(n10049)
         );
  NAND2_X1 U10784 ( .A1(n10049), .A2(n9972), .ZN(n9935) );
  AOI22_X1 U10785 ( .A1(n10786), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9933), 
        .B2(n10775), .ZN(n9934) );
  OAI211_X1 U10786 ( .C1(n10110), .C2(n9976), .A(n9935), .B(n9934), .ZN(n9936)
         );
  AOI21_X1 U10787 ( .B1(n10048), .B2(n10560), .A(n9936), .ZN(n9937) );
  OAI21_X1 U10788 ( .B1(n9938), .B2(n9979), .A(n9937), .ZN(P1_U3276) );
  OAI21_X1 U10789 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(n10053) );
  INV_X1 U10790 ( .A(n9942), .ZN(n9946) );
  AOI21_X1 U10791 ( .B1(n9963), .B2(n9944), .A(n9943), .ZN(n9945) );
  NOR2_X1 U10792 ( .A1(n9946), .A2(n9945), .ZN(n9947) );
  OAI222_X1 U10793 ( .A1(n10551), .A2(n9950), .B1(n9949), .B2(n9948), .C1(
        n10563), .C2(n9947), .ZN(n10054) );
  AOI211_X1 U10794 ( .C1(n9952), .C2(n9968), .A(n9915), .B(n9951), .ZN(n10055)
         );
  NAND2_X1 U10795 ( .A1(n10055), .A2(n9972), .ZN(n9955) );
  AOI22_X1 U10796 ( .A1(n10786), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9953), 
        .B2(n10775), .ZN(n9954) );
  OAI211_X1 U10797 ( .C1(n10114), .C2(n9976), .A(n9955), .B(n9954), .ZN(n9956)
         );
  AOI21_X1 U10798 ( .B1(n10054), .B2(n10560), .A(n9956), .ZN(n9957) );
  OAI21_X1 U10799 ( .B1(n10053), .B2(n9979), .A(n9957), .ZN(P1_U3277) );
  XNOR2_X1 U10800 ( .A(n9958), .B(n9960), .ZN(n10061) );
  INV_X1 U10801 ( .A(n10061), .ZN(n9980) );
  NAND3_X1 U10802 ( .A1(n9961), .A2(n9960), .A3(n9959), .ZN(n9962) );
  NAND3_X1 U10803 ( .A1(n9963), .A2(n10752), .A3(n9962), .ZN(n9967) );
  AOI22_X1 U10804 ( .A1(n10759), .A2(n9965), .B1(n9964), .B2(n10756), .ZN(
        n9966) );
  NAND2_X1 U10805 ( .A1(n9967), .A2(n9966), .ZN(n10059) );
  INV_X1 U10806 ( .A(n9968), .ZN(n9969) );
  AOI211_X1 U10807 ( .C1(n9971), .C2(n9970), .A(n9915), .B(n9969), .ZN(n10060)
         );
  NAND2_X1 U10808 ( .A1(n10060), .A2(n9972), .ZN(n9975) );
  AOI22_X1 U10809 ( .A1(n10786), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9973), 
        .B2(n10775), .ZN(n9974) );
  OAI211_X1 U10810 ( .C1(n10118), .C2(n9976), .A(n9975), .B(n9974), .ZN(n9977)
         );
  AOI21_X1 U10811 ( .B1(n10059), .B2(n10560), .A(n9977), .ZN(n9978) );
  OAI21_X1 U10812 ( .B1(n9980), .B2(n9979), .A(n9978), .ZN(P1_U3278) );
  INV_X1 U10813 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9983) );
  NOR2_X1 U10814 ( .A1(n9982), .A2(n9981), .ZN(n10070) );
  MUX2_X1 U10815 ( .A(n9983), .B(n10070), .S(n10770), .Z(n9984) );
  OAI21_X1 U10816 ( .B1(n10073), .B2(n10069), .A(n9984), .ZN(P1_U3553) );
  INV_X1 U10817 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9987) );
  AND2_X1 U10818 ( .A1(n9986), .A2(n9985), .ZN(n10074) );
  MUX2_X1 U10819 ( .A(n9987), .B(n10074), .S(n10770), .Z(n9988) );
  OAI21_X1 U10820 ( .B1(n10077), .B2(n10069), .A(n9988), .ZN(P1_U3552) );
  NAND2_X1 U10821 ( .A1(n9989), .A2(n10767), .ZN(n9992) );
  MUX2_X1 U10822 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10078), .S(n10770), .Z(
        P1_U3551) );
  AOI211_X1 U10823 ( .C1(n10619), .C2(n9995), .A(n9994), .B(n9993), .ZN(n9996)
         );
  OAI21_X1 U10824 ( .B1(n9997), .B2(n10623), .A(n9996), .ZN(n10079) );
  MUX2_X1 U10825 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10079), .S(n10770), .Z(
        P1_U3550) );
  INV_X1 U10826 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10001) );
  AOI211_X1 U10827 ( .C1(n10000), .C2(n10767), .A(n9999), .B(n9998), .ZN(
        n10080) );
  MUX2_X1 U10828 ( .A(n10001), .B(n10080), .S(n10770), .Z(n10002) );
  OAI21_X1 U10829 ( .B1(n10083), .B2(n10069), .A(n10002), .ZN(P1_U3549) );
  AOI211_X1 U10830 ( .C1(n10619), .C2(n10005), .A(n10004), .B(n10003), .ZN(
        n10006) );
  OAI21_X1 U10831 ( .B1(n10007), .B2(n10623), .A(n10006), .ZN(n10084) );
  MUX2_X1 U10832 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10084), .S(n10770), .Z(
        P1_U3548) );
  INV_X1 U10833 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10011) );
  AOI211_X1 U10834 ( .C1(n10010), .C2(n10767), .A(n10009), .B(n10008), .ZN(
        n10085) );
  MUX2_X1 U10835 ( .A(n10011), .B(n10085), .S(n10770), .Z(n10012) );
  OAI21_X1 U10836 ( .B1(n10088), .B2(n10069), .A(n10012), .ZN(P1_U3547) );
  AOI211_X1 U10837 ( .C1(n10619), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10016) );
  OAI21_X1 U10838 ( .B1(n10017), .B2(n10623), .A(n10016), .ZN(n10089) );
  MUX2_X1 U10839 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10089), .S(n10770), .Z(
        P1_U3546) );
  INV_X1 U10840 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10021) );
  AOI211_X1 U10841 ( .C1(n10020), .C2(n10767), .A(n10019), .B(n10018), .ZN(
        n10090) );
  MUX2_X1 U10842 ( .A(n10021), .B(n10090), .S(n10770), .Z(n10022) );
  OAI21_X1 U10843 ( .B1(n10093), .B2(n10069), .A(n10022), .ZN(P1_U3545) );
  AOI21_X1 U10844 ( .B1(n10619), .B2(n10024), .A(n10023), .ZN(n10025) );
  OAI211_X1 U10845 ( .C1(n10027), .C2(n10623), .A(n10026), .B(n10025), .ZN(
        n10094) );
  MUX2_X1 U10846 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10094), .S(n10770), .Z(
        P1_U3544) );
  AOI211_X1 U10847 ( .C1(n10619), .C2(n10030), .A(n10029), .B(n10028), .ZN(
        n10031) );
  OAI21_X1 U10848 ( .B1(n10032), .B2(n10623), .A(n10031), .ZN(n10095) );
  MUX2_X1 U10849 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10095), .S(n10770), .Z(
        P1_U3543) );
  INV_X1 U10850 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10036) );
  AOI211_X1 U10851 ( .C1(n10035), .C2(n10767), .A(n10034), .B(n10033), .ZN(
        n10096) );
  MUX2_X1 U10852 ( .A(n10036), .B(n10096), .S(n10770), .Z(n10037) );
  OAI21_X1 U10853 ( .B1(n10099), .B2(n10069), .A(n10037), .ZN(P1_U3542) );
  INV_X1 U10854 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10041) );
  AOI211_X1 U10855 ( .C1(n10040), .C2(n10767), .A(n10039), .B(n10038), .ZN(
        n10100) );
  MUX2_X1 U10856 ( .A(n10041), .B(n10100), .S(n10770), .Z(n10042) );
  OAI21_X1 U10857 ( .B1(n5120), .B2(n10069), .A(n10042), .ZN(P1_U3541) );
  AOI211_X1 U10858 ( .C1(n10045), .C2(n10767), .A(n10044), .B(n10043), .ZN(
        n10103) );
  MUX2_X1 U10859 ( .A(n10046), .B(n10103), .S(n10770), .Z(n10047) );
  OAI21_X1 U10860 ( .B1(n10106), .B2(n10069), .A(n10047), .ZN(P1_U3540) );
  AOI211_X1 U10861 ( .C1(n10050), .C2(n10767), .A(n10049), .B(n10048), .ZN(
        n10107) );
  MUX2_X1 U10862 ( .A(n10051), .B(n10107), .S(n10770), .Z(n10052) );
  OAI21_X1 U10863 ( .B1(n10110), .B2(n10069), .A(n10052), .ZN(P1_U3539) );
  INV_X1 U10864 ( .A(n10053), .ZN(n10056) );
  AOI211_X1 U10865 ( .C1(n10056), .C2(n10767), .A(n10055), .B(n10054), .ZN(
        n10111) );
  MUX2_X1 U10866 ( .A(n10057), .B(n10111), .S(n10770), .Z(n10058) );
  OAI21_X1 U10867 ( .B1(n10114), .B2(n10069), .A(n10058), .ZN(P1_U3538) );
  AOI211_X1 U10868 ( .C1(n10061), .C2(n10767), .A(n10060), .B(n10059), .ZN(
        n10115) );
  MUX2_X1 U10869 ( .A(n10062), .B(n10115), .S(n10770), .Z(n10063) );
  OAI21_X1 U10870 ( .B1(n10118), .B2(n10069), .A(n10063), .ZN(P1_U3537) );
  INV_X1 U10871 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10067) );
  AOI211_X1 U10872 ( .C1(n10066), .C2(n10767), .A(n10065), .B(n10064), .ZN(
        n10119) );
  MUX2_X1 U10873 ( .A(n10067), .B(n10119), .S(n10770), .Z(n10068) );
  OAI21_X1 U10874 ( .B1(n10123), .B2(n10069), .A(n10068), .ZN(P1_U3536) );
  INV_X1 U10875 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10071) );
  MUX2_X1 U10876 ( .A(n10071), .B(n10070), .S(n10774), .Z(n10072) );
  OAI21_X1 U10877 ( .B1(n10073), .B2(n10122), .A(n10072), .ZN(P1_U3521) );
  INV_X1 U10878 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10075) );
  MUX2_X1 U10879 ( .A(n10075), .B(n10074), .S(n10774), .Z(n10076) );
  OAI21_X1 U10880 ( .B1(n10077), .B2(n10122), .A(n10076), .ZN(P1_U3520) );
  MUX2_X1 U10881 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10078), .S(n10774), .Z(
        P1_U3519) );
  MUX2_X1 U10882 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10079), .S(n10774), .Z(
        P1_U3518) );
  INV_X1 U10883 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10081) );
  MUX2_X1 U10884 ( .A(n10081), .B(n10080), .S(n10774), .Z(n10082) );
  OAI21_X1 U10885 ( .B1(n10083), .B2(n10122), .A(n10082), .ZN(P1_U3517) );
  MUX2_X1 U10886 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10084), .S(n10774), .Z(
        P1_U3516) );
  INV_X1 U10887 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10086) );
  MUX2_X1 U10888 ( .A(n10086), .B(n10085), .S(n10774), .Z(n10087) );
  OAI21_X1 U10889 ( .B1(n10088), .B2(n10122), .A(n10087), .ZN(P1_U3515) );
  MUX2_X1 U10890 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10089), .S(n10774), .Z(
        P1_U3514) );
  INV_X1 U10891 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10091) );
  MUX2_X1 U10892 ( .A(n10091), .B(n10090), .S(n10774), .Z(n10092) );
  OAI21_X1 U10893 ( .B1(n10093), .B2(n10122), .A(n10092), .ZN(P1_U3513) );
  MUX2_X1 U10894 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10094), .S(n10774), .Z(
        P1_U3512) );
  MUX2_X1 U10895 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10095), .S(n10774), .Z(
        P1_U3511) );
  INV_X1 U10896 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10097) );
  MUX2_X1 U10897 ( .A(n10097), .B(n10096), .S(n10774), .Z(n10098) );
  OAI21_X1 U10898 ( .B1(n10099), .B2(n10122), .A(n10098), .ZN(P1_U3510) );
  INV_X1 U10899 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10101) );
  MUX2_X1 U10900 ( .A(n10101), .B(n10100), .S(n10774), .Z(n10102) );
  OAI21_X1 U10901 ( .B1(n5120), .B2(n10122), .A(n10102), .ZN(P1_U3509) );
  INV_X1 U10902 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10104) );
  MUX2_X1 U10903 ( .A(n10104), .B(n10103), .S(n10774), .Z(n10105) );
  OAI21_X1 U10904 ( .B1(n10106), .B2(n10122), .A(n10105), .ZN(P1_U3507) );
  INV_X1 U10905 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10108) );
  MUX2_X1 U10906 ( .A(n10108), .B(n10107), .S(n10774), .Z(n10109) );
  OAI21_X1 U10907 ( .B1(n10110), .B2(n10122), .A(n10109), .ZN(P1_U3504) );
  INV_X1 U10908 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10112) );
  MUX2_X1 U10909 ( .A(n10112), .B(n10111), .S(n10774), .Z(n10113) );
  OAI21_X1 U10910 ( .B1(n10114), .B2(n10122), .A(n10113), .ZN(P1_U3501) );
  INV_X1 U10911 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10116) );
  MUX2_X1 U10912 ( .A(n10116), .B(n10115), .S(n10774), .Z(n10117) );
  OAI21_X1 U10913 ( .B1(n10118), .B2(n10122), .A(n10117), .ZN(P1_U3498) );
  INV_X1 U10914 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10120) );
  MUX2_X1 U10915 ( .A(n10120), .B(n10119), .S(n10774), .Z(n10121) );
  OAI21_X1 U10916 ( .B1(n10123), .B2(n10122), .A(n10121), .ZN(P1_U3495) );
  NOR4_X1 U10917 ( .A1(n5554), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10124), .A4(
        P1_U3086), .ZN(n10125) );
  AOI21_X1 U10918 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n10126), .A(n10125), 
        .ZN(n10127) );
  OAI21_X1 U10919 ( .B1(n10128), .B2(n10138), .A(n10127), .ZN(P1_U3324) );
  OAI222_X1 U10920 ( .A1(n10132), .A2(n10131), .B1(P1_U3086), .B2(n10130), 
        .C1(n10138), .C2(n10129), .ZN(P1_U3326) );
  OAI222_X1 U10921 ( .A1(P1_U3086), .A2(n10135), .B1(n10138), .B2(n10134), 
        .C1(n10133), .C2(n10132), .ZN(P1_U3327) );
  OAI222_X1 U10922 ( .A1(P1_U3086), .A2(n10139), .B1(n10138), .B2(n10137), 
        .C1(n10136), .C2(n10132), .ZN(P1_U3328) );
  MUX2_X1 U10923 ( .A(n10140), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U10924 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10141), .ZN(P1_U3323) );
  AND2_X1 U10925 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10141), .ZN(P1_U3322) );
  AND2_X1 U10926 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10141), .ZN(P1_U3321) );
  AND2_X1 U10927 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10141), .ZN(P1_U3320) );
  AND2_X1 U10928 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10141), .ZN(P1_U3319) );
  AND2_X1 U10929 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10141), .ZN(P1_U3318) );
  AND2_X1 U10930 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10141), .ZN(P1_U3317) );
  AND2_X1 U10931 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10141), .ZN(P1_U3316) );
  AND2_X1 U10932 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10141), .ZN(P1_U3315) );
  AND2_X1 U10933 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10141), .ZN(P1_U3314) );
  AND2_X1 U10934 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10141), .ZN(P1_U3313) );
  AND2_X1 U10935 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10141), .ZN(P1_U3312) );
  AND2_X1 U10936 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10141), .ZN(P1_U3311) );
  AND2_X1 U10937 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10141), .ZN(P1_U3310) );
  AND2_X1 U10938 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10141), .ZN(P1_U3309) );
  AND2_X1 U10939 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10141), .ZN(P1_U3308) );
  AND2_X1 U10940 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10141), .ZN(P1_U3307) );
  AND2_X1 U10941 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10141), .ZN(P1_U3306) );
  AND2_X1 U10942 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10141), .ZN(P1_U3305) );
  AND2_X1 U10943 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10141), .ZN(P1_U3304) );
  AND2_X1 U10944 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10141), .ZN(P1_U3303) );
  AND2_X1 U10945 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10141), .ZN(P1_U3302) );
  AND2_X1 U10946 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10141), .ZN(P1_U3301) );
  AND2_X1 U10947 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10141), .ZN(P1_U3300) );
  AND2_X1 U10948 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10141), .ZN(P1_U3299) );
  AND2_X1 U10949 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10141), .ZN(P1_U3298) );
  AND2_X1 U10950 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10141), .ZN(P1_U3297) );
  AND2_X1 U10951 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10141), .ZN(P1_U3296) );
  AND2_X1 U10952 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10141), .ZN(P1_U3295) );
  AND2_X1 U10953 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10141), .ZN(P1_U3294) );
  OAI22_X1 U10954 ( .A1(n10364), .A2(keyinput_126), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_127), .ZN(n10142) );
  AOI221_X1 U10955 ( .B1(n10364), .B2(keyinput_126), .C1(keyinput_127), .C2(
        P2_REG3_REG_15__SCAN_IN), .A(n10142), .ZN(n10368) );
  INV_X1 U10956 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10361) );
  OAI22_X1 U10957 ( .A1(n10144), .A2(keyinput_124), .B1(n10597), .B2(
        keyinput_123), .ZN(n10143) );
  AOI221_X1 U10958 ( .B1(n10144), .B2(keyinput_124), .C1(keyinput_123), .C2(
        n10597), .A(n10143), .ZN(n10241) );
  AOI22_X1 U10959 ( .A1(n5947), .A2(keyinput_120), .B1(n10146), .B2(
        keyinput_119), .ZN(n10145) );
  OAI221_X1 U10960 ( .B1(n5947), .B2(keyinput_120), .C1(n10146), .C2(
        keyinput_119), .A(n10145), .ZN(n10239) );
  OAI22_X1 U10961 ( .A1(n6765), .A2(keyinput_118), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(keyinput_117), .ZN(n10147) );
  AOI221_X1 U10962 ( .B1(n6765), .B2(keyinput_118), .C1(keyinput_117), .C2(
        P2_REG3_REG_9__SCAN_IN), .A(n10147), .ZN(n10238) );
  XNOR2_X1 U10963 ( .A(n10346), .B(keyinput_115), .ZN(n10233) );
  INV_X1 U10964 ( .A(keyinput_114), .ZN(n10230) );
  INV_X1 U10965 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10337) );
  XOR2_X1 U10966 ( .A(n10337), .B(keyinput_109), .Z(n10227) );
  INV_X1 U10967 ( .A(keyinput_104), .ZN(n10216) );
  INV_X1 U10968 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10149) );
  OAI22_X1 U10969 ( .A1(n10149), .A2(keyinput_100), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .ZN(n10148) );
  AOI221_X1 U10970 ( .B1(n10149), .B2(keyinput_100), .C1(keyinput_101), .C2(
        P2_REG3_REG_14__SCAN_IN), .A(n10148), .ZN(n10214) );
  INV_X1 U10971 ( .A(keyinput_99), .ZN(n10210) );
  AOI22_X1 U10972 ( .A1(SI_5_), .A2(keyinput_91), .B1(n10151), .B2(keyinput_90), .ZN(n10150) );
  OAI221_X1 U10973 ( .B1(SI_5_), .B2(keyinput_91), .C1(n10151), .C2(
        keyinput_90), .A(n10150), .ZN(n10193) );
  OAI22_X1 U10974 ( .A1(n10298), .A2(keyinput_88), .B1(keyinput_89), .B2(SI_7_), .ZN(n10152) );
  AOI221_X1 U10975 ( .B1(n10298), .B2(keyinput_88), .C1(SI_7_), .C2(
        keyinput_89), .A(n10152), .ZN(n10190) );
  INV_X1 U10976 ( .A(SI_10_), .ZN(n10291) );
  INV_X1 U10977 ( .A(SI_13_), .ZN(n10288) );
  INV_X1 U10978 ( .A(keyinput_83), .ZN(n10183) );
  INV_X1 U10979 ( .A(keyinput_82), .ZN(n10181) );
  INV_X1 U10980 ( .A(keyinput_81), .ZN(n10179) );
  OAI22_X1 U10981 ( .A1(n10250), .A2(keyinput_80), .B1(SI_18_), .B2(
        keyinput_78), .ZN(n10153) );
  AOI221_X1 U10982 ( .B1(n10250), .B2(keyinput_80), .C1(keyinput_78), .C2(
        SI_18_), .A(n10153), .ZN(n10176) );
  AOI22_X1 U10983 ( .A1(SI_21_), .A2(keyinput_75), .B1(n10155), .B2(
        keyinput_76), .ZN(n10154) );
  OAI221_X1 U10984 ( .B1(SI_21_), .B2(keyinput_75), .C1(n10155), .C2(
        keyinput_76), .A(n10154), .ZN(n10174) );
  INV_X1 U10985 ( .A(SI_22_), .ZN(n10273) );
  INV_X1 U10986 ( .A(keyinput_74), .ZN(n10171) );
  INV_X1 U10987 ( .A(keyinput_67), .ZN(n10160) );
  INV_X1 U10988 ( .A(keyinput_66), .ZN(n10158) );
  OAI22_X1 U10989 ( .A1(SI_31_), .A2(keyinput_65), .B1(P2_WR_REG_SCAN_IN), 
        .B2(keyinput_64), .ZN(n10156) );
  AOI221_X1 U10990 ( .B1(SI_31_), .B2(keyinput_65), .C1(keyinput_64), .C2(
        P2_WR_REG_SCAN_IN), .A(n10156), .ZN(n10157) );
  AOI221_X1 U10991 ( .B1(SI_30_), .B2(keyinput_66), .C1(n10262), .C2(n10158), 
        .A(n10157), .ZN(n10159) );
  AOI221_X1 U10992 ( .B1(SI_29_), .B2(n10160), .C1(n10266), .C2(keyinput_67), 
        .A(n10159), .ZN(n10169) );
  INV_X1 U10993 ( .A(SI_25_), .ZN(n10258) );
  AOI22_X1 U10994 ( .A1(n10258), .A2(keyinput_71), .B1(n10256), .B2(
        keyinput_69), .ZN(n10161) );
  OAI221_X1 U10995 ( .B1(n10258), .B2(keyinput_71), .C1(n10256), .C2(
        keyinput_69), .A(n10161), .ZN(n10168) );
  AOI22_X1 U10996 ( .A1(SI_28_), .A2(keyinput_68), .B1(n10163), .B2(
        keyinput_72), .ZN(n10162) );
  OAI221_X1 U10997 ( .B1(SI_28_), .B2(keyinput_68), .C1(n10163), .C2(
        keyinput_72), .A(n10162), .ZN(n10167) );
  AOI22_X1 U10998 ( .A1(n10255), .A2(keyinput_73), .B1(n10165), .B2(
        keyinput_70), .ZN(n10164) );
  OAI221_X1 U10999 ( .B1(n10255), .B2(keyinput_73), .C1(n10165), .C2(
        keyinput_70), .A(n10164), .ZN(n10166) );
  NOR4_X1 U11000 ( .A1(n10169), .A2(n10168), .A3(n10167), .A4(n10166), .ZN(
        n10170) );
  AOI221_X1 U11001 ( .B1(SI_22_), .B2(keyinput_74), .C1(n10273), .C2(n10171), 
        .A(n10170), .ZN(n10173) );
  NAND2_X1 U11002 ( .A1(n10277), .A2(keyinput_77), .ZN(n10172) );
  OAI221_X1 U11003 ( .B1(n10174), .B2(n10173), .C1(n10277), .C2(keyinput_77), 
        .A(n10172), .ZN(n10175) );
  OAI211_X1 U11004 ( .C1(SI_17_), .C2(keyinput_79), .A(n10176), .B(n10175), 
        .ZN(n10177) );
  AOI21_X1 U11005 ( .B1(SI_17_), .B2(keyinput_79), .A(n10177), .ZN(n10178) );
  AOI221_X1 U11006 ( .B1(SI_15_), .B2(n10179), .C1(n10283), .C2(keyinput_81), 
        .A(n10178), .ZN(n10180) );
  AOI221_X1 U11007 ( .B1(SI_14_), .B2(n10181), .C1(n10286), .C2(keyinput_82), 
        .A(n10180), .ZN(n10182) );
  AOI221_X1 U11008 ( .B1(SI_13_), .B2(keyinput_83), .C1(n10288), .C2(n10183), 
        .A(n10182), .ZN(n10187) );
  AOI22_X1 U11009 ( .A1(SI_12_), .A2(keyinput_84), .B1(n10185), .B2(
        keyinput_85), .ZN(n10184) );
  OAI221_X1 U11010 ( .B1(SI_12_), .B2(keyinput_84), .C1(n10185), .C2(
        keyinput_85), .A(n10184), .ZN(n10186) );
  AOI211_X1 U11011 ( .C1(n10291), .C2(keyinput_86), .A(n10187), .B(n10186), 
        .ZN(n10188) );
  OAI21_X1 U11012 ( .B1(n10291), .B2(keyinput_86), .A(n10188), .ZN(n10189) );
  OAI211_X1 U11013 ( .C1(SI_9_), .C2(keyinput_87), .A(n10190), .B(n10189), 
        .ZN(n10191) );
  AOI21_X1 U11014 ( .B1(SI_9_), .B2(keyinput_87), .A(n10191), .ZN(n10192) );
  OAI22_X1 U11015 ( .A1(keyinput_92), .A2(n10195), .B1(n10193), .B2(n10192), 
        .ZN(n10194) );
  AOI21_X1 U11016 ( .B1(keyinput_92), .B2(n10195), .A(n10194), .ZN(n10198) );
  INV_X1 U11017 ( .A(keyinput_93), .ZN(n10196) );
  MUX2_X1 U11018 ( .A(keyinput_93), .B(n10196), .S(SI_3_), .Z(n10197) );
  NOR2_X1 U11019 ( .A1(n10198), .A2(n10197), .ZN(n10201) );
  INV_X1 U11020 ( .A(keyinput_94), .ZN(n10199) );
  MUX2_X1 U11021 ( .A(n10199), .B(keyinput_94), .S(SI_2_), .Z(n10200) );
  NOR2_X1 U11022 ( .A1(n10201), .A2(n10200), .ZN(n10206) );
  INV_X1 U11023 ( .A(keyinput_95), .ZN(n10202) );
  MUX2_X1 U11024 ( .A(n10202), .B(keyinput_95), .S(SI_1_), .Z(n10205) );
  INV_X1 U11025 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10530) );
  XOR2_X1 U11026 ( .A(n10530), .B(keyinput_97), .Z(n10204) );
  XNOR2_X1 U11027 ( .A(SI_0_), .B(keyinput_96), .ZN(n10203) );
  OAI211_X1 U11028 ( .C1(n10206), .C2(n10205), .A(n10204), .B(n10203), .ZN(
        n10208) );
  NAND2_X1 U11029 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_98), .ZN(n10207)
         );
  OAI211_X1 U11030 ( .C1(P2_STATE_REG_SCAN_IN), .C2(keyinput_98), .A(n10208), 
        .B(n10207), .ZN(n10209) );
  OAI221_X1 U11031 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_99), .C1(n10317), .C2(n10210), .A(n10209), .ZN(n10213) );
  AOI22_X1 U11032 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_103), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_102), .ZN(n10211) );
  OAI221_X1 U11033 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_103), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_102), .A(n10211), .ZN(n10212)
         );
  AOI21_X1 U11034 ( .B1(n10214), .B2(n10213), .A(n10212), .ZN(n10215) );
  AOI221_X1 U11035 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .C1(
        n10244), .C2(n10216), .A(n10215), .ZN(n10221) );
  AOI22_X1 U11036 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_105), .B1(
        n10325), .B2(keyinput_106), .ZN(n10217) );
  OAI221_X1 U11037 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .C1(
        n10325), .C2(keyinput_106), .A(n10217), .ZN(n10220) );
  XNOR2_X1 U11038 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_108), .ZN(n10219)
         );
  XNOR2_X1 U11039 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_107), .ZN(n10218)
         );
  OAI211_X1 U11040 ( .C1(n10221), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        n10226) );
  AOI22_X1 U11041 ( .A1(n5814), .A2(keyinput_113), .B1(n10340), .B2(
        keyinput_112), .ZN(n10222) );
  OAI221_X1 U11042 ( .B1(n5814), .B2(keyinput_113), .C1(n10340), .C2(
        keyinput_112), .A(n10222), .ZN(n10225) );
  AOI22_X1 U11043 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_110), .B1(
        P2_REG3_REG_25__SCAN_IN), .B2(keyinput_111), .ZN(n10223) );
  OAI221_X1 U11044 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput_111), .A(n10223), .ZN(n10224)
         );
  AOI211_X1 U11045 ( .C1(n10227), .C2(n10226), .A(n10225), .B(n10224), .ZN(
        n10228) );
  AOI221_X1 U11046 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(n10230), .C1(n10229), 
        .C2(keyinput_114), .A(n10228), .ZN(n10232) );
  INV_X1 U11047 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10350) );
  NAND2_X1 U11048 ( .A1(n10350), .A2(keyinput_116), .ZN(n10231) );
  OAI221_X1 U11049 ( .B1(n10233), .B2(n10232), .C1(n10350), .C2(keyinput_116), 
        .A(n10231), .ZN(n10237) );
  OAI22_X1 U11050 ( .A1(n10235), .A2(keyinput_121), .B1(keyinput_122), .B2(
        P2_REG3_REG_11__SCAN_IN), .ZN(n10234) );
  AOI221_X1 U11051 ( .B1(n10235), .B2(keyinput_121), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_122), .A(n10234), .ZN(n10236)
         );
  OAI221_X1 U11052 ( .B1(n10239), .B2(n10238), .C1(n10239), .C2(n10237), .A(
        n10236), .ZN(n10240) );
  AOI22_X1 U11053 ( .A1(keyinput_125), .A2(n10361), .B1(n10241), .B2(n10240), 
        .ZN(n10242) );
  OAI21_X1 U11054 ( .B1(n10361), .B2(keyinput_125), .A(n10242), .ZN(n10367) );
  AOI22_X1 U11055 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_60), .B1(n10597), .B2(keyinput_59), .ZN(n10243) );
  OAI221_X1 U11056 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .C1(
        n10597), .C2(keyinput_59), .A(n10243), .ZN(n10359) );
  INV_X1 U11057 ( .A(keyinput_52), .ZN(n10349) );
  INV_X1 U11058 ( .A(keyinput_51), .ZN(n10347) );
  XOR2_X1 U11059 ( .A(n10244), .B(keyinput_40), .Z(n10329) );
  INV_X1 U11060 ( .A(keyinput_35), .ZN(n10316) );
  AOI22_X1 U11061 ( .A1(SI_6_), .A2(keyinput_26), .B1(n10246), .B2(keyinput_27), .ZN(n10245) );
  OAI221_X1 U11062 ( .B1(SI_6_), .B2(keyinput_26), .C1(n10246), .C2(
        keyinput_27), .A(n10245), .ZN(n10300) );
  OAI22_X1 U11063 ( .A1(n10248), .A2(keyinput_23), .B1(keyinput_25), .B2(SI_7_), .ZN(n10247) );
  AOI221_X1 U11064 ( .B1(n10248), .B2(keyinput_23), .C1(SI_7_), .C2(
        keyinput_25), .A(n10247), .ZN(n10296) );
  INV_X1 U11065 ( .A(keyinput_19), .ZN(n10289) );
  INV_X1 U11066 ( .A(keyinput_18), .ZN(n10285) );
  INV_X1 U11067 ( .A(keyinput_17), .ZN(n10282) );
  OAI22_X1 U11068 ( .A1(n10251), .A2(keyinput_15), .B1(n10250), .B2(
        keyinput_16), .ZN(n10249) );
  AOI221_X1 U11069 ( .B1(n10251), .B2(keyinput_15), .C1(keyinput_16), .C2(
        n10250), .A(n10249), .ZN(n10279) );
  OAI22_X1 U11070 ( .A1(n10253), .A2(keyinput_11), .B1(SI_20_), .B2(
        keyinput_12), .ZN(n10252) );
  AOI221_X1 U11071 ( .B1(n10253), .B2(keyinput_11), .C1(keyinput_12), .C2(
        SI_20_), .A(n10252), .ZN(n10275) );
  INV_X1 U11072 ( .A(keyinput_10), .ZN(n10272) );
  OAI22_X1 U11073 ( .A1(n10256), .A2(keyinput_5), .B1(n10255), .B2(keyinput_9), 
        .ZN(n10254) );
  AOI221_X1 U11074 ( .B1(n10256), .B2(keyinput_5), .C1(keyinput_9), .C2(n10255), .A(n10254), .ZN(n10270) );
  OAI22_X1 U11075 ( .A1(n10258), .A2(keyinput_7), .B1(SI_26_), .B2(keyinput_6), 
        .ZN(n10257) );
  AOI221_X1 U11076 ( .B1(n10258), .B2(keyinput_7), .C1(keyinput_6), .C2(SI_26_), .A(n10257), .ZN(n10269) );
  OAI22_X1 U11077 ( .A1(SI_24_), .A2(keyinput_8), .B1(SI_28_), .B2(keyinput_4), 
        .ZN(n10259) );
  AOI221_X1 U11078 ( .B1(SI_24_), .B2(keyinput_8), .C1(keyinput_4), .C2(SI_28_), .A(n10259), .ZN(n10268) );
  INV_X1 U11079 ( .A(keyinput_3), .ZN(n10265) );
  INV_X1 U11080 ( .A(keyinput_2), .ZN(n10263) );
  AOI22_X1 U11081 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n10260) );
  OAI221_X1 U11082 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_31_), 
        .C2(keyinput_1), .A(n10260), .ZN(n10261) );
  OAI221_X1 U11083 ( .B1(SI_30_), .B2(n10263), .C1(n10262), .C2(keyinput_2), 
        .A(n10261), .ZN(n10264) );
  OAI221_X1 U11084 ( .B1(SI_29_), .B2(keyinput_3), .C1(n10266), .C2(n10265), 
        .A(n10264), .ZN(n10267) );
  NAND4_X1 U11085 ( .A1(n10270), .A2(n10269), .A3(n10268), .A4(n10267), .ZN(
        n10271) );
  OAI221_X1 U11086 ( .B1(SI_22_), .B2(keyinput_10), .C1(n10273), .C2(n10272), 
        .A(n10271), .ZN(n10274) );
  AOI22_X1 U11087 ( .A1(keyinput_13), .A2(n10277), .B1(n10275), .B2(n10274), 
        .ZN(n10276) );
  OAI21_X1 U11088 ( .B1(n10277), .B2(keyinput_13), .A(n10276), .ZN(n10278) );
  OAI211_X1 U11089 ( .C1(SI_18_), .C2(keyinput_14), .A(n10279), .B(n10278), 
        .ZN(n10280) );
  AOI21_X1 U11090 ( .B1(SI_18_), .B2(keyinput_14), .A(n10280), .ZN(n10281) );
  AOI221_X1 U11091 ( .B1(SI_15_), .B2(keyinput_17), .C1(n10283), .C2(n10282), 
        .A(n10281), .ZN(n10284) );
  AOI221_X1 U11092 ( .B1(SI_14_), .B2(keyinput_18), .C1(n10286), .C2(n10285), 
        .A(n10284), .ZN(n10287) );
  AOI221_X1 U11093 ( .B1(SI_13_), .B2(n10289), .C1(n10288), .C2(keyinput_19), 
        .A(n10287), .ZN(n10293) );
  AOI22_X1 U11094 ( .A1(SI_12_), .A2(keyinput_20), .B1(n10291), .B2(
        keyinput_22), .ZN(n10290) );
  OAI221_X1 U11095 ( .B1(SI_12_), .B2(keyinput_20), .C1(n10291), .C2(
        keyinput_22), .A(n10290), .ZN(n10292) );
  AOI211_X1 U11096 ( .C1(SI_11_), .C2(keyinput_21), .A(n10293), .B(n10292), 
        .ZN(n10294) );
  OAI21_X1 U11097 ( .B1(SI_11_), .B2(keyinput_21), .A(n10294), .ZN(n10295) );
  OAI211_X1 U11098 ( .C1(n10298), .C2(keyinput_24), .A(n10296), .B(n10295), 
        .ZN(n10297) );
  AOI21_X1 U11099 ( .B1(n10298), .B2(keyinput_24), .A(n10297), .ZN(n10299) );
  OAI22_X1 U11100 ( .A1(n10300), .A2(n10299), .B1(keyinput_28), .B2(SI_4_), 
        .ZN(n10301) );
  AOI21_X1 U11101 ( .B1(keyinput_28), .B2(SI_4_), .A(n10301), .ZN(n10304) );
  INV_X1 U11102 ( .A(keyinput_29), .ZN(n10302) );
  MUX2_X1 U11103 ( .A(n10302), .B(keyinput_29), .S(SI_3_), .Z(n10303) );
  NOR2_X1 U11104 ( .A1(n10304), .A2(n10303), .ZN(n10307) );
  INV_X1 U11105 ( .A(keyinput_30), .ZN(n10305) );
  MUX2_X1 U11106 ( .A(keyinput_30), .B(n10305), .S(SI_2_), .Z(n10306) );
  NOR2_X1 U11107 ( .A1(n10307), .A2(n10306), .ZN(n10310) );
  INV_X1 U11108 ( .A(keyinput_31), .ZN(n10308) );
  MUX2_X1 U11109 ( .A(keyinput_31), .B(n10308), .S(SI_1_), .Z(n10309) );
  NOR2_X1 U11110 ( .A1(n10310), .A2(n10309), .ZN(n10313) );
  AOI22_X1 U11111 ( .A1(SI_0_), .A2(keyinput_32), .B1(n10530), .B2(keyinput_33), .ZN(n10311) );
  OAI221_X1 U11112 ( .B1(SI_0_), .B2(keyinput_32), .C1(n10530), .C2(
        keyinput_33), .A(n10311), .ZN(n10312) );
  OAI22_X1 U11113 ( .A1(n10313), .A2(n10312), .B1(keyinput_34), .B2(P2_U3151), 
        .ZN(n10314) );
  AOI21_X1 U11114 ( .B1(keyinput_34), .B2(P2_U3151), .A(n10314), .ZN(n10315)
         );
  AOI221_X1 U11115 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_35), .C1(n10317), .C2(n10316), .A(n10315), .ZN(n10323) );
  AOI22_X1 U11116 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_37), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_36), .ZN(n10318) );
  OAI221_X1 U11117 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_36), .A(n10318), .ZN(n10322) );
  INV_X1 U11118 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10320) );
  OAI22_X1 U11119 ( .A1(n10320), .A2(keyinput_39), .B1(keyinput_38), .B2(
        P2_REG3_REG_23__SCAN_IN), .ZN(n10319) );
  AOI221_X1 U11120 ( .B1(n10320), .B2(keyinput_39), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_38), .A(n10319), .ZN(n10321) );
  OAI21_X1 U11121 ( .B1(n10323), .B2(n10322), .A(n10321), .ZN(n10328) );
  INV_X1 U11122 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U11123 ( .A1(n10326), .A2(keyinput_41), .B1(n10325), .B2(
        keyinput_42), .ZN(n10324) );
  OAI221_X1 U11124 ( .B1(n10326), .B2(keyinput_41), .C1(n10325), .C2(
        keyinput_42), .A(n10324), .ZN(n10327) );
  AOI21_X1 U11125 ( .B1(n10329), .B2(n10328), .A(n10327), .ZN(n10333) );
  XNOR2_X1 U11126 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .ZN(n10331)
         );
  XNOR2_X1 U11127 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_43), .ZN(n10330)
         );
  NAND2_X1 U11128 ( .A1(n10331), .A2(n10330), .ZN(n10332) );
  OAI22_X1 U11129 ( .A1(n10333), .A2(n10332), .B1(keyinput_45), .B2(n10337), 
        .ZN(n10338) );
  INV_X1 U11130 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10335) );
  OAI22_X1 U11131 ( .A1(n10335), .A2(keyinput_47), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(keyinput_49), .ZN(n10334) );
  AOI221_X1 U11132 ( .B1(n10335), .B2(keyinput_47), .C1(keyinput_49), .C2(
        P2_REG3_REG_5__SCAN_IN), .A(n10334), .ZN(n10336) );
  OAI221_X1 U11133 ( .B1(n10338), .B2(keyinput_45), .C1(n10338), .C2(n10337), 
        .A(n10336), .ZN(n10343) );
  AOI22_X1 U11134 ( .A1(n10341), .A2(keyinput_46), .B1(n10340), .B2(
        keyinput_48), .ZN(n10339) );
  OAI221_X1 U11135 ( .B1(n10341), .B2(keyinput_46), .C1(n10340), .C2(
        keyinput_48), .A(n10339), .ZN(n10342) );
  OAI22_X1 U11136 ( .A1(n10343), .A2(n10342), .B1(keyinput_50), .B2(
        P2_REG3_REG_17__SCAN_IN), .ZN(n10344) );
  AOI21_X1 U11137 ( .B1(keyinput_50), .B2(P2_REG3_REG_17__SCAN_IN), .A(n10344), 
        .ZN(n10345) );
  AOI221_X1 U11138 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n10347), .C1(n10346), 
        .C2(keyinput_51), .A(n10345), .ZN(n10348) );
  AOI221_X1 U11139 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_52), .C1(n10350), .C2(n10349), .A(n10348), .ZN(n10357) );
  OAI22_X1 U11140 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_55), .B1(
        keyinput_56), .B2(P2_REG3_REG_13__SCAN_IN), .ZN(n10351) );
  AOI221_X1 U11141 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_55), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_56), .A(n10351), .ZN(n10356) );
  AOI22_X1 U11142 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_53), .B1(n6765), 
        .B2(keyinput_54), .ZN(n10352) );
  OAI221_X1 U11143 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .C1(n6765), 
        .C2(keyinput_54), .A(n10352), .ZN(n10355) );
  AOI22_X1 U11144 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_58), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .ZN(n10353) );
  OAI221_X1 U11145 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_57), .A(n10353), .ZN(n10354) );
  AOI221_X1 U11146 ( .B1(n10357), .B2(n10356), .C1(n10355), .C2(n10356), .A(
        n10354), .ZN(n10358) );
  OAI22_X1 U11147 ( .A1(keyinput_61), .A2(n10361), .B1(n10359), .B2(n10358), 
        .ZN(n10360) );
  AOI21_X1 U11148 ( .B1(keyinput_61), .B2(n10361), .A(n10360), .ZN(n10366) );
  AOI22_X1 U11149 ( .A1(n10364), .A2(keyinput_62), .B1(keyinput_63), .B2(
        n10363), .ZN(n10362) );
  OAI221_X1 U11150 ( .B1(n10364), .B2(keyinput_62), .C1(n10363), .C2(
        keyinput_63), .A(n10362), .ZN(n10365) );
  AOI211_X1 U11151 ( .C1(n10368), .C2(n10367), .A(n10366), .B(n10365), .ZN(
        n10372) );
  MUX2_X1 U11152 ( .A(n10370), .B(n10369), .S(P1_U3973), .Z(n10371) );
  XNOR2_X1 U11153 ( .A(n10372), .B(n10371), .ZN(P1_U3583) );
  XOR2_X1 U11154 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI222_X1 U11155 ( .A1(n10377), .A2(n10376), .B1(n10377), .B2(n10375), .C1(
        n10374), .C2(n10373), .ZN(ADD_1068_U5) );
  AOI21_X1 U11156 ( .B1(n10380), .B2(n10379), .A(n10378), .ZN(ADD_1068_U54) );
  AOI21_X1 U11157 ( .B1(n10383), .B2(n10382), .A(n10381), .ZN(ADD_1068_U53) );
  OAI21_X1 U11158 ( .B1(n10386), .B2(n10385), .A(n10384), .ZN(ADD_1068_U52) );
  OAI21_X1 U11159 ( .B1(n10389), .B2(n10388), .A(n10387), .ZN(ADD_1068_U51) );
  OAI21_X1 U11160 ( .B1(n10392), .B2(n10391), .A(n10390), .ZN(ADD_1068_U50) );
  OAI21_X1 U11161 ( .B1(n10395), .B2(n10394), .A(n10393), .ZN(ADD_1068_U49) );
  OAI21_X1 U11162 ( .B1(n10398), .B2(n10397), .A(n10396), .ZN(ADD_1068_U48) );
  OAI21_X1 U11163 ( .B1(n10401), .B2(n10400), .A(n10399), .ZN(ADD_1068_U47) );
  OAI21_X1 U11164 ( .B1(n10404), .B2(n10403), .A(n10402), .ZN(ADD_1068_U63) );
  OAI21_X1 U11165 ( .B1(n10407), .B2(n10406), .A(n10405), .ZN(ADD_1068_U62) );
  OAI21_X1 U11166 ( .B1(n10410), .B2(n10409), .A(n10408), .ZN(ADD_1068_U61) );
  OAI21_X1 U11167 ( .B1(n10413), .B2(n10412), .A(n10411), .ZN(ADD_1068_U60) );
  OAI21_X1 U11168 ( .B1(n10416), .B2(n10415), .A(n10414), .ZN(ADD_1068_U59) );
  OAI21_X1 U11169 ( .B1(n10419), .B2(n10418), .A(n10417), .ZN(ADD_1068_U58) );
  OAI21_X1 U11170 ( .B1(n10422), .B2(n10421), .A(n10420), .ZN(ADD_1068_U57) );
  OAI21_X1 U11171 ( .B1(n10425), .B2(n10424), .A(n10423), .ZN(ADD_1068_U56) );
  OAI21_X1 U11172 ( .B1(n10428), .B2(n10427), .A(n10426), .ZN(ADD_1068_U55) );
  OAI21_X1 U11173 ( .B1(n10431), .B2(n10430), .A(n10429), .ZN(n10432) );
  AOI22_X1 U11174 ( .A1(n10525), .A2(n10432), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(P2_U3151), .ZN(n10442) );
  NAND2_X1 U11175 ( .A1(n10434), .A2(n10433), .ZN(n10441) );
  NAND2_X1 U11176 ( .A1(n10516), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n10440) );
  OAI21_X1 U11177 ( .B1(n10437), .B2(n10436), .A(n10435), .ZN(n10438) );
  NAND2_X1 U11178 ( .A1(n10492), .A2(n10438), .ZN(n10439) );
  AND4_X1 U11179 ( .A1(n10442), .A2(n10441), .A3(n10440), .A4(n10439), .ZN(
        n10447) );
  XOR2_X1 U11180 ( .A(n10444), .B(n10443), .Z(n10445) );
  NAND2_X1 U11181 ( .A1(n10445), .A2(n10519), .ZN(n10446) );
  NAND2_X1 U11182 ( .A1(n10447), .A2(n10446), .ZN(P2_U3184) );
  INV_X1 U11183 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10468) );
  AOI21_X1 U11184 ( .B1(n10449), .B2(n6316), .A(n10448), .ZN(n10452) );
  INV_X1 U11185 ( .A(n10450), .ZN(n10451) );
  OAI21_X1 U11186 ( .B1(n10496), .B2(n10452), .A(n10451), .ZN(n10453) );
  INV_X1 U11187 ( .A(n10453), .ZN(n10458) );
  AND2_X1 U11188 ( .A1(n10454), .A2(n6315), .ZN(n10455) );
  OAI21_X1 U11189 ( .B1(n10456), .B2(n10455), .A(n10492), .ZN(n10457) );
  OAI211_X1 U11190 ( .C1(n10511), .C2(n10459), .A(n10458), .B(n10457), .ZN(
        n10460) );
  INV_X1 U11191 ( .A(n10460), .ZN(n10467) );
  AOI21_X1 U11192 ( .B1(n10463), .B2(n10462), .A(n10461), .ZN(n10465) );
  OR2_X1 U11193 ( .A1(n10465), .A2(n10464), .ZN(n10466) );
  OAI211_X1 U11194 ( .C1(n10468), .C2(n10506), .A(n10467), .B(n10466), .ZN(
        P2_U3185) );
  AOI21_X1 U11195 ( .B1(n5041), .B2(n10470), .A(n10469), .ZN(n10472) );
  OAI22_X1 U11196 ( .A1(n10514), .A2(n10472), .B1(n10471), .B2(n10511), .ZN(
        n10473) );
  AOI21_X1 U11197 ( .B1(n10516), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n10473), .ZN(
        n10484) );
  OAI211_X1 U11198 ( .C1(n10476), .C2(n10475), .A(n10474), .B(n10519), .ZN(
        n10482) );
  AOI21_X1 U11199 ( .B1(n10479), .B2(n10478), .A(n10477), .ZN(n10480) );
  OR2_X1 U11200 ( .A1(n10496), .A2(n10480), .ZN(n10481) );
  NAND4_X1 U11201 ( .A1(n10484), .A2(n10483), .A3(n10482), .A4(n10481), .ZN(
        P2_U3186) );
  INV_X1 U11202 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10507) );
  AOI21_X1 U11203 ( .B1(n10486), .B2(n5816), .A(n10485), .ZN(n10497) );
  NAND2_X1 U11204 ( .A1(n10487), .A2(n5812), .ZN(n10490) );
  INV_X1 U11205 ( .A(n10488), .ZN(n10489) );
  NAND2_X1 U11206 ( .A1(n10490), .A2(n10489), .ZN(n10491) );
  NAND2_X1 U11207 ( .A1(n10492), .A2(n10491), .ZN(n10495) );
  INV_X1 U11208 ( .A(n10493), .ZN(n10494) );
  OAI211_X1 U11209 ( .C1(n10497), .C2(n10496), .A(n10495), .B(n10494), .ZN(
        n10500) );
  NOR2_X1 U11210 ( .A1(n10511), .A2(n10498), .ZN(n10499) );
  NOR2_X1 U11211 ( .A1(n10500), .A2(n10499), .ZN(n10505) );
  XOR2_X1 U11212 ( .A(n10501), .B(n10502), .Z(n10503) );
  NAND2_X1 U11213 ( .A1(n10503), .A2(n10519), .ZN(n10504) );
  OAI211_X1 U11214 ( .C1(n10507), .C2(n10506), .A(n10505), .B(n10504), .ZN(
        P2_U3187) );
  AOI21_X1 U11215 ( .B1(n10510), .B2(n10509), .A(n10508), .ZN(n10513) );
  OAI22_X1 U11216 ( .A1(n10514), .A2(n10513), .B1(n10512), .B2(n10511), .ZN(
        n10515) );
  AOI21_X1 U11217 ( .B1(n10516), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n10515), .ZN(
        n10529) );
  XOR2_X1 U11218 ( .A(n10517), .B(n10518), .Z(n10520) );
  NAND2_X1 U11219 ( .A1(n10520), .A2(n10519), .ZN(n10527) );
  OAI21_X1 U11220 ( .B1(n10523), .B2(n10522), .A(n10521), .ZN(n10524) );
  NAND2_X1 U11221 ( .A1(n10525), .A2(n10524), .ZN(n10526) );
  NAND4_X1 U11222 ( .A1(n10529), .A2(n10528), .A3(n10527), .A4(n10526), .ZN(
        P2_U3188) );
  XOR2_X1 U11223 ( .A(P1_RD_REG_SCAN_IN), .B(n10530), .Z(U126) );
  AOI21_X1 U11224 ( .B1(n10532), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n10531), .ZN(
        n10550) );
  OAI21_X1 U11225 ( .B1(n10535), .B2(n10534), .A(n10533), .ZN(n10545) );
  INV_X1 U11226 ( .A(n10536), .ZN(n10537) );
  OAI211_X1 U11227 ( .C1(n10540), .C2(n10539), .A(n10538), .B(n10537), .ZN(
        n10544) );
  NAND2_X1 U11228 ( .A1(n10542), .A2(n10541), .ZN(n10543) );
  OAI211_X1 U11229 ( .C1(n10546), .C2(n10545), .A(n10544), .B(n10543), .ZN(
        n10547) );
  INV_X1 U11230 ( .A(n10547), .ZN(n10549) );
  NAND3_X1 U11231 ( .A1(n10550), .A2(n10549), .A3(n10548), .ZN(P1_U3247) );
  NOR2_X1 U11232 ( .A1(n10552), .A2(n10551), .ZN(n10565) );
  NOR2_X1 U11233 ( .A1(n10554), .A2(n10553), .ZN(n10558) );
  NOR2_X1 U11234 ( .A1(n10562), .A2(n10555), .ZN(n10557) );
  MUX2_X1 U11235 ( .A(n10558), .B(n10557), .S(n10556), .Z(n10559) );
  AOI211_X1 U11236 ( .C1(n10775), .C2(P1_REG3_REG_0__SCAN_IN), .A(n10565), .B(
        n10559), .ZN(n10561) );
  AOI22_X1 U11237 ( .A1(n10786), .A2(n6477), .B1(n10561), .B2(n10560), .ZN(
        P1_U3293) );
  AOI21_X1 U11238 ( .B1(n10563), .B2(n10623), .A(n10562), .ZN(n10564) );
  AOI211_X1 U11239 ( .C1(n10567), .C2(n10566), .A(n10565), .B(n10564), .ZN(
        n10570) );
  AOI22_X1 U11240 ( .A1(n10770), .A2(n10570), .B1(n10568), .B2(n10768), .ZN(
        P1_U3522) );
  INV_X1 U11241 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U11242 ( .A1(n10774), .A2(n10570), .B1(n10569), .B2(n10771), .ZN(
        P1_U3453) );
  NOR2_X1 U11243 ( .A1(n10571), .A2(n10799), .ZN(n10573) );
  AOI211_X1 U11244 ( .C1(n10720), .C2(n10574), .A(n10573), .B(n10572), .ZN(
        n10576) );
  AOI22_X1 U11245 ( .A1(n10806), .A2(n10576), .B1(n10575), .B2(n10805), .ZN(
        P2_U3460) );
  AOI22_X1 U11246 ( .A1(n10810), .A2(n10576), .B1(n5750), .B2(n10807), .ZN(
        P2_U3393) );
  OAI21_X1 U11247 ( .B1(n10578), .B2(n10765), .A(n10577), .ZN(n10580) );
  AOI211_X1 U11248 ( .C1(n10767), .C2(n10581), .A(n10580), .B(n10579), .ZN(
        n10584) );
  INV_X1 U11249 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10582) );
  AOI22_X1 U11250 ( .A1(n10770), .A2(n10584), .B1(n10582), .B2(n10768), .ZN(
        P1_U3524) );
  INV_X1 U11251 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10583) );
  AOI22_X1 U11252 ( .A1(n10774), .A2(n10584), .B1(n10583), .B2(n10771), .ZN(
        P1_U3459) );
  XNOR2_X1 U11253 ( .A(n10585), .B(n10587), .ZN(n10603) );
  NAND3_X1 U11254 ( .A1(n10588), .A2(n10587), .A3(n10586), .ZN(n10589) );
  NAND2_X1 U11255 ( .A1(n10590), .A2(n10589), .ZN(n10593) );
  AOI222_X1 U11256 ( .A1(n10641), .A2(n10593), .B1(n10592), .B2(n6190), .C1(
        n10591), .C2(n10637), .ZN(n10600) );
  OAI21_X1 U11257 ( .B1(n10599), .B2(n10799), .A(n10600), .ZN(n10594) );
  AOI21_X1 U11258 ( .B1(n10603), .B2(n10720), .A(n10594), .ZN(n10596) );
  AOI22_X1 U11259 ( .A1(n10748), .A2(n10596), .B1(n6245), .B2(n10805), .ZN(
        P2_U3461) );
  INV_X1 U11260 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U11261 ( .A1(n10810), .A2(n10596), .B1(n10595), .B2(n10807), .ZN(
        P2_U3396) );
  OAI22_X1 U11262 ( .A1(n10599), .A2(n10598), .B1(n10597), .B2(n10650), .ZN(
        n10602) );
  INV_X1 U11263 ( .A(n10600), .ZN(n10601) );
  AOI211_X1 U11264 ( .C1(n10603), .C2(n10700), .A(n10602), .B(n10601), .ZN(
        n10604) );
  AOI22_X1 U11265 ( .A1(n9017), .A2(n6271), .B1(n10604), .B2(n10709), .ZN(
        P2_U3231) );
  NOR2_X1 U11266 ( .A1(n10605), .A2(n10799), .ZN(n10607) );
  AOI211_X1 U11267 ( .C1(n10608), .C2(n10720), .A(n10607), .B(n10606), .ZN(
        n10610) );
  AOI22_X1 U11268 ( .A1(n10748), .A2(n10610), .B1(n6315), .B2(n10805), .ZN(
        P2_U3462) );
  INV_X1 U11269 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U11270 ( .A1(n10810), .A2(n10610), .B1(n10609), .B2(n10807), .ZN(
        P2_U3399) );
  OAI21_X1 U11271 ( .B1(n10612), .B2(n10799), .A(n10611), .ZN(n10613) );
  AOI21_X1 U11272 ( .B1(n10720), .B2(n10614), .A(n10613), .ZN(n10616) );
  AOI22_X1 U11273 ( .A1(n10748), .A2(n10616), .B1(n10615), .B2(n10805), .ZN(
        P2_U3463) );
  AOI22_X1 U11274 ( .A1(n10810), .A2(n10616), .B1(n5798), .B2(n10807), .ZN(
        P2_U3402) );
  AOI21_X1 U11275 ( .B1(n10619), .B2(n10618), .A(n10617), .ZN(n10620) );
  OAI211_X1 U11276 ( .C1(n10623), .C2(n10622), .A(n10621), .B(n10620), .ZN(
        n10624) );
  INV_X1 U11277 ( .A(n10624), .ZN(n10627) );
  AOI22_X1 U11278 ( .A1(n10770), .A2(n10627), .B1(n10625), .B2(n10768), .ZN(
        P1_U3526) );
  INV_X1 U11279 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U11280 ( .A1(n10774), .A2(n10627), .B1(n10626), .B2(n10771), .ZN(
        P1_U3465) );
  NAND2_X1 U11281 ( .A1(n10629), .A2(n10628), .ZN(n10630) );
  XOR2_X1 U11282 ( .A(n10632), .B(n10630), .Z(n10642) );
  AOI21_X1 U11283 ( .B1(n10633), .B2(n10632), .A(n10631), .ZN(n10649) );
  INV_X1 U11284 ( .A(n10634), .ZN(n10639) );
  AOI22_X1 U11285 ( .A1(n10637), .A2(n10636), .B1(n10635), .B2(n6190), .ZN(
        n10638) );
  OAI21_X1 U11286 ( .B1(n10649), .B2(n10639), .A(n10638), .ZN(n10640) );
  AOI21_X1 U11287 ( .B1(n10642), .B2(n10641), .A(n10640), .ZN(n10657) );
  INV_X1 U11288 ( .A(n10657), .ZN(n10645) );
  OAI22_X1 U11289 ( .A1(n10649), .A2(n10643), .B1(n10652), .B2(n10799), .ZN(
        n10644) );
  NOR2_X1 U11290 ( .A1(n10645), .A2(n10644), .ZN(n10647) );
  AOI22_X1 U11291 ( .A1(n10748), .A2(n10647), .B1(n5812), .B2(n10805), .ZN(
        P2_U3464) );
  INV_X1 U11292 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U11293 ( .A1(n10810), .A2(n10647), .B1(n10646), .B2(n10807), .ZN(
        P2_U3405) );
  NOR3_X1 U11294 ( .A1(n10649), .A2(n9017), .A3(n10648), .ZN(n10655) );
  OAI22_X1 U11295 ( .A1(n10653), .A2(n10652), .B1(n10651), .B2(n10650), .ZN(
        n10654) );
  NOR2_X1 U11296 ( .A1(n10655), .A2(n10654), .ZN(n10656) );
  OAI221_X1 U11297 ( .B1(n9017), .B2(n10657), .C1(n10709), .C2(n5816), .A(
        n10656), .ZN(P2_U3228) );
  NOR2_X1 U11298 ( .A1(n10659), .A2(n10658), .ZN(n10664) );
  AOI22_X1 U11299 ( .A1(n10786), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n10660), 
        .B2(n10775), .ZN(n10661) );
  OAI21_X1 U11300 ( .B1(n10662), .B2(n9976), .A(n10661), .ZN(n10663) );
  AOI211_X1 U11301 ( .C1(n10665), .C2(n10781), .A(n10664), .B(n10663), .ZN(
        n10666) );
  OAI21_X1 U11302 ( .B1(n10786), .B2(n10667), .A(n10666), .ZN(P1_U3288) );
  OAI22_X1 U11303 ( .A1(n10669), .A2(n10801), .B1(n10668), .B2(n10799), .ZN(
        n10672) );
  INV_X1 U11304 ( .A(n10670), .ZN(n10671) );
  NOR2_X1 U11305 ( .A1(n10672), .A2(n10671), .ZN(n10674) );
  AOI22_X1 U11306 ( .A1(n10748), .A2(n10674), .B1(n6314), .B2(n10805), .ZN(
        P2_U3465) );
  INV_X1 U11307 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U11308 ( .A1(n10810), .A2(n10674), .B1(n10673), .B2(n10807), .ZN(
        P2_U3408) );
  OAI21_X1 U11309 ( .B1(n10676), .B2(n10765), .A(n10675), .ZN(n10678) );
  AOI211_X1 U11310 ( .C1(n10693), .C2(n10679), .A(n10678), .B(n10677), .ZN(
        n10682) );
  INV_X1 U11311 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U11312 ( .A1(n10770), .A2(n10682), .B1(n10680), .B2(n10768), .ZN(
        P1_U3528) );
  INV_X1 U11313 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U11314 ( .A1(n10774), .A2(n10682), .B1(n10681), .B2(n10771), .ZN(
        P1_U3471) );
  NOR3_X1 U11315 ( .A1(n10684), .A2(n10683), .A3(n10801), .ZN(n10686) );
  AOI211_X1 U11316 ( .C1(n10747), .C2(n10687), .A(n10686), .B(n10685), .ZN(
        n10689) );
  AOI22_X1 U11317 ( .A1(n10748), .A2(n10689), .B1(n6312), .B2(n10805), .ZN(
        P2_U3466) );
  INV_X1 U11318 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U11319 ( .A1(n10810), .A2(n10689), .B1(n10688), .B2(n10807), .ZN(
        P2_U3411) );
  OAI21_X1 U11320 ( .B1(n10691), .B2(n10765), .A(n10690), .ZN(n10692) );
  AOI21_X1 U11321 ( .B1(n10694), .B2(n10693), .A(n10692), .ZN(n10695) );
  AND2_X1 U11322 ( .A1(n10696), .A2(n10695), .ZN(n10699) );
  INV_X1 U11323 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U11324 ( .A1(n10770), .A2(n10699), .B1(n10697), .B2(n10768), .ZN(
        P1_U3530) );
  INV_X1 U11325 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U11326 ( .A1(n10774), .A2(n10699), .B1(n10698), .B2(n10771), .ZN(
        P1_U3477) );
  INV_X1 U11327 ( .A(n10700), .ZN(n10703) );
  OAI21_X1 U11328 ( .B1(n10703), .B2(n10702), .A(n10701), .ZN(n10708) );
  AOI222_X1 U11329 ( .A1(n10709), .A2(n10708), .B1(n10707), .B2(n10706), .C1(
        n10705), .C2(n10704), .ZN(n10710) );
  OAI21_X1 U11330 ( .B1(n10709), .B2(n6311), .A(n10710), .ZN(P2_U3225) );
  OAI211_X1 U11331 ( .C1(n10713), .C2(n10765), .A(n10712), .B(n10711), .ZN(
        n10714) );
  AOI21_X1 U11332 ( .B1(n10767), .B2(n10715), .A(n10714), .ZN(n10718) );
  AOI22_X1 U11333 ( .A1(n10770), .A2(n10718), .B1(n10716), .B2(n10768), .ZN(
        P1_U3531) );
  INV_X1 U11334 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U11335 ( .A1(n10774), .A2(n10718), .B1(n10717), .B2(n10771), .ZN(
        P1_U3480) );
  AND3_X1 U11336 ( .A1(n10721), .A2(n10720), .A3(n10719), .ZN(n10723) );
  AOI211_X1 U11337 ( .C1(n10747), .C2(n10724), .A(n10723), .B(n10722), .ZN(
        n10727) );
  AOI22_X1 U11338 ( .A1(n10748), .A2(n10727), .B1(n10725), .B2(n10805), .ZN(
        P2_U3468) );
  INV_X1 U11339 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U11340 ( .A1(n10810), .A2(n10727), .B1(n10726), .B2(n10807), .ZN(
        P2_U3417) );
  OAI21_X1 U11341 ( .B1(n10729), .B2(n10765), .A(n10728), .ZN(n10730) );
  AOI211_X1 U11342 ( .C1(n10732), .C2(n10767), .A(n10731), .B(n10730), .ZN(
        n10734) );
  AOI22_X1 U11343 ( .A1(n10770), .A2(n10734), .B1(n6665), .B2(n10768), .ZN(
        P1_U3532) );
  INV_X1 U11344 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U11345 ( .A1(n10774), .A2(n10734), .B1(n10733), .B2(n10771), .ZN(
        P1_U3483) );
  INV_X1 U11346 ( .A(n10735), .ZN(n10736) );
  NOR2_X1 U11347 ( .A1(n10736), .A2(n10799), .ZN(n10738) );
  AOI211_X1 U11348 ( .C1(n10740), .C2(n10739), .A(n10738), .B(n10737), .ZN(
        n10742) );
  AOI22_X1 U11349 ( .A1(n10806), .A2(n10742), .B1(n5903), .B2(n10805), .ZN(
        P2_U3469) );
  INV_X1 U11350 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U11351 ( .A1(n10810), .A2(n10742), .B1(n10741), .B2(n10807), .ZN(
        P2_U3420) );
  NOR2_X1 U11352 ( .A1(n10743), .A2(n10801), .ZN(n10744) );
  AOI211_X1 U11353 ( .C1(n10747), .C2(n10746), .A(n10745), .B(n10744), .ZN(
        n10750) );
  AOI22_X1 U11354 ( .A1(n10748), .A2(n10750), .B1(n5916), .B2(n10805), .ZN(
        P2_U3470) );
  INV_X1 U11355 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U11356 ( .A1(n10810), .A2(n10750), .B1(n10749), .B2(n10807), .ZN(
        P2_U3423) );
  XNOR2_X1 U11357 ( .A(n10751), .B(n10755), .ZN(n10782) );
  OAI211_X1 U11358 ( .C1(n10755), .C2(n10754), .A(n10753), .B(n10752), .ZN(
        n10761) );
  AOI22_X1 U11359 ( .A1(n10759), .A2(n10758), .B1(n10757), .B2(n10756), .ZN(
        n10760) );
  AND2_X1 U11360 ( .A1(n10761), .A2(n10760), .ZN(n10785) );
  OAI211_X1 U11361 ( .C1(n5540), .C2(n10764), .A(n10763), .B(n10762), .ZN(
        n10779) );
  OAI211_X1 U11362 ( .C1(n5540), .C2(n10765), .A(n10785), .B(n10779), .ZN(
        n10766) );
  AOI21_X1 U11363 ( .B1(n10782), .B2(n10767), .A(n10766), .ZN(n10773) );
  AOI22_X1 U11364 ( .A1(n10770), .A2(n10773), .B1(n10769), .B2(n10768), .ZN(
        P1_U3534) );
  INV_X1 U11365 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U11366 ( .A1(n10774), .A2(n10773), .B1(n10772), .B2(n10771), .ZN(
        P1_U3489) );
  AOI222_X1 U11367 ( .A1(n10778), .A2(n10777), .B1(n10776), .B2(n10775), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(n10786), .ZN(n10784) );
  INV_X1 U11368 ( .A(n10779), .ZN(n10780) );
  AOI22_X1 U11369 ( .A1(n10782), .A2(n10781), .B1(n10780), .B2(n9972), .ZN(
        n10783) );
  OAI211_X1 U11370 ( .C1(n10786), .C2(n10785), .A(n10784), .B(n10783), .ZN(
        P1_U3281) );
  OAI22_X1 U11371 ( .A1(n10788), .A2(n10801), .B1(n10787), .B2(n10799), .ZN(
        n10790) );
  NOR2_X1 U11372 ( .A1(n10790), .A2(n10789), .ZN(n10792) );
  AOI22_X1 U11373 ( .A1(n10806), .A2(n10792), .B1(n5946), .B2(n10805), .ZN(
        P2_U3472) );
  INV_X1 U11374 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U11375 ( .A1(n10810), .A2(n10792), .B1(n10791), .B2(n10807), .ZN(
        P2_U3429) );
  OAI22_X1 U11376 ( .A1(n10794), .A2(n10801), .B1(n10793), .B2(n10799), .ZN(
        n10796) );
  NOR2_X1 U11377 ( .A1(n10796), .A2(n10795), .ZN(n10798) );
  AOI22_X1 U11378 ( .A1(n10806), .A2(n10798), .B1(n5960), .B2(n10805), .ZN(
        P2_U3473) );
  INV_X1 U11379 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10797) );
  AOI22_X1 U11380 ( .A1(n10810), .A2(n10798), .B1(n10797), .B2(n10807), .ZN(
        P2_U3432) );
  OAI22_X1 U11381 ( .A1(n10802), .A2(n10801), .B1(n10800), .B2(n10799), .ZN(
        n10804) );
  NOR2_X1 U11382 ( .A1(n10804), .A2(n10803), .ZN(n10809) );
  AOI22_X1 U11383 ( .A1(n10806), .A2(n10809), .B1(n5977), .B2(n10805), .ZN(
        P2_U3474) );
  INV_X1 U11384 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U11385 ( .A1(n10810), .A2(n10809), .B1(n10808), .B2(n10807), .ZN(
        P2_U3435) );
  XNOR2_X1 U11386 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X1 U5025 ( .A(n7898), .Z(n8070) );
endmodule

