

module b22_C_SARLock_k_128_2 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628;

  OAI21_X1 U7317 ( .B1(n14980), .B2(n6913), .A(n6912), .ZN(n14759) );
  INV_X1 U7318 ( .A(n13292), .ZN(n13107) );
  AOI22_X1 U7319 ( .A1(n13223), .A2(n13049), .B1(n13078), .B2(n7531), .ZN(
        n13209) );
  NAND2_X1 U7320 ( .A1(n8426), .A2(n8425), .ZN(n13330) );
  INV_X2 U7321 ( .A(n12044), .ZN(n12070) );
  CLKBUF_X2 U7322 ( .A(n8795), .Z(n6570) );
  CLKBUF_X2 U7323 ( .A(n8795), .Z(n6569) );
  INV_X1 U7324 ( .A(n13850), .ZN(n13524) );
  NAND2_X1 U7325 ( .A1(n14564), .A2(n11694), .ZN(n10020) );
  NAND2_X1 U7326 ( .A1(n7919), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7253) );
  NAND2_X1 U7327 ( .A1(n7730), .A2(n7729), .ZN(n7728) );
  NAND2_X1 U7328 ( .A1(n13073), .A2(n13072), .ZN(n13245) );
  NAND2_X1 U7329 ( .A1(n13080), .A2(n13079), .ZN(n13197) );
  NAND2_X1 U7330 ( .A1(n11061), .A2(n11060), .ZN(n11190) );
  INV_X1 U7331 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7992) );
  NAND2_X2 U7332 ( .A1(n10020), .A2(n6568), .ZN(n13850) );
  CLKBUF_X2 U7333 ( .A(n10717), .Z(n13607) );
  NAND2_X1 U7334 ( .A1(n14672), .A2(n14673), .ZN(n14674) );
  INV_X1 U7335 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8709) );
  INV_X1 U7336 ( .A(n11315), .ZN(n12806) );
  BUF_X1 U7337 ( .A(n10289), .Z(n12824) );
  INV_X1 U7338 ( .A(n7965), .ZN(n8611) );
  NAND2_X1 U7339 ( .A1(n13268), .A2(n13267), .ZN(n13266) );
  INV_X1 U7340 ( .A(n10020), .ZN(n13523) );
  NAND2_X1 U7341 ( .A1(n9993), .A2(n11698), .ZN(n13842) );
  INV_X1 U7342 ( .A(n13844), .ZN(n13832) );
  XNOR2_X1 U7343 ( .A(n14674), .B(n7468), .ZN(n14710) );
  OR2_X1 U7344 ( .A1(n8758), .A2(n8709), .ZN(n8738) );
  NAND2_X1 U7345 ( .A1(n9991), .A2(n9993), .ZN(n13692) );
  INV_X1 U7346 ( .A(n15147), .ZN(n15076) );
  AOI21_X2 U7347 ( .B1(n9361), .B2(n12636), .A(n9360), .ZN(n11715) );
  OR2_X2 U7348 ( .A1(n6911), .A2(n14965), .ZN(n7454) );
  XNOR2_X2 U7349 ( .A(n7253), .B(P2_IR_REG_29__SCAN_IN), .ZN(n7906) );
  NOR2_X2 U7350 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n7934) );
  AND4_X4 U7351 ( .A1(n6622), .A2(n9395), .A3(n7810), .A4(n9448), .ZN(n10332)
         );
  NOR2_X2 U7352 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9448) );
  NAND2_X2 U7353 ( .A1(n13395), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7904) );
  NAND2_X2 U7354 ( .A1(n14776), .A2(n14742), .ZN(n14784) );
  AOI21_X1 U7355 ( .B1(n8280), .B2(n7758), .A(n7756), .ZN(n7277) );
  NAND2_X1 U7356 ( .A1(n10020), .A2(n10019), .ZN(n13836) );
  XNOR2_X2 U7357 ( .A(n8738), .B(n8757), .ZN(n9254) );
  XNOR2_X2 U7358 ( .A(n14726), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14727) );
  XNOR2_X2 U7359 ( .A(n14676), .B(n7466), .ZN(n14726) );
  OAI21_X4 U7360 ( .B1(n9376), .B2(n12079), .A(n8736), .ZN(n8804) );
  INV_X2 U7361 ( .A(n10019), .ZN(n6568) );
  INV_X4 U7362 ( .A(n7353), .ZN(n13436) );
  INV_X2 U7363 ( .A(n10019), .ZN(n8510) );
  NAND2_X1 U7364 ( .A1(n10163), .A2(n13436), .ZN(n8795) );
  INV_X1 U7365 ( .A(n8092), .ZN(n6571) );
  AND2_X1 U7366 ( .A1(n13402), .A2(n7907), .ZN(n7996) );
  OAI21_X2 U7367 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n14753), .A(n14976), .ZN(
        n14980) );
  NAND2_X1 U7368 ( .A1(n11309), .A2(n7536), .ZN(n11502) );
  INV_X2 U7369 ( .A(n8803), .ZN(n10473) );
  INV_X2 U7370 ( .A(n8804), .ZN(n8803) );
  INV_X2 U7371 ( .A(n8592), .ZN(n8617) );
  INV_X2 U7372 ( .A(n14021), .ZN(n14029) );
  INV_X4 U7373 ( .A(n8790), .ZN(n8962) );
  CLKBUF_X2 U7374 ( .A(n6603), .Z(n8586) );
  NAND2_X1 U7375 ( .A1(n9990), .A2(n9991), .ZN(n10037) );
  CLKBUF_X1 U7376 ( .A(n14564), .Z(n6573) );
  INV_X1 U7377 ( .A(n13436), .ZN(n10019) );
  NOR2_X2 U7378 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7966) );
  OR2_X1 U7379 ( .A1(n9389), .A2(n15601), .ZN(n9374) );
  OAI21_X1 U7380 ( .B1(n14910), .B2(n11716), .A(n11715), .ZN(n9389) );
  NOR2_X1 U7381 ( .A1(n8671), .A2(n9696), .ZN(n7167) );
  OAI21_X1 U7382 ( .B1(n6677), .B2(n6763), .A(n6589), .ZN(n8671) );
  NAND2_X1 U7383 ( .A1(n7162), .A2(n7161), .ZN(n6763) );
  XNOR2_X1 U7384 ( .A(n11877), .B(n9297), .ZN(n11716) );
  OAI21_X1 U7385 ( .B1(n7139), .B2(n7137), .A(n7140), .ZN(n7168) );
  OR2_X1 U7386 ( .A1(n12427), .A2(n12428), .ZN(n7203) );
  AOI21_X1 U7387 ( .B1(n7581), .B2(n6733), .A(n7579), .ZN(n7578) );
  NOR2_X1 U7388 ( .A1(n12457), .A2(n12052), .ZN(n12445) );
  OR2_X1 U7389 ( .A1(n12459), .A2(n12458), .ZN(n7011) );
  OAI211_X1 U7390 ( .C1(n12818), .C2(n6922), .A(n6921), .B(n12880), .ZN(n12883) );
  NAND2_X1 U7391 ( .A1(n14807), .A2(n14805), .ZN(n14811) );
  AOI21_X1 U7392 ( .B1(n7235), .B2(n7233), .A(n6697), .ZN(n7232) );
  NAND2_X1 U7393 ( .A1(n13161), .A2(n13146), .ZN(n13141) );
  AND2_X1 U7394 ( .A1(n7238), .A2(n6704), .ZN(n7235) );
  OAI21_X1 U7395 ( .B1(n9339), .B2(n7087), .A(n7085), .ZN(n12520) );
  XNOR2_X1 U7396 ( .A(n8560), .B(n8559), .ZN(n14560) );
  NAND2_X1 U7397 ( .A1(n13679), .A2(n13678), .ZN(n14452) );
  NAND2_X1 U7398 ( .A1(n7532), .A2(n7531), .ZN(n13217) );
  OR2_X1 U7399 ( .A1(n9147), .A2(n13416), .ZN(n9160) );
  XNOR2_X1 U7400 ( .A(n8569), .B(n8568), .ZN(n13676) );
  NAND2_X1 U7401 ( .A1(n8494), .A2(n8493), .ZN(n13313) );
  NAND2_X1 U7402 ( .A1(n11507), .A2(n11506), .ZN(n11509) );
  NAND2_X1 U7403 ( .A1(n13600), .A2(n13599), .ZN(n14472) );
  OR2_X1 U7404 ( .A1(n11307), .A2(n11306), .ZN(n11507) );
  AND2_X1 U7405 ( .A1(n7326), .A2(n7325), .ZN(n11576) );
  XNOR2_X1 U7406 ( .A(n7362), .B(n8486), .ZN(n13582) );
  OAI21_X1 U7407 ( .B1(n11190), .B2(n11195), .A(n11196), .ZN(n7330) );
  OAI21_X1 U7408 ( .B1(n9106), .B2(n13542), .A(n9109), .ZN(n9115) );
  OR2_X1 U7409 ( .A1(n13196), .A2(n7725), .ZN(n7724) );
  NAND2_X1 U7410 ( .A1(n7535), .A2(n7539), .ZN(n11585) );
  INV_X1 U7411 ( .A(n11502), .ZN(n7535) );
  NAND2_X1 U7412 ( .A1(n6698), .A2(n7296), .ZN(n11319) );
  NAND2_X1 U7413 ( .A1(n10987), .A2(n10986), .ZN(n11065) );
  NAND2_X1 U7414 ( .A1(n8462), .A2(n8461), .ZN(n8465) );
  AND2_X2 U7415 ( .A1(n7538), .A2(n7537), .ZN(n11309) );
  NAND2_X1 U7416 ( .A1(n8381), .A2(n8380), .ZN(n13343) );
  OR2_X1 U7417 ( .A1(n10747), .A2(n10984), .ZN(n10989) );
  OAI21_X1 U7418 ( .B1(n13437), .B2(n8440), .A(n8442), .ZN(n8462) );
  OAI21_X1 U7419 ( .B1(n11350), .B2(n11977), .A(n11609), .ZN(n9270) );
  XNOR2_X1 U7420 ( .A(n8441), .B(SI_22_), .ZN(n13437) );
  NAND2_X1 U7421 ( .A1(n8363), .A2(n8362), .ZN(n13348) );
  OAI21_X1 U7422 ( .B1(n7633), .B2(n8357), .A(n7631), .ZN(n8441) );
  CLKBUF_X2 U7423 ( .A(n12429), .Z(n6575) );
  OAI21_X1 U7424 ( .B1(n6615), .B2(n7633), .A(n8424), .ZN(n7632) );
  NAND2_X1 U7425 ( .A1(n7065), .A2(n7063), .ZN(n11275) );
  OR2_X1 U7426 ( .A1(n8353), .A2(n6997), .ZN(n8357) );
  OR2_X1 U7427 ( .A1(n10829), .A2(n6630), .ZN(n7065) );
  NAND2_X2 U7428 ( .A1(n8119), .A2(n8118), .ZN(n10647) );
  NOR2_X1 U7429 ( .A1(n9196), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9247) );
  OR2_X1 U7430 ( .A1(n9180), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9196) );
  NAND2_X1 U7431 ( .A1(n7185), .A2(n6659), .ZN(n7461) );
  NAND2_X1 U7432 ( .A1(n8130), .A2(n8114), .ZN(n10870) );
  NAND2_X1 U7433 ( .A1(n8138), .A2(n8137), .ZN(n10745) );
  OR2_X1 U7434 ( .A1(n14775), .A2(n14774), .ZN(n7185) );
  NAND2_X1 U7435 ( .A1(n8083), .A2(n8109), .ZN(n10857) );
  NAND2_X1 U7436 ( .A1(n8064), .A2(n8063), .ZN(n15365) );
  INV_X1 U7437 ( .A(n10252), .ZN(n6572) );
  NOR2_X1 U7438 ( .A1(n9364), .A2(n9260), .ZN(n11868) );
  AND4_X1 U7439 ( .A1(n8824), .A2(n8823), .A3(n8822), .A4(n8821), .ZN(n10964)
         );
  NAND2_X1 U7440 ( .A1(n7995), .A2(n7994), .ZN(n15348) );
  NOR2_X2 U7441 ( .A1(n7010), .A2(n6618), .ZN(n8812) );
  AND2_X1 U7442 ( .A1(n7607), .A2(n7359), .ZN(n7358) );
  AND4_X1 U7443 ( .A1(n8842), .A2(n8841), .A3(n8840), .A4(n8839), .ZN(n11206)
         );
  NAND4_X1 U7444 ( .A1(n8001), .A2(n8000), .A3(n7999), .A4(n7998), .ZN(n12991)
         );
  NAND2_X1 U7445 ( .A1(n7968), .A2(n7969), .ZN(n7166) );
  NAND2_X1 U7446 ( .A1(n6675), .A2(n8020), .ZN(n12990) );
  AOI21_X1 U7447 ( .B1(n7639), .B2(n7644), .A(SI_27_), .ZN(n7638) );
  INV_X2 U7448 ( .A(n7009), .ZN(n8788) );
  OAI21_X1 U7449 ( .B1(n6710), .B2(n7611), .A(n8307), .ZN(n7610) );
  CLKBUF_X1 U7450 ( .A(n10721), .Z(n13626) );
  OAI21_X1 U7451 ( .B1(n8848), .B2(n7386), .A(n7384), .ZN(n8879) );
  NAND2_X2 U7452 ( .A1(n14015), .A2(n13866), .ZN(n14021) );
  AOI21_X1 U7453 ( .B1(n8172), .B2(n7616), .A(n6692), .ZN(n7614) );
  INV_X2 U7454 ( .A(n10072), .ZN(n13627) );
  AND2_X2 U7455 ( .A1(n8766), .A2(n12781), .ZN(n9354) );
  NAND2_X1 U7456 ( .A1(n10163), .A2(n10019), .ZN(n8799) );
  NAND2_X2 U7457 ( .A1(n9254), .A2(n9255), .ZN(n10163) );
  NAND2_X1 U7458 ( .A1(n9986), .A2(n13856), .ZN(n10072) );
  INV_X1 U7459 ( .A(n10146), .ZN(n11403) );
  NOR2_X1 U7460 ( .A1(n7906), .A2(n7907), .ZN(n6603) );
  NAND2_X1 U7461 ( .A1(n9990), .A2(n11698), .ZN(n13844) );
  NAND2_X1 U7462 ( .A1(n9939), .A2(n7288), .ZN(n9712) );
  OR2_X2 U7463 ( .A1(n14022), .A2(n15139), .ZN(n15147) );
  XNOR2_X1 U7464 ( .A(n8760), .B(n12774), .ZN(n8766) );
  NAND2_X1 U7465 ( .A1(n7586), .A2(n7938), .ZN(n10146) );
  OAI21_X1 U7466 ( .B1(n6637), .B2(n8715), .A(n6846), .ZN(n11932) );
  CLKBUF_X1 U7467 ( .A(n8618), .Z(n9939) );
  INV_X1 U7468 ( .A(n8260), .ZN(n8284) );
  NAND2_X2 U7469 ( .A1(n7928), .A2(n7940), .ZN(n10945) );
  NAND2_X1 U7470 ( .A1(n8762), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8760) );
  INV_X2 U7471 ( .A(n14559), .ZN(n11699) );
  NOR2_X1 U7472 ( .A1(n6568), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14780) );
  AND3_X1 U7473 ( .A1(n8672), .A2(n7933), .A3(n7932), .ZN(n9938) );
  XNOR2_X1 U7474 ( .A(n14671), .B(n7187), .ZN(n14713) );
  INV_X1 U7475 ( .A(n7453), .ZN(n7098) );
  NOR2_X1 U7476 ( .A1(n7452), .A2(n7453), .ZN(n8758) );
  NAND2_X1 U7477 ( .A1(n14669), .A2(n7188), .ZN(n14671) );
  NOR2_X1 U7478 ( .A1(n7901), .A2(n7914), .ZN(n7902) );
  NAND2_X1 U7479 ( .A1(n10332), .A2(n6627), .ZN(n9664) );
  NAND4_X1 U7480 ( .A1(n6820), .A2(n6819), .A3(n8702), .A4(n6818), .ZN(n8703)
         );
  AND4_X1 U7481 ( .A1(n8716), .A2(n9223), .A3(n8715), .A4(n8714), .ZN(n8717)
         );
  AND2_X1 U7482 ( .A1(n8700), .A2(n8701), .ZN(n7863) );
  AND2_X1 U7483 ( .A1(n6910), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14717) );
  AND2_X2 U7484 ( .A1(n7966), .A2(n7896), .ZN(n8179) );
  AND4_X1 U7485 ( .A1(n9394), .A2(n9393), .A3(n9392), .A4(n7814), .ZN(n7810)
         );
  XNOR2_X1 U7486 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n14716) );
  NOR2_X1 U7487 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n8716) );
  INV_X1 U7488 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n12378) );
  INV_X1 U7489 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8693) );
  NOR2_X1 U7490 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n7889) );
  NOR2_X1 U7491 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7888) );
  INV_X1 U7492 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8920) );
  NOR2_X1 U7493 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n6819) );
  INV_X1 U7494 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8289) );
  NOR2_X1 U7495 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8773) );
  INV_X4 U7496 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7497 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8701) );
  XNOR2_X1 U7498 ( .A(n6793), .B(n9665), .ZN(n14564) );
  AOI21_X2 U7499 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(n14743), .A(n14783), .ZN(
        n14793) );
  XNOR2_X2 U7500 ( .A(n6791), .B(n9987), .ZN(n11694) );
  NOR2_X2 U7501 ( .A1(n13271), .A2(n13353), .ZN(n7534) );
  INV_X4 U7502 ( .A(n7997), .ZN(n8564) );
  CLKBUF_X2 U7503 ( .A(n8645), .Z(n6574) );
  OAI211_X1 U7504 ( .C1(n8611), .C2(n10021), .A(n7952), .B(n7951), .ZN(n8645)
         );
  NAND2_X1 U7505 ( .A1(n8617), .A2(n12986), .ZN(n7176) );
  NAND2_X1 U7506 ( .A1(n10647), .A2(n8615), .ZN(n7177) );
  INV_X1 U7507 ( .A(n8766), .ZN(n8764) );
  AOI21_X1 U7508 ( .B1(n6579), .B2(n6928), .A(n6694), .ZN(n6927) );
  INV_X1 U7509 ( .A(n7568), .ZN(n6928) );
  OR2_X1 U7510 ( .A1(n12938), .A2(n12941), .ZN(n12811) );
  NAND2_X1 U7511 ( .A1(n7732), .A2(n7731), .ZN(n7730) );
  INV_X1 U7512 ( .A(n13154), .ZN(n7731) );
  NAND2_X1 U7513 ( .A1(n14358), .A2(n14172), .ZN(n7698) );
  NAND2_X1 U7514 ( .A1(n7008), .A2(n8766), .ZN(n7009) );
  AND2_X1 U7515 ( .A1(n7855), .A2(n9345), .ZN(n7076) );
  INV_X1 U7516 ( .A(n8799), .ZN(n11887) );
  INV_X1 U7518 ( .A(n8586), .ZN(n8614) );
  INV_X1 U7519 ( .A(n8611), .ZN(n8400) );
  NOR2_X1 U7520 ( .A1(n6631), .A2(n7806), .ZN(n13268) );
  AND2_X1 U7521 ( .A1(n13069), .A2(n13065), .ZN(n7806) );
  NAND2_X1 U7522 ( .A1(n6950), .A2(n6948), .ZN(n14229) );
  OR2_X1 U7523 ( .A1(n6591), .A2(n6632), .ZN(n6950) );
  NOR2_X1 U7524 ( .A1(n6951), .A2(n6632), .ZN(n6949) );
  NAND2_X1 U7525 ( .A1(n7166), .A2(n8635), .ZN(n7975) );
  AOI22_X1 U7526 ( .A1(n7166), .A2(n8615), .B1(n12992), .B2(n8635), .ZN(n7982)
         );
  NAND2_X1 U7527 ( .A1(n8002), .A2(n8003), .ZN(n8006) );
  NOR2_X1 U7528 ( .A1(n7561), .A2(n13903), .ZN(n7560) );
  NAND2_X1 U7529 ( .A1(n13902), .A2(n13901), .ZN(n13905) );
  INV_X1 U7530 ( .A(n6777), .ZN(n6774) );
  AND2_X1 U7531 ( .A1(n8152), .A2(n6580), .ZN(n7165) );
  NAND2_X1 U7532 ( .A1(n7754), .A2(n7753), .ZN(n7752) );
  INV_X1 U7533 ( .A(n8327), .ZN(n7754) );
  INV_X1 U7534 ( .A(n8326), .ZN(n7753) );
  NAND2_X1 U7535 ( .A1(n13959), .A2(n13960), .ZN(n13958) );
  NAND2_X1 U7536 ( .A1(n13976), .A2(n6790), .ZN(n6789) );
  NOR2_X1 U7537 ( .A1(n13974), .A2(n13975), .ZN(n7224) );
  AND2_X1 U7538 ( .A1(n7281), .A2(n7282), .ZN(n7280) );
  INV_X1 U7539 ( .A(n6713), .ZN(n7281) );
  NAND2_X1 U7540 ( .A1(n8458), .A2(n6713), .ZN(n7279) );
  NAND2_X1 U7541 ( .A1(n13992), .A2(n7217), .ZN(n7216) );
  NAND2_X1 U7542 ( .A1(n7146), .A2(n6588), .ZN(n8481) );
  OR2_X1 U7543 ( .A1(n12516), .A2(n12522), .ZN(n12033) );
  AND2_X1 U7544 ( .A1(n11911), .A2(n11951), .ZN(n7431) );
  INV_X1 U7545 ( .A(n9087), .ZN(n7109) );
  OAI21_X1 U7546 ( .B1(n7283), .B2(n6605), .A(n8526), .ZN(n7141) );
  INV_X1 U7547 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U7548 ( .A1(n7355), .A2(n7354), .ZN(n8355) );
  AOI21_X1 U7549 ( .B1(n7356), .B2(n7610), .A(n6691), .ZN(n7354) );
  AND2_X1 U7550 ( .A1(n7358), .A2(n6705), .ZN(n7356) );
  INV_X1 U7551 ( .A(n8288), .ZN(n7611) );
  AOI21_X1 U7552 ( .B1(n7614), .B2(n7615), .A(n7613), .ZN(n7612) );
  INV_X1 U7553 ( .A(n8220), .ZN(n7613) );
  AND2_X1 U7554 ( .A1(n6703), .A2(n7680), .ZN(n7679) );
  NAND2_X1 U7555 ( .A1(n11782), .A2(n12557), .ZN(n7680) );
  AND2_X1 U7556 ( .A1(n11932), .A2(n9353), .ZN(n9228) );
  NAND2_X1 U7557 ( .A1(n10380), .A2(n15453), .ZN(n7052) );
  OR2_X1 U7558 ( .A1(n9349), .A2(n12094), .ZN(n9350) );
  OR2_X1 U7559 ( .A1(n11742), .A2(n12495), .ZN(n12042) );
  NOR2_X1 U7560 ( .A1(n12611), .A2(n7440), .ZN(n7439) );
  NAND2_X1 U7561 ( .A1(n9327), .A2(n7095), .ZN(n7094) );
  NAND2_X1 U7562 ( .A1(n8812), .A2(n10704), .ZN(n11942) );
  NAND2_X1 U7563 ( .A1(n8806), .A2(n9302), .ZN(n11935) );
  AND2_X1 U7564 ( .A1(n10403), .A2(n14638), .ZN(n9382) );
  NAND2_X1 U7565 ( .A1(n8741), .A2(n8740), .ZN(n9255) );
  NAND2_X1 U7566 ( .A1(n8737), .A2(n6801), .ZN(n8741) );
  NOR2_X1 U7567 ( .A1(n7202), .A2(n8709), .ZN(n6801) );
  INV_X1 U7568 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8714) );
  INV_X1 U7569 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8708) );
  INV_X1 U7570 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7875) );
  AND2_X1 U7571 ( .A1(n7878), .A2(n6638), .ZN(n7683) );
  INV_X1 U7572 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U7573 ( .A1(n7582), .A2(n10283), .ZN(n7583) );
  NAND2_X1 U7574 ( .A1(n7164), .A2(n7163), .ZN(n7162) );
  INV_X1 U7575 ( .A(n8598), .ZN(n7163) );
  NAND2_X1 U7576 ( .A1(n8600), .A2(n8599), .ZN(n7164) );
  AND2_X1 U7577 ( .A1(n13318), .A2(n13052), .ZN(n7798) );
  INV_X1 U7578 ( .A(n7244), .ZN(n7241) );
  AND2_X1 U7579 ( .A1(n6702), .A2(n11067), .ZN(n7245) );
  NAND2_X1 U7580 ( .A1(n15358), .A2(n12990), .ZN(n7332) );
  AND2_X1 U7581 ( .A1(n7923), .A2(n6568), .ZN(n7965) );
  NAND2_X1 U7582 ( .A1(n13197), .A2(n13196), .ZN(n7723) );
  OR2_X1 U7583 ( .A1(n13353), .A2(n13042), .ZN(n7805) );
  AND2_X1 U7584 ( .A1(n7897), .A2(n6644), .ZN(n7319) );
  NAND2_X1 U7585 ( .A1(n7486), .A2(n7485), .ZN(n7484) );
  NAND2_X1 U7586 ( .A1(n7487), .A2(n7490), .ZN(n7485) );
  NAND2_X1 U7587 ( .A1(n7488), .A2(n13742), .ZN(n7486) );
  INV_X1 U7588 ( .A(n13714), .ZN(n7487) );
  AND2_X1 U7589 ( .A1(n7515), .A2(n11681), .ZN(n7514) );
  INV_X1 U7590 ( .A(n9990), .ZN(n9993) );
  INV_X1 U7591 ( .A(n11698), .ZN(n9991) );
  AND2_X1 U7592 ( .A1(n14323), .A2(n14196), .ZN(n7829) );
  INV_X1 U7593 ( .A(n6968), .ZN(n6967) );
  OAI21_X1 U7594 ( .B1(n6614), .B2(n6969), .A(n14185), .ZN(n6968) );
  AND2_X1 U7595 ( .A1(n7876), .A2(n11147), .ZN(n7714) );
  INV_X1 U7596 ( .A(n15060), .ZN(n13925) );
  INV_X1 U7597 ( .A(n10228), .ZN(n7819) );
  AND2_X1 U7598 ( .A1(n10026), .A2(n13856), .ZN(n13517) );
  NAND2_X1 U7599 ( .A1(n9981), .A2(n11298), .ZN(n14022) );
  NOR2_X1 U7600 ( .A1(n9660), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U7601 ( .A1(n7630), .A2(n8377), .ZN(n8420) );
  NAND2_X1 U7602 ( .A1(n8357), .A2(n6615), .ZN(n7630) );
  INV_X1 U7603 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9398) );
  NOR2_X1 U7604 ( .A1(n8990), .A2(n9329), .ZN(n7663) );
  OAI21_X1 U7605 ( .B1(n11864), .B2(n6833), .A(n6830), .ZN(n11745) );
  AOI21_X1 U7606 ( .B1(n6832), .B2(n6831), .A(n6636), .ZN(n6830) );
  NAND2_X1 U7607 ( .A1(n6840), .A2(n11756), .ZN(n6839) );
  AOI21_X1 U7608 ( .B1(n11562), .B2(n6576), .A(n6740), .ZN(n6845) );
  NAND2_X1 U7609 ( .A1(n8843), .A2(n11206), .ZN(n6828) );
  AND2_X1 U7610 ( .A1(n7409), .A2(n7408), .ZN(n12072) );
  AOI21_X1 U7611 ( .B1(n14899), .B2(n11898), .A(n11895), .ZN(n7408) );
  INV_X1 U7612 ( .A(n14638), .ZN(n11927) );
  OR2_X1 U7613 ( .A1(n12735), .A2(n12487), .ZN(n7886) );
  AOI21_X1 U7614 ( .B1(n12497), .B2(n11908), .A(n12039), .ZN(n12481) );
  NOR2_X1 U7615 ( .A1(n7884), .A2(n7860), .ZN(n7859) );
  INV_X1 U7616 ( .A(n7439), .ZN(n7438) );
  AOI21_X1 U7617 ( .B1(n7439), .B2(n7437), .A(n7436), .ZN(n7435) );
  INV_X1 U7618 ( .A(n7442), .ZN(n7437) );
  INV_X1 U7619 ( .A(n12001), .ZN(n7436) );
  AOI21_X1 U7620 ( .B1(n7070), .B2(n7072), .A(n6738), .ZN(n7068) );
  AOI21_X1 U7621 ( .B1(n6989), .B2(n11959), .A(n11912), .ZN(n6987) );
  INV_X1 U7622 ( .A(n11909), .ZN(n6989) );
  AND2_X1 U7623 ( .A1(n9420), .A2(n12772), .ZN(n10160) );
  INV_X1 U7624 ( .A(n11402), .ZN(n8724) );
  NAND2_X1 U7625 ( .A1(n7403), .A2(n7402), .ZN(n11725) );
  AND2_X1 U7626 ( .A1(n11722), .A2(n9289), .ZN(n7402) );
  INV_X1 U7627 ( .A(n9255), .ZN(n10182) );
  OAI21_X1 U7628 ( .B1(n9159), .B2(n7401), .A(n7398), .ZN(n9190) );
  NAND2_X1 U7629 ( .A1(n9175), .A2(n14572), .ZN(n7401) );
  NAND2_X1 U7630 ( .A1(n7873), .A2(n7098), .ZN(n8737) );
  INV_X1 U7631 ( .A(n9059), .ZN(n7115) );
  AND3_X1 U7632 ( .A1(n7683), .A2(n8919), .A3(n6662), .ZN(n8718) );
  NOR2_X1 U7633 ( .A1(n8750), .A2(n8703), .ZN(n8919) );
  NAND2_X1 U7634 ( .A1(n6926), .A2(n6927), .ZN(n12813) );
  INV_X1 U7635 ( .A(n6749), .ZN(n7302) );
  INV_X1 U7636 ( .A(n13087), .ZN(n13088) );
  OR2_X1 U7637 ( .A1(n10970), .A2(n10969), .ZN(n6932) );
  INV_X2 U7638 ( .A(n8160), .ZN(n8585) );
  NAND2_X1 U7639 ( .A1(n13126), .A2(n13292), .ZN(n13115) );
  NAND2_X1 U7640 ( .A1(n13299), .A2(n6660), .ZN(n13106) );
  INV_X1 U7641 ( .A(n8611), .ZN(n8532) );
  AOI21_X1 U7642 ( .B1(n7344), .B2(n7722), .A(n7343), .ZN(n7342) );
  INV_X1 U7643 ( .A(n13085), .ZN(n7343) );
  OR2_X1 U7644 ( .A1(n13325), .A2(n13051), .ZN(n7799) );
  NAND2_X1 U7645 ( .A1(n13197), .A2(n7721), .ZN(n7347) );
  NAND2_X1 U7646 ( .A1(n8316), .A2(n8315), .ZN(n13069) );
  NAND2_X1 U7647 ( .A1(n7807), .A2(n7231), .ZN(n7230) );
  AOI21_X1 U7648 ( .B1(n7808), .B2(n11575), .A(n7809), .ZN(n7807) );
  NAND2_X1 U7649 ( .A1(n11509), .A2(n7808), .ZN(n7231) );
  NAND2_X1 U7650 ( .A1(n7329), .A2(n6656), .ZN(n7325) );
  NAND2_X1 U7651 ( .A1(n10532), .A2(n10629), .ZN(n10751) );
  NOR2_X2 U7652 ( .A1(n10450), .A2(n10647), .ZN(n10532) );
  OAI211_X1 U7653 ( .C1(n8064), .C2(n12988), .A(n7769), .B(n7768), .ZN(n10344)
         );
  NAND2_X1 U7654 ( .A1(n10350), .A2(n7771), .ZN(n7768) );
  NAND2_X1 U7655 ( .A1(n7770), .A2(n8064), .ZN(n7769) );
  NOR2_X1 U7656 ( .A1(n10350), .A2(n7771), .ZN(n7770) );
  INV_X1 U7657 ( .A(n13063), .ZN(n13289) );
  NAND2_X1 U7658 ( .A1(n13100), .A2(n13099), .ZN(n13101) );
  INV_X1 U7659 ( .A(n15376), .ZN(n15366) );
  OR2_X1 U7660 ( .A1(n7929), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n7940) );
  NAND2_X1 U7661 ( .A1(n7017), .A2(n6611), .ZN(n10673) );
  INV_X2 U7662 ( .A(n10721), .ZN(n13680) );
  NAND2_X1 U7663 ( .A1(n7032), .A2(n6640), .ZN(n13703) );
  NAND2_X2 U7664 ( .A1(n9986), .A2(n10229), .ZN(n13681) );
  AND2_X1 U7665 ( .A1(n14179), .A2(n13805), .ZN(n14248) );
  NAND2_X1 U7666 ( .A1(n14258), .A2(n6891), .ZN(n6883) );
  OR2_X1 U7667 ( .A1(n14258), .A2(n14199), .ZN(n6887) );
  NAND2_X1 U7668 ( .A1(n7688), .A2(n6629), .ZN(n7015) );
  NAND2_X1 U7669 ( .A1(n14386), .A2(n7688), .ZN(n7016) );
  NAND2_X1 U7670 ( .A1(n13526), .A2(n13525), .ZN(n14375) );
  AOI22_X1 U7671 ( .A1(n14405), .A2(n14404), .B1(n14414), .B2(n14170), .ZN(
        n14388) );
  AOI21_X1 U7672 ( .B1(n6941), .B2(n6943), .A(n6736), .ZN(n6939) );
  NAND2_X1 U7673 ( .A1(n14797), .A2(n14058), .ZN(n7707) );
  NAND2_X1 U7674 ( .A1(n10893), .A2(n10892), .ZN(n11023) );
  OAI21_X1 U7675 ( .B1(n6869), .B2(n6866), .A(n6863), .ZN(n10893) );
  INV_X1 U7676 ( .A(n6872), .ZN(n6866) );
  AOI21_X1 U7677 ( .B1(n13885), .B2(n7818), .A(n7822), .ZN(n7817) );
  NOR2_X1 U7678 ( .A1(n13891), .A2(n13892), .ZN(n7822) );
  NAND2_X1 U7679 ( .A1(n10500), .A2(n10777), .ZN(n13888) );
  OR2_X1 U7680 ( .A1(n15147), .A2(n14265), .ZN(n10769) );
  INV_X1 U7681 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9987) );
  AND3_X1 U7682 ( .A1(n9406), .A2(n9405), .A3(n9404), .ZN(n9410) );
  AND4_X1 U7683 ( .A1(n9098), .A2(n9097), .A3(n9096), .A4(n9095), .ZN(n12509)
         );
  NAND2_X1 U7684 ( .A1(n14637), .A2(n6757), .ZN(n6812) );
  NAND2_X1 U7685 ( .A1(n9079), .A2(n9078), .ZN(n12755) );
  NOR2_X1 U7686 ( .A1(n12841), .A2(n7311), .ZN(n7310) );
  INV_X1 U7687 ( .A(n12834), .ZN(n7311) );
  OAI21_X1 U7688 ( .B1(n7581), .B2(n12968), .A(n12957), .ZN(n6915) );
  NAND2_X1 U7689 ( .A1(n12789), .A2(n12788), .ZN(n12893) );
  INV_X1 U7690 ( .A(n7574), .ZN(n7573) );
  OAI21_X1 U7691 ( .B1(n7577), .B2(n7575), .A(n12907), .ZN(n7574) );
  OAI21_X1 U7692 ( .B1(n13291), .B2(n15352), .A(n7787), .ZN(n7254) );
  NAND2_X1 U7693 ( .A1(n7503), .A2(n7504), .ZN(n13664) );
  NAND2_X1 U7694 ( .A1(n13733), .A2(n7507), .ZN(n7503) );
  XNOR2_X1 U7695 ( .A(n7012), .B(n6962), .ZN(n7595) );
  AOI21_X1 U7696 ( .B1(n7014), .B2(n6645), .A(n7013), .ZN(n7012) );
  NOR2_X1 U7697 ( .A1(n14182), .A2(n14233), .ZN(n7013) );
  AND2_X1 U7698 ( .A1(n6898), .A2(n6896), .ZN(n14462) );
  OR2_X1 U7699 ( .A1(n14235), .A2(n15178), .ZN(n6898) );
  AOI21_X1 U7700 ( .B1(n14458), .B2(n15074), .A(n6897), .ZN(n6896) );
  AND3_X1 U7701 ( .A1(n7943), .A2(n7942), .A3(n7941), .ZN(n7123) );
  AND2_X1 U7702 ( .A1(n13875), .A2(n13876), .ZN(n13879) );
  OR2_X1 U7703 ( .A1(n8074), .A2(n7127), .ZN(n7124) );
  NAND2_X1 U7704 ( .A1(n8074), .A2(n7127), .ZN(n7126) );
  NAND2_X1 U7705 ( .A1(n7560), .A2(n7559), .ZN(n7558) );
  NAND2_X1 U7706 ( .A1(n7561), .A2(n13903), .ZN(n7559) );
  NAND2_X1 U7707 ( .A1(n13916), .A2(n6772), .ZN(n6771) );
  NAND2_X1 U7708 ( .A1(n6774), .A2(n6773), .ZN(n6772) );
  INV_X1 U7709 ( .A(n6775), .ZN(n6773) );
  AND2_X1 U7710 ( .A1(n6770), .A2(n6769), .ZN(n6768) );
  NAND2_X1 U7711 ( .A1(n7564), .A2(n6775), .ZN(n6769) );
  NAND2_X1 U7712 ( .A1(n6780), .A2(n6777), .ZN(n6770) );
  AOI21_X1 U7713 ( .B1(n8169), .B2(n8168), .A(n8167), .ZN(n8171) );
  OAI22_X1 U7714 ( .A1(n13932), .A2(n13931), .B1(n13937), .B2(n13936), .ZN(
        n6782) );
  AOI21_X1 U7715 ( .B1(n7160), .B2(n7158), .A(n7157), .ZN(n7156) );
  INV_X1 U7716 ( .A(n6688), .ZN(n7160) );
  INV_X1 U7717 ( .A(n13965), .ZN(n6798) );
  INV_X1 U7718 ( .A(n13959), .ZN(n13962) );
  INV_X1 U7719 ( .A(n7752), .ZN(n7191) );
  NAND2_X1 U7720 ( .A1(n8350), .A2(n7751), .ZN(n7750) );
  NAND2_X1 U7721 ( .A1(n7755), .A2(n7752), .ZN(n7751) );
  AND2_X1 U7722 ( .A1(n8326), .A2(n8327), .ZN(n7755) );
  NOR2_X1 U7723 ( .A1(n6790), .A2(n13976), .ZN(n7567) );
  OR2_X1 U7724 ( .A1(n7567), .A2(n6788), .ZN(n6787) );
  INV_X1 U7725 ( .A(n6786), .ZN(n6785) );
  OAI21_X1 U7726 ( .B1(n6789), .B2(n6788), .A(n13978), .ZN(n6786) );
  NOR2_X1 U7727 ( .A1(n7224), .A2(n14192), .ZN(n7223) );
  OR2_X1 U7728 ( .A1(n7224), .A2(n7225), .ZN(n7222) );
  AOI21_X1 U7729 ( .B1(n13974), .B2(n13975), .A(n7226), .ZN(n7225) );
  INV_X1 U7730 ( .A(n13973), .ZN(n7226) );
  NAND2_X1 U7731 ( .A1(n7766), .A2(n7764), .ZN(n7763) );
  AOI21_X1 U7732 ( .B1(n8376), .B2(n8375), .A(n8374), .ZN(n7290) );
  NAND2_X1 U7733 ( .A1(n8437), .A2(n8438), .ZN(n7762) );
  NAND2_X1 U7734 ( .A1(n7280), .A2(n7279), .ZN(n7278) );
  NAND2_X1 U7735 ( .A1(n7154), .A2(n7153), .ZN(n7152) );
  INV_X1 U7736 ( .A(n8437), .ZN(n7153) );
  INV_X1 U7737 ( .A(n8438), .ZN(n7154) );
  NAND2_X1 U7738 ( .A1(n13991), .A2(n7215), .ZN(n7214) );
  NAND2_X1 U7739 ( .A1(n13993), .A2(n13995), .ZN(n7550) );
  NAND2_X1 U7740 ( .A1(n7285), .A2(n6605), .ZN(n7284) );
  INV_X1 U7741 ( .A(n12029), .ZN(n7449) );
  INV_X1 U7742 ( .A(n7285), .ZN(n6765) );
  NOR2_X1 U7743 ( .A1(n7184), .A2(n8527), .ZN(n7183) );
  INV_X1 U7744 ( .A(n6605), .ZN(n7184) );
  NAND2_X1 U7745 ( .A1(n8485), .A2(n7138), .ZN(n7137) );
  INV_X1 U7746 ( .A(n7283), .ZN(n7138) );
  INV_X1 U7747 ( .A(n12990), .ZN(n8021) );
  XNOR2_X1 U7748 ( .A(n13861), .B(n14265), .ZN(n13865) );
  INV_X1 U7749 ( .A(n13998), .ZN(n14001) );
  OR2_X1 U7750 ( .A1(n7636), .A2(n7634), .ZN(n7633) );
  INV_X1 U7751 ( .A(n8377), .ZN(n7634) );
  NAND2_X1 U7752 ( .A1(n6741), .A2(n6598), .ZN(n7636) );
  INV_X1 U7753 ( .A(n8378), .ZN(n7635) );
  NOR2_X1 U7754 ( .A1(n8199), .A2(n7617), .ZN(n7616) );
  INV_X1 U7755 ( .A(n8175), .ZN(n7617) );
  NAND4_X1 U7756 ( .A1(n7910), .A2(n7911), .A3(n7909), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7604) );
  NAND2_X1 U7757 ( .A1(n10191), .A2(n10357), .ZN(n6808) );
  NAND2_X1 U7758 ( .A1(n10554), .A2(n6971), .ZN(n12392) );
  NAND2_X1 U7759 ( .A1(n10547), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n6971) );
  NAND2_X1 U7760 ( .A1(n15551), .A2(n14652), .ZN(n14653) );
  INV_X1 U7761 ( .A(n14839), .ZN(n7060) );
  INV_X1 U7762 ( .A(n14592), .ZN(n7059) );
  OR2_X1 U7763 ( .A1(n12652), .A2(n6575), .ZN(n12063) );
  INV_X1 U7764 ( .A(n12025), .ZN(n7001) );
  AOI21_X1 U7765 ( .B1(n7447), .B2(n7449), .A(n7445), .ZN(n7444) );
  INV_X1 U7766 ( .A(n12033), .ZN(n7445) );
  OR2_X1 U7767 ( .A1(n12550), .A2(n9274), .ZN(n12018) );
  INV_X1 U7768 ( .A(n9314), .ZN(n7066) );
  NAND3_X1 U7769 ( .A1(n7683), .A2(n7007), .A3(n7006), .ZN(n7453) );
  INV_X1 U7770 ( .A(n8703), .ZN(n7007) );
  NOR2_X1 U7771 ( .A1(n8750), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n7006) );
  AND2_X1 U7772 ( .A1(n7686), .A2(n9223), .ZN(n7685) );
  AND2_X1 U7773 ( .A1(n8714), .A2(n8715), .ZN(n7686) );
  NOR2_X1 U7774 ( .A1(n8871), .A2(n7388), .ZN(n7387) );
  INV_X1 U7775 ( .A(n8850), .ZN(n7388) );
  INV_X1 U7776 ( .A(n8847), .ZN(n7385) );
  INV_X1 U7777 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8844) );
  INV_X1 U7778 ( .A(n9919), .ZN(n9899) );
  NAND2_X1 U7779 ( .A1(n7306), .A2(n10615), .ZN(n7304) );
  INV_X1 U7780 ( .A(n12876), .ZN(n6929) );
  INV_X1 U7781 ( .A(n7737), .ZN(n7735) );
  OR3_X1 U7782 ( .A1(n8248), .A2(n11225), .A3(n11321), .ZN(n8271) );
  OR2_X1 U7783 ( .A1(n8185), .A2(n8184), .ZN(n8209) );
  NOR2_X1 U7784 ( .A1(n10742), .A2(n7323), .ZN(n7322) );
  INV_X1 U7785 ( .A(n10528), .ZN(n7323) );
  AND2_X1 U7786 ( .A1(n10988), .A2(n8640), .ZN(n10746) );
  NAND2_X1 U7787 ( .A1(n8642), .A2(n10121), .ZN(n10112) );
  OR2_X1 U7788 ( .A1(n9939), .A2(n11403), .ZN(n9711) );
  NOR2_X1 U7789 ( .A1(n7940), .A2(n7939), .ZN(n7588) );
  AND3_X2 U7790 ( .A1(n7228), .A2(n8179), .A3(n8178), .ZN(n7122) );
  NOR2_X1 U7791 ( .A1(n8176), .A2(n7892), .ZN(n7228) );
  INV_X1 U7792 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7891) );
  INV_X1 U7793 ( .A(n11645), .ZN(n7029) );
  AND2_X1 U7794 ( .A1(n7518), .A2(n7516), .ZN(n7515) );
  NAND2_X1 U7795 ( .A1(n7519), .A2(n6626), .ZN(n7518) );
  NAND2_X1 U7796 ( .A1(n13647), .A2(n7520), .ZN(n7519) );
  INV_X1 U7797 ( .A(n13479), .ZN(n7520) );
  AND2_X1 U7798 ( .A1(n6626), .A2(n13480), .ZN(n7521) );
  NAND2_X1 U7799 ( .A1(n14158), .A2(n14021), .ZN(n14030) );
  NAND2_X1 U7800 ( .A1(n6891), .A2(n14199), .ZN(n6890) );
  NOR2_X1 U7801 ( .A1(n7702), .A2(n7706), .ZN(n7701) );
  AND2_X1 U7802 ( .A1(n14304), .A2(n14176), .ZN(n7706) );
  INV_X1 U7803 ( .A(n7704), .ZN(n7702) );
  AND2_X1 U7804 ( .A1(n6977), .A2(n6851), .ZN(n6850) );
  NAND2_X1 U7805 ( .A1(n14334), .A2(n6852), .ZN(n6851) );
  AND2_X1 U7806 ( .A1(n6711), .A2(n6586), .ZN(n6977) );
  INV_X1 U7807 ( .A(n14174), .ZN(n6852) );
  NOR2_X1 U7808 ( .A1(n6876), .A2(n11623), .ZN(n6875) );
  INV_X1 U7809 ( .A(n6610), .ZN(n6876) );
  INV_X1 U7810 ( .A(n11238), .ZN(n6878) );
  AND2_X1 U7811 ( .A1(n6607), .A2(n10894), .ZN(n6860) );
  NAND2_X1 U7812 ( .A1(n6861), .A2(n13815), .ZN(n6856) );
  NAND2_X1 U7813 ( .A1(n6619), .A2(n10894), .ZN(n6861) );
  NAND2_X1 U7814 ( .A1(n7817), .A2(n7821), .ZN(n6936) );
  XNOR2_X1 U7815 ( .A(n14434), .B(n13880), .ZN(n13809) );
  OR2_X1 U7816 ( .A1(n14460), .A2(n14246), .ZN(n7828) );
  NAND2_X1 U7817 ( .A1(n6944), .A2(n6945), .ZN(n14300) );
  AOI21_X1 U7818 ( .B1(n14309), .B2(n6946), .A(n6671), .ZN(n6945) );
  NAND2_X1 U7819 ( .A1(n8465), .A2(n8464), .ZN(n8487) );
  INV_X1 U7820 ( .A(n8354), .ZN(n6997) );
  NAND2_X1 U7821 ( .A1(n6981), .A2(n6979), .ZN(n8244) );
  AOI21_X1 U7822 ( .B1(n6982), .B2(n6984), .A(n6980), .ZN(n6979) );
  INV_X1 U7823 ( .A(n8239), .ZN(n6980) );
  NAND2_X1 U7824 ( .A1(n7609), .A2(n7360), .ZN(n7359) );
  AOI21_X1 U7825 ( .B1(n7609), .B2(n7611), .A(n6684), .ZN(n7607) );
  INV_X1 U7826 ( .A(n8243), .ZN(n7360) );
  NAND2_X1 U7827 ( .A1(n8244), .A2(n8243), .ZN(n8283) );
  XNOR2_X1 U7828 ( .A(n8283), .B(n9676), .ZN(n8262) );
  NAND2_X1 U7829 ( .A1(n8154), .A2(n8153), .ZN(n8174) );
  NAND2_X1 U7830 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7189), .ZN(n7188) );
  INV_X1 U7831 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7189) );
  INV_X1 U7832 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14691) );
  AOI21_X1 U7833 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n15017), .A(n14692), .ZN(
        n14749) );
  AND2_X1 U7834 ( .A1(n11204), .A2(n6828), .ZN(n6821) );
  NAND2_X1 U7835 ( .A1(n6839), .A2(n6843), .ZN(n9135) );
  NAND2_X1 U7836 ( .A1(n10594), .A2(n10595), .ZN(n7674) );
  NOR2_X1 U7837 ( .A1(n8810), .A2(n8808), .ZN(n10476) );
  AND2_X1 U7838 ( .A1(n8806), .A2(n8807), .ZN(n8808) );
  OR2_X1 U7839 ( .A1(n11561), .A2(n11562), .ZN(n11559) );
  NAND2_X1 U7840 ( .A1(n6842), .A2(n6841), .ZN(n6840) );
  NAND2_X1 U7841 ( .A1(n9120), .A2(n9121), .ZN(n6843) );
  AND3_X1 U7842 ( .A1(n8777), .A2(n8776), .A3(n8775), .ZN(n10704) );
  NAND2_X1 U7843 ( .A1(n10958), .A2(n6665), .ZN(n6827) );
  INV_X1 U7844 ( .A(n7661), .ZN(n7659) );
  NOR2_X1 U7845 ( .A1(n7880), .A2(n8991), .ZN(n7661) );
  AND2_X1 U7846 ( .A1(n11901), .A2(n11900), .ZN(n11906) );
  NAND2_X1 U7847 ( .A1(n12072), .A2(n7407), .ZN(n7406) );
  NOR2_X1 U7848 ( .A1(n11926), .A2(n12066), .ZN(n7407) );
  AND4_X1 U7849 ( .A1(n8989), .A2(n8988), .A3(n8987), .A4(n8986), .ZN(n9329)
         );
  OAI21_X1 U7850 ( .B1(n10279), .B2(n15396), .A(n6606), .ZN(n10266) );
  OAI21_X1 U7851 ( .B1(n10182), .B2(n10605), .A(n6811), .ZN(n6810) );
  NAND2_X1 U7852 ( .A1(n10182), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n6811) );
  AND3_X1 U7853 ( .A1(n6583), .A2(n6726), .A3(n7365), .ZN(n10379) );
  OAI21_X1 U7854 ( .B1(n7049), .B2(n7047), .A(n7048), .ZN(n7045) );
  OR2_X1 U7855 ( .A1(n7367), .A2(n14642), .ZN(n7048) );
  NOR2_X1 U7856 ( .A1(n12382), .A2(n12383), .ZN(n12385) );
  OR2_X1 U7857 ( .A1(n15477), .A2(n7364), .ZN(n7363) );
  AND2_X1 U7858 ( .A1(n15485), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7364) );
  OR2_X1 U7859 ( .A1(n15511), .A2(n7042), .ZN(n7041) );
  NOR2_X1 U7860 ( .A1(n14648), .A2(n14583), .ZN(n7042) );
  XNOR2_X1 U7861 ( .A(n14622), .B(n14827), .ZN(n14831) );
  OR2_X1 U7862 ( .A1(n14831), .A2(n14832), .ZN(n6815) );
  NAND2_X1 U7863 ( .A1(n7375), .A2(n7374), .ZN(n14587) );
  AOI21_X1 U7864 ( .B1(n14585), .B2(n7376), .A(n7377), .ZN(n7374) );
  XNOR2_X1 U7865 ( .A(n14653), .B(n14623), .ZN(n14824) );
  NAND2_X1 U7866 ( .A1(n14824), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n14823) );
  AND2_X1 U7867 ( .A1(n9247), .A2(n9246), .ZN(n12408) );
  OAI21_X1 U7868 ( .B1(n12452), .B2(n7083), .A(n7078), .ZN(n12427) );
  AND2_X1 U7869 ( .A1(n7079), .A2(n7081), .ZN(n7078) );
  NAND2_X1 U7870 ( .A1(n6680), .A2(n7084), .ZN(n7081) );
  NAND2_X1 U7871 ( .A1(n7082), .A2(n7080), .ZN(n7079) );
  NAND2_X1 U7872 ( .A1(n12426), .A2(n9350), .ZN(n12412) );
  NAND2_X1 U7873 ( .A1(n12427), .A2(n12428), .ZN(n12426) );
  AND2_X1 U7874 ( .A1(n9203), .A2(n9202), .ZN(n12443) );
  AND2_X1 U7875 ( .A1(n9186), .A2(n9185), .ZN(n12456) );
  AOI21_X1 U7876 ( .B1(n12461), .B2(n8789), .A(n9169), .ZN(n12473) );
  NAND2_X1 U7877 ( .A1(n7075), .A2(n7073), .ZN(n12482) );
  NOR2_X1 U7878 ( .A1(n7879), .A2(n7074), .ZN(n7073) );
  INV_X1 U7879 ( .A(n12483), .ZN(n7074) );
  NAND2_X1 U7880 ( .A1(n7857), .A2(n7856), .ZN(n7855) );
  INV_X1 U7881 ( .A(n7884), .ZN(n7856) );
  INV_X1 U7882 ( .A(n7862), .ZN(n7857) );
  OR2_X1 U7883 ( .A1(n12039), .A2(n12038), .ZN(n12496) );
  NOR2_X1 U7884 ( .A1(n12519), .A2(n7451), .ZN(n7450) );
  INV_X1 U7885 ( .A(n12024), .ZN(n7451) );
  AND2_X1 U7886 ( .A1(n9105), .A2(n9104), .ZN(n12522) );
  INV_X1 U7887 ( .A(n7086), .ZN(n7085) );
  OAI21_X1 U7888 ( .B1(n6613), .B2(n7087), .A(n9343), .ZN(n7086) );
  NAND2_X1 U7889 ( .A1(n7002), .A2(n12025), .ZN(n9275) );
  INV_X1 U7890 ( .A(n12530), .ZN(n7002) );
  NAND2_X1 U7891 ( .A1(n9339), .A2(n6613), .ZN(n12543) );
  AND2_X1 U7892 ( .A1(n12018), .A2(n12019), .ZN(n12546) );
  INV_X1 U7893 ( .A(n7435), .ZN(n7005) );
  AND2_X1 U7894 ( .A1(n7433), .A2(n7004), .ZN(n7003) );
  NAND2_X1 U7895 ( .A1(n7435), .A2(n12642), .ZN(n7004) );
  NOR2_X1 U7896 ( .A1(n11998), .A2(n7443), .ZN(n7442) );
  INV_X1 U7897 ( .A(n11993), .ZN(n7443) );
  NAND2_X1 U7898 ( .A1(n12643), .A2(n12630), .ZN(n9273) );
  AOI21_X1 U7899 ( .B1(n7852), .B2(n7854), .A(n6732), .ZN(n7850) );
  NAND2_X1 U7900 ( .A1(n11275), .A2(n7852), .ZN(n7849) );
  NAND2_X1 U7901 ( .A1(n11275), .A2(n9317), .ZN(n7851) );
  AND4_X1 U7902 ( .A1(n8930), .A2(n8929), .A3(n8928), .A4(n8927), .ZN(n11836)
         );
  NAND2_X1 U7903 ( .A1(n11117), .A2(n11909), .ZN(n11119) );
  AND4_X1 U7904 ( .A1(n8859), .A2(n8858), .A3(n8857), .A4(n8856), .ZN(n11288)
         );
  NAND2_X1 U7905 ( .A1(n10824), .A2(n11948), .ZN(n10823) );
  OR2_X1 U7906 ( .A1(n9258), .A2(n12044), .ZN(n12587) );
  OR2_X1 U7907 ( .A1(n11932), .A2(n14790), .ZN(n12044) );
  NAND2_X1 U7908 ( .A1(n9195), .A2(n9194), .ZN(n9349) );
  NAND2_X1 U7909 ( .A1(n7120), .A2(n9179), .ZN(n9348) );
  NAND2_X1 U7910 ( .A1(n11399), .A2(n11887), .ZN(n7120) );
  NAND2_X1 U7911 ( .A1(n9164), .A2(n9163), .ZN(n9301) );
  INV_X1 U7912 ( .A(n6570), .ZN(n9063) );
  NAND2_X1 U7913 ( .A1(n9258), .A2(n12070), .ZN(n12589) );
  OAI21_X1 U7914 ( .B1(n9209), .B2(P3_D_REG_0__SCAN_IN), .A(n8727), .ZN(n9376)
         );
  NOR2_X1 U7915 ( .A1(n9287), .A2(n7405), .ZN(n7404) );
  INV_X1 U7916 ( .A(n9282), .ZN(n7405) );
  NAND2_X1 U7917 ( .A1(n8717), .A2(n6662), .ZN(n7874) );
  NAND2_X1 U7918 ( .A1(n9160), .A2(n9148), .ZN(n9159) );
  AOI21_X1 U7919 ( .B1(n7104), .B2(n7106), .A(n6753), .ZN(n7102) );
  NAND2_X1 U7920 ( .A1(n8718), .A2(n7686), .ZN(n9222) );
  AND2_X1 U7921 ( .A1(n9089), .A2(n9076), .ZN(n9087) );
  AOI21_X1 U7922 ( .B1(n7114), .B2(n9057), .A(n7112), .ZN(n7111) );
  INV_X1 U7923 ( .A(n9075), .ZN(n7112) );
  AND2_X1 U7924 ( .A1(n9075), .A2(n9060), .ZN(n9072) );
  INV_X1 U7925 ( .A(n9058), .ZN(n7118) );
  NAND2_X1 U7926 ( .A1(n7100), .A2(n9029), .ZN(n9042) );
  INV_X1 U7927 ( .A(n8955), .ZN(n7394) );
  NAND2_X1 U7928 ( .A1(n7397), .A2(n7396), .ZN(n7395) );
  INV_X1 U7929 ( .A(n8954), .ZN(n7397) );
  NAND2_X1 U7930 ( .A1(n7099), .A2(n8918), .ZN(n8936) );
  NAND2_X1 U7931 ( .A1(n8879), .A2(n8878), .ZN(n8881) );
  NAND2_X1 U7932 ( .A1(n8831), .A2(n8830), .ZN(n8848) );
  XNOR2_X1 U7933 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8847) );
  NOR2_X1 U7934 ( .A1(n13411), .A2(n13412), .ZN(n9419) );
  OAI21_X1 U7935 ( .B1(n10094), .B2(n7583), .A(n6590), .ZN(n10293) );
  OR2_X1 U7936 ( .A1(n11011), .A2(n11012), .ZN(n7301) );
  OR2_X1 U7937 ( .A1(n9704), .A2(n9708), .ZN(n13031) );
  INV_X1 U7938 ( .A(n12894), .ZN(n7577) );
  OR2_X1 U7939 ( .A1(n8317), .A2(n12902), .ZN(n8338) );
  INV_X1 U7940 ( .A(n12991), .ZN(n9920) );
  AND3_X1 U7941 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_27__SCAN_IN), .ZN(n7922) );
  NAND2_X1 U7942 ( .A1(n7300), .A2(n7299), .ZN(n7295) );
  INV_X1 U7943 ( .A(n7301), .ZN(n7299) );
  NAND2_X1 U7944 ( .A1(n6932), .A2(n6642), .ZN(n7296) );
  NAND2_X1 U7945 ( .A1(n8160), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7134) );
  NAND2_X1 U7946 ( .A1(n13313), .A2(n13086), .ZN(n7729) );
  INV_X1 U7947 ( .A(n7730), .ZN(n13153) );
  INV_X1 U7948 ( .A(n7797), .ZN(n7793) );
  AND2_X1 U7949 ( .A1(n7789), .A2(n7239), .ZN(n7238) );
  NAND2_X1 U7950 ( .A1(n7790), .A2(n7791), .ZN(n7789) );
  NAND2_X1 U7951 ( .A1(n7792), .A2(n13196), .ZN(n7239) );
  INV_X1 U7952 ( .A(n7798), .ZN(n7791) );
  NOR2_X1 U7953 ( .A1(n13184), .A2(n7801), .ZN(n7797) );
  NOR2_X1 U7954 ( .A1(n7346), .A2(n7795), .ZN(n7794) );
  INV_X1 U7955 ( .A(n7799), .ZN(n7795) );
  AND2_X1 U7956 ( .A1(n7720), .A2(n6722), .ZN(n7719) );
  INV_X1 U7957 ( .A(n13084), .ZN(n7346) );
  NAND2_X1 U7958 ( .A1(n13209), .A2(n13208), .ZN(n13207) );
  NAND2_X1 U7959 ( .A1(n7334), .A2(n7333), .ZN(n13080) );
  AOI21_X1 U7960 ( .B1(n7335), .B2(n7338), .A(n6653), .ZN(n7333) );
  NOR2_X1 U7961 ( .A1(n7804), .A2(n7251), .ZN(n7250) );
  INV_X1 U7962 ( .A(n7805), .ZN(n7251) );
  NOR2_X1 U7963 ( .A1(n13348), .A2(n13043), .ZN(n7804) );
  NAND2_X1 U7964 ( .A1(n7534), .A2(n7533), .ZN(n13250) );
  NOR2_X1 U7965 ( .A1(n7740), .A2(n11590), .ZN(n7739) );
  INV_X1 U7966 ( .A(n11578), .ZN(n7740) );
  NAND2_X1 U7967 ( .A1(n7738), .A2(n12978), .ZN(n7737) );
  INV_X1 U7968 ( .A(n11595), .ZN(n7229) );
  AND2_X1 U7969 ( .A1(n11570), .A2(n11572), .ZN(n7808) );
  OR2_X1 U7970 ( .A1(n11509), .A2(n11575), .ZN(n11571) );
  AOI21_X1 U7971 ( .B1(n7245), .B2(n11064), .A(n6689), .ZN(n7244) );
  NAND2_X1 U7972 ( .A1(n11065), .A2(n7245), .ZN(n7242) );
  INV_X1 U7973 ( .A(n13264), .ZN(n13247) );
  OAI21_X2 U7974 ( .B1(n10857), .B2(n8611), .A(n8087), .ZN(n10564) );
  NOR2_X1 U7975 ( .A1(n10302), .A2(n7777), .ZN(n7776) );
  INV_X1 U7976 ( .A(n10116), .ZN(n7777) );
  AND2_X1 U7977 ( .A1(n8641), .A2(n10304), .ZN(n10124) );
  NOR2_X2 U7978 ( .A1(n10397), .A2(n15348), .ZN(n10440) );
  INV_X1 U7979 ( .A(n10112), .ZN(n10204) );
  NAND2_X1 U7980 ( .A1(n8647), .A2(n10118), .ZN(n10252) );
  INV_X1 U7981 ( .A(n13294), .ZN(n13270) );
  NAND2_X1 U7982 ( .A1(n7288), .A2(n8618), .ZN(n7287) );
  XNOR2_X1 U7983 ( .A(n9712), .B(n11403), .ZN(n7585) );
  NAND2_X1 U7984 ( .A1(n8648), .A2(n10129), .ZN(n8649) );
  INV_X1 U7985 ( .A(n13040), .ZN(n13287) );
  NAND2_X1 U7986 ( .A1(n13092), .A2(n7784), .ZN(n7783) );
  INV_X1 U7987 ( .A(n7788), .ZN(n7784) );
  NAND2_X1 U7988 ( .A1(n13107), .A2(n13096), .ZN(n7788) );
  AND2_X1 U7989 ( .A1(n9679), .A2(n9693), .ZN(n15314) );
  INV_X1 U7990 ( .A(n7929), .ZN(n7169) );
  AND2_X1 U7991 ( .A1(n7915), .A2(n7916), .ZN(n7526) );
  INV_X1 U7992 ( .A(n7929), .ZN(n7925) );
  OR2_X1 U7993 ( .A1(n8085), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8116) );
  INV_X1 U7994 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8742) );
  OR2_X1 U7995 ( .A1(n7484), .A2(n13775), .ZN(n7483) );
  INV_X1 U7996 ( .A(n13658), .ZN(n7479) );
  OAI21_X1 U7997 ( .B1(n7483), .B2(n7037), .A(n7480), .ZN(n7476) );
  INV_X1 U7998 ( .A(n7481), .ZN(n7480) );
  OAI21_X1 U7999 ( .B1(n7484), .B2(n7482), .A(n7489), .ZN(n7481) );
  OR2_X1 U8000 ( .A1(n13633), .A2(n13632), .ZN(n7489) );
  AND2_X1 U8001 ( .A1(n7502), .A2(n7504), .ZN(n7501) );
  INV_X1 U8002 ( .A(n13665), .ZN(n7502) );
  NAND2_X1 U8003 ( .A1(n11266), .A2(n7522), .ZN(n11451) );
  NOR2_X1 U8004 ( .A1(n11269), .A2(n7523), .ZN(n7522) );
  INV_X1 U8005 ( .A(n11265), .ZN(n7523) );
  XNOR2_X1 U8006 ( .A(n7021), .B(n13517), .ZN(n10027) );
  OAI22_X1 U8007 ( .A1(n14428), .A2(n13681), .B1(n10072), .B2(n14423), .ZN(
        n7021) );
  NAND2_X1 U8008 ( .A1(n10673), .A2(n10672), .ZN(n10729) );
  AND3_X1 U8009 ( .A1(n10002), .A2(n10001), .A3(n10000), .ZN(n10030) );
  OR2_X1 U8010 ( .A1(n10006), .A2(n10030), .ZN(n10032) );
  INV_X1 U8011 ( .A(n13752), .ZN(n7031) );
  NAND2_X1 U8012 ( .A1(n13733), .A2(n7498), .ZN(n7497) );
  NOR2_X1 U8013 ( .A1(n7500), .A2(n7499), .ZN(n7498) );
  INV_X1 U8014 ( .A(n7509), .ZN(n7499) );
  INV_X1 U8015 ( .A(n7507), .ZN(n7500) );
  NAND2_X1 U8016 ( .A1(n7025), .A2(n7023), .ZN(n11669) );
  NAND2_X1 U8017 ( .A1(n11483), .A2(n7026), .ZN(n7025) );
  INV_X1 U8018 ( .A(n7024), .ZN(n7023) );
  NOR2_X1 U8019 ( .A1(n7029), .A2(n7027), .ZN(n7026) );
  OAI21_X1 U8020 ( .B1(n13876), .B2(n13681), .A(n7524), .ZN(n10073) );
  NAND2_X1 U8021 ( .A1(n13880), .A2(n13627), .ZN(n7524) );
  NAND2_X1 U8022 ( .A1(n7033), .A2(n13494), .ZN(n13786) );
  NAND2_X1 U8023 ( .A1(n7517), .A2(n7518), .ZN(n7033) );
  NAND2_X1 U8024 ( .A1(n13481), .A2(n7521), .ZN(n7517) );
  AND4_X1 U8025 ( .A1(n11430), .A2(n11429), .A3(n11428), .A4(n11427), .ZN(
        n13485) );
  AND4_X1 U8026 ( .A1(n11138), .A2(n11137), .A3(n11136), .A4(n11135), .ZN(
        n13929) );
  INV_X1 U8027 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14668) );
  NAND2_X1 U8028 ( .A1(n7351), .A2(n7350), .ZN(n7014) );
  NAND2_X1 U8029 ( .A1(n14460), .A2(n14180), .ZN(n7350) );
  INV_X1 U8030 ( .A(n14452), .ZN(n14182) );
  INV_X1 U8031 ( .A(n14233), .ZN(n14181) );
  INV_X1 U8032 ( .A(n7014), .ZN(n14214) );
  NAND2_X1 U8033 ( .A1(n14246), .A2(n15049), .ZN(n7196) );
  NAND2_X1 U8034 ( .A1(n14229), .A2(n14231), .ZN(n14228) );
  NOR2_X1 U8035 ( .A1(n7832), .A2(n6625), .ZN(n7831) );
  INV_X1 U8036 ( .A(n7837), .ZN(n7832) );
  INV_X1 U8037 ( .A(n14248), .ZN(n6952) );
  OR2_X1 U8038 ( .A1(n7833), .A2(n6625), .ZN(n7830) );
  NOR2_X1 U8039 ( .A1(n14276), .A2(n7838), .ZN(n7837) );
  INV_X1 U8040 ( .A(n14198), .ZN(n7838) );
  NOR2_X1 U8041 ( .A1(n14260), .A2(n7834), .ZN(n7833) );
  INV_X1 U8042 ( .A(n7836), .ZN(n7834) );
  OR2_X1 U8043 ( .A1(n14284), .A2(n14295), .ZN(n7836) );
  NAND2_X1 U8044 ( .A1(n14275), .A2(n7352), .ZN(n14258) );
  OR2_X1 U8045 ( .A1(n13806), .A2(n14326), .ZN(n14292) );
  NAND2_X1 U8046 ( .A1(n14338), .A2(n7829), .ZN(n14331) );
  INV_X1 U8047 ( .A(n7698), .ZN(n7690) );
  INV_X1 U8048 ( .A(n7695), .ZN(n7694) );
  NAND2_X1 U8049 ( .A1(n7689), .A2(n7698), .ZN(n7688) );
  NAND2_X1 U8050 ( .A1(n7692), .A2(n14356), .ZN(n7689) );
  NAND2_X1 U8051 ( .A1(n7695), .A2(n7693), .ZN(n7692) );
  INV_X1 U8052 ( .A(n7697), .ZN(n7693) );
  NAND2_X1 U8053 ( .A1(n13464), .A2(n13463), .ZN(n14358) );
  AND2_X1 U8054 ( .A1(n7699), .A2(n7700), .ZN(n7697) );
  NAND2_X1 U8055 ( .A1(n7696), .A2(n7699), .ZN(n7695) );
  INV_X1 U8056 ( .A(n14368), .ZN(n7696) );
  NAND2_X1 U8057 ( .A1(n6963), .A2(n6964), .ZN(n14355) );
  AOI21_X1 U8058 ( .B1(n6577), .B2(n6969), .A(n7839), .ZN(n6964) );
  NAND2_X1 U8059 ( .A1(n7843), .A2(n14189), .ZN(n14366) );
  NAND2_X1 U8060 ( .A1(n14187), .A2(n7844), .ZN(n7843) );
  NAND2_X1 U8061 ( .A1(n14388), .A2(n14387), .ZN(n14386) );
  NAND2_X1 U8062 ( .A1(n6965), .A2(n6967), .ZN(n14187) );
  NAND2_X1 U8063 ( .A1(n6966), .A2(n14183), .ZN(n6965) );
  INV_X1 U8064 ( .A(n14934), .ZN(n6966) );
  AOI21_X1 U8065 ( .B1(n14169), .B2(n14168), .A(n14167), .ZN(n14405) );
  NAND2_X1 U8066 ( .A1(n13821), .A2(n6880), .ZN(n6879) );
  INV_X1 U8067 ( .A(n7707), .ZN(n6880) );
  NAND2_X1 U8068 ( .A1(n6878), .A2(n6610), .ZN(n6877) );
  NAND2_X1 U8069 ( .A1(n7824), .A2(n7823), .ZN(n11420) );
  OR2_X1 U8070 ( .A1(n7825), .A2(n7826), .ZN(n7823) );
  AOI21_X1 U8071 ( .B1(n14952), .B2(n13925), .A(n7827), .ZN(n7826) );
  OR2_X1 U8072 ( .A1(n11238), .A2(n13820), .ZN(n7708) );
  NAND2_X1 U8073 ( .A1(n11146), .A2(n11145), .ZN(n15057) );
  NAND2_X1 U8074 ( .A1(n15053), .A2(n15054), .ZN(n15052) );
  NAND2_X1 U8075 ( .A1(n11023), .A2(n6860), .ZN(n6859) );
  NAND2_X1 U8076 ( .A1(n6856), .A2(n6607), .ZN(n6858) );
  NOR2_X1 U8077 ( .A1(n6868), .A2(n10890), .ZN(n6867) );
  INV_X1 U8078 ( .A(n10413), .ZN(n6868) );
  OR2_X1 U8079 ( .A1(n15095), .A2(n14063), .ZN(n6872) );
  NAND2_X1 U8080 ( .A1(n7816), .A2(n7818), .ZN(n7815) );
  NOR2_X1 U8081 ( .A1(n10411), .A2(n6871), .ZN(n6870) );
  INV_X1 U8082 ( .A(n13888), .ZN(n6871) );
  AOI22_X1 U8083 ( .A1(n13524), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n13523), 
        .B2(n14102), .ZN(n6933) );
  NAND2_X1 U8084 ( .A1(n11615), .A2(n10215), .ZN(n6800) );
  OR2_X1 U8085 ( .A1(n13517), .A2(n10231), .ZN(n10844) );
  OR2_X1 U8086 ( .A1(n14300), .A2(n14299), .ZN(n14485) );
  NAND2_X1 U8087 ( .A1(n11619), .A2(n11618), .ZN(n14534) );
  OR2_X1 U8088 ( .A1(n10012), .A2(n10011), .ZN(n10248) );
  NAND2_X1 U8089 ( .A1(n7625), .A2(n6752), .ZN(n8609) );
  NAND2_X1 U8090 ( .A1(n7626), .A2(n8553), .ZN(n8582) );
  XNOR2_X1 U8091 ( .A(n9417), .B(n9416), .ZN(n9663) );
  NOR2_X1 U8092 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n9397) );
  NOR2_X1 U8093 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9396) );
  INV_X1 U8094 ( .A(n7209), .ZN(n7208) );
  OAI21_X1 U8095 ( .B1(n8081), .B2(n7210), .A(n8112), .ZN(n7209) );
  OAI211_X1 U8096 ( .C1(n8024), .C2(n6919), .A(n8029), .B(n6917), .ZN(n8053)
         );
  AND2_X1 U8097 ( .A1(n8026), .A2(n8011), .ZN(n6918) );
  INV_X1 U8098 ( .A(n7961), .ZN(n7963) );
  XNOR2_X1 U8099 ( .A(n14716), .B(n6909), .ZN(n14720) );
  INV_X1 U8100 ( .A(n14717), .ZN(n6909) );
  INV_X1 U8101 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14712) );
  AND2_X1 U8102 ( .A1(n6905), .A2(n6904), .ZN(n14728) );
  OAI21_X1 U8103 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14685), .A(n14684), .ZN(
        n14708) );
  AOI21_X1 U8104 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n14689), .A(n14688), .ZN(
        n14746) );
  AOI21_X1 U8105 ( .B1(n14966), .B2(n14967), .A(n7455), .ZN(n6911) );
  OR2_X1 U8106 ( .A1(n8799), .A2(n9428), .ZN(n8800) );
  OAI21_X1 U8107 ( .B1(n11808), .B2(n11807), .A(n9101), .ZN(n11753) );
  AOI21_X1 U8108 ( .B1(n12474), .B2(n8789), .A(n9155), .ZN(n12487) );
  NAND2_X1 U8109 ( .A1(n11864), .A2(n9025), .ZN(n11784) );
  NAND2_X1 U8110 ( .A1(n9092), .A2(n9091), .ZN(n12524) );
  OAI21_X1 U8111 ( .B1(n11760), .B2(n8975), .A(n8974), .ZN(n11817) );
  NAND2_X1 U8112 ( .A1(n9119), .A2(n9118), .ZN(n11829) );
  AND4_X1 U8113 ( .A1(n9056), .A2(n9055), .A3(n9054), .A4(n9053), .ZN(n12548)
         );
  NAND2_X1 U8114 ( .A1(n6834), .A2(n7676), .ZN(n11844) );
  NAND2_X1 U8115 ( .A1(n11864), .A2(n6835), .ZN(n6834) );
  AND2_X1 U8116 ( .A1(n9237), .A2(n12639), .ZN(n11875) );
  AND2_X1 U8117 ( .A1(n9233), .A2(n10160), .ZN(n11863) );
  INV_X1 U8118 ( .A(n12587), .ZN(n12631) );
  INV_X1 U8119 ( .A(n12456), .ZN(n12095) );
  INV_X1 U8120 ( .A(n12548), .ZN(n12570) );
  INV_X1 U8121 ( .A(n9329), .ZN(n12634) );
  NOR2_X1 U8122 ( .A1(n10185), .A2(n6809), .ZN(n10264) );
  AND2_X1 U8123 ( .A1(n6810), .A2(n10279), .ZN(n6809) );
  XNOR2_X1 U8124 ( .A(n7363), .B(n15501), .ZN(n15496) );
  NOR2_X1 U8125 ( .A1(n15496), .A2(n11417), .ZN(n15495) );
  OAI21_X1 U8126 ( .B1(n14858), .B2(n7371), .A(n7369), .ZN(n14875) );
  OR2_X1 U8127 ( .A1(n14876), .A2(n14859), .ZN(n7371) );
  INV_X1 U8128 ( .A(n14876), .ZN(n7370) );
  XNOR2_X1 U8129 ( .A(n14636), .B(n14635), .ZN(n6813) );
  NOR2_X1 U8130 ( .A1(n14875), .A2(n7372), .ZN(n14597) );
  NOR2_X1 U8131 ( .A1(n14660), .A2(n14595), .ZN(n7372) );
  AND3_X1 U8132 ( .A1(n8756), .A2(n8755), .A3(n8754), .ZN(n10831) );
  NAND2_X1 U8133 ( .A1(n10658), .A2(n12639), .ZN(n14895) );
  AOI21_X1 U8134 ( .B1(n12780), .B2(n11887), .A(n9290), .ZN(n11718) );
  INV_X1 U8135 ( .A(n9349), .ZN(n12723) );
  INV_X1 U8136 ( .A(n9348), .ZN(n12727) );
  OR2_X1 U8137 ( .A1(n15601), .A2(n12621), .ZN(n12770) );
  AND2_X1 U8138 ( .A1(n9211), .A2(n9210), .ZN(n12771) );
  OR2_X1 U8139 ( .A1(n9209), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U8140 ( .A1(n7098), .A2(n7097), .ZN(n8762) );
  AND2_X1 U8141 ( .A1(n7873), .A2(n7870), .ZN(n7097) );
  NOR2_X1 U8142 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(n7871), .ZN(n7870) );
  NAND2_X1 U8143 ( .A1(n8759), .A2(n7202), .ZN(n7871) );
  NAND2_X1 U8144 ( .A1(n8735), .A2(n8734), .ZN(n14638) );
  XNOR2_X1 U8145 ( .A(n6916), .B(n6730), .ZN(n7581) );
  NAND2_X1 U8146 ( .A1(n12868), .A2(n12867), .ZN(n6916) );
  OR2_X1 U8147 ( .A1(n10870), .A2(n8611), .ZN(n8119) );
  AOI21_X1 U8148 ( .B1(n11013), .B2(n11011), .A(n7302), .ZN(n11015) );
  NOR2_X1 U8149 ( .A1(n7302), .A2(n6747), .ZN(n7300) );
  NAND2_X1 U8150 ( .A1(n11013), .A2(n7301), .ZN(n7297) );
  NAND2_X1 U8151 ( .A1(n8206), .A2(n8205), .ZN(n11195) );
  NAND2_X1 U8152 ( .A1(n7576), .A2(n7577), .ZN(n12912) );
  INV_X1 U8153 ( .A(n12893), .ZN(n7576) );
  NAND2_X1 U8154 ( .A1(n12893), .A2(n12791), .ZN(n7570) );
  NOR2_X1 U8155 ( .A1(n6628), .A2(n7318), .ZN(n7317) );
  INV_X1 U8156 ( .A(n12950), .ZN(n7318) );
  OR2_X1 U8157 ( .A1(n12800), .A2(n6628), .ZN(n7569) );
  NAND2_X1 U8158 ( .A1(n6932), .A2(n10975), .ZN(n11013) );
  NAND2_X1 U8159 ( .A1(n8182), .A2(n8181), .ZN(n11066) );
  NAND2_X1 U8160 ( .A1(n7571), .A2(n6587), .ZN(n12951) );
  NOR2_X1 U8161 ( .A1(n7575), .A2(n6729), .ZN(n7572) );
  NAND2_X1 U8162 ( .A1(n8513), .A2(n8512), .ZN(n13307) );
  OR2_X1 U8163 ( .A1(n8663), .A2(n9939), .ZN(n7194) );
  NAND2_X1 U8164 ( .A1(n8671), .A2(n8668), .ZN(n8669) );
  NAND2_X1 U8165 ( .A1(n8541), .A2(n8540), .ZN(n13089) );
  NAND2_X1 U8166 ( .A1(n8522), .A2(n8521), .ZN(n13087) );
  NAND2_X1 U8167 ( .A1(n8453), .A2(n8452), .ZN(n13051) );
  OR2_X1 U8168 ( .A1(n7997), .A2(n9578), .ZN(n7255) );
  NOR2_X1 U8169 ( .A1(n13288), .A2(n6650), .ZN(n7348) );
  INV_X1 U8170 ( .A(n7783), .ZN(n7781) );
  NAND2_X1 U8171 ( .A1(n7779), .A2(n13092), .ZN(n7778) );
  INV_X1 U8172 ( .A(n13105), .ZN(n7779) );
  AND4_X1 U8173 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n13891) );
  AND2_X1 U8174 ( .A1(n11234), .A2(n11233), .ZN(n14797) );
  NAND2_X1 U8175 ( .A1(n10010), .A2(n10009), .ZN(n13784) );
  NAND2_X1 U8176 ( .A1(n7488), .A2(n7037), .ZN(n7036) );
  NAND2_X1 U8177 ( .A1(n7488), .A2(n7035), .ZN(n7034) );
  INV_X1 U8178 ( .A(n13775), .ZN(n7038) );
  AND2_X1 U8179 ( .A1(n13772), .A2(n15200), .ZN(n13782) );
  AOI21_X1 U8180 ( .B1(n14048), .B2(n14049), .A(n7212), .ZN(n7211) );
  NAND2_X1 U8181 ( .A1(n14047), .A2(n14046), .ZN(n7212) );
  INV_X1 U8182 ( .A(n13929), .ZN(n14058) );
  NAND2_X1 U8183 ( .A1(n13616), .A2(n13615), .ZN(n14254) );
  NAND2_X1 U8184 ( .A1(n13498), .A2(n13497), .ZN(n14414) );
  NAND2_X1 U8185 ( .A1(n14934), .A2(n11620), .ZN(n11622) );
  OR2_X1 U8186 ( .A1(n15105), .A2(n10776), .ZN(n15096) );
  INV_X1 U8187 ( .A(n14379), .ZN(n15105) );
  INV_X1 U8188 ( .A(n14418), .ZN(n15065) );
  AND2_X1 U8189 ( .A1(n7596), .A2(n7594), .ZN(n7204) );
  NAND2_X1 U8190 ( .A1(n7595), .A2(n15196), .ZN(n7361) );
  NAND2_X1 U8191 ( .A1(n7713), .A2(n15207), .ZN(n7712) );
  NAND2_X1 U8192 ( .A1(n14462), .A2(n6894), .ZN(n14541) );
  INV_X1 U8193 ( .A(n6895), .ZN(n6894) );
  OAI21_X1 U8194 ( .B1(n14463), .B2(n14795), .A(n14461), .ZN(n6895) );
  NAND2_X1 U8195 ( .A1(n7847), .A2(n6668), .ZN(n14557) );
  INV_X1 U8196 ( .A(n9664), .ZN(n7847) );
  INV_X1 U8197 ( .A(n7848), .ZN(n7846) );
  XNOR2_X1 U8198 ( .A(n8609), .B(n8608), .ZN(n13837) );
  NAND2_X1 U8199 ( .A1(n9413), .A2(n9664), .ZN(n14567) );
  INV_X1 U8200 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9399) );
  OAI21_X1 U8201 ( .B1(n9401), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9400) );
  XNOR2_X1 U8202 ( .A(n9403), .B(n9402), .ZN(n14574) );
  INV_X1 U8203 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9402) );
  XNOR2_X1 U8204 ( .A(n14720), .B(n6908), .ZN(n15627) );
  OAI21_X1 U8205 ( .B1(n14770), .B2(n14771), .A(n6907), .ZN(n6906) );
  INV_X1 U8206 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6907) );
  NOR2_X1 U8207 ( .A1(n15623), .A2(n15624), .ZN(n15622) );
  XNOR2_X1 U8208 ( .A(n14730), .B(n7462), .ZN(n14775) );
  NAND2_X1 U8209 ( .A1(n14778), .A2(n14777), .ZN(n14776) );
  XNOR2_X1 U8210 ( .A(n7454), .B(n14750), .ZN(n14971) );
  NAND2_X1 U8211 ( .A1(n14971), .A2(n14970), .ZN(n14969) );
  OAI21_X1 U8212 ( .B1(n14811), .B2(n14810), .A(n11338), .ZN(n7465) );
  AOI21_X1 U8213 ( .B1(n15365), .B2(n8615), .A(n7128), .ZN(n7127) );
  NOR2_X1 U8214 ( .A1(n10350), .A2(n8615), .ZN(n7128) );
  NAND2_X1 U8215 ( .A1(n8128), .A2(n7744), .ZN(n7743) );
  NAND2_X1 U8216 ( .A1(n7747), .A2(n7746), .ZN(n7745) );
  INV_X1 U8217 ( .A(n8128), .ZN(n7746) );
  AND2_X1 U8218 ( .A1(n7558), .A2(n13909), .ZN(n7557) );
  OAI21_X1 U8219 ( .B1(n13905), .B2(n7560), .A(n6685), .ZN(n13911) );
  AOI21_X1 U8220 ( .B1(n6779), .B2(n13914), .A(n6778), .ZN(n6777) );
  INV_X1 U8221 ( .A(n13918), .ZN(n6778) );
  NOR2_X1 U8222 ( .A1(n13915), .A2(n13920), .ZN(n6779) );
  NAND2_X1 U8223 ( .A1(n7565), .A2(n13919), .ZN(n6780) );
  NOR2_X1 U8224 ( .A1(n6776), .A2(n13919), .ZN(n6775) );
  NOR2_X1 U8225 ( .A1(n7566), .A2(n13915), .ZN(n6776) );
  OAI22_X1 U8226 ( .A1(n13922), .A2(n7554), .B1(n13923), .B2(n7555), .ZN(
        n13928) );
  AND2_X1 U8227 ( .A1(n13923), .A2(n7555), .ZN(n7554) );
  NAND2_X1 U8228 ( .A1(n6771), .A2(n6768), .ZN(n13922) );
  INV_X1 U8229 ( .A(n8195), .ZN(n7291) );
  NOR2_X1 U8230 ( .A1(n8195), .A2(n7741), .ZN(n7292) );
  AND2_X1 U8231 ( .A1(n8278), .A2(n8279), .ZN(n7761) );
  NAND2_X1 U8232 ( .A1(n6781), .A2(n6647), .ZN(n13959) );
  NAND2_X1 U8233 ( .A1(n6782), .A2(n6646), .ZN(n6781) );
  NAND2_X1 U8234 ( .A1(n8258), .A2(n6688), .ZN(n7159) );
  AND2_X1 U8235 ( .A1(n8236), .A2(n8237), .ZN(n7767) );
  NAND2_X1 U8236 ( .A1(n7757), .A2(n8305), .ZN(n7756) );
  NAND2_X1 U8237 ( .A1(n7761), .A2(n7758), .ZN(n7757) );
  NAND2_X1 U8238 ( .A1(n7760), .A2(n7759), .ZN(n7758) );
  INV_X1 U8239 ( .A(n8278), .ZN(n7759) );
  INV_X1 U8240 ( .A(n8279), .ZN(n7760) );
  NAND2_X1 U8241 ( .A1(n13965), .A2(n13808), .ZN(n6799) );
  NAND2_X1 U8242 ( .A1(n14189), .A2(n6798), .ZN(n6797) );
  NAND2_X1 U8243 ( .A1(n8393), .A2(n8394), .ZN(n7765) );
  OAI21_X1 U8244 ( .B1(n8328), .B2(n7755), .A(n7190), .ZN(n8351) );
  NOR2_X1 U8245 ( .A1(n7191), .A2(n8350), .ZN(n7190) );
  INV_X1 U8246 ( .A(n8394), .ZN(n7766) );
  INV_X1 U8247 ( .A(n8393), .ZN(n7764) );
  NAND2_X1 U8248 ( .A1(n13986), .A2(n7546), .ZN(n7545) );
  NAND2_X1 U8249 ( .A1(n6634), .A2(n7547), .ZN(n7546) );
  OAI21_X1 U8250 ( .B1(n6686), .B2(n6784), .A(n6783), .ZN(n13982) );
  NOR2_X1 U8251 ( .A1(n6785), .A2(n6620), .ZN(n6784) );
  AOI22_X1 U8252 ( .A1(n6785), .A2(n6787), .B1(n6620), .B2(n7567), .ZN(n6783)
         );
  NAND2_X1 U8253 ( .A1(n13980), .A2(n7548), .ZN(n7547) );
  INV_X1 U8254 ( .A(n13981), .ZN(n7548) );
  INV_X1 U8255 ( .A(n8505), .ZN(n7286) );
  INV_X1 U8256 ( .A(n7142), .ZN(n7150) );
  NOR2_X1 U8257 ( .A1(n8416), .A2(n7144), .ZN(n7143) );
  INV_X1 U8258 ( .A(n8418), .ZN(n7144) );
  NAND2_X1 U8259 ( .A1(n7279), .A2(n7149), .ZN(n7145) );
  INV_X1 U8260 ( .A(n7152), .ZN(n7149) );
  INV_X1 U8261 ( .A(n8329), .ZN(n8330) );
  AND2_X1 U8262 ( .A1(n8506), .A2(n7286), .ZN(n7285) );
  AND2_X1 U8263 ( .A1(n6767), .A2(n6766), .ZN(n13998) );
  NAND2_X1 U8264 ( .A1(n6593), .A2(n7550), .ZN(n6766) );
  AND2_X1 U8265 ( .A1(n8507), .A2(SI_26_), .ZN(n7647) );
  INV_X1 U8266 ( .A(n11959), .ZN(n6990) );
  NOR2_X1 U8267 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8739) );
  NOR2_X1 U8268 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8706) );
  NOR2_X1 U8269 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8707) );
  AOI21_X1 U8270 ( .B1(n13076), .B2(n13074), .A(n7341), .ZN(n7340) );
  INV_X1 U8271 ( .A(n13213), .ZN(n7341) );
  INV_X1 U8272 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7890) );
  INV_X1 U8273 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7273) );
  INV_X1 U8274 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7893) );
  NAND2_X1 U8275 ( .A1(n14019), .A2(n13863), .ZN(n14015) );
  INV_X1 U8276 ( .A(n14197), .ZN(n6946) );
  INV_X1 U8277 ( .A(n11026), .ZN(n7593) );
  INV_X1 U8278 ( .A(n7647), .ZN(n7641) );
  AOI21_X1 U8279 ( .B1(n8508), .B2(n7647), .A(n7646), .ZN(n7645) );
  INV_X1 U8280 ( .A(n8529), .ZN(n7646) );
  AOI21_X1 U8281 ( .B1(n8508), .B2(n8507), .A(SI_26_), .ZN(n7648) );
  INV_X1 U8282 ( .A(SI_16_), .ZN(n8309) );
  INV_X1 U8283 ( .A(n6835), .ZN(n6831) );
  AND2_X1 U8284 ( .A1(n12417), .A2(n11907), .ZN(n12058) );
  NAND2_X1 U8285 ( .A1(n12394), .A2(n12395), .ZN(n12397) );
  NAND2_X1 U8286 ( .A1(n15480), .A2(n6751), .ZN(n14645) );
  NAND2_X1 U8287 ( .A1(n15514), .A2(n6970), .ZN(n14649) );
  OR2_X1 U8288 ( .A1(n14648), .A2(n14912), .ZN(n6970) );
  INV_X1 U8289 ( .A(n15549), .ZN(n7376) );
  NAND2_X1 U8290 ( .A1(n9348), .A2(n12095), .ZN(n7084) );
  INV_X1 U8291 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12199) );
  NAND2_X1 U8292 ( .A1(n9102), .A2(n12199), .ZN(n9122) );
  AND2_X1 U8293 ( .A1(n12503), .A2(n6592), .ZN(n7862) );
  NAND2_X1 U8294 ( .A1(n12520), .A2(n12519), .ZN(n7861) );
  INV_X1 U8295 ( .A(n7088), .ZN(n7087) );
  NOR2_X1 U8296 ( .A1(n12531), .A2(n7089), .ZN(n7088) );
  INV_X1 U8297 ( .A(n9341), .ZN(n7089) );
  AOI21_X1 U8298 ( .B1(n7435), .B2(n7438), .A(n7434), .ZN(n7433) );
  INV_X1 U8299 ( .A(n12591), .ZN(n7434) );
  INV_X1 U8300 ( .A(n7071), .ZN(n7070) );
  OAI21_X1 U8301 ( .B1(n11980), .B2(n7072), .A(n11917), .ZN(n7071) );
  INV_X1 U8302 ( .A(n9325), .ZN(n7072) );
  AND2_X1 U8303 ( .A1(n7853), .A2(n11352), .ZN(n7852) );
  OR2_X1 U8304 ( .A1(n9317), .A2(n7854), .ZN(n7853) );
  INV_X1 U8305 ( .A(n9324), .ZN(n7854) );
  NAND2_X1 U8306 ( .A1(n7430), .A2(n7432), .ZN(n7428) );
  INV_X1 U8307 ( .A(n11951), .ZN(n7432) );
  NAND2_X1 U8308 ( .A1(n10706), .A2(n9305), .ZN(n9308) );
  NAND2_X1 U8309 ( .A1(n10315), .A2(n11935), .ZN(n9267) );
  NAND2_X1 U8310 ( .A1(n11109), .A2(n9314), .ZN(n11120) );
  INV_X1 U8311 ( .A(n9175), .ZN(n7400) );
  INV_X1 U8312 ( .A(n9116), .ZN(n7106) );
  INV_X1 U8313 ( .A(n7105), .ZN(n7104) );
  OAI21_X1 U8314 ( .B1(n9114), .B2(n7106), .A(n9127), .ZN(n7105) );
  INV_X1 U8315 ( .A(n7111), .ZN(n7110) );
  AOI21_X1 U8316 ( .B1(n7111), .B2(n7113), .A(n7109), .ZN(n7108) );
  AOI21_X1 U8317 ( .B1(n7393), .B2(n8953), .A(n7392), .ZN(n7391) );
  INV_X1 U8318 ( .A(n8976), .ZN(n7392) );
  INV_X1 U8319 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7684) );
  NOR2_X1 U8320 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n6820) );
  INV_X1 U8321 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n12307) );
  INV_X1 U8322 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8917) );
  OR2_X1 U8323 ( .A1(n8882), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8896) );
  XNOR2_X1 U8324 ( .A(n10564), .B(n11315), .ZN(n10614) );
  NOR2_X1 U8325 ( .A1(n8597), .A2(n8637), .ZN(n7161) );
  NAND2_X1 U8326 ( .A1(n6764), .A2(n7183), .ZN(n8528) );
  INV_X1 U8327 ( .A(n7141), .ZN(n7140) );
  NAND2_X1 U8328 ( .A1(n6582), .A2(n7742), .ZN(n7619) );
  INV_X1 U8329 ( .A(n7792), .ZN(n7233) );
  INV_X1 U8330 ( .A(n7794), .ZN(n7790) );
  INV_X1 U8331 ( .A(n13082), .ZN(n7725) );
  AOI21_X1 U8332 ( .B1(n7340), .B2(n7337), .A(n7336), .ZN(n7335) );
  INV_X1 U8333 ( .A(n13076), .ZN(n7337) );
  INV_X1 U8334 ( .A(n13077), .ZN(n7336) );
  INV_X1 U8335 ( .A(n7340), .ZN(n7338) );
  NOR2_X2 U8336 ( .A1(n13250), .A2(n13343), .ZN(n7532) );
  INV_X1 U8337 ( .A(n11301), .ZN(n7327) );
  OR2_X1 U8338 ( .A1(n7536), .A2(n12980), .ZN(n7329) );
  INV_X1 U8339 ( .A(n8063), .ZN(n7771) );
  AOI22_X1 U8340 ( .A1(n7803), .A2(n7802), .B1(n13088), .B2(n13146), .ZN(
        n13128) );
  NAND2_X1 U8341 ( .A1(n13307), .A2(n13087), .ZN(n7802) );
  NAND2_X1 U8342 ( .A1(n12378), .A2(n8693), .ZN(n7920) );
  INV_X1 U8343 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7917) );
  INV_X1 U8344 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8673) );
  INV_X1 U8345 ( .A(n8672), .ZN(n8675) );
  INV_X1 U8346 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U8347 ( .A1(n8672), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7926) );
  INV_X1 U8348 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n12329) );
  INV_X1 U8349 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7887) );
  INV_X1 U8350 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7896) );
  OR2_X1 U8351 ( .A1(n13775), .A2(n7488), .ZN(n7482) );
  NOR2_X1 U8352 ( .A1(n10072), .A2(n15076), .ZN(n10721) );
  NAND2_X1 U8353 ( .A1(n13539), .A2(n13540), .ZN(n7509) );
  INV_X1 U8354 ( .A(n11481), .ZN(n7027) );
  NOR2_X1 U8355 ( .A1(n11653), .A2(n7493), .ZN(n7492) );
  INV_X1 U8356 ( .A(n11650), .ZN(n7493) );
  NAND2_X1 U8357 ( .A1(n14004), .A2(n14006), .ZN(n7220) );
  INV_X1 U8358 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n12306) );
  INV_X1 U8359 ( .A(n7831), .ZN(n6951) );
  NAND2_X1 U8360 ( .A1(n6882), .A2(n6663), .ZN(n7351) );
  INV_X1 U8361 ( .A(n14231), .ZN(n6881) );
  NAND2_X1 U8362 ( .A1(n6889), .A2(n14179), .ZN(n6884) );
  NAND2_X1 U8363 ( .A1(n14258), .A2(n6885), .ZN(n6882) );
  NOR2_X1 U8364 ( .A1(n6892), .A2(n6886), .ZN(n6885) );
  INV_X1 U8365 ( .A(n14179), .ZN(n6886) );
  NOR2_X1 U8366 ( .A1(n14358), .A2(n7270), .ZN(n7269) );
  INV_X1 U8367 ( .A(n7271), .ZN(n7270) );
  NOR2_X1 U8368 ( .A1(n14375), .A2(n14522), .ZN(n7271) );
  NOR2_X1 U8369 ( .A1(n14188), .A2(n7845), .ZN(n7844) );
  INV_X1 U8370 ( .A(n14186), .ZN(n7845) );
  OR2_X1 U8371 ( .A1(n14534), .A2(n13726), .ZN(n14166) );
  INV_X1 U8372 ( .A(n6942), .ZN(n6941) );
  OAI21_X1 U8373 ( .B1(n13820), .B2(n6943), .A(n11520), .ZN(n6942) );
  INV_X1 U8374 ( .A(n11421), .ZN(n6943) );
  NOR2_X1 U8375 ( .A1(n11434), .A2(n13934), .ZN(n7599) );
  NOR2_X1 U8376 ( .A1(n14952), .A2(n13925), .ZN(n7825) );
  INV_X1 U8377 ( .A(n11162), .ZN(n7827) );
  AOI21_X1 U8378 ( .B1(n6865), .B2(n6872), .A(n6864), .ZN(n6863) );
  INV_X1 U8379 ( .A(n6867), .ZN(n6865) );
  NOR2_X1 U8380 ( .A1(n7259), .A2(n10777), .ZN(n7260) );
  NOR2_X1 U8381 ( .A1(n14219), .A2(n6961), .ZN(n6960) );
  INV_X1 U8382 ( .A(n7828), .ZN(n6961) );
  NAND2_X1 U8383 ( .A1(n7593), .A2(n7592), .ZN(n11052) );
  NAND2_X1 U8384 ( .A1(n8581), .A2(n7628), .ZN(n7627) );
  INV_X1 U8385 ( .A(n8553), .ZN(n7628) );
  INV_X1 U8386 ( .A(n8568), .ZN(n7629) );
  AND2_X1 U8387 ( .A1(n7642), .A2(n7640), .ZN(n7639) );
  NAND2_X1 U8388 ( .A1(n7648), .A2(n7643), .ZN(n7642) );
  NAND2_X1 U8389 ( .A1(n7645), .A2(n7641), .ZN(n7640) );
  INV_X1 U8390 ( .A(n8507), .ZN(n7643) );
  NOR2_X1 U8391 ( .A1(n7648), .A2(n7645), .ZN(n7644) );
  NAND2_X1 U8392 ( .A1(n8509), .A2(n7639), .ZN(n7637) );
  OR2_X1 U8393 ( .A1(n8464), .A2(n7624), .ZN(n7622) );
  INV_X1 U8394 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9416) );
  INV_X1 U8395 ( .A(n7632), .ZN(n7631) );
  NOR2_X1 U8396 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7813) );
  NOR2_X1 U8397 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n7812) );
  NOR2_X1 U8398 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7811) );
  INV_X1 U8399 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9393) );
  INV_X1 U8400 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9394) );
  INV_X1 U8401 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9469) );
  OR2_X1 U8402 ( .A1(n10463), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n10788) );
  AND2_X1 U8403 ( .A1(n10332), .A2(n10333), .ZN(n10337) );
  INV_X1 U8404 ( .A(n7612), .ZN(n6984) );
  AOI21_X1 U8405 ( .B1(n7612), .B2(n6983), .A(n6683), .ZN(n6982) );
  INV_X1 U8406 ( .A(n7614), .ZN(n6983) );
  INV_X1 U8407 ( .A(n7616), .ZN(n7615) );
  INV_X1 U8408 ( .A(n8129), .ZN(n7207) );
  NAND2_X1 U8409 ( .A1(n8075), .A2(n8078), .ZN(n6994) );
  INV_X1 U8410 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U8411 ( .A1(n7988), .A2(n7987), .ZN(n7205) );
  NAND2_X1 U8412 ( .A1(n7605), .A2(n7218), .ZN(n7944) );
  NAND2_X1 U8413 ( .A1(n7353), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7218) );
  INV_X1 U8414 ( .A(n14724), .ZN(n6904) );
  NAND2_X1 U8415 ( .A1(n7467), .A2(n14675), .ZN(n14676) );
  NAND2_X1 U8416 ( .A1(n14710), .A2(n14711), .ZN(n7467) );
  INV_X1 U8417 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7466) );
  AOI22_X1 U8418 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14731), .B1(n14733), .B2(
        n14679), .ZN(n14681) );
  OR2_X1 U8419 ( .A1(n8854), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8861) );
  OR2_X1 U8420 ( .A1(n9066), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U8421 ( .A1(n7650), .A2(n7649), .ZN(n9207) );
  AOI21_X1 U8422 ( .B1(n7651), .B2(n7654), .A(n9188), .ZN(n7649) );
  NAND2_X1 U8423 ( .A1(n9173), .A2(n7651), .ZN(n7650) );
  AND3_X1 U8424 ( .A1(n8886), .A2(n8885), .A3(n8884), .ZN(n11971) );
  INV_X1 U8425 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U8426 ( .A1(n8827), .A2(n11106), .ZN(n6829) );
  NAND2_X1 U8427 ( .A1(n6817), .A2(n6816), .ZN(n11770) );
  INV_X1 U8428 ( .A(n11799), .ZN(n7668) );
  NAND2_X1 U8429 ( .A1(n9135), .A2(n9134), .ZN(n11798) );
  OR2_X1 U8430 ( .A1(n9137), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9151) );
  NOR2_X1 U8431 ( .A1(n9151), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9165) );
  AND2_X1 U8432 ( .A1(n8888), .A2(n8887), .ZN(n8906) );
  AND2_X1 U8433 ( .A1(n9093), .A2(n11809), .ZN(n9102) );
  NOR2_X1 U8434 ( .A1(n9080), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9093) );
  AOI21_X1 U8435 ( .B1(n6673), .B2(n7679), .A(n6585), .ZN(n7676) );
  NOR2_X1 U8436 ( .A1(n7677), .A2(n6836), .ZN(n6835) );
  INV_X1 U8437 ( .A(n9025), .ZN(n6836) );
  INV_X1 U8438 ( .A(n7679), .ZN(n7677) );
  AND2_X1 U8439 ( .A1(n11856), .A2(n7652), .ZN(n7651) );
  NAND2_X1 U8440 ( .A1(n7653), .A2(n9174), .ZN(n7652) );
  INV_X1 U8441 ( .A(n11772), .ZN(n7653) );
  INV_X1 U8442 ( .A(n9174), .ZN(n7654) );
  NAND2_X1 U8443 ( .A1(n11770), .A2(n11771), .ZN(n9173) );
  NOR2_X1 U8444 ( .A1(n9017), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9034) );
  NAND2_X1 U8445 ( .A1(n7381), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10268) );
  INV_X1 U8446 ( .A(n10266), .ZN(n7381) );
  NAND2_X1 U8447 ( .A1(n10173), .A2(n10174), .ZN(n10365) );
  NAND2_X1 U8448 ( .A1(n6804), .A2(n6667), .ZN(n15415) );
  NOR2_X1 U8449 ( .A1(n15412), .A2(n10185), .ZN(n6807) );
  NAND2_X1 U8450 ( .A1(n15430), .A2(n15429), .ZN(n15428) );
  OR2_X1 U8451 ( .A1(n15408), .A2(n7366), .ZN(n7365) );
  OR2_X1 U8452 ( .A1(n15426), .A2(n8820), .ZN(n7366) );
  OR2_X1 U8453 ( .A1(n15408), .A2(n8820), .ZN(n15406) );
  NAND2_X1 U8454 ( .A1(n6975), .A2(n6974), .ZN(n6973) );
  NAND2_X1 U8455 ( .A1(n15433), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6974) );
  INV_X1 U8456 ( .A(n15439), .ZN(n6975) );
  XNOR2_X1 U8457 ( .A(n6973), .B(n15453), .ZN(n15456) );
  INV_X1 U8458 ( .A(n7052), .ZN(n7051) );
  NAND2_X1 U8459 ( .A1(n7053), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7050) );
  XNOR2_X1 U8460 ( .A(n12392), .B(n12381), .ZN(n10556) );
  NAND2_X1 U8461 ( .A1(n10556), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n12394) );
  INV_X1 U8462 ( .A(n7368), .ZN(n14578) );
  NAND2_X1 U8463 ( .A1(n15471), .A2(n14643), .ZN(n15481) );
  NAND2_X1 U8464 ( .A1(n15481), .A2(n15482), .ZN(n15480) );
  NAND2_X1 U8465 ( .A1(n14601), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7367) );
  OR2_X1 U8466 ( .A1(n12385), .A2(n12384), .ZN(n7368) );
  XNOR2_X1 U8467 ( .A(n14645), .B(n14646), .ZN(n15498) );
  NAND2_X1 U8468 ( .A1(n15504), .A2(n14612), .ZN(n15523) );
  NAND2_X1 U8469 ( .A1(n15515), .A2(n15516), .ZN(n15514) );
  AND2_X1 U8470 ( .A1(n15524), .A2(n14614), .ZN(n15542) );
  NAND2_X1 U8471 ( .A1(n15542), .A2(n15541), .ZN(n15540) );
  XNOR2_X1 U8472 ( .A(n14649), .B(n14650), .ZN(n15533) );
  NAND2_X1 U8473 ( .A1(n15533), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n15532) );
  INV_X1 U8474 ( .A(n7041), .ZN(n14584) );
  NAND2_X1 U8475 ( .A1(n7055), .A2(n7054), .ZN(n7061) );
  INV_X1 U8476 ( .A(n14588), .ZN(n7054) );
  INV_X1 U8477 ( .A(n14820), .ZN(n7055) );
  NAND2_X1 U8478 ( .A1(n6815), .A2(n6814), .ZN(n14626) );
  NAND2_X1 U8479 ( .A1(n14624), .A2(n14623), .ZN(n6814) );
  NAND2_X1 U8480 ( .A1(n14823), .A2(n14654), .ZN(n14842) );
  NAND2_X1 U8481 ( .A1(n7061), .A2(n7060), .ZN(n14837) );
  AND2_X1 U8482 ( .A1(n14864), .A2(n14863), .ZN(n14865) );
  XNOR2_X1 U8483 ( .A(n14630), .B(n14877), .ZN(n14885) );
  INV_X1 U8484 ( .A(n7058), .ZN(n7057) );
  OR2_X1 U8485 ( .A1(n14588), .A2(n7059), .ZN(n7056) );
  OAI21_X1 U8486 ( .B1(n7060), .B2(n7059), .A(n14868), .ZN(n7058) );
  OR2_X1 U8487 ( .A1(n14858), .A2(n14859), .ZN(n7373) );
  NOR2_X1 U8488 ( .A1(n14865), .A2(n14629), .ZN(n14630) );
  AOI21_X1 U8489 ( .B1(n7867), .B2(n11907), .A(n6672), .ZN(n7866) );
  AOI21_X1 U8490 ( .B1(n7417), .B2(n7419), .A(n12062), .ZN(n7416) );
  NOR2_X1 U8491 ( .A1(n7869), .A2(n7422), .ZN(n7417) );
  INV_X1 U8492 ( .A(n7420), .ZN(n7419) );
  AOI21_X1 U8493 ( .B1(n7121), .B2(n11907), .A(n12064), .ZN(n7420) );
  NAND2_X1 U8494 ( .A1(n7423), .A2(n12057), .ZN(n7121) );
  OR2_X1 U8495 ( .A1(n12408), .A2(n9248), .ZN(n12419) );
  OAI21_X1 U8496 ( .B1(n7011), .B2(n12057), .A(n7423), .ZN(n12425) );
  AND2_X1 U8497 ( .A1(n7444), .A2(n7000), .ZN(n6999) );
  NAND2_X1 U8498 ( .A1(n7447), .A2(n7001), .ZN(n7000) );
  AND2_X1 U8499 ( .A1(n7861), .A2(n7862), .ZN(n12506) );
  OAI21_X1 U8500 ( .B1(n12542), .B2(n9340), .A(n12018), .ZN(n12530) );
  AND2_X1 U8501 ( .A1(n12543), .A2(n9341), .ZN(n12533) );
  NAND2_X1 U8502 ( .A1(n12543), .A2(n7088), .ZN(n12532) );
  NAND2_X1 U8503 ( .A1(n12560), .A2(n12020), .ZN(n12542) );
  NAND2_X1 U8504 ( .A1(n9051), .A2(n12256), .ZN(n9066) );
  AND2_X1 U8505 ( .A1(n9034), .A2(n9033), .ZN(n9051) );
  INV_X1 U8506 ( .A(n12013), .ZN(n12561) );
  NAND2_X1 U8507 ( .A1(n12590), .A2(n12004), .ZN(n12574) );
  INV_X1 U8508 ( .A(n9335), .ZN(n12573) );
  NOR2_X1 U8509 ( .A1(n12600), .A2(n7093), .ZN(n7092) );
  INV_X1 U8510 ( .A(n9330), .ZN(n7093) );
  INV_X1 U8511 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11818) );
  NOR2_X1 U8512 ( .A1(n8963), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8984) );
  AND3_X1 U8513 ( .A1(n8945), .A2(n8944), .A3(n8943), .ZN(n11414) );
  OR2_X1 U8514 ( .A1(n8925), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8946) );
  OR2_X1 U8515 ( .A1(n8946), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U8516 ( .A1(n11470), .A2(n11980), .ZN(n7069) );
  AND4_X1 U8517 ( .A1(n8968), .A2(n8967), .A3(n8966), .A4(n8965), .ZN(n11820)
         );
  AND3_X1 U8518 ( .A1(n8924), .A2(n8923), .A3(n8922), .ZN(n11472) );
  NAND2_X1 U8519 ( .A1(n11987), .A2(n11410), .ZN(n11980) );
  INV_X1 U8520 ( .A(n7064), .ZN(n7063) );
  OAI21_X1 U8521 ( .B1(n6581), .B2(n6630), .A(n9316), .ZN(n7064) );
  AND4_X1 U8522 ( .A1(n8893), .A2(n8892), .A3(n8891), .A4(n8890), .ZN(n11564)
         );
  NAND2_X1 U8523 ( .A1(n10829), .A2(n6581), .ZN(n11109) );
  NAND2_X1 U8524 ( .A1(n10829), .A2(n9313), .ZN(n11107) );
  INV_X1 U8525 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n11099) );
  AND3_X1 U8526 ( .A1(n8836), .A2(n8835), .A3(n8834), .ZN(n11112) );
  NAND2_X1 U8527 ( .A1(n9308), .A2(n9307), .ZN(n7865) );
  NAND2_X1 U8528 ( .A1(n7410), .A2(n11942), .ZN(n10663) );
  AND2_X1 U8529 ( .A1(n10403), .A2(n11927), .ZN(n10705) );
  NAND2_X1 U8530 ( .A1(n10581), .A2(n10580), .ZN(n10658) );
  INV_X1 U8531 ( .A(n12621), .ZN(n14898) );
  AND3_X1 U8532 ( .A1(n8819), .A2(n8818), .A3(n8817), .ZN(n9311) );
  INV_X1 U8533 ( .A(n8806), .ZN(n10708) );
  INV_X1 U8534 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U8535 ( .A1(n7873), .A2(n7202), .ZN(n7452) );
  OAI21_X1 U8536 ( .B1(n9190), .B2(n9189), .A(n9191), .ZN(n9279) );
  XNOR2_X1 U8537 ( .A(n9232), .B(n8710), .ZN(n10161) );
  NAND2_X1 U8538 ( .A1(n6748), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9232) );
  NOR2_X1 U8539 ( .A1(n8730), .A2(n8728), .ZN(n9353) );
  NAND2_X1 U8540 ( .A1(n7383), .A2(n9011), .ZN(n9028) );
  NAND2_X1 U8541 ( .A1(n8903), .A2(n8902), .ZN(n8916) );
  INV_X1 U8542 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8901) );
  XNOR2_X1 U8543 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8899) );
  AOI21_X1 U8544 ( .B1(n7387), .B2(n7385), .A(n6693), .ZN(n7384) );
  INV_X1 U8545 ( .A(n7387), .ZN(n7386) );
  XNOR2_X1 U8546 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8828) );
  NAND2_X1 U8547 ( .A1(n8742), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8797) );
  INV_X1 U8548 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11321) );
  NAND2_X1 U8549 ( .A1(n9901), .A2(n9919), .ZN(n9902) );
  AOI21_X1 U8550 ( .B1(n7568), .B2(n7316), .A(n6687), .ZN(n7315) );
  INV_X1 U8551 ( .A(n7317), .ZN(n7316) );
  NAND2_X1 U8552 ( .A1(n6931), .A2(n7568), .ZN(n6930) );
  INV_X1 U8553 ( .A(n12951), .ZN(n6931) );
  NAND2_X1 U8554 ( .A1(n8382), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8404) );
  INV_X1 U8555 ( .A(n8384), .ZN(n8382) );
  NAND2_X1 U8556 ( .A1(n12818), .A2(n6923), .ZN(n12918) );
  XNOR2_X1 U8557 ( .A(n12806), .B(n15348), .ZN(n9919) );
  OR2_X1 U8558 ( .A1(n9904), .A2(n9903), .ZN(n9914) );
  OAI21_X1 U8559 ( .B1(n10293), .B2(n6678), .A(n7305), .ZN(n10620) );
  INV_X1 U8560 ( .A(n7303), .ZN(n7305) );
  OAI21_X1 U8561 ( .B1(n10637), .B2(n7304), .A(n10641), .ZN(n7303) );
  NAND2_X1 U8562 ( .A1(n10620), .A2(n10621), .ZN(n10682) );
  NAND2_X1 U8563 ( .A1(n8207), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8248) );
  OR2_X1 U8564 ( .A1(n8427), .A2(n12942), .ZN(n8447) );
  NAND2_X1 U8565 ( .A1(n6930), .A2(n6579), .ZN(n12937) );
  NAND2_X1 U8566 ( .A1(n10284), .A2(n7584), .ZN(n10324) );
  AND2_X1 U8567 ( .A1(n8574), .A2(n8536), .ZN(n13129) );
  AND2_X1 U8568 ( .A1(n13307), .A2(n13088), .ZN(n7349) );
  NAND2_X1 U8569 ( .A1(n13146), .A2(n13087), .ZN(n7727) );
  INV_X1 U8570 ( .A(n13055), .ZN(n13127) );
  NOR2_X2 U8571 ( .A1(n13313), .A2(n6602), .ZN(n13161) );
  NOR2_X2 U8572 ( .A1(n13217), .A2(n13330), .ZN(n13200) );
  NOR2_X1 U8573 ( .A1(n7249), .A2(n6682), .ZN(n7247) );
  INV_X1 U8574 ( .A(n7532), .ZN(n13234) );
  NAND2_X1 U8575 ( .A1(n7339), .A2(n13076), .ZN(n13230) );
  OR2_X1 U8576 ( .A1(n13245), .A2(n13074), .ZN(n7339) );
  NAND2_X1 U8577 ( .A1(n8337), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8365) );
  INV_X1 U8578 ( .A(n8338), .ZN(n8337) );
  NOR2_X1 U8579 ( .A1(n7734), .A2(n6734), .ZN(n7733) );
  NOR2_X1 U8580 ( .A1(n7739), .A2(n6616), .ZN(n7734) );
  NOR2_X2 U8581 ( .A1(n11585), .A2(n13364), .ZN(n11597) );
  NOR2_X1 U8582 ( .A1(n7241), .A2(n11303), .ZN(n7240) );
  INV_X1 U8583 ( .A(n7538), .ZN(n11193) );
  INV_X1 U8584 ( .A(n7322), .ZN(n7321) );
  OR2_X1 U8585 ( .A1(n8120), .A2(n10633), .ZN(n8141) );
  NAND2_X1 U8586 ( .A1(n10352), .A2(n10351), .ZN(n10452) );
  AOI21_X1 U8587 ( .B1(n10344), .B2(n7773), .A(n6655), .ZN(n7772) );
  INV_X1 U8588 ( .A(n10301), .ZN(n7773) );
  XNOR2_X1 U8589 ( .A(n10564), .B(n10455), .ZN(n10446) );
  AOI21_X1 U8590 ( .B1(n10435), .B2(n7718), .A(n7717), .ZN(n7716) );
  INV_X1 U8591 ( .A(n10122), .ZN(n7717) );
  INV_X1 U8592 ( .A(n10121), .ZN(n7718) );
  AOI22_X1 U8593 ( .A1(n8561), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n8334), .B2(
        n9531), .ZN(n7968) );
  NAND2_X1 U8594 ( .A1(n6572), .A2(n6762), .ZN(n10254) );
  NOR2_X1 U8595 ( .A1(n9711), .A2(n9696), .ZN(n9701) );
  NAND2_X1 U8596 ( .A1(n13128), .A2(n13127), .ZN(n13299) );
  NAND2_X1 U8597 ( .A1(n7723), .A2(n13082), .ZN(n13186) );
  NAND2_X1 U8598 ( .A1(n13266), .A2(n7805), .ZN(n13254) );
  NAND2_X1 U8599 ( .A1(n8336), .A2(n8335), .ZN(n13353) );
  NAND2_X1 U8600 ( .A1(n11579), .A2(n11578), .ZN(n11591) );
  NAND2_X1 U8601 ( .A1(n9945), .A2(n9707), .ZN(n15376) );
  XNOR2_X1 U8602 ( .A(n8692), .B(P2_IR_REG_28__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U8603 ( .A1(n8678), .A2(n8677), .ZN(n8681) );
  INV_X1 U8604 ( .A(n8690), .ZN(n9475) );
  NOR2_X1 U8605 ( .A1(n7588), .A2(n7587), .ZN(n7586) );
  INV_X1 U8606 ( .A(n7937), .ZN(n7587) );
  OR2_X1 U8607 ( .A1(n8116), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8156) );
  AND2_X1 U8608 ( .A1(n8062), .A2(n8085), .ZN(n9634) );
  OR2_X1 U8609 ( .A1(n8032), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8055) );
  NOR2_X1 U8610 ( .A1(n13768), .A2(n7508), .ZN(n7507) );
  INV_X1 U8611 ( .A(n13731), .ZN(n7508) );
  INV_X1 U8612 ( .A(n7505), .ZN(n7504) );
  OAI21_X1 U8613 ( .B1(n13768), .B2(n7506), .A(n7510), .ZN(n7505) );
  OR2_X1 U8614 ( .A1(n13597), .A2(n13596), .ZN(n7491) );
  INV_X1 U8615 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n12184) );
  OR2_X1 U8616 ( .A1(n11530), .A2(n11529), .ZN(n11625) );
  NAND2_X1 U8617 ( .A1(n7028), .A2(n7030), .ZN(n11479) );
  NAND2_X1 U8618 ( .A1(n7496), .A2(n7509), .ZN(n7495) );
  INV_X1 U8619 ( .A(n7501), .ZN(n7496) );
  OR2_X1 U8620 ( .A1(n13529), .A2(n13667), .ZN(n13546) );
  NAND2_X1 U8621 ( .A1(n10028), .A2(n10027), .ZN(n10074) );
  AND3_X1 U8622 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n10415) );
  INV_X1 U8623 ( .A(n10726), .ZN(n7474) );
  AND2_X1 U8624 ( .A1(n7490), .A2(n7491), .ZN(n7488) );
  NOR2_X1 U8625 ( .A1(n6597), .A2(n13658), .ZN(n7035) );
  INV_X1 U8626 ( .A(n7484), .ZN(n7040) );
  NAND2_X1 U8627 ( .A1(n7515), .A2(n7513), .ZN(n7512) );
  INV_X1 U8628 ( .A(n7521), .ZN(n7513) );
  INV_X1 U8629 ( .A(n13692), .ZN(n13553) );
  INV_X1 U8630 ( .A(n13842), .ZN(n13831) );
  INV_X1 U8631 ( .A(n10037), .ZN(n13688) );
  OAI22_X1 U8632 ( .A1(n13692), .A2(n7471), .B1(n13842), .B2(n14435), .ZN(
        n7470) );
  NAND2_X1 U8633 ( .A1(n13840), .A2(n13839), .ZN(n14162) );
  OR2_X1 U8634 ( .A1(n13837), .A2(n13836), .ZN(n13840) );
  NAND2_X1 U8635 ( .A1(n14201), .A2(n6959), .ZN(n6958) );
  OR2_X1 U8636 ( .A1(n6960), .A2(n6958), .ZN(n6955) );
  NAND2_X1 U8637 ( .A1(n14200), .A2(n6962), .ZN(n6957) );
  AND2_X1 U8638 ( .A1(n6960), .A2(n6962), .ZN(n6956) );
  NOR2_X1 U8639 ( .A1(n14236), .A2(n14452), .ZN(n14218) );
  INV_X1 U8640 ( .A(n7351), .ZN(n14230) );
  NAND2_X1 U8641 ( .A1(n6882), .A2(n6884), .ZN(n14232) );
  INV_X1 U8642 ( .A(n14234), .ZN(n6897) );
  NOR2_X1 U8643 ( .A1(n14282), .A2(n14472), .ZN(n14261) );
  NAND2_X1 U8644 ( .A1(n14261), .A2(n14465), .ZN(n14250) );
  NAND2_X1 U8645 ( .A1(n7601), .A2(n7600), .ZN(n14282) );
  NAND2_X1 U8646 ( .A1(n6850), .A2(n14323), .ZN(n6848) );
  AND2_X1 U8647 ( .A1(n7703), .A2(n7701), .ZN(n14277) );
  INV_X1 U8648 ( .A(n7601), .ZN(n14297) );
  NAND2_X1 U8649 ( .A1(n14299), .A2(n7705), .ZN(n7704) );
  INV_X1 U8650 ( .A(n14292), .ZN(n7705) );
  AND2_X1 U8651 ( .A1(n6978), .A2(n6586), .ZN(n14317) );
  NAND2_X1 U8652 ( .A1(n14324), .A2(n14334), .ZN(n6978) );
  NAND2_X1 U8653 ( .A1(n14317), .A2(n6947), .ZN(n14291) );
  NAND2_X1 U8654 ( .A1(n7602), .A2(n13806), .ZN(n14311) );
  NAND2_X1 U8655 ( .A1(n14340), .A2(n14174), .ZN(n14324) );
  NAND2_X1 U8656 ( .A1(n14393), .A2(n7267), .ZN(n14344) );
  NOR2_X1 U8657 ( .A1(n7272), .A2(n7268), .ZN(n7267) );
  INV_X1 U8658 ( .A(n7269), .ZN(n7268) );
  NAND2_X1 U8659 ( .A1(n14393), .A2(n7271), .ZN(n14373) );
  AND2_X1 U8660 ( .A1(n13511), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13527) );
  NAND2_X1 U8661 ( .A1(n14393), .A2(n14397), .ZN(n14394) );
  NAND2_X1 U8662 ( .A1(n6874), .A2(n6873), .ZN(n14169) );
  NAND2_X1 U8663 ( .A1(n6701), .A2(n13942), .ZN(n6873) );
  NAND2_X1 U8664 ( .A1(n6878), .A2(n6875), .ZN(n6874) );
  NAND2_X1 U8665 ( .A1(n7599), .A2(n7598), .ZN(n11634) );
  INV_X1 U8666 ( .A(n7599), .ZN(n11518) );
  NAND2_X1 U8667 ( .A1(n7264), .A2(n7263), .ZN(n11251) );
  NOR2_X1 U8668 ( .A1(n13924), .A2(n15201), .ZN(n7263) );
  OR2_X1 U8669 ( .A1(n10897), .A2(n10896), .ZN(n11040) );
  OR2_X1 U8670 ( .A1(n11040), .A2(n12362), .ZN(n11153) );
  NAND2_X1 U8671 ( .A1(n6700), .A2(n6856), .ZN(n6853) );
  AND2_X1 U8672 ( .A1(n6855), .A2(n11140), .ZN(n6854) );
  NOR2_X1 U8673 ( .A1(n15075), .A2(n15084), .ZN(n15079) );
  NAND2_X1 U8674 ( .A1(n15079), .A2(n15177), .ZN(n11026) );
  INV_X1 U8675 ( .A(n6936), .ZN(n6937) );
  NAND2_X1 U8676 ( .A1(n10424), .A2(n15095), .ZN(n15075) );
  AND3_X1 U8677 ( .A1(n13892), .A2(n15156), .A3(n7260), .ZN(n10424) );
  AND4_X1 U8678 ( .A1(n10043), .A2(n10042), .A3(n10041), .A4(n10040), .ZN(
        n13876) );
  OR2_X1 U8679 ( .A1(n10037), .A2(n9754), .ZN(n10043) );
  NAND2_X1 U8680 ( .A1(n10768), .A2(n10767), .ZN(n14206) );
  AND2_X1 U8681 ( .A1(n13868), .A2(n13871), .ZN(n10948) );
  NAND2_X1 U8682 ( .A1(n15156), .A2(n14425), .ZN(n10949) );
  NAND2_X1 U8683 ( .A1(n14419), .A2(n10224), .ZN(n10954) );
  AND3_X1 U8684 ( .A1(n10024), .A2(n10023), .A3(n10022), .ZN(n14423) );
  OR2_X1 U8685 ( .A1(n14444), .A2(n15147), .ZN(n7596) );
  INV_X1 U8686 ( .A(n14448), .ZN(n7594) );
  NAND2_X1 U8687 ( .A1(n14228), .A2(n7828), .ZN(n14220) );
  NAND2_X1 U8688 ( .A1(n14386), .A2(n7700), .ZN(n14367) );
  NAND2_X1 U8689 ( .A1(n10769), .A2(n10776), .ZN(n15200) );
  INV_X1 U8690 ( .A(n15200), .ZN(n15191) );
  NAND2_X1 U8691 ( .A1(n9617), .A2(n9616), .ZN(n9979) );
  INV_X1 U8692 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9989) );
  NAND2_X1 U8693 ( .A1(n9665), .A2(n9987), .ZN(n7848) );
  OAI21_X1 U8694 ( .B1(n8509), .B2(n8508), .A(n8507), .ZN(n8530) );
  NOR2_X1 U8695 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7562) );
  XNOR2_X1 U8696 ( .A(n9662), .B(P1_IR_REG_21__SCAN_IN), .ZN(n15139) );
  XNOR2_X1 U8697 ( .A(n8399), .B(n8398), .ZN(n13450) );
  NAND2_X1 U8698 ( .A1(n8357), .A2(n8356), .ZN(n8379) );
  NAND2_X1 U8699 ( .A1(n7357), .A2(n7358), .ZN(n8331) );
  OR2_X1 U8700 ( .A1(n8244), .A2(n7610), .ZN(n7357) );
  NAND2_X1 U8701 ( .A1(n7608), .A2(n8288), .ZN(n8308) );
  NAND2_X1 U8702 ( .A1(n8283), .A2(n6710), .ZN(n7608) );
  OR2_X1 U8703 ( .A1(n10332), .A2(n10335), .ZN(n10513) );
  INV_X1 U8704 ( .A(n8262), .ZN(n8259) );
  NAND2_X1 U8705 ( .A1(n7618), .A2(n8175), .ZN(n8200) );
  NAND2_X1 U8706 ( .A1(n8174), .A2(n8173), .ZN(n7618) );
  NAND2_X1 U8707 ( .A1(n6996), .A2(n7206), .ZN(n8134) );
  OAI211_X1 U8708 ( .C1(n8077), .C2(n6995), .A(n6994), .B(n7208), .ZN(n6996)
         );
  AOI21_X1 U8709 ( .B1(n7208), .B2(n7210), .A(n7207), .ZN(n7206) );
  INV_X1 U8710 ( .A(n8078), .ZN(n6995) );
  INV_X1 U8711 ( .A(n8108), .ZN(n7210) );
  INV_X1 U8712 ( .A(n8080), .ZN(n8081) );
  NAND2_X1 U8713 ( .A1(n6993), .A2(n8078), .ZN(n8082) );
  NAND2_X1 U8714 ( .A1(n8082), .A2(n8081), .ZN(n8109) );
  NOR2_X1 U8715 ( .A1(n6992), .A2(n9962), .ZN(n7946) );
  NAND2_X1 U8716 ( .A1(n7460), .A2(n7459), .ZN(n14715) );
  NAND2_X1 U8717 ( .A1(n14668), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7459) );
  NOR2_X1 U8718 ( .A1(n15619), .A2(n14737), .ZN(n14740) );
  INV_X1 U8719 ( .A(n7461), .ZN(n14736) );
  AOI21_X1 U8720 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14687), .A(n14686), .ZN(
        n14706) );
  OAI21_X1 U8721 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14691), .A(n14690), .ZN(
        n14704) );
  OAI21_X1 U8722 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14696), .A(n14695), .ZN(
        n14700) );
  OR2_X1 U8723 ( .A1(n14981), .A2(n6914), .ZN(n6912) );
  AND2_X1 U8724 ( .A1(n14981), .A2(n6914), .ZN(n6913) );
  INV_X1 U8725 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6914) );
  OAI21_X1 U8726 ( .B1(n6827), .B2(n6824), .A(n6823), .ZN(n11287) );
  AOI21_X1 U8727 ( .B1(n6822), .B2(n6821), .A(n6652), .ZN(n6823) );
  NAND2_X1 U8728 ( .A1(n7664), .A2(n7662), .ZN(n11731) );
  INV_X1 U8729 ( .A(n7663), .ZN(n7662) );
  NAND2_X1 U8730 ( .A1(n7666), .A2(n7665), .ZN(n7664) );
  NAND2_X1 U8731 ( .A1(n9131), .A2(n9130), .ZN(n11742) );
  NAND2_X1 U8732 ( .A1(n11559), .A2(n8913), .ZN(n11605) );
  NAND2_X1 U8733 ( .A1(n11559), .A2(n6576), .ZN(n11606) );
  AND2_X1 U8734 ( .A1(n7674), .A2(n7675), .ZN(n10782) );
  INV_X1 U8735 ( .A(n7673), .ZN(n7672) );
  NAND2_X1 U8736 ( .A1(n9207), .A2(n9206), .ZN(n11713) );
  NAND2_X1 U8737 ( .A1(n10473), .A2(n7090), .ZN(n10474) );
  NAND2_X1 U8738 ( .A1(n10958), .A2(n6829), .ZN(n11098) );
  NAND2_X1 U8739 ( .A1(n7681), .A2(n7682), .ZN(n11792) );
  NAND2_X1 U8740 ( .A1(n11784), .A2(n11782), .ZN(n7682) );
  NAND2_X1 U8741 ( .A1(n7678), .A2(n12557), .ZN(n7681) );
  OR2_X1 U8742 ( .A1(n11784), .A2(n11782), .ZN(n7678) );
  AOI21_X1 U8743 ( .B1(n11745), .B2(n11746), .A(n6837), .ZN(n11808) );
  INV_X1 U8744 ( .A(n6839), .ZN(n6838) );
  NAND2_X1 U8745 ( .A1(n6843), .A2(n6840), .ZN(n11825) );
  AND4_X1 U8746 ( .A1(n8951), .A2(n8950), .A3(n8949), .A4(n8948), .ZN(n11832)
         );
  NAND2_X1 U8747 ( .A1(n10475), .A2(n8811), .ZN(n10594) );
  XNOR2_X1 U8748 ( .A(n8813), .B(n12106), .ZN(n10595) );
  OR2_X1 U8749 ( .A1(n6826), .A2(n11097), .ZN(n6825) );
  INV_X1 U8750 ( .A(n6828), .ZN(n6826) );
  NAND2_X1 U8751 ( .A1(n11202), .A2(n11204), .ZN(n11203) );
  AND4_X1 U8752 ( .A1(n9039), .A2(n9038), .A3(n9037), .A4(n9036), .ZN(n12588)
         );
  AOI21_X1 U8753 ( .B1(n7660), .B2(n7659), .A(n7658), .ZN(n7657) );
  INV_X1 U8754 ( .A(n11865), .ZN(n7658) );
  NAND2_X1 U8755 ( .A1(n7656), .A2(n7660), .ZN(n11866) );
  NAND2_X1 U8756 ( .A1(n7666), .A2(n7661), .ZN(n7656) );
  NOR2_X1 U8757 ( .A1(n12071), .A2(n7406), .ZN(n11928) );
  INV_X1 U8758 ( .A(n12509), .ZN(n12534) );
  INV_X1 U8759 ( .A(n9274), .ZN(n12558) );
  INV_X1 U8760 ( .A(n11820), .ZN(n12616) );
  INV_X1 U8761 ( .A(n11832), .ZN(n12632) );
  INV_X1 U8762 ( .A(n11836), .ZN(n12099) );
  INV_X1 U8763 ( .A(n11564), .ZN(n12101) );
  INV_X1 U8764 ( .A(n11288), .ZN(n12103) );
  AND2_X1 U8765 ( .A1(n6806), .A2(n6805), .ZN(n15413) );
  INV_X1 U8766 ( .A(n10191), .ZN(n6806) );
  NAND2_X1 U8767 ( .A1(n10263), .A2(n10192), .ZN(n6805) );
  NAND2_X1 U8768 ( .A1(n6583), .A2(n7365), .ZN(n15425) );
  AND2_X1 U8769 ( .A1(n15406), .A2(n10374), .ZN(n15427) );
  XNOR2_X1 U8770 ( .A(n10379), .B(n10378), .ZN(n15444) );
  NOR2_X1 U8771 ( .A1(n15444), .A2(n15445), .ZN(n15443) );
  OAI22_X1 U8772 ( .A1(n15456), .A2(n10367), .B1(n6972), .B2(n10378), .ZN(
        n10369) );
  INV_X1 U8773 ( .A(n6973), .ZN(n6972) );
  INV_X1 U8774 ( .A(n7045), .ZN(n7044) );
  NAND2_X1 U8775 ( .A1(n6803), .A2(n6802), .ZN(n15524) );
  INV_X1 U8776 ( .A(n15522), .ZN(n6802) );
  INV_X1 U8777 ( .A(n15523), .ZN(n6803) );
  NOR2_X1 U8778 ( .A1(n14582), .A2(n15495), .ZN(n15513) );
  INV_X1 U8779 ( .A(n7363), .ZN(n14581) );
  NOR2_X1 U8780 ( .A1(n15513), .A2(n15512), .ZN(n15511) );
  NOR2_X1 U8781 ( .A1(n15530), .A2(n15531), .ZN(n15529) );
  XNOR2_X1 U8782 ( .A(n7041), .B(n15537), .ZN(n15530) );
  NOR2_X1 U8783 ( .A1(n15529), .A2(n14585), .ZN(n15550) );
  NOR2_X1 U8784 ( .A1(n15550), .A2(n15549), .ZN(n15548) );
  OR2_X1 U8785 ( .A1(n15566), .A2(n15565), .ZN(n15567) );
  INV_X1 U8786 ( .A(n6815), .ZN(n14830) );
  NOR2_X1 U8787 ( .A1(n14821), .A2(n14822), .ZN(n14820) );
  XNOR2_X1 U8788 ( .A(n14587), .B(n14827), .ZN(n14821) );
  INV_X1 U8789 ( .A(n14626), .ZN(n14853) );
  MUX2_X1 U8790 ( .A(n10178), .B(n12107), .S(n12083), .Z(n15555) );
  XNOR2_X1 U8791 ( .A(n14593), .B(n14628), .ZN(n14858) );
  AND2_X1 U8792 ( .A1(n14837), .A2(n14592), .ZN(n14593) );
  NAND2_X1 U8793 ( .A1(n12426), .A2(n7867), .ZN(n12415) );
  NAND2_X1 U8794 ( .A1(n12451), .A2(n6617), .ZN(n12441) );
  NAND2_X1 U8795 ( .A1(n9150), .A2(n9149), .ZN(n12478) );
  AND2_X1 U8796 ( .A1(n7075), .A2(n7077), .ZN(n12484) );
  NAND2_X1 U8797 ( .A1(n7858), .A2(n7855), .ZN(n12493) );
  NAND2_X1 U8798 ( .A1(n9275), .A2(n7450), .ZN(n7446) );
  NAND2_X1 U8799 ( .A1(n9111), .A2(n9110), .ZN(n12516) );
  NAND2_X1 U8800 ( .A1(n9275), .A2(n12024), .ZN(n12523) );
  NAND2_X1 U8801 ( .A1(n9339), .A2(n9338), .ZN(n12545) );
  OAI21_X1 U8802 ( .B1(n9273), .B2(n7438), .A(n7435), .ZN(n12592) );
  NAND2_X1 U8803 ( .A1(n7441), .A2(n11916), .ZN(n12612) );
  NAND2_X1 U8804 ( .A1(n9273), .A2(n7442), .ZN(n7441) );
  NAND2_X1 U8805 ( .A1(n11119), .A2(n11959), .ZN(n11279) );
  NAND2_X1 U8806 ( .A1(n10823), .A2(n11951), .ZN(n11105) );
  AND2_X1 U8807 ( .A1(n10160), .A2(n9236), .ZN(n12624) );
  NAND2_X1 U8808 ( .A1(n11357), .A2(n10584), .ZN(n12627) );
  INV_X1 U8809 ( .A(n12624), .ZN(n12639) );
  INV_X1 U8810 ( .A(n12478), .ZN(n12735) );
  INV_X1 U8811 ( .A(n11829), .ZN(n12743) );
  NAND2_X1 U8812 ( .A1(n9002), .A2(n9001), .ZN(n12769) );
  INV_X1 U8813 ( .A(n9311), .ZN(n10934) );
  AND2_X1 U8814 ( .A1(n10161), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12772) );
  OAI21_X1 U8815 ( .B1(n11884), .B2(n11883), .A(n11882), .ZN(n11886) );
  MUX2_X1 U8816 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8761), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8763) );
  NAND2_X1 U8817 ( .A1(n8757), .A2(n7202), .ZN(n7201) );
  NAND2_X1 U8818 ( .A1(n7403), .A2(n9289), .ZN(n11723) );
  XNOR2_X1 U8819 ( .A(n9190), .B(n9178), .ZN(n11399) );
  NAND2_X1 U8820 ( .A1(n8737), .A2(n8723), .ZN(n11402) );
  OAI21_X1 U8821 ( .B1(n9159), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n9160), .ZN(
        n9176) );
  NAND2_X1 U8822 ( .A1(n8720), .A2(n6604), .ZN(n11297) );
  XNOR2_X1 U8823 ( .A(n8713), .B(n8712), .ZN(n8726) );
  INV_X1 U8824 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8712) );
  INV_X1 U8825 ( .A(n8711), .ZN(n8713) );
  XNOR2_X1 U8826 ( .A(n9224), .B(n9223), .ZN(n14790) );
  NAND2_X1 U8827 ( .A1(n9222), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9224) );
  NAND2_X1 U8828 ( .A1(n7103), .A2(n9116), .ZN(n9128) );
  NAND2_X1 U8829 ( .A1(n9115), .A2(n9114), .ZN(n7103) );
  AOI21_X1 U8830 ( .B1(n8709), .B2(n8715), .A(n6847), .ZN(n6846) );
  INV_X1 U8831 ( .A(n9222), .ZN(n6847) );
  INV_X1 U8832 ( .A(n9353), .ZN(n10403) );
  INV_X1 U8833 ( .A(SI_19_), .ZN(n10139) );
  NAND2_X1 U8834 ( .A1(n7107), .A2(n7111), .ZN(n9088) );
  NAND2_X1 U8835 ( .A1(n9058), .A2(n7114), .ZN(n7107) );
  NAND2_X1 U8836 ( .A1(n7116), .A2(n9059), .ZN(n9074) );
  NAND2_X1 U8837 ( .A1(n7118), .A2(n7117), .ZN(n7116) );
  INV_X1 U8838 ( .A(SI_13_), .ZN(n9614) );
  NAND2_X1 U8839 ( .A1(n7395), .A2(n7393), .ZN(n8977) );
  NAND2_X1 U8840 ( .A1(n7395), .A2(n8955), .ZN(n8958) );
  INV_X1 U8841 ( .A(SI_12_), .ZN(n9474) );
  INV_X1 U8842 ( .A(SI_11_), .ZN(n9460) );
  INV_X1 U8843 ( .A(n15485), .ZN(n14644) );
  NAND2_X1 U8844 ( .A1(n7389), .A2(n8850), .ZN(n8872) );
  NAND2_X1 U8845 ( .A1(n8848), .A2(n8847), .ZN(n7389) );
  AND2_X1 U8846 ( .A1(n8753), .A2(n8832), .ZN(n10375) );
  AND3_X1 U8847 ( .A1(n8774), .A2(n7379), .A3(n7378), .ZN(n10371) );
  NAND2_X1 U8848 ( .A1(n8709), .A2(n8700), .ZN(n7378) );
  INV_X1 U8849 ( .A(n8773), .ZN(n7380) );
  XNOR2_X1 U8850 ( .A(n7382), .B(n8794), .ZN(n10279) );
  INV_X1 U8851 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7382) );
  NAND2_X1 U8852 ( .A1(n10293), .A2(n10292), .ZN(n10616) );
  NAND2_X1 U8853 ( .A1(n12969), .A2(n12834), .ZN(n12840) );
  NAND2_X1 U8854 ( .A1(n8159), .A2(n8158), .ZN(n11003) );
  NAND2_X1 U8855 ( .A1(n10616), .A2(n10615), .ZN(n10642) );
  NAND2_X1 U8856 ( .A1(n6930), .A2(n7315), .ZN(n12875) );
  INV_X1 U8857 ( .A(n12823), .ZN(n6922) );
  NAND2_X1 U8858 ( .A1(n10094), .A2(n10100), .ZN(n10284) );
  NAND2_X1 U8859 ( .A1(n12818), .A2(n12817), .ZN(n12920) );
  INV_X1 U8860 ( .A(n10129), .ZN(n10260) );
  NOR2_X1 U8861 ( .A1(n11221), .A2(n7298), .ZN(n7294) );
  NAND2_X1 U8862 ( .A1(n7296), .A2(n6600), .ZN(n11222) );
  NAND2_X1 U8863 ( .A1(n12951), .A2(n12950), .ZN(n12949) );
  NAND2_X1 U8864 ( .A1(n10284), .A2(n10283), .ZN(n10326) );
  NAND2_X1 U8865 ( .A1(n11551), .A2(n11550), .ZN(n12789) );
  XNOR2_X1 U8866 ( .A(n12785), .B(n12786), .ZN(n11551) );
  NAND2_X1 U8867 ( .A1(n6603), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7954) );
  NAND2_X1 U8868 ( .A1(n8160), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U8869 ( .A1(n6603), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7133) );
  OR2_X1 U8870 ( .A1(n7997), .A2(n7908), .ZN(n7132) );
  NAND2_X1 U8871 ( .A1(n13030), .A2(n13294), .ZN(n13283) );
  AND2_X1 U8872 ( .A1(n8584), .A2(n8583), .ZN(n13063) );
  NAND2_X1 U8873 ( .A1(n8534), .A2(n8533), .ZN(n13301) );
  INV_X1 U8874 ( .A(n13307), .ZN(n13146) );
  INV_X1 U8875 ( .A(n7728), .ZN(n13137) );
  INV_X1 U8876 ( .A(n7732), .ZN(n13155) );
  NAND2_X1 U8877 ( .A1(n7236), .A2(n7238), .ZN(n13152) );
  NAND2_X1 U8878 ( .A1(n7237), .A2(n7792), .ZN(n7236) );
  AND2_X1 U8879 ( .A1(n7796), .A2(n7794), .ZN(n13173) );
  NAND2_X1 U8880 ( .A1(n7796), .A2(n7799), .ZN(n13174) );
  NAND2_X1 U8881 ( .A1(n13207), .A2(n7797), .ZN(n7796) );
  NAND2_X1 U8882 ( .A1(n7347), .A2(n7344), .ZN(n13170) );
  NAND2_X1 U8883 ( .A1(n13207), .A2(n7800), .ZN(n13183) );
  AND2_X1 U8884 ( .A1(n7248), .A2(n7252), .ZN(n13227) );
  NAND2_X1 U8885 ( .A1(n7736), .A2(n7737), .ZN(n13067) );
  NAND2_X1 U8886 ( .A1(n11579), .A2(n7739), .ZN(n7736) );
  INV_X1 U8887 ( .A(n7230), .ZN(n11596) );
  AND2_X1 U8888 ( .A1(n11571), .A2(n7808), .ZN(n11594) );
  NAND2_X1 U8889 ( .A1(n11571), .A2(n11570), .ZN(n11573) );
  NAND2_X1 U8890 ( .A1(n7328), .A2(n11301), .ZN(n11498) );
  NAND2_X1 U8891 ( .A1(n6739), .A2(n7330), .ZN(n7328) );
  NAND2_X1 U8892 ( .A1(n7242), .A2(n7244), .ZN(n11304) );
  NAND2_X1 U8893 ( .A1(n7330), .A2(n11191), .ZN(n11299) );
  NAND2_X1 U8894 ( .A1(n7243), .A2(n11067), .ZN(n11197) );
  OR2_X1 U8895 ( .A1(n11065), .A2(n11064), .ZN(n7243) );
  INV_X1 U8896 ( .A(n10532), .ZN(n10534) );
  NAND2_X1 U8897 ( .A1(n7324), .A2(n10528), .ZN(n10743) );
  NAND2_X1 U8898 ( .A1(n10526), .A2(n10525), .ZN(n7324) );
  NAND2_X1 U8899 ( .A1(n7775), .A2(n10301), .ZN(n10345) );
  NAND2_X1 U8900 ( .A1(n10117), .A2(n10116), .ZN(n10303) );
  NAND2_X1 U8901 ( .A1(n10434), .A2(n10435), .ZN(n10433) );
  NAND2_X1 U8902 ( .A1(n10202), .A2(n10121), .ZN(n10434) );
  INV_X1 U8903 ( .A(n13277), .ZN(n13240) );
  NAND2_X1 U8904 ( .A1(n15327), .A2(n9701), .ZN(n13236) );
  OR2_X1 U8905 ( .A1(n13335), .A2(n13334), .ZN(n13386) );
  AND2_X1 U8906 ( .A1(n7902), .A2(n7905), .ZN(n7170) );
  NAND2_X1 U8907 ( .A1(n8683), .A2(n8686), .ZN(n13411) );
  INV_X1 U8908 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13413) );
  NAND2_X1 U8909 ( .A1(n7925), .A2(n7915), .ZN(n8687) );
  INV_X1 U8910 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13416) );
  XNOR2_X1 U8911 ( .A(n8682), .B(P2_IR_REG_24__SCAN_IN), .ZN(n13414) );
  NAND2_X1 U8912 ( .A1(n8681), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8682) );
  INV_X1 U8913 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10947) );
  MUX2_X1 U8914 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7927), .S(
        P2_IR_REG_19__SCAN_IN), .Z(n7928) );
  NAND2_X1 U8915 ( .A1(n7929), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7927) );
  INV_X1 U8916 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10466) );
  INV_X1 U8917 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10331) );
  INV_X1 U8918 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10572) );
  INV_X1 U8919 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n12254) );
  INV_X1 U8920 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9927) );
  AND2_X1 U8921 ( .A1(n8086), .A2(n8116), .ZN(n15232) );
  INV_X1 U8922 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9549) );
  NOR2_X1 U8923 ( .A1(n8510), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13397) );
  INV_X1 U8924 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9467) );
  INV_X1 U8925 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9447) );
  CLKBUF_X1 U8926 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n15229) );
  NAND2_X1 U8927 ( .A1(n11088), .A2(n11087), .ZN(n11266) );
  NAND2_X1 U8928 ( .A1(n7477), .A2(n7475), .ZN(n13675) );
  INV_X1 U8929 ( .A(n7476), .ZN(n7475) );
  NOR2_X1 U8930 ( .A1(n7483), .A2(n7479), .ZN(n7478) );
  NAND2_X1 U8931 ( .A1(n13422), .A2(n13421), .ZN(n14460) );
  AOI21_X1 U8932 ( .B1(n13481), .B2(n13480), .A(n13479), .ZN(n13646) );
  NAND2_X1 U8933 ( .A1(n11478), .A2(n11479), .ZN(n11646) );
  NAND2_X1 U8934 ( .A1(n11266), .A2(n11265), .ZN(n11268) );
  AND2_X1 U8935 ( .A1(n13650), .A2(n15059), .ZN(n13776) );
  AND2_X1 U8936 ( .A1(n13650), .A2(n15049), .ZN(n13777) );
  NAND2_X1 U8937 ( .A1(n10030), .A2(n13682), .ZN(n10031) );
  NAND2_X1 U8938 ( .A1(n10034), .A2(n10033), .ZN(n10075) );
  AND2_X1 U8939 ( .A1(n7032), .A2(n6624), .ZN(n13704) );
  OAI21_X1 U8940 ( .B1(n13741), .B2(n13742), .A(n7491), .ZN(n13713) );
  NAND2_X1 U8941 ( .A1(n13720), .A2(n13506), .ZN(n13733) );
  XNOR2_X1 U8942 ( .A(n10729), .B(n10674), .ZN(n10727) );
  NAND2_X1 U8943 ( .A1(n7497), .A2(n7495), .ZN(n13753) );
  NAND2_X1 U8944 ( .A1(n7494), .A2(n11650), .ZN(n11652) );
  NAND2_X1 U8945 ( .A1(n11646), .A2(n11645), .ZN(n7494) );
  NAND2_X1 U8946 ( .A1(n10076), .A2(n10077), .ZN(n7017) );
  NOR2_X1 U8947 ( .A1(n10248), .A2(n10013), .ZN(n13650) );
  AOI21_X1 U8948 ( .B1(n13733), .B2(n13731), .A(n13730), .ZN(n13767) );
  NAND2_X1 U8949 ( .A1(n7019), .A2(n7018), .ZN(n10920) );
  INV_X1 U8950 ( .A(n7020), .ZN(n7019) );
  NAND2_X1 U8951 ( .A1(n10727), .A2(n6654), .ZN(n7018) );
  OAI21_X1 U8952 ( .B1(n10730), .B2(n7473), .A(n10913), .ZN(n7020) );
  NAND2_X1 U8953 ( .A1(n10920), .A2(n10919), .ZN(n11081) );
  OR2_X1 U8954 ( .A1(n13788), .A2(n13787), .ZN(n13792) );
  INV_X1 U8955 ( .A(n13784), .ZN(n13790) );
  NOR2_X1 U8956 ( .A1(n14034), .A2(n14044), .ZN(n7552) );
  AOI21_X1 U8957 ( .B1(n14216), .B2(n15196), .A(n7195), .ZN(n14457) );
  NAND2_X1 U8958 ( .A1(n7197), .A2(n7196), .ZN(n7195) );
  NAND2_X1 U8959 ( .A1(n14215), .A2(n15059), .ZN(n7197) );
  NAND2_X1 U8960 ( .A1(n6953), .A2(n7830), .ZN(n14249) );
  NAND2_X1 U8961 ( .A1(n14485), .A2(n7831), .ZN(n6953) );
  NAND2_X1 U8962 ( .A1(n6887), .A2(n6891), .ZN(n14245) );
  NAND2_X1 U8963 ( .A1(n6883), .A2(n6888), .ZN(n14244) );
  NAND2_X1 U8964 ( .A1(n7835), .A2(n7836), .ZN(n14259) );
  NAND2_X1 U8965 ( .A1(n14485), .A2(n7837), .ZN(n7835) );
  NAND2_X1 U8966 ( .A1(n14485), .A2(n14198), .ZN(n14274) );
  NAND2_X1 U8967 ( .A1(n13567), .A2(n13566), .ZN(n14304) );
  NAND2_X1 U8968 ( .A1(n14331), .A2(n14197), .ZN(n14310) );
  NAND2_X1 U8969 ( .A1(n14338), .A2(n14196), .ZN(n14333) );
  NAND2_X1 U8970 ( .A1(n7687), .A2(n7688), .ZN(n14342) );
  OR2_X1 U8971 ( .A1(n14386), .A2(n6629), .ZN(n7687) );
  NAND2_X1 U8972 ( .A1(n7691), .A2(n7695), .ZN(n14357) );
  NAND2_X1 U8973 ( .A1(n14386), .A2(n7697), .ZN(n7691) );
  NAND2_X1 U8974 ( .A1(n14187), .A2(n14186), .ZN(n14385) );
  NAND2_X1 U8975 ( .A1(n14184), .A2(n14183), .ZN(n14403) );
  NAND2_X1 U8976 ( .A1(n11523), .A2(n11522), .ZN(n14934) );
  INV_X1 U8977 ( .A(n13951), .ZN(n11522) );
  AND2_X1 U8978 ( .A1(n6877), .A2(n6633), .ZN(n11624) );
  NAND2_X1 U8979 ( .A1(n6877), .A2(n6879), .ZN(n11513) );
  NAND2_X1 U8980 ( .A1(n11420), .A2(n13820), .ZN(n6940) );
  NAND2_X1 U8981 ( .A1(n15057), .A2(n11147), .ZN(n11235) );
  NAND2_X1 U8982 ( .A1(n15052), .A2(n11162), .ZN(n11231) );
  INV_X1 U8983 ( .A(n15087), .ZN(n15063) );
  NAND2_X1 U8984 ( .A1(n6858), .A2(n6859), .ZN(n11139) );
  OAI21_X1 U8985 ( .B1(n11023), .B2(n6619), .A(n10894), .ZN(n11039) );
  NAND2_X1 U8986 ( .A1(n6862), .A2(n6872), .ZN(n15071) );
  NAND2_X1 U8987 ( .A1(n6869), .A2(n6867), .ZN(n6862) );
  NAND2_X1 U8988 ( .A1(n6869), .A2(n10413), .ZN(n10891) );
  NAND2_X1 U8989 ( .A1(n10763), .A2(n10227), .ZN(n7820) );
  NAND2_X1 U8990 ( .A1(n7715), .A2(n13888), .ZN(n10412) );
  INV_X1 U8991 ( .A(n7589), .ZN(n7257) );
  NAND2_X1 U8992 ( .A1(n11615), .A2(n10071), .ZN(n7256) );
  OAI21_X1 U8993 ( .B1(n13850), .B2(n7591), .A(n7590), .ZN(n7589) );
  AND2_X2 U8994 ( .A1(n10211), .A2(n10768), .ZN(n15224) );
  NAND2_X1 U8995 ( .A1(n14557), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9988) );
  XNOR2_X1 U8996 ( .A(n7525), .B(n9989), .ZN(n11698) );
  OAI21_X1 U8997 ( .B1(n9664), .B2(n7848), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7525) );
  NAND2_X1 U8998 ( .A1(n6792), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U8999 ( .A1(n9664), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6793) );
  XNOR2_X1 U9000 ( .A(n9661), .B(P1_IR_REG_22__SCAN_IN), .ZN(n13861) );
  NAND2_X1 U9001 ( .A1(n9660), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9661) );
  XNOR2_X1 U9002 ( .A(n9980), .B(n7563), .ZN(n11298) );
  INV_X1 U9003 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10944) );
  NAND2_X1 U9004 ( .A1(n9983), .A2(n9409), .ZN(n14265) );
  INV_X1 U9005 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n12269) );
  INV_X1 U9006 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n12347) );
  INV_X1 U9007 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10340) );
  INV_X1 U9008 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10342) );
  INV_X1 U9009 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9933) );
  INV_X1 U9010 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9809) );
  INV_X1 U9011 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9553) );
  INV_X1 U9012 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9547) );
  NAND2_X1 U9013 ( .A1(n6920), .A2(n8026), .ZN(n8030) );
  NAND2_X1 U9014 ( .A1(n8025), .A2(n8024), .ZN(n6920) );
  INV_X1 U9015 ( .A(P2_RD_REG_SCAN_IN), .ZN(n14767) );
  INV_X1 U9016 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14718) );
  NOR2_X1 U9017 ( .A1(n15626), .A2(n14721), .ZN(n14770) );
  AOI21_X1 U9018 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14722), .A(n15622), .ZN(
        n15614) );
  NAND2_X1 U9019 ( .A1(n6900), .A2(n6902), .ZN(n15617) );
  NAND2_X1 U9020 ( .A1(n6905), .A2(n6901), .ZN(n6900) );
  NAND2_X1 U9021 ( .A1(n6903), .A2(n14727), .ZN(n6902) );
  NOR2_X1 U9022 ( .A1(n14727), .A2(n14724), .ZN(n6901) );
  XNOR2_X1 U9023 ( .A(n7461), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15620) );
  NOR2_X1 U9024 ( .A1(n15620), .A2(n15621), .ZN(n15619) );
  XNOR2_X1 U9025 ( .A(n14740), .B(n7458), .ZN(n14778) );
  INV_X1 U9026 ( .A(n14741), .ZN(n7458) );
  AND2_X1 U9027 ( .A1(n7456), .A2(n7457), .ZN(n14966) );
  NAND2_X1 U9028 ( .A1(n14969), .A2(n14752), .ZN(n14973) );
  INV_X1 U9029 ( .A(n7454), .ZN(n14751) );
  NAND2_X1 U9030 ( .A1(n14973), .A2(n14974), .ZN(n14972) );
  NAND2_X1 U9031 ( .A1(n6899), .A2(n14972), .ZN(n14978) );
  OAI21_X1 U9032 ( .B1(n14973), .B2(n14974), .A(n7186), .ZN(n6899) );
  INV_X1 U9033 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7186) );
  NOR2_X1 U9034 ( .A1(n14759), .A2(n14758), .ZN(n14806) );
  OAI21_X1 U9035 ( .B1(n11775), .B2(n11776), .A(n11863), .ZN(n11781) );
  INV_X1 U9036 ( .A(n7173), .ZN(n7172) );
  OAI21_X1 U9037 ( .B1(n12727), .B2(n11875), .A(n11861), .ZN(n7173) );
  AOI21_X1 U9038 ( .B1(n6813), .B2(n15543), .A(n6812), .ZN(n14665) );
  NOR2_X1 U9039 ( .A1(n7200), .A2(n7199), .ZN(n7198) );
  NOR2_X1 U9040 ( .A1(n15599), .A2(n12722), .ZN(n7199) );
  NOR2_X1 U9041 ( .A1(n12723), .A2(n12770), .ZN(n7200) );
  NAND2_X1 U9042 ( .A1(n7580), .A2(n7578), .ZN(P2_U3192) );
  OAI21_X1 U9043 ( .B1(n13111), .B2(n12967), .A(n12872), .ZN(n7579) );
  NAND2_X1 U9044 ( .A1(n7297), .A2(n7300), .ZN(n11216) );
  NAND2_X1 U9045 ( .A1(n7570), .A2(n7573), .ZN(n12915) );
  NAND2_X1 U9046 ( .A1(n7314), .A2(n7568), .ZN(n12935) );
  NAND2_X1 U9047 ( .A1(n12951), .A2(n7317), .ZN(n7314) );
  OR2_X1 U9048 ( .A1(n15392), .A2(n7529), .ZN(n7528) );
  NAND2_X1 U9049 ( .A1(n7254), .A2(n15392), .ZN(n7530) );
  INV_X1 U9050 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7529) );
  OAI211_X1 U9051 ( .C1(n7787), .C2(n15381), .A(n7785), .B(n7786), .ZN(
        P2_U3496) );
  NOR2_X1 U9052 ( .A1(n7781), .A2(n6760), .ZN(n7780) );
  OAI21_X1 U9053 ( .B1(n13837), .B2(n13399), .A(n7748), .ZN(P2_U3297) );
  INV_X1 U9054 ( .A(n7749), .ZN(n7748) );
  INV_X1 U9055 ( .A(n9618), .ZN(n9418) );
  XNOR2_X1 U9056 ( .A(n7039), .B(n7038), .ZN(n13785) );
  INV_X1 U9057 ( .A(n7595), .ZN(n14449) );
  AOI211_X1 U9058 ( .C1(n7713), .C2(n15065), .A(n14211), .B(n14210), .ZN(
        n14212) );
  OR2_X1 U9059 ( .A1(n15224), .A2(n7710), .ZN(n7709) );
  NAND2_X1 U9060 ( .A1(n14539), .A2(n15224), .ZN(n7711) );
  INV_X1 U9061 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7710) );
  NAND2_X1 U9062 ( .A1(n14539), .A2(n15209), .ZN(n7262) );
  NAND2_X1 U9063 ( .A1(n6893), .A2(n6745), .ZN(P1_U3523) );
  NAND2_X1 U9064 ( .A1(n14541), .A2(n15209), .ZN(n6893) );
  INV_X1 U9065 ( .A(n7185), .ZN(n14773) );
  XNOR2_X1 U9066 ( .A(n14819), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n7463) );
  XNOR2_X1 U9067 ( .A(n14818), .B(n14817), .ZN(n14819) );
  INV_X1 U9068 ( .A(n8635), .ZN(n8592) );
  AND2_X1 U9069 ( .A1(n8931), .A2(n8913), .ZN(n6576) );
  AND2_X1 U9070 ( .A1(n6967), .A2(n7841), .ZN(n6577) );
  AND2_X1 U9071 ( .A1(n7592), .A2(n7265), .ZN(n6578) );
  INV_X1 U9072 ( .A(n7309), .ZN(n15362) );
  NAND2_X2 U9073 ( .A1(n7906), .A2(n7907), .ZN(n7997) );
  AND2_X1 U9074 ( .A1(n7315), .A2(n6929), .ZN(n6579) );
  INV_X1 U9075 ( .A(n8645), .ZN(n10130) );
  AND2_X1 U9076 ( .A1(n8150), .A2(n8149), .ZN(n6580) );
  INV_X1 U9077 ( .A(n13895), .ZN(n7821) );
  NAND2_X1 U9078 ( .A1(n7497), .A2(n6664), .ZN(n7032) );
  NAND2_X1 U9079 ( .A1(n11425), .A2(n11424), .ZN(n13934) );
  INV_X1 U9080 ( .A(n10344), .ZN(n7774) );
  AND2_X1 U9081 ( .A1(n7426), .A2(n9313), .ZN(n6581) );
  NAND2_X1 U9082 ( .A1(n11144), .A2(n11143), .ZN(n15201) );
  OAI21_X1 U9083 ( .B1(n14340), .B2(n14323), .A(n6850), .ZN(n7703) );
  OR2_X1 U9084 ( .A1(n8628), .A2(n8627), .ZN(n6582) );
  INV_X1 U9085 ( .A(n8416), .ZN(n7175) );
  AOI21_X1 U9086 ( .B1(n11753), .B2(n11752), .A(n9113), .ZN(n9120) );
  INV_X1 U9087 ( .A(n7610), .ZN(n7609) );
  NOR2_X1 U9088 ( .A1(n7819), .A2(n10406), .ZN(n7818) );
  INV_X1 U9089 ( .A(n12417), .ZN(n7869) );
  OR2_X1 U9090 ( .A1(n10374), .A2(n15426), .ZN(n6583) );
  NAND2_X1 U9091 ( .A1(n8919), .A2(n6638), .ZN(n6584) );
  XNOR2_X1 U9092 ( .A(n9988), .B(n14554), .ZN(n9990) );
  INV_X1 U9093 ( .A(n13977), .ZN(n6790) );
  AND2_X1 U9094 ( .A1(n11790), .A2(n12548), .ZN(n6585) );
  OR2_X1 U9095 ( .A1(n14496), .A2(n14175), .ZN(n6586) );
  INV_X1 U9096 ( .A(n10615), .ZN(n7307) );
  OR2_X1 U9097 ( .A1(n7573), .A2(n6729), .ZN(n6587) );
  INV_X1 U9098 ( .A(n8991), .ZN(n7665) );
  AND2_X1 U9099 ( .A1(n6699), .A2(n7145), .ZN(n6588) );
  INV_X1 U9100 ( .A(n10327), .ZN(n7582) );
  AND2_X1 U9101 ( .A1(n7619), .A2(n8636), .ZN(n6589) );
  AND2_X1 U9102 ( .A1(n7312), .A2(n10291), .ZN(n6590) );
  AND2_X1 U9103 ( .A1(n7830), .A2(n6952), .ZN(n6591) );
  NAND2_X1 U9104 ( .A1(n12524), .A2(n12534), .ZN(n6592) );
  NAND2_X1 U9105 ( .A1(n6717), .A2(n7214), .ZN(n6593) );
  INV_X1 U9106 ( .A(n8458), .ZN(n7282) );
  OR2_X1 U9107 ( .A1(n7029), .A2(n11457), .ZN(n6594) );
  AND3_X1 U9108 ( .A1(n7279), .A2(n7762), .A3(n6709), .ZN(n6595) );
  OR2_X1 U9109 ( .A1(n13934), .A2(n13935), .ZN(n6596) );
  INV_X1 U9110 ( .A(n10555), .ZN(n10547) );
  AND2_X1 U9111 ( .A1(n13581), .A2(n13580), .ZN(n6597) );
  NAND2_X1 U9112 ( .A1(n7367), .A2(n14642), .ZN(n7047) );
  OR2_X1 U9113 ( .A1(n8422), .A2(SI_21_), .ZN(n6598) );
  INV_X1 U9114 ( .A(n12384), .ZN(n7049) );
  OR2_X1 U9115 ( .A1(n12384), .A2(n14642), .ZN(n6599) );
  INV_X1 U9116 ( .A(n7266), .ZN(n7264) );
  NAND2_X1 U9117 ( .A1(n11037), .A2(n11036), .ZN(n13917) );
  INV_X1 U9118 ( .A(n13917), .ZN(n7265) );
  AND2_X1 U9119 ( .A1(n7295), .A2(n11215), .ZN(n6600) );
  AND2_X1 U9120 ( .A1(n7264), .A2(n11163), .ZN(n6601) );
  NAND2_X1 U9121 ( .A1(n11905), .A2(n9383), .ZN(n12636) );
  INV_X1 U9122 ( .A(n12636), .ZN(n12584) );
  OR2_X1 U9123 ( .A1(n13189), .A2(n13318), .ZN(n6602) );
  NAND2_X1 U9124 ( .A1(n9286), .A2(n9285), .ZN(n12652) );
  AND2_X1 U9125 ( .A1(n10218), .A2(n10217), .ZN(n13892) );
  NAND2_X1 U9126 ( .A1(n7309), .A2(n9712), .ZN(n11315) );
  OR2_X1 U9127 ( .A1(n9061), .A2(n7872), .ZN(n6604) );
  OR2_X1 U9128 ( .A1(n7286), .A2(n8506), .ZN(n6605) );
  OR3_X1 U9129 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n10184), .ZN(n6606) );
  INV_X1 U9130 ( .A(n13092), .ZN(n13093) );
  NAND4_X1 U9131 ( .A1(n9996), .A2(n9997), .A3(n9998), .A4(n9995), .ZN(n10212)
         );
  OR2_X1 U9132 ( .A1(n13913), .A2(n11260), .ZN(n6607) );
  INV_X1 U9133 ( .A(n8592), .ZN(n8616) );
  XNOR2_X1 U9134 ( .A(n14358), .B(n14345), .ZN(n14356) );
  AND2_X1 U9135 ( .A1(n9408), .A2(n9398), .ZN(n6608) );
  NAND2_X1 U9136 ( .A1(n13374), .A2(n11300), .ZN(n6609) );
  INV_X1 U9137 ( .A(n14183), .ZN(n6969) );
  NOR2_X1 U9138 ( .A1(n7798), .A2(n7793), .ZN(n7792) );
  NOR2_X1 U9139 ( .A1(n11520), .A2(n13820), .ZN(n6610) );
  AND2_X1 U9140 ( .A1(n7569), .A2(n12930), .ZN(n7568) );
  OR2_X1 U9141 ( .A1(n12524), .A2(n12509), .ZN(n12029) );
  AND2_X1 U9142 ( .A1(n10505), .A2(n10504), .ZN(n6611) );
  NAND2_X1 U9143 ( .A1(n14228), .A2(n6960), .ZN(n6612) );
  AND2_X1 U9144 ( .A1(n9340), .A2(n9338), .ZN(n6613) );
  AND2_X1 U9145 ( .A1(n13823), .A2(n11620), .ZN(n6614) );
  AND2_X1 U9146 ( .A1(n8356), .A2(n7635), .ZN(n6615) );
  OR2_X1 U9147 ( .A1(n7735), .A2(n13066), .ZN(n6616) );
  OR2_X1 U9148 ( .A1(n12731), .A2(n12473), .ZN(n6617) );
  AND2_X1 U9149 ( .A1(n8789), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n6618) );
  OR3_X1 U9150 ( .A1(n14570), .A2(n14574), .A3(n14567), .ZN(n9986) );
  NAND2_X1 U9151 ( .A1(n7863), .A2(n8773), .ZN(n8750) );
  AND2_X1 U9152 ( .A1(n13906), .A2(n11085), .ZN(n6619) );
  INV_X1 U9153 ( .A(n13885), .ZN(n10227) );
  XNOR2_X1 U9154 ( .A(n10500), .B(n15163), .ZN(n13885) );
  AND2_X1 U9155 ( .A1(n6789), .A2(n6788), .ZN(n6620) );
  OR2_X1 U9156 ( .A1(n13844), .A2(n10014), .ZN(n6621) );
  INV_X1 U9157 ( .A(n12519), .ZN(n7860) );
  AND4_X1 U9158 ( .A1(n7811), .A2(n7812), .A3(n7813), .A4(n9469), .ZN(n6622)
         );
  INV_X1 U9159 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14670) );
  NAND2_X1 U9160 ( .A1(n14028), .A2(n14027), .ZN(n6623) );
  INV_X1 U9161 ( .A(n12458), .ZN(n7080) );
  NAND2_X1 U9162 ( .A1(n6933), .A2(n6800), .ZN(n10777) );
  INV_X1 U9163 ( .A(n10777), .ZN(n15163) );
  NAND2_X1 U9164 ( .A1(n13556), .A2(n13555), .ZN(n6624) );
  NAND2_X1 U9165 ( .A1(n10332), .A2(n6608), .ZN(n9409) );
  AND2_X1 U9166 ( .A1(n14472), .A2(n14278), .ZN(n6625) );
  NAND2_X1 U9167 ( .A1(n13489), .A2(n13488), .ZN(n6626) );
  AND3_X1 U9168 ( .A1(n9410), .A2(n9408), .A3(n9407), .ZN(n6627) );
  INV_X1 U9169 ( .A(n13348), .ZN(n7533) );
  AND2_X1 U9170 ( .A1(n12802), .A2(n12801), .ZN(n6628) );
  INV_X1 U9171 ( .A(n13979), .ZN(n6788) );
  OR2_X1 U9172 ( .A1(n7694), .A2(n7690), .ZN(n6629) );
  OR2_X1 U9173 ( .A1(n11909), .A2(n7066), .ZN(n6630) );
  AND2_X1 U9174 ( .A1(n7230), .A2(n7229), .ZN(n6631) );
  NAND2_X1 U9175 ( .A1(n7412), .A2(n8792), .ZN(n8806) );
  AND2_X1 U9176 ( .A1(n14254), .A2(n14262), .ZN(n6632) );
  AND2_X1 U9177 ( .A1(n6879), .A2(n6596), .ZN(n6633) );
  NAND3_X1 U9178 ( .A1(n7469), .A2(n6621), .A3(n10016), .ZN(n14066) );
  INV_X1 U9179 ( .A(n14066), .ZN(n14428) );
  AND2_X1 U9180 ( .A1(n7549), .A2(n13981), .ZN(n6634) );
  AND2_X1 U9181 ( .A1(n7446), .A2(n12029), .ZN(n6635) );
  NAND2_X1 U9182 ( .A1(n8247), .A2(n8246), .ZN(n11505) );
  INV_X1 U9183 ( .A(n11505), .ZN(n7536) );
  NAND4_X1 U9184 ( .A1(n10084), .A2(n10083), .A3(n10082), .A4(n10081), .ZN(
        n14065) );
  NAND2_X1 U9185 ( .A1(n8402), .A2(n8401), .ZN(n13337) );
  INV_X1 U9186 ( .A(n13337), .ZN(n7531) );
  XNOR2_X1 U9187 ( .A(n7926), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8618) );
  AND2_X1 U9188 ( .A1(n11842), .A2(n12558), .ZN(n6636) );
  NAND2_X1 U9189 ( .A1(n11151), .A2(n11150), .ZN(n13924) );
  INV_X1 U9190 ( .A(n14201), .ZN(n6962) );
  OR2_X1 U9191 ( .A1(n8728), .A2(n8709), .ZN(n6637) );
  NOR2_X1 U9192 ( .A1(n9061), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8731) );
  OAI21_X1 U9193 ( .B1(n9173), .B2(n7654), .A(n7651), .ZN(n11854) );
  AND2_X1 U9194 ( .A1(n8920), .A2(n7684), .ZN(n6638) );
  OR2_X1 U9195 ( .A1(n11842), .A2(n12558), .ZN(n6639) );
  NAND2_X1 U9196 ( .A1(n13453), .A2(n13452), .ZN(n14496) );
  NAND4_X2 U9197 ( .A1(n7956), .A2(n7955), .A3(n7954), .A4(n7953), .ZN(n12994)
         );
  AND2_X1 U9198 ( .A1(n13705), .A2(n6624), .ZN(n6640) );
  AND2_X1 U9199 ( .A1(n7669), .A2(n12495), .ZN(n6641) );
  AND2_X1 U9200 ( .A1(n7300), .A2(n10975), .ZN(n6642) );
  NAND3_X1 U9201 ( .A1(n10332), .A2(n6608), .A3(n7563), .ZN(n6643) );
  AOI21_X1 U9202 ( .B1(n13657), .B2(n13658), .A(n6597), .ZN(n13741) );
  AND2_X1 U9203 ( .A1(n12329), .A2(n7924), .ZN(n6644) );
  OR2_X1 U9204 ( .A1(n14452), .A2(n14181), .ZN(n6645) );
  INV_X1 U9205 ( .A(n13904), .ZN(n7561) );
  AND3_X1 U9206 ( .A1(n13953), .A2(n13943), .A3(n13947), .ZN(n6646) );
  INV_X1 U9207 ( .A(n13821), .ZN(n11520) );
  AND3_X1 U9208 ( .A1(n13954), .A2(n13955), .A3(n13956), .ZN(n6647) );
  INV_X1 U9209 ( .A(n6892), .ZN(n6891) );
  AND2_X1 U9210 ( .A1(n14575), .A2(n10020), .ZN(n14314) );
  NAND2_X1 U9211 ( .A1(n8826), .A2(n9268), .ZN(n6648) );
  NOR2_X1 U9212 ( .A1(n11729), .A2(n12586), .ZN(n6649) );
  AND2_X1 U9213 ( .A1(n13289), .A2(n15366), .ZN(n6650) );
  OR2_X1 U9214 ( .A1(n9061), .A2(n7874), .ZN(n6651) );
  AND2_X1 U9215 ( .A1(n13544), .A2(n13543), .ZN(n14502) );
  INV_X1 U9216 ( .A(n14502), .ZN(n7272) );
  AND2_X1 U9217 ( .A1(n8860), .A2(n12103), .ZN(n6652) );
  NAND2_X1 U9218 ( .A1(n13510), .A2(n13509), .ZN(n14522) );
  AND2_X1 U9219 ( .A1(n13337), .A2(n13078), .ZN(n6653) );
  NOR2_X1 U9220 ( .A1(n7473), .A2(n7474), .ZN(n6654) );
  AND2_X1 U9221 ( .A1(n15365), .A2(n12988), .ZN(n6655) );
  INV_X1 U9222 ( .A(n13914), .ZN(n7566) );
  OR2_X1 U9223 ( .A1(n11497), .A2(n7327), .ZN(n6656) );
  NOR2_X1 U9224 ( .A1(n6810), .A2(n10279), .ZN(n10185) );
  INV_X1 U9225 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n6818) );
  INV_X1 U9226 ( .A(n7258), .ZN(n14236) );
  NOR2_X1 U9227 ( .A1(n14250), .A2(n14460), .ZN(n7258) );
  AND2_X1 U9228 ( .A1(n9310), .A2(n9307), .ZN(n6657) );
  AND2_X1 U9229 ( .A1(n7347), .A2(n7719), .ZN(n6658) );
  OR2_X1 U9230 ( .A1(n14730), .A2(n7462), .ZN(n6659) );
  INV_X1 U9231 ( .A(n7424), .ZN(n7423) );
  OAI21_X1 U9232 ( .B1(n12057), .B2(n9278), .A(n12055), .ZN(n7424) );
  OR2_X1 U9233 ( .A1(n13090), .A2(n13056), .ZN(n6660) );
  INV_X1 U9234 ( .A(n7722), .ZN(n7721) );
  NAND2_X1 U9235 ( .A1(n13184), .A2(n7724), .ZN(n7722) );
  AND2_X1 U9236 ( .A1(n7503), .A2(n7501), .ZN(n6661) );
  AND2_X1 U9237 ( .A1(n8708), .A2(n7875), .ZN(n6662) );
  INV_X1 U9238 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6908) );
  INV_X1 U9239 ( .A(n7062), .ZN(n14594) );
  OAI21_X1 U9240 ( .B1(n14820), .B2(n7056), .A(n7057), .ZN(n7062) );
  AND2_X1 U9241 ( .A1(n6884), .A2(n6881), .ZN(n6663) );
  AND2_X1 U9242 ( .A1(n7495), .A2(n7031), .ZN(n6664) );
  AND2_X1 U9243 ( .A1(n6829), .A2(n6828), .ZN(n6665) );
  INV_X1 U9244 ( .A(n7841), .ZN(n7840) );
  NOR2_X1 U9245 ( .A1(n14191), .A2(n7842), .ZN(n7841) );
  OR2_X1 U9246 ( .A1(n8219), .A2(n8218), .ZN(n6666) );
  AND2_X1 U9247 ( .A1(n6808), .A2(n15411), .ZN(n6667) );
  INV_X1 U9248 ( .A(n12600), .ZN(n12611) );
  AND2_X1 U9249 ( .A1(n12001), .A2(n12002), .ZN(n12600) );
  INV_X1 U9250 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8700) );
  AND2_X1 U9251 ( .A1(n7846), .A2(n9989), .ZN(n6668) );
  AND2_X1 U9252 ( .A1(n12024), .A2(n12025), .ZN(n12531) );
  AND2_X1 U9253 ( .A1(n7835), .A2(n7833), .ZN(n6669) );
  INV_X1 U9254 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7202) );
  AND2_X1 U9255 ( .A1(n6953), .A2(n6591), .ZN(n6670) );
  NOR2_X1 U9256 ( .A1(n14314), .A2(n14326), .ZN(n6671) );
  INV_X1 U9257 ( .A(n7880), .ZN(n7667) );
  AND2_X1 U9258 ( .A1(n12652), .A2(n12093), .ZN(n6672) );
  NAND2_X1 U9259 ( .A1(n7284), .A2(n8527), .ZN(n7283) );
  NAND2_X1 U9260 ( .A1(n8763), .A2(n8762), .ZN(n12781) );
  INV_X1 U9261 ( .A(n12781), .ZN(n7008) );
  NOR2_X1 U9262 ( .A1(n11782), .A2(n12557), .ZN(n6673) );
  AND3_X1 U9263 ( .A1(n8069), .A2(n8070), .A3(n7255), .ZN(n6674) );
  AND3_X1 U9264 ( .A1(n8017), .A2(n8018), .A3(n8019), .ZN(n6675) );
  INV_X1 U9265 ( .A(n7422), .ZN(n7421) );
  NOR2_X1 U9266 ( .A1(n7424), .A2(n12064), .ZN(n7422) );
  INV_X1 U9267 ( .A(n12988), .ZN(n10350) );
  NAND2_X1 U9268 ( .A1(n6674), .A2(n8071), .ZN(n12988) );
  INV_X1 U9269 ( .A(n7331), .ZN(n10435) );
  NAND2_X1 U9270 ( .A1(n10122), .A2(n7332), .ZN(n7331) );
  AND2_X1 U9271 ( .A1(n7703), .A2(n7704), .ZN(n6676) );
  NOR2_X1 U9272 ( .A1(n8600), .A2(n8599), .ZN(n6677) );
  OR2_X1 U9273 ( .A1(n10637), .A2(n7307), .ZN(n6678) );
  INV_X1 U9274 ( .A(n14200), .ZN(n6959) );
  NAND2_X1 U9275 ( .A1(n10332), .A2(n9408), .ZN(n6679) );
  AND2_X1 U9276 ( .A1(n12727), .A2(n12456), .ZN(n6680) );
  INV_X1 U9277 ( .A(n7801), .ZN(n7800) );
  NOR2_X1 U9278 ( .A1(n13050), .A2(n13081), .ZN(n7801) );
  OR2_X1 U9279 ( .A1(n6990), .A2(n6991), .ZN(n6681) );
  INV_X1 U9280 ( .A(n14309), .ZN(n6947) );
  NOR2_X1 U9281 ( .A1(n13045), .A2(n13044), .ZN(n6682) );
  AND2_X1 U9282 ( .A1(n8222), .A2(n9474), .ZN(n6683) );
  AND2_X1 U9283 ( .A1(n8310), .A2(n8309), .ZN(n6684) );
  AND2_X1 U9284 ( .A1(n13910), .A2(n7559), .ZN(n6685) );
  AND2_X1 U9285 ( .A1(n7221), .A2(n7222), .ZN(n6686) );
  AND2_X1 U9286 ( .A1(n12805), .A2(n12804), .ZN(n6687) );
  AND2_X1 U9287 ( .A1(n8256), .A2(n8255), .ZN(n6688) );
  INV_X1 U9288 ( .A(n7345), .ZN(n7344) );
  NAND2_X1 U9289 ( .A1(n7719), .A2(n7346), .ZN(n7345) );
  NOR2_X1 U9290 ( .A1(n14927), .A2(n11196), .ZN(n6689) );
  NAND2_X1 U9291 ( .A1(n8992), .A2(n7119), .ZN(n6690) );
  AND2_X1 U9292 ( .A1(n8330), .A2(SI_17_), .ZN(n6691) );
  AND2_X1 U9293 ( .A1(n8198), .A2(n9460), .ZN(n6692) );
  AND2_X1 U9294 ( .A1(n9547), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U9295 ( .A1(n12936), .A2(n12811), .ZN(n6694) );
  INV_X1 U9296 ( .A(n7083), .ZN(n7082) );
  NAND2_X1 U9297 ( .A1(n6617), .A2(n7084), .ZN(n7083) );
  INV_X1 U9298 ( .A(n6833), .ZN(n6832) );
  NAND2_X1 U9299 ( .A1(n7676), .A2(n6639), .ZN(n6833) );
  OR2_X1 U9300 ( .A1(n6649), .A2(n7663), .ZN(n6695) );
  OAI21_X1 U9301 ( .B1(n7840), .B2(n7844), .A(n14190), .ZN(n7839) );
  OR2_X1 U9302 ( .A1(n11902), .A2(n12407), .ZN(n7409) );
  AND2_X1 U9303 ( .A1(n7701), .A2(n14276), .ZN(n6696) );
  INV_X1 U9304 ( .A(n7873), .ZN(n7872) );
  NOR2_X1 U9305 ( .A1(n7874), .A2(P3_IR_REG_25__SCAN_IN), .ZN(n7873) );
  NOR2_X1 U9306 ( .A1(n13054), .A2(n13086), .ZN(n6697) );
  AND2_X1 U9307 ( .A1(n7295), .A2(n7294), .ZN(n6698) );
  AND2_X1 U9308 ( .A1(n7278), .A2(n8482), .ZN(n6699) );
  AND2_X1 U9309 ( .A1(n13817), .A2(n6607), .ZN(n6700) );
  INV_X1 U9310 ( .A(n13980), .ZN(n7549) );
  INV_X1 U9311 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U9312 ( .A1(n7177), .A2(n7176), .ZN(n7747) );
  INV_X1 U9313 ( .A(n7747), .ZN(n7744) );
  INV_X1 U9314 ( .A(n6889), .ZN(n6888) );
  NAND2_X1 U9315 ( .A1(n6890), .A2(n14248), .ZN(n6889) );
  INV_X1 U9316 ( .A(n7565), .ZN(n7564) );
  NAND2_X1 U9317 ( .A1(n7566), .A2(n13915), .ZN(n7565) );
  INV_X1 U9318 ( .A(n13992), .ZN(n7215) );
  NAND2_X1 U9319 ( .A1(n6633), .A2(n13933), .ZN(n6701) );
  OR2_X1 U9320 ( .A1(n11195), .A2(n12982), .ZN(n6702) );
  OR2_X1 U9321 ( .A1(n11790), .A2(n12548), .ZN(n6703) );
  OR2_X1 U9322 ( .A1(n13313), .A2(n13053), .ZN(n6704) );
  INV_X1 U9323 ( .A(n10381), .ZN(n7053) );
  OR2_X1 U9324 ( .A1(n8330), .A2(SI_17_), .ZN(n6705) );
  AND3_X1 U9325 ( .A1(n6794), .A2(n7211), .A3(n7213), .ZN(n6706) );
  AND2_X1 U9326 ( .A1(n11955), .A2(n11956), .ZN(n7430) );
  INV_X1 U9327 ( .A(n7430), .ZN(n7426) );
  NOR2_X1 U9328 ( .A1(n7825), .A2(n11145), .ZN(n6707) );
  AND2_X1 U9329 ( .A1(n12063), .A2(n12061), .ZN(n12417) );
  NOR2_X1 U9330 ( .A1(n14980), .A2(n14981), .ZN(n6708) );
  OR2_X1 U9331 ( .A1(n7175), .A2(n8418), .ZN(n6709) );
  AND2_X1 U9332 ( .A1(n8282), .A2(n8286), .ZN(n6710) );
  AND2_X1 U9333 ( .A1(n14299), .A2(n6947), .ZN(n6711) );
  AND2_X1 U9334 ( .A1(n7685), .A2(n8710), .ZN(n6712) );
  AND2_X1 U9335 ( .A1(n8455), .A2(n8454), .ZN(n6713) );
  OR2_X1 U9336 ( .A1(n14006), .A2(n14004), .ZN(n6714) );
  AND2_X1 U9337 ( .A1(n7368), .A2(n7367), .ZN(n6715) );
  AND2_X1 U9338 ( .A1(n7329), .A2(n6609), .ZN(n6716) );
  NAND2_X1 U9339 ( .A1(n13994), .A2(n7551), .ZN(n6717) );
  AND2_X1 U9340 ( .A1(n7373), .A2(n7062), .ZN(n6718) );
  NAND2_X1 U9341 ( .A1(n6695), .A2(n7667), .ZN(n7660) );
  AND2_X1 U9342 ( .A1(n7040), .A2(n7034), .ZN(n6719) );
  AND2_X1 U9343 ( .A1(n7216), .A2(n7550), .ZN(n6720) );
  AND2_X1 U9344 ( .A1(n14309), .A2(n7829), .ZN(n6721) );
  OR2_X1 U9345 ( .A1(n13325), .A2(n13083), .ZN(n6722) );
  OR2_X1 U9346 ( .A1(n7009), .A2(n10186), .ZN(n6723) );
  INV_X1 U9347 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7905) );
  INV_X1 U9348 ( .A(n7448), .ZN(n7447) );
  OAI21_X1 U9349 ( .B1(n7450), .B2(n7449), .A(n12034), .ZN(n7448) );
  AND2_X1 U9350 ( .A1(n6955), .A2(n6957), .ZN(n6724) );
  INV_X1 U9351 ( .A(n7868), .ZN(n7867) );
  NAND2_X1 U9352 ( .A1(n7869), .A2(n9350), .ZN(n7868) );
  OR2_X1 U9353 ( .A1(n10745), .A2(n10744), .ZN(n6725) );
  NAND2_X1 U9354 ( .A1(n8773), .A2(n8700), .ZN(n8774) );
  INV_X1 U9355 ( .A(n6924), .ZN(n6923) );
  NAND2_X1 U9356 ( .A1(n12817), .A2(n6925), .ZN(n6924) );
  NAND2_X1 U9357 ( .A1(n15433), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6726) );
  INV_X1 U9358 ( .A(n13817), .ZN(n6857) );
  INV_X1 U9359 ( .A(n15467), .ZN(n14642) );
  OAI211_X1 U9360 ( .C1(n8962), .C2(n9126), .A(n9125), .B(n9124), .ZN(n12507)
         );
  AND2_X1 U9361 ( .A1(n12949), .A2(n12800), .ZN(n6727) );
  AND2_X1 U9362 ( .A1(n14393), .A2(n7269), .ZN(n6728) );
  INV_X1 U9363 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8715) );
  INV_X1 U9364 ( .A(n13494), .ZN(n7516) );
  AND2_X1 U9365 ( .A1(n12794), .A2(n12793), .ZN(n6729) );
  INV_X1 U9366 ( .A(n11916), .ZN(n7440) );
  INV_X1 U9367 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7606) );
  XOR2_X1 U9368 ( .A(n12870), .B(n12869), .Z(n6730) );
  NAND2_X1 U9369 ( .A1(n6940), .A2(n11421), .ZN(n11521) );
  NAND2_X1 U9370 ( .A1(n9273), .A2(n11993), .ZN(n12619) );
  INV_X1 U9371 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7563) );
  NAND2_X1 U9372 ( .A1(n13584), .A2(n13583), .ZN(n14284) );
  INV_X1 U9373 ( .A(n14284), .ZN(n7600) );
  OR2_X1 U9374 ( .A1(n12723), .A2(n12715), .ZN(n6731) );
  AND2_X1 U9375 ( .A1(n12100), .A2(n11977), .ZN(n6732) );
  NAND2_X1 U9376 ( .A1(n7257), .A2(n7256), .ZN(n13880) );
  INV_X1 U9377 ( .A(n13880), .ZN(n15156) );
  NAND2_X1 U9378 ( .A1(n7094), .A2(n9330), .ZN(n12599) );
  AND2_X1 U9379 ( .A1(n13292), .A2(n12961), .ZN(n6733) );
  INV_X1 U9380 ( .A(n9121), .ZN(n6841) );
  NAND2_X1 U9381 ( .A1(n8919), .A2(n8920), .ZN(n8940) );
  AND2_X1 U9382 ( .A1(n13069), .A2(n13068), .ZN(n6734) );
  AND2_X1 U9383 ( .A1(n8580), .A2(n8579), .ZN(n13058) );
  INV_X1 U9384 ( .A(n13058), .ZN(n13096) );
  INV_X1 U9385 ( .A(n7602), .ZN(n14327) );
  NOR2_X1 U9386 ( .A1(n14344), .A2(n14496), .ZN(n7602) );
  INV_X1 U9387 ( .A(n7534), .ZN(n13269) );
  INV_X1 U9388 ( .A(n11106), .ZN(n12105) );
  AND4_X1 U9389 ( .A1(n8770), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(n11106)
         );
  AND2_X1 U9390 ( .A1(n14194), .A2(n14193), .ZN(n6735) );
  INV_X1 U9391 ( .A(n7597), .ZN(n14406) );
  NOR2_X1 U9392 ( .A1(n14534), .A2(n11634), .ZN(n7597) );
  INV_X1 U9393 ( .A(n8953), .ZN(n7396) );
  AND2_X1 U9394 ( .A1(n9809), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8953) );
  AND2_X1 U9395 ( .A1(n11894), .A2(n11893), .ZN(n12407) );
  NAND3_X1 U9396 ( .A1(n7992), .A2(n8056), .A3(n7273), .ZN(n8176) );
  NOR2_X1 U9397 ( .A1(n13934), .A2(n14057), .ZN(n6736) );
  NAND2_X1 U9398 ( .A1(n14934), .A2(n6614), .ZN(n14184) );
  AND2_X1 U9399 ( .A1(n6838), .A2(n6843), .ZN(n6737) );
  INV_X1 U9400 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10048) );
  AND2_X1 U9401 ( .A1(n12632), .A2(n11414), .ZN(n6738) );
  AND2_X1 U9402 ( .A1(n8571), .A2(n8570), .ZN(n13292) );
  AND2_X1 U9403 ( .A1(n11191), .A2(n6609), .ZN(n6739) );
  AND2_X1 U9404 ( .A1(n8933), .A2(n12099), .ZN(n6740) );
  INV_X1 U9405 ( .A(n6597), .ZN(n7037) );
  OR2_X1 U9406 ( .A1(n8419), .A2(SI_20_), .ZN(n6741) );
  INV_X1 U9407 ( .A(n14189), .ZN(n7842) );
  AND2_X1 U9408 ( .A1(n7391), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n6742) );
  AND3_X1 U9409 ( .A1(n9394), .A2(n9392), .A3(n9469), .ZN(n6743) );
  NOR2_X1 U9410 ( .A1(n8957), .A2(n7394), .ZN(n7393) );
  AND2_X1 U9411 ( .A1(n7708), .A2(n7707), .ZN(n6744) );
  INV_X1 U9412 ( .A(n7252), .ZN(n7249) );
  NAND2_X1 U9413 ( .A1(n13348), .A2(n13043), .ZN(n7252) );
  INV_X1 U9414 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9223) );
  INV_X1 U9415 ( .A(n7879), .ZN(n7077) );
  INV_X1 U9416 ( .A(n7047), .ZN(n7046) );
  NAND2_X1 U9417 ( .A1(n7585), .A2(n10945), .ZN(n7309) );
  INV_X1 U9418 ( .A(n7996), .ZN(n8092) );
  INV_X1 U9419 ( .A(n13913), .ZN(n7592) );
  OR2_X1 U9420 ( .A1(n15209), .A2(n13428), .ZN(n6745) );
  NAND2_X1 U9421 ( .A1(n8294), .A2(n8293), .ZN(n13364) );
  INV_X1 U9422 ( .A(n13364), .ZN(n7738) );
  NAND2_X1 U9423 ( .A1(n7851), .A2(n9324), .ZN(n11351) );
  NAND2_X1 U9424 ( .A1(n7069), .A2(n9325), .ZN(n11406) );
  NAND2_X1 U9425 ( .A1(n8268), .A2(n8267), .ZN(n13369) );
  INV_X1 U9426 ( .A(n13369), .ZN(n7539) );
  INV_X1 U9427 ( .A(n14648), .ZN(n15519) );
  NAND2_X1 U9428 ( .A1(n11517), .A2(n11516), .ZN(n13648) );
  INV_X1 U9429 ( .A(n13648), .ZN(n7598) );
  OR2_X1 U9430 ( .A1(n15209), .A2(n13693), .ZN(n6746) );
  XOR2_X1 U9431 ( .A(n11212), .B(n11213), .Z(n6747) );
  NAND2_X1 U9432 ( .A1(n8725), .A2(n8724), .ZN(n9209) );
  NAND2_X1 U9433 ( .A1(n8718), .A2(n7685), .ZN(n6748) );
  NAND2_X1 U9434 ( .A1(n8919), .A2(n7683), .ZN(n9061) );
  NAND2_X1 U9435 ( .A1(n6827), .A2(n6825), .ZN(n11202) );
  NAND2_X1 U9436 ( .A1(n11011), .A2(n11012), .ZN(n6749) );
  AND2_X1 U9437 ( .A1(n7815), .A2(n7817), .ZN(n6750) );
  INV_X1 U9438 ( .A(n7114), .ZN(n7113) );
  NOR2_X1 U9439 ( .A1(n9073), .A2(n7115), .ZN(n7114) );
  OR2_X1 U9440 ( .A1(n14644), .A2(n15609), .ZN(n6751) );
  INV_X1 U9441 ( .A(n13730), .ZN(n7506) );
  INV_X1 U9442 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7462) );
  INV_X1 U9443 ( .A(n9057), .ZN(n7117) );
  AND2_X1 U9444 ( .A1(n12347), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9057) );
  INV_X1 U9445 ( .A(n12791), .ZN(n7575) );
  INV_X1 U9446 ( .A(n11215), .ZN(n7298) );
  AND2_X1 U9447 ( .A1(n7627), .A2(n8555), .ZN(n6752) );
  AND2_X1 U9448 ( .A1(n9129), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6753) );
  AND2_X1 U9449 ( .A1(n8464), .A2(n7624), .ZN(n6754) );
  AND2_X1 U9450 ( .A1(n7622), .A2(n8486), .ZN(n6755) );
  INV_X1 U9451 ( .A(n7583), .ZN(n7584) );
  NAND2_X1 U9452 ( .A1(n8229), .A2(n8228), .ZN(n13374) );
  INV_X1 U9453 ( .A(n13374), .ZN(n7537) );
  INV_X1 U9454 ( .A(n15196), .ZN(n15178) );
  AND2_X1 U9455 ( .A1(n7260), .A2(n15156), .ZN(n6756) );
  INV_X1 U9456 ( .A(n12968), .ZN(n12961) );
  NAND4_X1 U9457 ( .A1(n8787), .A2(n8786), .A3(n8785), .A4(n8784), .ZN(n12108)
         );
  INV_X1 U9458 ( .A(n12108), .ZN(n7415) );
  INV_X1 U9459 ( .A(n15365), .ZN(n7527) );
  OR2_X1 U9460 ( .A1(n15555), .A2(n14638), .ZN(n6757) );
  NAND2_X1 U9461 ( .A1(n10131), .A2(n10135), .ZN(n10311) );
  NOR2_X1 U9462 ( .A1(n15443), .A2(n7051), .ZN(n6758) );
  AND2_X1 U9463 ( .A1(n11946), .A2(n11945), .ZN(n9309) );
  INV_X1 U9464 ( .A(n10253), .ZN(n6762) );
  NAND2_X1 U9465 ( .A1(n7672), .A2(n7674), .ZN(n6759) );
  NAND2_X1 U9466 ( .A1(n15383), .A2(n15373), .ZN(n6760) );
  INV_X1 U9467 ( .A(n11956), .ZN(n6991) );
  INV_X1 U9468 ( .A(SI_24_), .ZN(n7624) );
  INV_X1 U9469 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7910) );
  INV_X1 U9470 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7911) );
  INV_X1 U9471 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7468) );
  NOR2_X1 U9472 ( .A1(n11694), .A2(n9670), .ZN(n6761) );
  INV_X1 U9473 ( .A(n15369), .ZN(n7308) );
  NOR2_X1 U9474 ( .A1(n10945), .A2(n9938), .ZN(n10147) );
  NAND2_X1 U9475 ( .A1(n7169), .A2(n7170), .ZN(n13395) );
  OR2_X1 U9476 ( .A1(n15614), .A2(n15613), .ZN(n6905) );
  INV_X1 U9477 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7455) );
  INV_X1 U9478 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7912) );
  INV_X1 U9479 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7591) );
  INV_X1 U9480 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7471) );
  INV_X1 U9481 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6910) );
  INV_X1 U9482 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7187) );
  INV_X1 U9483 ( .A(n15352), .ZN(n15373) );
  NOR2_X2 U9484 ( .A1(n15362), .A2(n7308), .ZN(n15352) );
  NOR2_X1 U9485 ( .A1(n14966), .A2(n14967), .ZN(n14965) );
  NAND2_X1 U9486 ( .A1(n15617), .A2(n15616), .ZN(n15615) );
  NOR2_X1 U9487 ( .A1(n14784), .A2(n14785), .ZN(n14783) );
  NOR2_X2 U9488 ( .A1(n13115), .A2(n13289), .ZN(n13059) );
  INV_X1 U9489 ( .A(n7235), .ZN(n7234) );
  INV_X1 U9490 ( .A(n8465), .ZN(n7620) );
  INV_X1 U9491 ( .A(n13147), .ZN(n7803) );
  XNOR2_X1 U9492 ( .A(n8355), .B(SI_18_), .ZN(n8353) );
  NAND2_X1 U9493 ( .A1(n14715), .A2(n14714), .ZN(n14669) );
  NAND2_X1 U9494 ( .A1(n14759), .A2(n14758), .ZN(n14808) );
  NAND2_X1 U9495 ( .A1(n10390), .A2(n10120), .ZN(n10203) );
  OAI22_X2 U9496 ( .A1(n13122), .A2(n13127), .B1(n13090), .B2(n13089), .ZN(
        n13109) );
  OAI21_X2 U9497 ( .B1(n11579), .B2(n6616), .A(n7733), .ZN(n13261) );
  NAND2_X1 U9498 ( .A1(n7530), .A2(n7528), .ZN(P2_U3528) );
  OAI211_X1 U9499 ( .C1(n10526), .C2(n7321), .A(n7320), .B(n6725), .ZN(n10747)
         );
  XNOR2_X1 U9500 ( .A(n13094), .B(n13093), .ZN(n7726) );
  AOI21_X1 U9501 ( .B1(n7726), .B2(n13264), .A(n13101), .ZN(n13290) );
  OR2_X1 U9502 ( .A1(n7151), .A2(n7175), .ZN(n7148) );
  OR2_X1 U9503 ( .A1(n8171), .A2(n8170), .ZN(n7293) );
  NAND3_X1 U9504 ( .A1(n8484), .A2(n8485), .A3(n6765), .ZN(n6764) );
  OAI22_X2 U9505 ( .A1(n8151), .A2(n7165), .B1(n8152), .B2(n6580), .ZN(n8169)
         );
  NAND2_X1 U9506 ( .A1(n7125), .A2(n7124), .ZN(n8103) );
  NOR2_X1 U9507 ( .A1(n7123), .A2(n7976), .ZN(n7980) );
  OR2_X1 U9508 ( .A1(n8008), .A2(n8004), .ZN(n7131) );
  NAND2_X1 U9509 ( .A1(n7155), .A2(n7159), .ZN(n8280) );
  NAND3_X1 U9510 ( .A1(n13989), .A2(n13990), .A3(n6720), .ZN(n6767) );
  NAND3_X1 U9511 ( .A1(n10332), .A2(n6627), .A3(n9665), .ZN(n6792) );
  NAND2_X1 U9512 ( .A1(n6795), .A2(n7553), .ZN(n6794) );
  NAND2_X1 U9513 ( .A1(n14014), .A2(n14013), .ZN(n6795) );
  NAND2_X1 U9514 ( .A1(n14012), .A2(n14011), .ZN(n14013) );
  NAND2_X1 U9515 ( .A1(n14008), .A2(n14007), .ZN(n14014) );
  NAND2_X1 U9516 ( .A1(n6796), .A2(n6799), .ZN(n13968) );
  NAND3_X1 U9517 ( .A1(n13964), .A2(n6797), .A3(n13963), .ZN(n6796) );
  NAND2_X1 U9518 ( .A1(n6807), .A2(n10263), .ZN(n6804) );
  NAND2_X1 U9519 ( .A1(n15415), .A2(n10362), .ZN(n15430) );
  INV_X2 U9520 ( .A(n10182), .ZN(n14633) );
  AOI21_X1 U9521 ( .B1(n11798), .B2(n9346), .A(n7668), .ZN(n6816) );
  NAND2_X1 U9522 ( .A1(n11738), .A2(n11798), .ZN(n6817) );
  INV_X1 U9523 ( .A(n11097), .ZN(n6822) );
  INV_X1 U9524 ( .A(n11204), .ZN(n6824) );
  AND2_X1 U9525 ( .A1(n9086), .A2(n12098), .ZN(n6837) );
  INV_X1 U9526 ( .A(n9120), .ZN(n6842) );
  NAND2_X1 U9527 ( .A1(n11561), .A2(n6576), .ZN(n6844) );
  NAND2_X1 U9528 ( .A1(n6844), .A2(n6845), .ZN(n11760) );
  NAND2_X1 U9529 ( .A1(n14340), .A2(n6850), .ZN(n6849) );
  NAND3_X1 U9530 ( .A1(n6849), .A2(n6696), .A3(n6848), .ZN(n14275) );
  NAND2_X1 U9531 ( .A1(n6854), .A2(n6853), .ZN(n15055) );
  NAND3_X1 U9532 ( .A1(n11023), .A2(n6860), .A3(n13817), .ZN(n6855) );
  INV_X1 U9533 ( .A(n13814), .ZN(n6864) );
  NAND2_X1 U9534 ( .A1(n6870), .A2(n7715), .ZN(n6869) );
  NOR2_X1 U9535 ( .A1(n14178), .A2(n14278), .ZN(n6892) );
  NAND2_X1 U9536 ( .A1(n6905), .A2(n6904), .ZN(n6903) );
  INV_X1 U9537 ( .A(n6905), .ZN(n15612) );
  NAND2_X1 U9538 ( .A1(n14769), .A2(n6906), .ZN(n15623) );
  NAND2_X1 U9539 ( .A1(n11549), .A2(n11548), .ZN(n12785) );
  NAND2_X1 U9540 ( .A1(n6915), .A2(n13107), .ZN(n7580) );
  NAND2_X1 U9541 ( .A1(n6976), .A2(n8011), .ZN(n8025) );
  NAND2_X1 U9542 ( .A1(n6976), .A2(n6918), .ZN(n6917) );
  INV_X1 U9543 ( .A(n8026), .ZN(n6919) );
  NAND2_X1 U9544 ( .A1(n6924), .A2(n12823), .ZN(n6921) );
  INV_X1 U9545 ( .A(n12921), .ZN(n6925) );
  NAND2_X1 U9546 ( .A1(n6579), .A2(n12951), .ZN(n6926) );
  NAND2_X1 U9547 ( .A1(n6936), .A2(n10850), .ZN(n6934) );
  NAND3_X1 U9548 ( .A1(n6864), .A2(n6935), .A3(n6934), .ZN(n15069) );
  NAND3_X1 U9549 ( .A1(n7816), .A2(n7818), .A3(n10850), .ZN(n6935) );
  NAND2_X1 U9550 ( .A1(n10851), .A2(n10850), .ZN(n15070) );
  NAND2_X1 U9551 ( .A1(n7815), .A2(n6937), .ZN(n10851) );
  NAND2_X1 U9552 ( .A1(n11420), .A2(n6941), .ZN(n6938) );
  NAND2_X1 U9553 ( .A1(n6938), .A2(n6939), .ZN(n11524) );
  NAND2_X1 U9554 ( .A1(n14338), .A2(n6721), .ZN(n6944) );
  NAND2_X1 U9555 ( .A1(n14485), .A2(n6949), .ZN(n6948) );
  NAND2_X1 U9556 ( .A1(n14228), .A2(n6956), .ZN(n6954) );
  OAI211_X1 U9557 ( .C1(n14228), .C2(n6958), .A(n6724), .B(n6954), .ZN(n14451)
         );
  NAND2_X1 U9558 ( .A1(n14934), .A2(n6577), .ZN(n6963) );
  MUX2_X1 U9559 ( .A(n10186), .B(P3_REG1_REG_2__SCAN_IN), .S(n10371), .Z(
        n10174) );
  NAND2_X1 U9560 ( .A1(n7205), .A2(n8010), .ZN(n6976) );
  NAND2_X1 U9561 ( .A1(n7960), .A2(n7961), .ZN(n7988) );
  NAND2_X1 U9562 ( .A1(n7711), .A2(n7709), .ZN(P1_U3557) );
  NAND2_X1 U9563 ( .A1(n8174), .A2(n6982), .ZN(n6981) );
  OAI21_X1 U9564 ( .B1(n8174), .B2(n6984), .A(n6982), .ZN(n8240) );
  NAND2_X1 U9565 ( .A1(n7429), .A2(n6985), .ZN(n6988) );
  NOR2_X1 U9566 ( .A1(n6986), .A2(n6681), .ZN(n6985) );
  INV_X1 U9567 ( .A(n7427), .ZN(n6986) );
  NAND2_X1 U9568 ( .A1(n6988), .A2(n6987), .ZN(n11278) );
  NAND3_X1 U9569 ( .A1(n7427), .A2(n7429), .A3(n11956), .ZN(n11117) );
  NAND2_X1 U9570 ( .A1(n7945), .A2(n7946), .ZN(n7958) );
  MUX2_X1 U9571 ( .A(n8742), .B(n8780), .S(n7353), .Z(n6992) );
  NAND2_X2 U9572 ( .A1(n7603), .A2(n7604), .ZN(n7353) );
  NAND2_X1 U9573 ( .A1(n8077), .A2(n8076), .ZN(n6993) );
  NAND2_X1 U9574 ( .A1(n12530), .A2(n7447), .ZN(n6998) );
  NAND2_X1 U9575 ( .A1(n6998), .A2(n6999), .ZN(n12497) );
  OAI21_X1 U9576 ( .B1(n12643), .B2(n7005), .A(n7003), .ZN(n12590) );
  NAND3_X1 U9577 ( .A1(n8779), .A2(n6723), .A3(n8778), .ZN(n7010) );
  INV_X2 U9578 ( .A(n7011), .ZN(n12457) );
  NOR2_X2 U9579 ( .A1(n12466), .A2(n12046), .ZN(n12459) );
  NAND3_X1 U9580 ( .A1(n7016), .A2(n14341), .A3(n7015), .ZN(n14340) );
  NAND2_X1 U9581 ( .A1(n7017), .A2(n10504), .ZN(n10507) );
  OAI21_X1 U9582 ( .B1(n10076), .B2(n10077), .A(n7017), .ZN(n10078) );
  NOR2_X1 U9583 ( .A1(n10025), .A2(n7022), .ZN(n10028) );
  AND2_X1 U9584 ( .A1(n10721), .A2(n14066), .ZN(n7022) );
  INV_X1 U9585 ( .A(n11458), .ZN(n7028) );
  NAND2_X1 U9586 ( .A1(n11483), .A2(n11481), .ZN(n11478) );
  OAI21_X1 U9587 ( .B1(n11458), .B2(n6594), .A(n7492), .ZN(n7024) );
  INV_X1 U9588 ( .A(n11457), .ZN(n7030) );
  INV_X1 U9589 ( .A(n7032), .ZN(n13751) );
  NAND3_X1 U9590 ( .A1(n13792), .A2(n13721), .A3(n13786), .ZN(n13720) );
  OAI21_X1 U9591 ( .B1(n13657), .B2(n7036), .A(n6719), .ZN(n7039) );
  NAND3_X1 U9592 ( .A1(n10332), .A2(n6608), .A3(n7562), .ZN(n9660) );
  NOR2_X1 U9593 ( .A1(n15479), .A2(n15478), .ZN(n15477) );
  NAND2_X1 U9594 ( .A1(n12385), .A2(n7046), .ZN(n7043) );
  OAI211_X1 U9595 ( .C1(n12385), .C2(n6599), .A(n7043), .B(n7044), .ZN(n15462)
         );
  NOR2_X1 U9596 ( .A1(n15462), .A2(n11359), .ZN(n15461) );
  OAI22_X1 U9597 ( .A1(n15444), .A2(n7050), .B1(n7052), .B2(n10381), .ZN(
        n10544) );
  INV_X1 U9598 ( .A(n7061), .ZN(n14840) );
  NAND2_X1 U9599 ( .A1(n11470), .A2(n7070), .ZN(n7067) );
  NAND2_X1 U9600 ( .A1(n7067), .A2(n7068), .ZN(n12629) );
  AND2_X1 U9601 ( .A1(n8789), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7413) );
  AND2_X2 U9602 ( .A1(n8764), .A2(n7008), .ZN(n8789) );
  NAND2_X1 U9603 ( .A1(n7858), .A2(n7076), .ZN(n7075) );
  NAND2_X1 U9604 ( .A1(n12452), .A2(n12458), .ZN(n12451) );
  NAND2_X1 U9605 ( .A1(n11936), .A2(n11935), .ZN(n7091) );
  NAND2_X1 U9606 ( .A1(n7091), .A2(n10586), .ZN(n9304) );
  INV_X1 U9607 ( .A(n7091), .ZN(n11930) );
  XNOR2_X1 U9608 ( .A(n7091), .B(n10586), .ZN(n10589) );
  XNOR2_X1 U9609 ( .A(n10585), .B(n7091), .ZN(n10602) );
  AND2_X1 U9610 ( .A1(n10585), .A2(n7091), .ZN(n7090) );
  NAND2_X1 U9611 ( .A1(n7094), .A2(n7092), .ZN(n12602) );
  NAND2_X1 U9612 ( .A1(n9327), .A2(n9326), .ZN(n12615) );
  NOR2_X1 U9613 ( .A1(n9328), .A2(n7096), .ZN(n7095) );
  INV_X1 U9614 ( .A(n9326), .ZN(n7096) );
  NAND2_X1 U9615 ( .A1(n8936), .A2(n8935), .ZN(n8938) );
  NAND2_X1 U9616 ( .A1(n8916), .A2(n8915), .ZN(n7099) );
  NAND2_X1 U9617 ( .A1(n9042), .A2(n9041), .ZN(n9044) );
  NAND2_X1 U9618 ( .A1(n9028), .A2(n9027), .ZN(n7100) );
  NAND2_X1 U9619 ( .A1(n9115), .A2(n7104), .ZN(n7101) );
  NAND2_X1 U9620 ( .A1(n7101), .A2(n7102), .ZN(n9143) );
  OAI21_X1 U9621 ( .B1(n9058), .B2(n7110), .A(n7108), .ZN(n9090) );
  NAND2_X1 U9622 ( .A1(n7390), .A2(n7391), .ZN(n8978) );
  NAND3_X1 U9623 ( .A1(n8992), .A2(n7119), .A3(P1_DATAO_REG_13__SCAN_IN), .ZN(
        n8993) );
  NAND2_X1 U9624 ( .A1(n7390), .A2(n6742), .ZN(n7119) );
  OAI21_X1 U9625 ( .B1(n9389), .B2(n15608), .A(n9390), .ZN(n9391) );
  NAND2_X2 U9626 ( .A1(n7122), .A2(n7897), .ZN(n7929) );
  NAND2_X1 U9627 ( .A1(n7319), .A2(n7122), .ZN(n8672) );
  NAND2_X1 U9628 ( .A1(n7976), .A2(n7123), .ZN(n7977) );
  OAI211_X1 U9629 ( .C1(n7130), .C2(n7129), .A(n7126), .B(n8051), .ZN(n7125)
         );
  AOI21_X1 U9630 ( .B1(n7131), .B2(n8048), .A(n8047), .ZN(n7129) );
  OAI22_X1 U9631 ( .A1(n7131), .A2(n8048), .B1(n8050), .B2(n8049), .ZN(n7130)
         );
  NAND4_X1 U9632 ( .A1(n7136), .A2(n7134), .A3(n7133), .A4(n7132), .ZN(n8648)
         );
  AND2_X2 U9633 ( .A1(n7135), .A2(n7906), .ZN(n8160) );
  INV_X1 U9634 ( .A(n7907), .ZN(n7135) );
  NAND2_X1 U9635 ( .A1(n7996), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7136) );
  INV_X1 U9636 ( .A(n7906), .ZN(n13402) );
  INV_X1 U9637 ( .A(n8484), .ZN(n7139) );
  AND2_X1 U9638 ( .A1(n8417), .A2(n8418), .ZN(n7151) );
  OAI21_X1 U9639 ( .B1(n8417), .B2(n8418), .A(n7762), .ZN(n7142) );
  OAI21_X1 U9640 ( .B1(n8417), .B2(n7143), .A(n6595), .ZN(n7146) );
  NAND2_X1 U9641 ( .A1(n7147), .A2(n7152), .ZN(n8459) );
  NAND2_X1 U9642 ( .A1(n7148), .A2(n7150), .ZN(n7147) );
  OAI21_X1 U9643 ( .B1(n8238), .B2(n7767), .A(n7156), .ZN(n7155) );
  NOR2_X1 U9644 ( .A1(n8237), .A2(n8236), .ZN(n7157) );
  INV_X1 U9645 ( .A(n8258), .ZN(n7158) );
  OAI22_X1 U9646 ( .A1(n7293), .A2(n7292), .B1(n8196), .B2(n7291), .ZN(n8219)
         );
  OAI22_X1 U9647 ( .A1(n7277), .A2(n7276), .B1(n7275), .B2(n7274), .ZN(n8328)
         );
  OAI21_X1 U9648 ( .B1(n7290), .B2(n7289), .A(n7763), .ZN(n8417) );
  NAND2_X1 U9649 ( .A1(n7168), .A2(n8528), .ZN(n8600) );
  NOR2_X1 U9650 ( .A1(n7167), .A2(n7194), .ZN(n7193) );
  OAI21_X1 U9651 ( .B1(n8376), .B2(n8375), .A(n7765), .ZN(n7289) );
  INV_X1 U9652 ( .A(n8217), .ZN(n7179) );
  NAND2_X1 U9653 ( .A1(n7169), .A2(n7902), .ZN(n7919) );
  NAND3_X1 U9654 ( .A1(n8107), .A2(n7171), .A3(n7743), .ZN(n7192) );
  NAND2_X1 U9655 ( .A1(n8106), .A2(n8105), .ZN(n7171) );
  NAND3_X1 U9656 ( .A1(n10594), .A2(n6648), .A3(n10595), .ZN(n7670) );
  NAND2_X1 U9657 ( .A1(n8791), .A2(n8793), .ZN(n7414) );
  NAND2_X1 U9658 ( .A1(n11774), .A2(n9174), .ZN(n11855) );
  NAND2_X1 U9659 ( .A1(n7174), .A2(n7172), .ZN(P3_U3180) );
  NAND2_X1 U9660 ( .A1(n11857), .A2(n11863), .ZN(n7174) );
  NAND3_X1 U9661 ( .A1(n10476), .A2(n8809), .A3(n10586), .ZN(n10475) );
  NAND2_X1 U9662 ( .A1(n7671), .A2(n7670), .ZN(n10959) );
  NAND2_X1 U9663 ( .A1(n7655), .A2(n7657), .ZN(n11864) );
  NAND2_X1 U9664 ( .A1(n11393), .A2(n11392), .ZN(n11391) );
  NAND2_X1 U9665 ( .A1(n7944), .A2(SI_1_), .ZN(n7957) );
  OAI211_X1 U9666 ( .C1(n8459), .C2(n7280), .A(n7279), .B(n8483), .ZN(n8484)
         );
  NAND2_X1 U9667 ( .A1(n6666), .A2(n7178), .ZN(n8238) );
  NAND2_X1 U9668 ( .A1(n7180), .A2(n7179), .ZN(n7178) );
  NAND2_X1 U9669 ( .A1(n8219), .A2(n8218), .ZN(n7180) );
  AOI21_X1 U9670 ( .B1(n8007), .B2(n8006), .A(n8005), .ZN(n8008) );
  NAND2_X1 U9671 ( .A1(n7181), .A2(n8349), .ZN(n8352) );
  INV_X1 U9672 ( .A(n7182), .ZN(n7181) );
  AOI21_X1 U9673 ( .B1(n8328), .B2(n7752), .A(n7750), .ZN(n7182) );
  NAND2_X1 U9674 ( .A1(n7986), .A2(n7985), .ZN(n8007) );
  AOI21_X2 U9675 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(n14744), .A(n14791), .ZN(
        n14963) );
  NAND2_X1 U9676 ( .A1(n14812), .A2(n7465), .ZN(n7464) );
  XNOR2_X1 U9677 ( .A(n7464), .B(n7463), .ZN(SUB_1596_U4) );
  NAND2_X1 U9678 ( .A1(n10132), .A2(n7527), .ZN(n10347) );
  OR2_X1 U9679 ( .A1(n10396), .A2(n7166), .ZN(n10397) );
  NOR2_X2 U9680 ( .A1(n10751), .A2(n11003), .ZN(n10995) );
  OAI21_X1 U9681 ( .B1(n8680), .B2(n7193), .A(n11491), .ZN(n8699) );
  NAND2_X1 U9682 ( .A1(n8109), .A2(n8108), .ZN(n8113) );
  NAND2_X1 U9683 ( .A1(n7192), .A2(n7745), .ZN(n8151) );
  NAND2_X1 U9684 ( .A1(n8103), .A2(n8104), .ZN(n8102) );
  NAND2_X2 U9685 ( .A1(n10146), .A2(n10197), .ZN(n8635) );
  OAI21_X2 U9686 ( .B1(n12481), .B2(n12483), .A(n12042), .ZN(n12467) );
  INV_X1 U9687 ( .A(n9228), .ZN(n12079) );
  XNOR2_X1 U9688 ( .A(n9107), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n9106) );
  NAND2_X1 U9689 ( .A1(n9044), .A2(n9043), .ZN(n9058) );
  NAND2_X1 U9690 ( .A1(n8993), .A2(n8992), .ZN(n9010) );
  OAI21_X1 U9691 ( .B1(n9160), .B2(n7400), .A(n9177), .ZN(n7399) );
  NAND2_X1 U9692 ( .A1(n9283), .A2(n9282), .ZN(n9288) );
  NAND2_X1 U9693 ( .A1(n12556), .A2(n12013), .ZN(n9339) );
  NAND2_X1 U9694 ( .A1(n12470), .A2(n12469), .ZN(n12468) );
  AOI21_X1 U9695 ( .B1(n12431), .B2(n12636), .A(n12430), .ZN(n12432) );
  NAND2_X1 U9696 ( .A1(n7673), .A2(n6648), .ZN(n7671) );
  NAND2_X1 U9697 ( .A1(n10959), .A2(n10960), .ZN(n10958) );
  NAND2_X1 U9698 ( .A1(n8813), .A2(n8812), .ZN(n7675) );
  NAND2_X1 U9699 ( .A1(n10771), .A2(n13885), .ZN(n7715) );
  NAND4_X1 U9700 ( .A1(n14457), .A2(n14455), .A3(n14454), .A4(n14456), .ZN(
        n14540) );
  NOR2_X1 U9701 ( .A1(n7414), .A2(n7413), .ZN(n7412) );
  OAI21_X1 U9702 ( .B1(n12721), .B2(n15601), .A(n7198), .ZN(P3_U3454) );
  NAND2_X1 U9703 ( .A1(n11409), .A2(n11983), .ZN(n11412) );
  NAND2_X1 U9704 ( .A1(n12660), .A2(n6731), .ZN(P3_U3486) );
  NAND2_X1 U9705 ( .A1(n12602), .A2(n9331), .ZN(n12583) );
  OAI21_X1 U9706 ( .B1(n8737), .B2(n7201), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8761) );
  NAND2_X1 U9707 ( .A1(n12426), .A2(n7203), .ZN(n12431) );
  INV_X1 U9708 ( .A(n14451), .ZN(n7713) );
  NAND2_X1 U9709 ( .A1(n7262), .A2(n6746), .ZN(P1_U3525) );
  NAND3_X1 U9710 ( .A1(n7712), .A2(n7361), .A3(n7204), .ZN(n14539) );
  NAND2_X1 U9711 ( .A1(n14716), .A2(n14717), .ZN(n7460) );
  INV_X1 U9712 ( .A(n14961), .ZN(n7457) );
  NAND2_X1 U9713 ( .A1(n14747), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7456) );
  OAI21_X1 U9714 ( .B1(n12433), .B2(n12434), .A(n12432), .ZN(n12657) );
  XNOR2_X1 U9715 ( .A(n7205), .B(n8009), .ZN(n10215) );
  OAI21_X1 U9716 ( .B1(n8082), .B2(n7210), .A(n7208), .ZN(n8130) );
  NAND3_X1 U9717 ( .A1(n14014), .A2(n14013), .A3(n7552), .ZN(n7213) );
  INV_X1 U9718 ( .A(n13991), .ZN(n7217) );
  NAND2_X1 U9719 ( .A1(n7219), .A2(n7220), .ZN(n14009) );
  NAND3_X1 U9720 ( .A1(n14003), .A2(n6714), .A3(n14002), .ZN(n7219) );
  NAND3_X1 U9721 ( .A1(n13970), .A2(n7223), .A3(n13969), .ZN(n7221) );
  NAND2_X1 U9722 ( .A1(n10738), .A2(n10739), .ZN(n10741) );
  NAND2_X1 U9723 ( .A1(n7227), .A2(n10540), .ZN(n10738) );
  NAND2_X1 U9724 ( .A1(n10539), .A2(n10538), .ZN(n7227) );
  NAND2_X1 U9725 ( .A1(n10449), .A2(n10448), .ZN(n10539) );
  AND3_X2 U9726 ( .A1(n7894), .A2(n7895), .A3(n7893), .ZN(n8178) );
  INV_X1 U9727 ( .A(n13209), .ZN(n7237) );
  OAI21_X2 U9728 ( .B1(n7237), .B2(n7234), .A(n7232), .ZN(n13147) );
  NAND2_X1 U9729 ( .A1(n7242), .A2(n7240), .ZN(n7246) );
  NAND2_X1 U9730 ( .A1(n7246), .A2(n11305), .ZN(n11306) );
  NAND2_X1 U9731 ( .A1(n13266), .A2(n7250), .ZN(n7248) );
  NAND2_X1 U9732 ( .A1(n7248), .A2(n7247), .ZN(n13046) );
  INV_X2 U9733 ( .A(n13836), .ZN(n11615) );
  INV_X1 U9734 ( .A(n14425), .ZN(n7259) );
  INV_X1 U9735 ( .A(n13892), .ZN(n7261) );
  NAND2_X1 U9736 ( .A1(n7593), .A2(n6578), .ZN(n7266) );
  INV_X2 U9737 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8056) );
  NAND2_X1 U9738 ( .A1(n7758), .A2(n8306), .ZN(n7274) );
  NOR2_X1 U9739 ( .A1(n8280), .A2(n7761), .ZN(n7275) );
  INV_X1 U9740 ( .A(n8304), .ZN(n7276) );
  NOR2_X2 U9741 ( .A1(n10945), .A2(n7287), .ZN(n10197) );
  INV_X2 U9742 ( .A(n9938), .ZN(n7288) );
  INV_X1 U9743 ( .A(n10292), .ZN(n7306) );
  NAND2_X1 U9744 ( .A1(n7309), .A2(n10198), .ZN(n10199) );
  NOR2_X1 U9745 ( .A1(n10151), .A2(n7309), .ZN(n10125) );
  NOR2_X1 U9746 ( .A1(n15370), .A2(n7309), .ZN(n10308) );
  NAND2_X1 U9747 ( .A1(n12969), .A2(n7310), .ZN(n12868) );
  NAND3_X1 U9748 ( .A1(n7582), .A2(n7313), .A3(n10283), .ZN(n7312) );
  INV_X1 U9749 ( .A(n10100), .ZN(n7313) );
  XNOR2_X1 U9750 ( .A(n10280), .B(n10281), .ZN(n10100) );
  NAND2_X1 U9751 ( .A1(n10538), .A2(n7322), .ZN(n7320) );
  NAND3_X1 U9752 ( .A1(n7330), .A2(n11191), .A3(n6716), .ZN(n7326) );
  NAND2_X1 U9753 ( .A1(n13245), .A2(n7335), .ZN(n7334) );
  OAI21_X2 U9754 ( .B1(n13197), .B2(n7345), .A(n7342), .ZN(n7732) );
  AND2_X2 U9755 ( .A1(n13290), .A2(n7348), .ZN(n7787) );
  AOI21_X2 U9756 ( .B1(n7728), .B2(n7727), .A(n7349), .ZN(n13122) );
  OR2_X1 U9757 ( .A1(n14284), .A2(n14177), .ZN(n7352) );
  NAND2_X1 U9758 ( .A1(n8244), .A2(n7356), .ZN(n7355) );
  NAND3_X1 U9759 ( .A1(n7621), .A2(n7622), .A3(n7623), .ZN(n7362) );
  NAND2_X1 U9760 ( .A1(n14594), .A2(n7370), .ZN(n7369) );
  INV_X1 U9761 ( .A(n7373), .ZN(n14857) );
  NAND2_X1 U9762 ( .A1(n15529), .A2(n7376), .ZN(n7375) );
  INV_X1 U9763 ( .A(n14620), .ZN(n7377) );
  NAND3_X1 U9764 ( .A1(n7380), .A2(P3_IR_REG_2__SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n7379) );
  NAND2_X1 U9765 ( .A1(n9010), .A2(n9009), .ZN(n7383) );
  NAND2_X1 U9766 ( .A1(n8954), .A2(n7393), .ZN(n7390) );
  INV_X1 U9767 ( .A(n7399), .ZN(n7398) );
  NAND2_X1 U9768 ( .A1(n9283), .A2(n7404), .ZN(n7403) );
  NAND2_X1 U9769 ( .A1(n7411), .A2(n7410), .ZN(n15578) );
  NAND2_X1 U9770 ( .A1(n10703), .A2(n10707), .ZN(n7410) );
  OR2_X1 U9771 ( .A1(n10703), .A2(n10707), .ZN(n7411) );
  INV_X1 U9772 ( .A(n10317), .ZN(n10316) );
  AND2_X1 U9773 ( .A1(n7415), .A2(n10317), .ZN(n10315) );
  OAI211_X1 U9774 ( .C1(n15402), .C2(n10163), .A(n8783), .B(n8782), .ZN(n10317) );
  OAI21_X1 U9775 ( .B1(n12457), .B2(n7421), .A(n7419), .ZN(n12418) );
  NAND2_X1 U9776 ( .A1(n7418), .A2(n7416), .ZN(n11877) );
  NAND3_X1 U9777 ( .A1(n12457), .A2(n7419), .A3(n12417), .ZN(n7418) );
  NOR2_X1 U9778 ( .A1(n7426), .A2(n7431), .ZN(n7425) );
  NAND2_X1 U9779 ( .A1(n10824), .A2(n7425), .ZN(n7429) );
  OR2_X1 U9780 ( .A1(n7431), .A2(n7428), .ZN(n7427) );
  NAND3_X1 U9781 ( .A1(n9270), .A2(n9271), .A3(n9269), .ZN(n11409) );
  NAND2_X1 U9782 ( .A1(n9270), .A2(n9269), .ZN(n11475) );
  INV_X1 U9783 ( .A(n7470), .ZN(n7469) );
  NAND2_X1 U9784 ( .A1(n7472), .A2(n10730), .ZN(n10912) );
  NAND2_X1 U9785 ( .A1(n10727), .A2(n10726), .ZN(n7472) );
  INV_X1 U9786 ( .A(n10911), .ZN(n7473) );
  NAND2_X1 U9787 ( .A1(n13657), .A2(n7478), .ZN(n7477) );
  NAND2_X1 U9788 ( .A1(n13613), .A2(n13612), .ZN(n7490) );
  OR2_X1 U9789 ( .A1(n13537), .A2(n13536), .ZN(n7510) );
  NAND2_X1 U9790 ( .A1(n11682), .A2(n7514), .ZN(n7511) );
  NAND2_X1 U9791 ( .A1(n7511), .A2(n7512), .ZN(n13788) );
  NAND2_X1 U9792 ( .A1(n11682), .A2(n11681), .ZN(n13481) );
  NAND3_X1 U9793 ( .A1(n6573), .A2(n11694), .A3(n14088), .ZN(n7590) );
  NAND2_X1 U9794 ( .A1(n7925), .A2(n7526), .ZN(n8684) );
  INV_X1 U9795 ( .A(n8684), .ZN(n7918) );
  AND2_X1 U9796 ( .A1(n10440), .A2(n15358), .ZN(n10131) );
  NOR2_X2 U9797 ( .A1(n13141), .A2(n13301), .ZN(n13126) );
  NOR2_X2 U9798 ( .A1(n11069), .A2(n11195), .ZN(n7538) );
  NAND2_X1 U9799 ( .A1(n13890), .A2(n13889), .ZN(n7543) );
  NAND2_X1 U9800 ( .A1(n7540), .A2(n13893), .ZN(n13897) );
  NAND2_X1 U9801 ( .A1(n13890), .A2(n7541), .ZN(n7540) );
  NOR2_X1 U9802 ( .A1(n7542), .A2(n13894), .ZN(n7541) );
  INV_X1 U9803 ( .A(n13889), .ZN(n7542) );
  NAND2_X1 U9804 ( .A1(n7543), .A2(n13894), .ZN(n13896) );
  AOI21_X1 U9805 ( .B1(n13982), .B2(n7547), .A(n7545), .ZN(n7544) );
  OAI21_X1 U9806 ( .B1(n13982), .B2(n6634), .A(n7547), .ZN(n13985) );
  INV_X1 U9807 ( .A(n7544), .ZN(n13984) );
  INV_X1 U9808 ( .A(n13993), .ZN(n7551) );
  AND2_X1 U9809 ( .A1(n14026), .A2(n6623), .ZN(n7553) );
  NOR2_X1 U9810 ( .A1(n13928), .A2(n13927), .ZN(n13931) );
  INV_X1 U9811 ( .A(n13921), .ZN(n7555) );
  NAND2_X1 U9812 ( .A1(n7556), .A2(n7557), .ZN(n13908) );
  NAND2_X1 U9813 ( .A1(n13905), .A2(n7559), .ZN(n7556) );
  AOI21_X1 U9814 ( .B1(n13928), .B2(n13927), .A(n13926), .ZN(n13932) );
  NAND2_X1 U9815 ( .A1(n13912), .A2(n13911), .ZN(n13916) );
  NAND2_X1 U9816 ( .A1(n9090), .A2(n9089), .ZN(n9107) );
  NAND2_X1 U9817 ( .A1(n9146), .A2(n9145), .ZN(n9147) );
  NAND2_X1 U9818 ( .A1(n12893), .A2(n7572), .ZN(n7571) );
  NAND2_X1 U9819 ( .A1(n10682), .A2(n10681), .ZN(n10970) );
  INV_X2 U9820 ( .A(n12806), .ZN(n12869) );
  NOR2_X2 U9821 ( .A1(n14406), .A2(n14414), .ZN(n14393) );
  NOR2_X2 U9822 ( .A1(n14311), .A2(n14304), .ZN(n7601) );
  NAND4_X1 U9823 ( .A1(n7912), .A2(n14767), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7603) );
  NAND3_X1 U9824 ( .A1(n7604), .A2(P1_DATAO_REG_1__SCAN_IN), .A3(n7603), .ZN(
        n7605) );
  OAI21_X1 U9825 ( .B1(n8174), .B2(n7615), .A(n7614), .ZN(n8221) );
  NAND3_X1 U9826 ( .A1(n7621), .A2(n6755), .A3(n7623), .ZN(n8489) );
  NAND2_X1 U9827 ( .A1(n8465), .A2(n6754), .ZN(n7623) );
  NAND2_X1 U9828 ( .A1(n7620), .A2(SI_24_), .ZN(n7621) );
  NAND2_X1 U9829 ( .A1(n8550), .A2(n8549), .ZN(n8569) );
  NAND4_X1 U9830 ( .A1(n8550), .A2(n8549), .A3(n7629), .A4(n8581), .ZN(n7625)
         );
  NAND3_X1 U9831 ( .A1(n8550), .A2(n8549), .A3(n7629), .ZN(n7626) );
  OAI21_X1 U9832 ( .B1(n8509), .B2(n7644), .A(n7639), .ZN(n8547) );
  NAND2_X1 U9833 ( .A1(n7637), .A2(n7638), .ZN(n8546) );
  NAND2_X1 U9834 ( .A1(n9173), .A2(n11772), .ZN(n11774) );
  INV_X1 U9835 ( .A(n11817), .ZN(n7666) );
  NAND2_X1 U9836 ( .A1(n11817), .A2(n7660), .ZN(n7655) );
  INV_X1 U9837 ( .A(n11738), .ZN(n7669) );
  NAND2_X1 U9838 ( .A1(n7675), .A2(n10783), .ZN(n7673) );
  AOI21_X1 U9839 ( .B1(n8718), .B2(n6712), .A(n8709), .ZN(n8711) );
  AND2_X1 U9840 ( .A1(n8718), .A2(n8714), .ZN(n8728) );
  NAND2_X1 U9841 ( .A1(n14376), .A2(n14390), .ZN(n7699) );
  OR2_X1 U9842 ( .A1(n14522), .A2(n14171), .ZN(n7700) );
  INV_X1 U9843 ( .A(n7708), .ZN(n11426) );
  NAND2_X1 U9844 ( .A1(n15057), .A2(n7714), .ZN(n11237) );
  OAI21_X1 U9845 ( .B1(n10202), .B2(n7331), .A(n7716), .ZN(n10123) );
  NAND2_X1 U9846 ( .A1(n10203), .A2(n10204), .ZN(n10202) );
  NAND3_X1 U9847 ( .A1(n13184), .A2(n7724), .A3(n7725), .ZN(n7720) );
  INV_X1 U9848 ( .A(n8196), .ZN(n7741) );
  INV_X1 U9849 ( .A(n8637), .ZN(n7742) );
  OAI22_X1 U9850 ( .A1(n7907), .A2(P2_U3088), .B1(n11726), .B2(n13417), .ZN(
        n7749) );
  NAND2_X1 U9851 ( .A1(n10117), .A2(n7776), .ZN(n7775) );
  OAI21_X1 U9852 ( .B1(n7775), .B2(n7774), .A(n7772), .ZN(n10447) );
  NAND3_X1 U9853 ( .A1(n7782), .A2(n7783), .A3(n7778), .ZN(n13291) );
  NAND3_X1 U9854 ( .A1(n7782), .A2(n7780), .A3(n7778), .ZN(n7785) );
  NAND3_X1 U9855 ( .A1(n13105), .A2(n7788), .A3(n13093), .ZN(n7782) );
  OR2_X1 U9856 ( .A1(n15383), .A2(n12257), .ZN(n7786) );
  INV_X1 U9857 ( .A(n7923), .ZN(n8334) );
  AND2_X2 U9858 ( .A1(n7923), .A2(n10019), .ZN(n8561) );
  MUX2_X1 U9859 ( .A(n9518), .B(n13418), .S(n7923), .Z(n10129) );
  AND2_X1 U9860 ( .A1(n13364), .A2(n12978), .ZN(n7809) );
  NAND4_X1 U9861 ( .A1(n6743), .A2(n9448), .A3(n9393), .A4(n7814), .ZN(n9545)
         );
  NAND2_X1 U9862 ( .A1(n9448), .A2(n9392), .ZN(n9452) );
  INV_X1 U9863 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7814) );
  INV_X1 U9864 ( .A(n10763), .ZN(n7816) );
  NAND2_X1 U9865 ( .A1(n7820), .A2(n10228), .ZN(n10407) );
  NAND2_X1 U9866 ( .A1(n15053), .A2(n6707), .ZN(n7824) );
  INV_X1 U9867 ( .A(n14427), .ZN(n13810) );
  NAND2_X1 U9868 ( .A1(n14420), .A2(n14427), .ZN(n14419) );
  NAND2_X1 U9869 ( .A1(n13872), .A2(n13871), .ZN(n14427) );
  NAND2_X1 U9870 ( .A1(n7849), .A2(n7850), .ZN(n11470) );
  NAND2_X1 U9871 ( .A1(n12520), .A2(n7859), .ZN(n7858) );
  AND2_X1 U9872 ( .A1(n7861), .A2(n6592), .ZN(n12504) );
  NAND2_X1 U9873 ( .A1(n9308), .A2(n6657), .ZN(n10664) );
  NAND2_X1 U9874 ( .A1(n10664), .A2(n7864), .ZN(n10666) );
  AOI21_X1 U9875 ( .B1(n7865), .B2(n9309), .A(n12584), .ZN(n7864) );
  OAI21_X1 U9876 ( .B1(n12427), .B2(n7868), .A(n7866), .ZN(n9352) );
  NAND2_X1 U9877 ( .A1(n10826), .A2(n11911), .ZN(n10829) );
  NAND2_X1 U9878 ( .A1(n10147), .A2(n10146), .ZN(n15369) );
  OR2_X1 U9879 ( .A1(n13861), .A2(n14032), .ZN(n10776) );
  NAND2_X1 U9880 ( .A1(n10741), .A2(n10740), .ZN(n10985) );
  NAND2_X1 U9881 ( .A1(n8684), .A2(n8689), .ZN(n13412) );
  OAI21_X1 U9882 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(n7920), .A(n7919), .ZN(
        n7921) );
  AOI22_X1 U9883 ( .A1(n6574), .A2(n8592), .B1(n12994), .B2(n8635), .ZN(n7976)
         );
  NAND4_X2 U9884 ( .A1(n7973), .A2(n7972), .A3(n7971), .A4(n7970), .ZN(n12992)
         );
  NAND2_X1 U9885 ( .A1(n9267), .A2(n11936), .ZN(n10703) );
  AOI21_X1 U9886 ( .B1(n11936), .B2(n8805), .A(n8807), .ZN(n8810) );
  INV_X1 U9887 ( .A(n8796), .ZN(n8801) );
  INV_X1 U9888 ( .A(n9305), .ZN(n10707) );
  NOR2_X1 U9889 ( .A1(n8758), .A2(n8739), .ZN(n8740) );
  OR2_X1 U9890 ( .A1(n13924), .A2(n13925), .ZN(n7876) );
  OR2_X1 U9891 ( .A1(n11718), .A2(n12770), .ZN(n7877) );
  AND2_X1 U9892 ( .A1(n9371), .A2(n9370), .ZN(n15601) );
  INV_X2 U9893 ( .A(n15608), .ZN(n15611) );
  AND4_X1 U9894 ( .A1(n8707), .A2(n8706), .A3(n8705), .A4(n8704), .ZN(n7878)
         );
  AND2_X1 U9895 ( .A1(n12743), .A2(n11756), .ZN(n7879) );
  AND2_X1 U9896 ( .A1(n11729), .A2(n12586), .ZN(n7880) );
  OR2_X1 U9897 ( .A1(n8021), .A2(n8635), .ZN(n7881) );
  OR2_X1 U9898 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10172), .ZN(n7882) );
  AND2_X1 U9899 ( .A1(n13436), .A2(P2_U3088), .ZN(n13404) );
  INV_X1 U9900 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7991) );
  AND2_X1 U9901 ( .A1(n14206), .A2(n15080), .ZN(n15093) );
  INV_X1 U9902 ( .A(n15093), .ZN(n14379) );
  INV_X1 U9903 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9033) );
  INV_X1 U9904 ( .A(n13256), .ZN(n13280) );
  INV_X1 U9905 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14725) );
  OAI21_X1 U9906 ( .B1(n13707), .B2(n13692), .A(n13459), .ZN(n14347) );
  OR2_X1 U9907 ( .A1(n11718), .A2(n12715), .ZN(n7883) );
  INV_X1 U9908 ( .A(n11742), .ZN(n12739) );
  INV_X1 U9909 ( .A(n13823), .ZN(n14168) );
  NAND2_X2 U9910 ( .A1(n9936), .A2(n13236), .ZN(n13252) );
  AND2_X1 U9911 ( .A1(n12747), .A2(n12522), .ZN(n7884) );
  OR2_X1 U9912 ( .A1(n11906), .A2(n12719), .ZN(n7885) );
  AND3_X1 U9913 ( .A1(n9141), .A2(n9140), .A3(n9139), .ZN(n12495) );
  INV_X1 U9914 ( .A(n12495), .ZN(n9346) );
  OR2_X1 U9915 ( .A1(n10248), .A2(n10247), .ZN(n15208) );
  INV_X2 U9916 ( .A(n15208), .ZN(n15209) );
  AND2_X1 U9917 ( .A1(n13858), .A2(n13871), .ZN(n13859) );
  OR2_X1 U9918 ( .A1(n14021), .A2(n15156), .ZN(n13875) );
  NAND2_X1 U9919 ( .A1(n8302), .A2(n8301), .ZN(n8305) );
  INV_X1 U9920 ( .A(n8305), .ZN(n8306) );
  NAND2_X1 U9921 ( .A1(n13962), .A2(n13961), .ZN(n13963) );
  NAND2_X1 U9922 ( .A1(n8352), .A2(n8351), .ZN(n8376) );
  NAND2_X1 U9923 ( .A1(n13988), .A2(n13987), .ZN(n13989) );
  INV_X1 U9924 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8704) );
  INV_X1 U9925 ( .A(n8594), .ZN(n8595) );
  OR4_X1 U9926 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n9217) );
  INV_X1 U9927 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8702) );
  INV_X1 U9928 ( .A(n12546), .ZN(n9340) );
  INV_X1 U9929 ( .A(n7914), .ZN(n7915) );
  INV_X1 U9930 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7924) );
  INV_X1 U9931 ( .A(n13681), .ZN(n10717) );
  INV_X1 U9932 ( .A(n14347), .ZN(n14175) );
  OAI22_X1 U9933 ( .A1(n6569), .A2(n9427), .B1(n10163), .B2(n10279), .ZN(n8796) );
  INV_X1 U9934 ( .A(n12531), .ZN(n9342) );
  INV_X1 U9935 ( .A(n11971), .ZN(n9320) );
  INV_X1 U9936 ( .A(n9309), .ZN(n9310) );
  INV_X1 U9937 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8403) );
  INV_X1 U9938 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7916) );
  INV_X1 U9939 ( .A(n10508), .ZN(n10505) );
  OAI211_X1 U9940 ( .C1(n14158), .C2(n14157), .A(n14031), .B(n14030), .ZN(
        n14038) );
  INV_X1 U9941 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13545) );
  INV_X1 U9942 ( .A(n14195), .ZN(n14173) );
  AND2_X1 U9943 ( .A1(n9397), .A2(n9396), .ZN(n9408) );
  INV_X1 U9944 ( .A(n9206), .ZN(n9204) );
  OR2_X1 U9945 ( .A1(n9122), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9137) );
  INV_X1 U9946 ( .A(n15501), .ZN(n14646) );
  INV_X1 U9947 ( .A(n12503), .ZN(n9344) );
  NAND2_X1 U9948 ( .A1(n11984), .A2(n11990), .ZN(n11917) );
  NAND2_X1 U9949 ( .A1(n11368), .A2(n11973), .ZN(n11350) );
  AND2_X1 U9950 ( .A1(n11959), .A2(n11960), .ZN(n11909) );
  OR2_X1 U9951 ( .A1(n12771), .A2(n9227), .ZN(n9364) );
  OR2_X1 U9952 ( .A1(n8535), .A2(n12843), .ZN(n8574) );
  OR2_X1 U9953 ( .A1(n8495), .A2(n12887), .ZN(n8516) );
  OR2_X1 U9954 ( .A1(n8404), .A2(n8403), .ZN(n8427) );
  OR2_X1 U9955 ( .A1(n15250), .A2(n15249), .ZN(n15252) );
  INV_X1 U9956 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8364) );
  AND2_X1 U9957 ( .A1(n9939), .A2(n11403), .ZN(n9703) );
  NAND2_X1 U9958 ( .A1(n13098), .A2(n13097), .ZN(n13099) );
  INV_X1 U9959 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7903) );
  NOR2_X1 U9960 ( .A1(n13546), .A2(n13545), .ZN(n13547) );
  INV_X1 U9961 ( .A(n14797), .ZN(n13930) );
  NAND2_X1 U9962 ( .A1(n13861), .A2(n15139), .ZN(n14023) );
  OR2_X1 U9963 ( .A1(n10212), .A2(n15140), .ZN(n13857) );
  INV_X1 U9964 ( .A(n14059), .ZN(n11654) );
  NAND2_X1 U9965 ( .A1(n8548), .A2(SI_27_), .ZN(n8549) );
  OR2_X1 U9966 ( .A1(n14731), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14679) );
  NOR2_X1 U9967 ( .A1(n8861), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8888) );
  OR2_X1 U9968 ( .A1(n9003), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9017) );
  INV_X1 U9969 ( .A(n11604), .ZN(n8931) );
  NAND2_X1 U9970 ( .A1(n8801), .A2(n8800), .ZN(n8802) );
  INV_X1 U9971 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n11777) );
  INV_X1 U9972 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n11809) );
  NAND3_X1 U9973 ( .A1(n12773), .A2(n12771), .A3(n9377), .ZN(n9367) );
  NAND2_X1 U9974 ( .A1(n10373), .A2(n10372), .ZN(n10374) );
  AOI21_X1 U9975 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10547), .A(n10544), .ZN(
        n12380) );
  INV_X1 U9976 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11563) );
  INV_X1 U9977 ( .A(n14655), .ZN(n14845) );
  INV_X1 U9978 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12256) );
  AND2_X1 U9979 ( .A1(n12005), .A2(n12004), .ZN(n12591) );
  OR2_X1 U9980 ( .A1(n10658), .A2(n10705), .ZN(n12641) );
  INV_X1 U9981 ( .A(n11911), .ZN(n11948) );
  AND2_X1 U9982 ( .A1(n9377), .A2(n10160), .ZN(n9378) );
  AND2_X1 U9983 ( .A1(n9300), .A2(n9380), .ZN(n12433) );
  NOR2_X1 U9984 ( .A1(n9259), .A2(n12044), .ZN(n9368) );
  INV_X1 U9985 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12887) );
  INV_X1 U9986 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n12902) );
  INV_X1 U9987 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11225) );
  NOR2_X1 U9988 ( .A1(n15326), .A2(n10144), .ZN(n9935) );
  INV_X1 U9989 ( .A(n8666), .ZN(n8670) );
  AND2_X1 U9990 ( .A1(n8516), .A2(n8496), .ZN(n13162) );
  INV_X1 U9991 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10633) );
  INV_X1 U9992 ( .A(n13053), .ZN(n13086) );
  OR2_X1 U9993 ( .A1(n8365), .A2(n8364), .ZN(n8384) );
  NAND2_X1 U9994 ( .A1(n9704), .A2(n9703), .ZN(n12916) );
  NAND2_X1 U9995 ( .A1(n13252), .A2(n10133), .ZN(n13277) );
  AND2_X1 U9996 ( .A1(n8679), .A2(n8681), .ZN(n8690) );
  NOR2_X1 U9997 ( .A1(n8203), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8226) );
  INV_X1 U9998 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13667) );
  NOR2_X1 U9999 ( .A1(n11625), .A2(n12184), .ZN(n13511) );
  OR2_X1 U10000 ( .A1(n13505), .A2(n13504), .ZN(n13506) );
  OR2_X1 U10001 ( .A1(n10764), .A2(n10765), .ZN(n10013) );
  NAND2_X1 U10002 ( .A1(n15196), .A2(n10036), .ZN(n14050) );
  AND2_X1 U10003 ( .A1(n13547), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n13455) );
  INV_X1 U10004 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14685) );
  INV_X1 U10005 ( .A(n14151), .ZN(n14447) );
  NAND2_X1 U10006 ( .A1(n6735), .A2(n14339), .ZN(n14338) );
  AND2_X1 U10007 ( .A1(n10766), .A2(n10765), .ZN(n10767) );
  INV_X1 U10008 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n12362) );
  INV_X1 U10009 ( .A(n13899), .ZN(n15095) );
  INV_X1 U10010 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14554) );
  AND2_X1 U10011 ( .A1(n9752), .A2(n12306), .ZN(n9931) );
  INV_X1 U10012 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14711) );
  NAND2_X1 U10013 ( .A1(n9231), .A2(n9230), .ZN(n9420) );
  OAI21_X1 U10014 ( .B1(n12723), .B2(n11875), .A(n9263), .ZN(n9264) );
  INV_X1 U10015 ( .A(n11875), .ZN(n11850) );
  NAND2_X1 U10016 ( .A1(n9245), .A2(n9244), .ZN(n11872) );
  AOI21_X1 U10017 ( .B1(n12419), .B2(n8789), .A(n9253), .ZN(n12429) );
  AND4_X1 U10018 ( .A1(n9071), .A2(n9070), .A3(n9069), .A4(n9068), .ZN(n9274)
         );
  INV_X1 U10019 ( .A(n10964), .ZN(n9268) );
  INV_X1 U10020 ( .A(n15406), .ZN(n15407) );
  NOR2_X1 U10021 ( .A1(n14579), .A2(n15461), .ZN(n15479) );
  AND2_X1 U10022 ( .A1(P3_U3897), .A2(n9254), .ZN(n15543) );
  INV_X1 U10023 ( .A(n12589), .ZN(n12633) );
  NAND2_X1 U10024 ( .A1(n15608), .A2(n9293), .ZN(n9390) );
  AND2_X1 U10025 ( .A1(n9379), .A2(n9378), .ZN(n10581) );
  AND2_X1 U10026 ( .A1(n12433), .A2(n12656), .ZN(n14910) );
  INV_X1 U10027 ( .A(n14910), .ZN(n15595) );
  NAND2_X1 U10028 ( .A1(n11932), .A2(n14790), .ZN(n12621) );
  OR2_X1 U10029 ( .A1(n9013), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n9047) );
  INV_X1 U10030 ( .A(n12393), .ZN(n12381) );
  INV_X1 U10031 ( .A(n12916), .ZN(n13095) );
  AND2_X1 U10032 ( .A1(n9890), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12965) );
  NAND2_X1 U10033 ( .A1(n9702), .A2(n13236), .ZN(n12972) );
  AND2_X1 U10034 ( .A1(n8591), .A2(n8590), .ZN(n8593) );
  INV_X1 U10035 ( .A(n15270), .ZN(n15306) );
  AND2_X1 U10036 ( .A1(n15277), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15305) );
  NAND2_X1 U10037 ( .A1(n9941), .A2(n9940), .ZN(n13264) );
  AND2_X1 U10038 ( .A1(n13252), .A2(n10945), .ZN(n13272) );
  INV_X1 U10039 ( .A(n8631), .ZN(n13284) );
  AND2_X1 U10040 ( .A1(n10145), .A2(n15326), .ZN(n10155) );
  AOI21_X1 U10041 ( .B1(n13414), .B2(n9419), .A(n8690), .ZN(n9697) );
  AND2_X1 U10042 ( .A1(n9663), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9618) );
  AND2_X1 U10043 ( .A1(n10494), .A2(n14052), .ZN(n13772) );
  AND4_X1 U10044 ( .A1(n11535), .A2(n11534), .A3(n11533), .A4(n11532), .ZN(
        n13726) );
  AND2_X1 U10045 ( .A1(n9669), .A2(n9668), .ZN(n9767) );
  INV_X1 U10046 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14731) );
  INV_X1 U10047 ( .A(n15043), .ZN(n15012) );
  INV_X1 U10048 ( .A(n9767), .ZN(n9765) );
  INV_X1 U10049 ( .A(n14199), .ZN(n14260) );
  INV_X1 U10050 ( .A(n10844), .ZN(n15074) );
  NOR2_X1 U10051 ( .A1(n15093), .A2(n14024), .ZN(n15100) );
  INV_X1 U10052 ( .A(n15096), .ZN(n15085) );
  INV_X1 U10053 ( .A(n10248), .ZN(n10768) );
  INV_X1 U10054 ( .A(n15207), .ZN(n14450) );
  OR2_X1 U10055 ( .A1(n14022), .A2(n14265), .ZN(n14795) );
  NAND2_X1 U10056 ( .A1(n9985), .A2(n13863), .ZN(n15196) );
  NAND2_X1 U10057 ( .A1(n10844), .A2(n14795), .ZN(n15207) );
  AND2_X1 U10058 ( .A1(n9986), .A2(n9618), .ZN(n14052) );
  INV_X1 U10059 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9665) );
  AND2_X1 U10060 ( .A1(n9932), .A2(n10050), .ZN(n15013) );
  AND2_X1 U10061 ( .A1(n9454), .A2(n9468), .ZN(n14102) );
  NOR2_X1 U10062 ( .A1(n8510), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14559) );
  AND2_X1 U10063 ( .A1(n10171), .A2(n10170), .ZN(n15535) );
  INV_X1 U10064 ( .A(n11863), .ZN(n11852) );
  INV_X1 U10065 ( .A(n11872), .ZN(n11613) );
  INV_X1 U10066 ( .A(n12443), .ZN(n12094) );
  INV_X1 U10067 ( .A(n15543), .ZN(n15564) );
  NAND2_X1 U10068 ( .A1(n10166), .A2(n10165), .ZN(n15571) );
  NAND2_X1 U10069 ( .A1(n11415), .A2(n14898), .ZN(n12595) );
  AND2_X1 U10070 ( .A1(n12605), .A2(n12604), .ZN(n12712) );
  INV_X2 U10071 ( .A(n14895), .ZN(n12648) );
  INV_X1 U10072 ( .A(n12627), .ZN(n12644) );
  NAND2_X1 U10073 ( .A1(n10581), .A2(n9388), .ZN(n15608) );
  NAND2_X1 U10074 ( .A1(n15611), .A2(n14898), .ZN(n12715) );
  INV_X1 U10075 ( .A(n9301), .ZN(n12731) );
  OR3_X1 U10076 ( .A1(n12705), .A2(n12704), .A3(n12703), .ZN(n12761) );
  INV_X2 U10077 ( .A(n15601), .ZN(n15599) );
  INV_X1 U10078 ( .A(n9724), .ZN(n9889) );
  NAND2_X1 U10079 ( .A1(n9209), .A2(n12772), .ZN(n9724) );
  INV_X1 U10080 ( .A(SI_26_), .ZN(n11401) );
  INV_X1 U10081 ( .A(SI_15_), .ZN(n12360) );
  INV_X1 U10082 ( .A(n14640), .ZN(n14601) );
  NAND2_X1 U10083 ( .A1(n13436), .A2(P3_U3151), .ZN(n12784) );
  INV_X1 U10084 ( .A(n12965), .ZN(n12928) );
  INV_X1 U10085 ( .A(n12972), .ZN(n12957) );
  INV_X1 U10086 ( .A(n8593), .ZN(n12976) );
  CLKBUF_X2 U10087 ( .A(P2_U3947), .Z(n12993) );
  OR2_X1 U10088 ( .A1(n9493), .A2(P2_U3088), .ZN(n15260) );
  INV_X1 U10089 ( .A(n15305), .ZN(n15262) );
  INV_X1 U10090 ( .A(n13272), .ZN(n13206) );
  OR2_X1 U10091 ( .A1(n11594), .A2(n11574), .ZN(n13367) );
  NAND2_X1 U10092 ( .A1(n13252), .A2(n10199), .ZN(n13256) );
  INV_X1 U10093 ( .A(n15392), .ZN(n15390) );
  INV_X1 U10094 ( .A(n15383), .ZN(n15381) );
  NOR2_X1 U10095 ( .A1(n15324), .A2(n15314), .ZN(n15320) );
  NAND2_X1 U10096 ( .A1(n9681), .A2(n9680), .ZN(n15326) );
  INV_X1 U10097 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13410) );
  INV_X1 U10098 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10792) );
  INV_X1 U10099 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9811) );
  AND2_X1 U10100 ( .A1(n10496), .A2(n14055), .ZN(n13780) );
  NAND2_X1 U10101 ( .A1(n13446), .A2(n13445), .ZN(n14326) );
  INV_X1 U10102 ( .A(n13485), .ZN(n14056) );
  INV_X1 U10103 ( .A(n13876), .ZN(n14434) );
  OR2_X1 U10104 ( .A1(n9765), .A2(n14079), .ZN(n15043) );
  INV_X1 U10105 ( .A(n15018), .ZN(n15047) );
  OR2_X1 U10106 ( .A1(n14206), .A2(n13462), .ZN(n15087) );
  OR2_X1 U10107 ( .A1(n15105), .A2(n10845), .ZN(n14418) );
  NAND2_X1 U10108 ( .A1(n14052), .A2(n10770), .ZN(n15080) );
  INV_X1 U10109 ( .A(n15224), .ZN(n15221) );
  AND2_X2 U10110 ( .A1(n9979), .A2(n14052), .ZN(n15136) );
  INV_X1 U10111 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14565) );
  INV_X1 U10112 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13542) );
  INV_X1 U10113 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10573) );
  AND2_X2 U10114 ( .A1(n9421), .A2(n12772), .ZN(P3_U3897) );
  NOR2_X1 U10115 ( .A1(P2_U3088), .A2(n9479), .ZN(P2_U3947) );
  NOR2_X1 U10116 ( .A1(n9986), .A2(n9418), .ZN(P1_U4016) );
  NAND4_X1 U10117 ( .A1(n7889), .A2(n7888), .A3(n7887), .A4(n8289), .ZN(n8312)
         );
  INV_X1 U10118 ( .A(n8312), .ZN(n7897) );
  NAND2_X1 U10119 ( .A1(n7891), .A2(n7890), .ZN(n7892) );
  NOR2_X2 U10120 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7895) );
  NOR2_X2 U10121 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n7894) );
  INV_X1 U10122 ( .A(n7920), .ZN(n7898) );
  NAND3_X1 U10123 ( .A1(n7898), .A2(n7917), .A3(n7916), .ZN(n7901) );
  NOR2_X1 U10124 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n7900) );
  NOR2_X1 U10125 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n7899) );
  NAND3_X1 U10126 ( .A1(n7934), .A2(n7900), .A3(n7899), .ZN(n7914) );
  XNOR2_X2 U10127 ( .A(n7904), .B(n7903), .ZN(n7907) );
  INV_X1 U10128 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7908) );
  INV_X1 U10129 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U10130 ( .A1(n8510), .A2(SI_0_), .ZN(n7913) );
  XNOR2_X1 U10131 ( .A(n7913), .B(n8742), .ZN(n13418) );
  INV_X1 U10132 ( .A(n15229), .ZN(n9518) );
  NAND2_X1 U10133 ( .A1(n7918), .A2(n7917), .ZN(n8683) );
  AOI21_X2 U10134 ( .B1(n8683), .B2(n7922), .A(n7921), .ZN(n7923) );
  NAND3_X1 U10135 ( .A1(n7929), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .ZN(n7933) );
  NAND2_X1 U10136 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n7930) );
  NAND2_X1 U10137 ( .A1(n7930), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7931) );
  OAI21_X1 U10138 ( .B1(n12329), .B2(P2_IR_REG_31__SCAN_IN), .A(n7931), .ZN(
        n7932) );
  NAND2_X1 U10139 ( .A1(n7934), .A2(n8674), .ZN(n7939) );
  NAND3_X1 U10140 ( .A1(n7940), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_22__SCAN_IN), .ZN(n7938) );
  INV_X1 U10141 ( .A(n7934), .ZN(n7936) );
  XNOR2_X1 U10142 ( .A(P2_IR_REG_22__SCAN_IN), .B(P2_IR_REG_31__SCAN_IN), .ZN(
        n7935) );
  OAI21_X1 U10143 ( .B1(n7936), .B2(n8674), .A(n7935), .ZN(n7937) );
  NAND2_X1 U10144 ( .A1(n8649), .A2(n8592), .ZN(n7943) );
  NAND2_X1 U10145 ( .A1(n10129), .A2(n9712), .ZN(n7942) );
  OAI211_X1 U10146 ( .C1(n10129), .C2(n9712), .A(n8648), .B(n8635), .ZN(n7941)
         );
  OAI21_X1 U10147 ( .B1(SI_1_), .B2(n7944), .A(n7957), .ZN(n7948) );
  INV_X1 U10148 ( .A(n7948), .ZN(n7945) );
  INV_X1 U10149 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8780) );
  INV_X1 U10150 ( .A(SI_0_), .ZN(n9962) );
  INV_X1 U10151 ( .A(n7946), .ZN(n7947) );
  NAND2_X1 U10152 ( .A1(n7948), .A2(n7947), .ZN(n7949) );
  NAND2_X1 U10153 ( .A1(n7958), .A2(n7949), .ZN(n10021) );
  NAND2_X1 U10154 ( .A1(n8561), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U10155 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n15229), .ZN(n7950) );
  XNOR2_X1 U10156 ( .A(n7950), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U10157 ( .A1(n8334), .A2(n9515), .ZN(n7951) );
  NAND2_X1 U10158 ( .A1(n7996), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7956) );
  NAND2_X1 U10159 ( .A1(n8564), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7953) );
  AOI22_X1 U10160 ( .A1(n6574), .A2(n8635), .B1(n12994), .B2(n8592), .ZN(n7979) );
  NAND2_X1 U10161 ( .A1(n7958), .A2(n7957), .ZN(n7961) );
  MUX2_X1 U10162 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n13436), .Z(n7959) );
  NAND2_X1 U10163 ( .A1(n7959), .A2(SI_2_), .ZN(n7987) );
  OAI21_X1 U10164 ( .B1(n7959), .B2(SI_2_), .A(n7987), .ZN(n7962) );
  INV_X1 U10165 ( .A(n7962), .ZN(n7960) );
  NAND2_X1 U10166 ( .A1(n7963), .A2(n7962), .ZN(n7964) );
  AND2_X1 U10167 ( .A1(n7988), .A2(n7964), .ZN(n10071) );
  NAND2_X1 U10168 ( .A1(n10071), .A2(n7965), .ZN(n7969) );
  OR2_X1 U10169 ( .A1(n7966), .A2(n7991), .ZN(n7967) );
  XNOR2_X1 U10170 ( .A(n7967), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9531) );
  NAND2_X1 U10171 ( .A1(n6603), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U10172 ( .A1(n8160), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U10173 ( .A1(n7996), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U10174 ( .A1(n8564), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U10175 ( .A1(n12992), .A2(n8592), .ZN(n7974) );
  NAND2_X1 U10176 ( .A1(n7975), .A2(n7974), .ZN(n7981) );
  NAND2_X1 U10177 ( .A1(n7981), .A2(n7982), .ZN(n7978) );
  OAI211_X1 U10178 ( .C1(n7980), .C2(n7979), .A(n7978), .B(n7977), .ZN(n7986)
         );
  INV_X1 U10179 ( .A(n7981), .ZN(n7984) );
  INV_X1 U10180 ( .A(n7982), .ZN(n7983) );
  NAND2_X1 U10181 ( .A1(n7984), .A2(n7983), .ZN(n7985) );
  MUX2_X1 U10182 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n13436), .Z(n7989) );
  NAND2_X1 U10183 ( .A1(n7989), .A2(SI_3_), .ZN(n8011) );
  OAI21_X1 U10184 ( .B1(n7989), .B2(SI_3_), .A(n8011), .ZN(n8009) );
  NAND2_X1 U10185 ( .A1(n10215), .A2(n8532), .ZN(n7995) );
  NOR2_X1 U10186 ( .A1(n8179), .A2(n7991), .ZN(n7990) );
  MUX2_X1 U10187 ( .A(n7991), .B(n7990), .S(P2_IR_REG_3__SCAN_IN), .Z(n7993)
         );
  AND2_X1 U10188 ( .A1(n8179), .A2(n7992), .ZN(n8013) );
  NOR2_X1 U10189 ( .A1(n7993), .A2(n8013), .ZN(n9562) );
  AOI22_X1 U10190 ( .A1(n8561), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n9562), .B2(
        n8334), .ZN(n7994) );
  INV_X4 U10191 ( .A(n8635), .ZN(n8615) );
  NAND2_X1 U10192 ( .A1(n15348), .A2(n8615), .ZN(n8003) );
  OR2_X1 U10193 ( .A1(n8585), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8001) );
  NAND2_X1 U10194 ( .A1(n7996), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10195 ( .A1(n8586), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U10196 ( .A1(n8564), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U10197 ( .A1(n12991), .A2(n8617), .ZN(n8002) );
  NOR2_X1 U10198 ( .A1(n8007), .A2(n8006), .ZN(n8004) );
  AOI22_X1 U10199 ( .A1(n15348), .A2(n8617), .B1(n8615), .B2(n12991), .ZN(
        n8005) );
  INV_X1 U10200 ( .A(n8009), .ZN(n8010) );
  MUX2_X1 U10201 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n13436), .Z(n8012) );
  NAND2_X1 U10202 ( .A1(n8012), .A2(SI_4_), .ZN(n8026) );
  OAI21_X1 U10203 ( .B1(n8012), .B2(SI_4_), .A(n8026), .ZN(n8023) );
  XNOR2_X1 U10204 ( .A(n8025), .B(n8023), .ZN(n10216) );
  NAND2_X1 U10205 ( .A1(n10216), .A2(n8532), .ZN(n8016) );
  INV_X1 U10206 ( .A(n8013), .ZN(n8032) );
  NAND2_X1 U10207 ( .A1(n8032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8014) );
  XNOR2_X1 U10208 ( .A(n8014), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9599) );
  AOI22_X1 U10209 ( .A1(n8561), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9599), .B2(
        n8334), .ZN(n8015) );
  NAND2_X1 U10210 ( .A1(n8016), .A2(n8015), .ZN(n10115) );
  NAND2_X1 U10211 ( .A1(n10115), .A2(n8617), .ZN(n8022) );
  AND2_X1 U10212 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8036) );
  INV_X1 U10213 ( .A(n8036), .ZN(n8038) );
  OAI21_X1 U10214 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8038), .ZN(n10441) );
  OR2_X1 U10215 ( .A1(n8585), .A2(n10441), .ZN(n8020) );
  NAND2_X1 U10216 ( .A1(n8564), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U10217 ( .A1(n7996), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U10218 ( .A1(n8586), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8017) );
  NAND2_X1 U10219 ( .A1(n8022), .A2(n7881), .ZN(n8048) );
  INV_X1 U10220 ( .A(n8023), .ZN(n8024) );
  MUX2_X1 U10221 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6568), .Z(n8027) );
  NAND2_X1 U10222 ( .A1(n8027), .A2(SI_5_), .ZN(n8052) );
  OAI21_X1 U10223 ( .B1(n8027), .B2(SI_5_), .A(n8052), .ZN(n8028) );
  INV_X1 U10224 ( .A(n8028), .ZN(n8029) );
  OR2_X1 U10225 ( .A1(n8030), .A2(n8029), .ZN(n8031) );
  NAND2_X1 U10226 ( .A1(n8053), .A2(n8031), .ZN(n9461) );
  OR2_X1 U10227 ( .A1(n9461), .A2(n8611), .ZN(n8035) );
  INV_X1 U10228 ( .A(n8561), .ZN(n8610) );
  INV_X2 U10229 ( .A(n8610), .ZN(n8361) );
  NAND2_X1 U10230 ( .A1(n8055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8033) );
  XNOR2_X1 U10231 ( .A(n8033), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9583) );
  AOI22_X1 U10232 ( .A1(n8361), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9583), .B2(
        n8334), .ZN(n8034) );
  NAND2_X2 U10233 ( .A1(n8035), .A2(n8034), .ZN(n10300) );
  NAND2_X1 U10234 ( .A1(n8036), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8067) );
  INV_X1 U10235 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U10236 ( .A1(n8038), .A2(n8037), .ZN(n8039) );
  NAND2_X1 U10237 ( .A1(n8067), .A2(n8039), .ZN(n10134) );
  OR2_X1 U10238 ( .A1(n8585), .A2(n10134), .ZN(n8043) );
  NAND2_X1 U10239 ( .A1(n8564), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8042) );
  NAND2_X1 U10240 ( .A1(n7996), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8041) );
  NAND2_X1 U10241 ( .A1(n8586), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8040) );
  NAND4_X1 U10242 ( .A1(n8043), .A2(n8042), .A3(n8041), .A4(n8040), .ZN(n12989) );
  AND2_X1 U10243 ( .A1(n12989), .A2(n8617), .ZN(n8044) );
  AOI21_X1 U10244 ( .B1(n10300), .B2(n8615), .A(n8044), .ZN(n8050) );
  NAND2_X1 U10245 ( .A1(n10300), .A2(n8617), .ZN(n8046) );
  NAND2_X1 U10246 ( .A1(n12989), .A2(n8615), .ZN(n8045) );
  NAND2_X1 U10247 ( .A1(n8046), .A2(n8045), .ZN(n8049) );
  AOI22_X1 U10248 ( .A1(n10115), .A2(n8615), .B1(n12990), .B2(n8616), .ZN(
        n8047) );
  NAND2_X1 U10249 ( .A1(n8050), .A2(n8049), .ZN(n8051) );
  NAND2_X1 U10250 ( .A1(n8053), .A2(n8052), .ZN(n8077) );
  MUX2_X1 U10251 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n8510), .Z(n8054) );
  NAND2_X1 U10252 ( .A1(n8054), .A2(SI_6_), .ZN(n8078) );
  OAI21_X1 U10253 ( .B1(SI_6_), .B2(n8054), .A(n8078), .ZN(n8075) );
  XNOR2_X1 U10254 ( .A(n8077), .B(n8075), .ZN(n10852) );
  NAND2_X1 U10255 ( .A1(n10852), .A2(n8532), .ZN(n8064) );
  INV_X1 U10256 ( .A(n8055), .ZN(n8057) );
  NAND2_X1 U10257 ( .A1(n8057), .A2(n8056), .ZN(n8059) );
  NAND2_X1 U10258 ( .A1(n8059), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8058) );
  MUX2_X1 U10259 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8058), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n8062) );
  INV_X1 U10260 ( .A(n8059), .ZN(n8061) );
  INV_X1 U10261 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U10262 ( .A1(n8061), .A2(n8060), .ZN(n8085) );
  AOI22_X1 U10263 ( .A1(n8361), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9634), .B2(
        n9476), .ZN(n8063) );
  NAND2_X1 U10264 ( .A1(n15365), .A2(n8616), .ZN(n8073) );
  INV_X1 U10265 ( .A(n8067), .ZN(n8065) );
  NAND2_X1 U10266 ( .A1(n8065), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8090) );
  INV_X1 U10267 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8066) );
  NAND2_X1 U10268 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  NAND2_X1 U10269 ( .A1(n8090), .A2(n8068), .ZN(n10323) );
  OR2_X1 U10270 ( .A1(n8585), .A2(n10323), .ZN(n8071) );
  NAND2_X1 U10271 ( .A1(n7996), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8070) );
  NAND2_X1 U10272 ( .A1(n8586), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U10273 ( .A1(n12988), .A2(n8615), .ZN(n8072) );
  NAND2_X1 U10274 ( .A1(n8073), .A2(n8072), .ZN(n8074) );
  INV_X1 U10275 ( .A(n8075), .ZN(n8076) );
  MUX2_X1 U10276 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6568), .Z(n8079) );
  NAND2_X1 U10277 ( .A1(n8079), .A2(SI_7_), .ZN(n8108) );
  OAI21_X1 U10278 ( .B1(n8079), .B2(SI_7_), .A(n8108), .ZN(n8080) );
  OR2_X1 U10279 ( .A1(n8082), .A2(n8081), .ZN(n8083) );
  NAND2_X1 U10280 ( .A1(n8085), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8084) );
  MUX2_X1 U10281 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8084), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n8086) );
  AOI22_X1 U10282 ( .A1(n8361), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n15232), 
        .B2(n9476), .ZN(n8087) );
  NAND2_X1 U10283 ( .A1(n10564), .A2(n8615), .ZN(n8098) );
  INV_X1 U10284 ( .A(n8090), .ZN(n8088) );
  NAND2_X1 U10285 ( .A1(n8088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8120) );
  INV_X1 U10286 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10287 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  NAND2_X1 U10288 ( .A1(n8120), .A2(n8091), .ZN(n10296) );
  OR2_X1 U10289 ( .A1(n8585), .A2(n10296), .ZN(n8096) );
  NAND2_X1 U10290 ( .A1(n8564), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U10291 ( .A1(n6571), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10292 ( .A1(n8586), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8093) );
  NAND4_X1 U10293 ( .A1(n8096), .A2(n8095), .A3(n8094), .A4(n8093), .ZN(n12987) );
  NAND2_X1 U10294 ( .A1(n12987), .A2(n8616), .ZN(n8097) );
  NAND2_X1 U10295 ( .A1(n8098), .A2(n8097), .ZN(n8104) );
  NAND2_X1 U10296 ( .A1(n10564), .A2(n8616), .ZN(n8100) );
  NAND2_X1 U10297 ( .A1(n12987), .A2(n8615), .ZN(n8099) );
  NAND2_X1 U10298 ( .A1(n8100), .A2(n8099), .ZN(n8101) );
  NAND2_X1 U10299 ( .A1(n8102), .A2(n8101), .ZN(n8107) );
  INV_X1 U10300 ( .A(n8103), .ZN(n8106) );
  INV_X1 U10301 ( .A(n8104), .ZN(n8105) );
  MUX2_X1 U10302 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n8510), .Z(n8110) );
  NAND2_X1 U10303 ( .A1(n8110), .A2(SI_8_), .ZN(n8129) );
  OAI21_X1 U10304 ( .B1(SI_8_), .B2(n8110), .A(n8129), .ZN(n8111) );
  INV_X1 U10305 ( .A(n8111), .ZN(n8112) );
  OR2_X1 U10306 ( .A1(n8113), .A2(n8112), .ZN(n8114) );
  NAND2_X1 U10307 ( .A1(n8116), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8115) );
  MUX2_X1 U10308 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8115), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8117) );
  NAND2_X1 U10309 ( .A1(n8117), .A2(n8156), .ZN(n13001) );
  INV_X1 U10310 ( .A(n13001), .ZN(n9640) );
  AOI22_X1 U10311 ( .A1(n9640), .A2(n9476), .B1(n8361), .B2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n8118) );
  NAND2_X1 U10312 ( .A1(n10647), .A2(n8616), .ZN(n8127) );
  NAND2_X1 U10313 ( .A1(n8120), .A2(n10633), .ZN(n8121) );
  NAND2_X1 U10314 ( .A1(n8141), .A2(n8121), .ZN(n10636) );
  OR2_X1 U10315 ( .A1(n8585), .A2(n10636), .ZN(n8125) );
  NAND2_X1 U10316 ( .A1(n6571), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8124) );
  NAND2_X1 U10317 ( .A1(n8586), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U10318 ( .A1(n8564), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8122) );
  NAND4_X1 U10319 ( .A1(n8125), .A2(n8124), .A3(n8123), .A4(n8122), .ZN(n12986) );
  NAND2_X1 U10320 ( .A1(n12986), .A2(n8615), .ZN(n8126) );
  NAND2_X1 U10321 ( .A1(n8127), .A2(n8126), .ZN(n8128) );
  MUX2_X1 U10322 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n8510), .Z(n8131) );
  NAND2_X1 U10323 ( .A1(n8131), .A2(SI_9_), .ZN(n8153) );
  OAI21_X1 U10324 ( .B1(n8131), .B2(SI_9_), .A(n8153), .ZN(n8132) );
  INV_X1 U10325 ( .A(n8132), .ZN(n8133) );
  NAND2_X1 U10326 ( .A1(n8134), .A2(n8133), .ZN(n8154) );
  OR2_X1 U10327 ( .A1(n8134), .A2(n8133), .ZN(n8135) );
  NAND2_X1 U10328 ( .A1(n8154), .A2(n8135), .ZN(n11035) );
  OR2_X1 U10329 ( .A1(n11035), .A2(n8611), .ZN(n8138) );
  NAND2_X1 U10330 ( .A1(n8156), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8136) );
  XNOR2_X1 U10331 ( .A(n8136), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9650) );
  AOI22_X1 U10332 ( .A1(n9650), .A2(n9476), .B1(n8361), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U10333 ( .A1(n10745), .A2(n8615), .ZN(n8148) );
  INV_X1 U10334 ( .A(n8141), .ZN(n8139) );
  NAND2_X1 U10335 ( .A1(n8139), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8185) );
  INV_X1 U10336 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U10337 ( .A1(n8141), .A2(n8140), .ZN(n8142) );
  NAND2_X1 U10338 ( .A1(n8185), .A2(n8142), .ZN(n10623) );
  OR2_X1 U10339 ( .A1(n8585), .A2(n10623), .ZN(n8146) );
  NAND2_X1 U10340 ( .A1(n6571), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U10341 ( .A1(n8586), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8144) );
  NAND2_X1 U10342 ( .A1(n8564), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8143) );
  NAND4_X1 U10343 ( .A1(n8146), .A2(n8145), .A3(n8144), .A4(n8143), .ZN(n12985) );
  NAND2_X1 U10344 ( .A1(n12985), .A2(n8617), .ZN(n8147) );
  NAND2_X1 U10345 ( .A1(n8148), .A2(n8147), .ZN(n8152) );
  NAND2_X1 U10346 ( .A1(n10745), .A2(n8617), .ZN(n8150) );
  NAND2_X1 U10347 ( .A1(n12985), .A2(n8615), .ZN(n8149) );
  MUX2_X1 U10348 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8510), .Z(n8155) );
  NAND2_X1 U10349 ( .A1(n8155), .A2(SI_10_), .ZN(n8175) );
  OAI21_X1 U10350 ( .B1(n8155), .B2(SI_10_), .A(n8175), .ZN(n8172) );
  XNOR2_X1 U10351 ( .A(n8174), .B(n8172), .ZN(n11141) );
  NAND2_X1 U10352 ( .A1(n11141), .A2(n8532), .ZN(n8159) );
  OAI21_X1 U10353 ( .B1(n8156), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8157) );
  XNOR2_X1 U10354 ( .A(n8157), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9817) );
  AOI22_X1 U10355 ( .A1(n9817), .A2(n9476), .B1(P1_DATAO_REG_10__SCAN_IN), 
        .B2(n8361), .ZN(n8158) );
  NAND2_X1 U10356 ( .A1(n11003), .A2(n8616), .ZN(n8166) );
  NAND2_X1 U10357 ( .A1(n8564), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10358 ( .A1(n6571), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8163) );
  XNOR2_X1 U10359 ( .A(n8185), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n10752) );
  NAND2_X1 U10360 ( .A1(n8160), .A2(n10752), .ZN(n8162) );
  NAND2_X1 U10361 ( .A1(n8586), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8161) );
  NAND4_X1 U10362 ( .A1(n8164), .A2(n8163), .A3(n8162), .A4(n8161), .ZN(n12984) );
  NAND2_X1 U10363 ( .A1(n12984), .A2(n8615), .ZN(n8165) );
  NAND2_X1 U10364 ( .A1(n8166), .A2(n8165), .ZN(n8168) );
  AOI22_X1 U10365 ( .A1(n11003), .A2(n8615), .B1(n12984), .B2(n8617), .ZN(
        n8167) );
  NOR2_X1 U10366 ( .A1(n8169), .A2(n8168), .ZN(n8170) );
  INV_X1 U10367 ( .A(n8172), .ZN(n8173) );
  MUX2_X1 U10368 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n8510), .Z(n8197) );
  XNOR2_X1 U10369 ( .A(n8197), .B(SI_11_), .ZN(n8199) );
  XNOR2_X1 U10370 ( .A(n8200), .B(n8199), .ZN(n11148) );
  NAND2_X1 U10371 ( .A1(n11148), .A2(n8532), .ZN(n8182) );
  INV_X1 U10372 ( .A(n8176), .ZN(n8177) );
  NAND3_X1 U10373 ( .A1(n8179), .A2(n8178), .A3(n8177), .ZN(n8313) );
  NAND2_X1 U10374 ( .A1(n8313), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8180) );
  XNOR2_X1 U10375 ( .A(n8180), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U10376 ( .A1(n8361), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n10806), 
        .B2(n9476), .ZN(n8181) );
  NAND2_X1 U10377 ( .A1(n11066), .A2(n8615), .ZN(n8192) );
  INV_X1 U10378 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9740) );
  INV_X1 U10379 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8183) );
  OAI21_X1 U10380 ( .B1(n8185), .B2(n9740), .A(n8183), .ZN(n8186) );
  NAND2_X1 U10381 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n8184) );
  NAND2_X1 U10382 ( .A1(n8186), .A2(n8209), .ZN(n10996) );
  OR2_X1 U10383 ( .A1(n8585), .A2(n10996), .ZN(n8190) );
  NAND2_X1 U10384 ( .A1(n6571), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U10385 ( .A1(n8586), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8188) );
  NAND2_X1 U10386 ( .A1(n8564), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8187) );
  NAND4_X1 U10387 ( .A1(n8190), .A2(n8189), .A3(n8188), .A4(n8187), .ZN(n12983) );
  NAND2_X1 U10388 ( .A1(n12983), .A2(n8617), .ZN(n8191) );
  NAND2_X1 U10389 ( .A1(n8192), .A2(n8191), .ZN(n8196) );
  NAND2_X1 U10390 ( .A1(n11066), .A2(n8617), .ZN(n8194) );
  NAND2_X1 U10391 ( .A1(n12983), .A2(n8615), .ZN(n8193) );
  NAND2_X1 U10392 ( .A1(n8194), .A2(n8193), .ZN(n8195) );
  INV_X1 U10393 ( .A(n8197), .ZN(n8198) );
  MUX2_X1 U10394 ( .A(n9933), .B(n9927), .S(n6568), .Z(n8222) );
  XNOR2_X1 U10395 ( .A(n8222), .B(SI_12_), .ZN(n8220) );
  XNOR2_X1 U10396 ( .A(n8221), .B(n8220), .ZN(n11232) );
  NAND2_X1 U10397 ( .A1(n11232), .A2(n8532), .ZN(n8206) );
  OR2_X1 U10398 ( .A1(n8313), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U10399 ( .A1(n8203), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8201) );
  MUX2_X1 U10400 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8201), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8202) );
  INV_X1 U10401 ( .A(n8202), .ZN(n8204) );
  NOR2_X1 U10402 ( .A1(n8204), .A2(n8226), .ZN(n10810) );
  AOI22_X1 U10403 ( .A1(n8361), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n10810), 
        .B2(n9476), .ZN(n8205) );
  NAND2_X1 U10404 ( .A1(n11195), .A2(n8617), .ZN(n8216) );
  INV_X1 U10405 ( .A(n8209), .ZN(n8207) );
  INV_X1 U10406 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8208) );
  NAND2_X1 U10407 ( .A1(n8209), .A2(n8208), .ZN(n8210) );
  NAND2_X1 U10408 ( .A1(n8248), .A2(n8210), .ZN(n11071) );
  OR2_X1 U10409 ( .A1(n8585), .A2(n11071), .ZN(n8214) );
  NAND2_X1 U10410 ( .A1(n8564), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8213) );
  NAND2_X1 U10411 ( .A1(n6571), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U10412 ( .A1(n8586), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8211) );
  NAND4_X1 U10413 ( .A1(n8214), .A2(n8213), .A3(n8212), .A4(n8211), .ZN(n12982) );
  NAND2_X1 U10414 ( .A1(n12982), .A2(n8615), .ZN(n8215) );
  NAND2_X1 U10415 ( .A1(n8216), .A2(n8215), .ZN(n8218) );
  AOI22_X1 U10416 ( .A1(n11195), .A2(n8615), .B1(n12982), .B2(n8617), .ZN(
        n8217) );
  MUX2_X1 U10417 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n13436), .Z(n8241) );
  XNOR2_X1 U10418 ( .A(n8241), .B(n9614), .ZN(n8239) );
  XNOR2_X1 U10419 ( .A(n8240), .B(n8239), .ZN(n11422) );
  NAND2_X1 U10420 ( .A1(n11422), .A2(n8400), .ZN(n8229) );
  INV_X1 U10421 ( .A(n8226), .ZN(n8223) );
  NAND2_X1 U10422 ( .A1(n8223), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8224) );
  MUX2_X1 U10423 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8224), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8227) );
  INV_X1 U10424 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U10425 ( .A1(n8226), .A2(n8225), .ZN(n8265) );
  NAND2_X1 U10426 ( .A1(n8227), .A2(n8265), .ZN(n15261) );
  INV_X1 U10427 ( .A(n15261), .ZN(n10811) );
  AOI22_X1 U10428 ( .A1(n8361), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n10811), 
        .B2(n8334), .ZN(n8228) );
  NAND2_X1 U10429 ( .A1(n13374), .A2(n8615), .ZN(n8235) );
  XNOR2_X1 U10430 ( .A(n8248), .B(P2_REG3_REG_13__SCAN_IN), .ZN(n11228) );
  NAND2_X1 U10431 ( .A1(n11228), .A2(n8160), .ZN(n8233) );
  NAND2_X1 U10432 ( .A1(n8564), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8232) );
  NAND2_X1 U10433 ( .A1(n6571), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8231) );
  NAND2_X1 U10434 ( .A1(n8586), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8230) );
  NAND4_X1 U10435 ( .A1(n8233), .A2(n8232), .A3(n8231), .A4(n8230), .ZN(n12981) );
  NAND2_X1 U10436 ( .A1(n12981), .A2(n8617), .ZN(n8234) );
  NAND2_X1 U10437 ( .A1(n8235), .A2(n8234), .ZN(n8237) );
  AOI22_X1 U10438 ( .A1(n13374), .A2(n8617), .B1(n8615), .B2(n12981), .ZN(
        n8236) );
  INV_X1 U10439 ( .A(n8241), .ZN(n8242) );
  NAND2_X1 U10440 ( .A1(n8242), .A2(n9614), .ZN(n8243) );
  MUX2_X1 U10441 ( .A(n10342), .B(n12254), .S(n13436), .Z(n8260) );
  XNOR2_X1 U10442 ( .A(n8259), .B(n8260), .ZN(n11514) );
  NAND2_X1 U10443 ( .A1(n11514), .A2(n8400), .ZN(n8247) );
  NAND2_X1 U10444 ( .A1(n8265), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8245) );
  XNOR2_X1 U10445 ( .A(n8245), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U10446 ( .A1(n8361), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n10812), 
        .B2(n9476), .ZN(n8246) );
  NAND2_X1 U10447 ( .A1(n11505), .A2(n8616), .ZN(n8256) );
  INV_X1 U10448 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8254) );
  OAI21_X1 U10449 ( .B1(n8248), .B2(n11225), .A(n11321), .ZN(n8249) );
  AND2_X1 U10450 ( .A1(n8249), .A2(n8271), .ZN(n11324) );
  NAND2_X1 U10451 ( .A1(n11324), .A2(n8160), .ZN(n8253) );
  NAND2_X1 U10452 ( .A1(n8564), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8251) );
  NAND2_X1 U10453 ( .A1(n6571), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8250) );
  AND2_X1 U10454 ( .A1(n8251), .A2(n8250), .ZN(n8252) );
  OAI211_X1 U10455 ( .C1(n8614), .C2(n8254), .A(n8253), .B(n8252), .ZN(n12980)
         );
  NAND2_X1 U10456 ( .A1(n12980), .A2(n8615), .ZN(n8255) );
  INV_X1 U10457 ( .A(n12980), .ZN(n11499) );
  NAND2_X1 U10458 ( .A1(n11505), .A2(n8615), .ZN(n8257) );
  OAI21_X1 U10459 ( .B1(n11499), .B2(n8592), .A(n8257), .ZN(n8258) );
  INV_X1 U10460 ( .A(n8283), .ZN(n8261) );
  OAI22_X1 U10461 ( .A1(n8262), .A2(n8284), .B1(n8261), .B2(SI_14_), .ZN(n8264) );
  MUX2_X1 U10462 ( .A(n10573), .B(n10572), .S(n13436), .Z(n8285) );
  XNOR2_X1 U10463 ( .A(n8285), .B(SI_15_), .ZN(n8263) );
  XNOR2_X1 U10464 ( .A(n8264), .B(n8263), .ZN(n11616) );
  NAND2_X1 U10465 ( .A1(n11616), .A2(n8400), .ZN(n8268) );
  OR2_X1 U10466 ( .A1(n8265), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U10467 ( .A1(n8266), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8290) );
  XNOR2_X1 U10468 ( .A(n8290), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15290) );
  AOI22_X1 U10469 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n8361), .B1(n15290), 
        .B2(n8334), .ZN(n8267) );
  NAND2_X1 U10470 ( .A1(n13369), .A2(n8615), .ZN(n8277) );
  INV_X1 U10471 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8275) );
  INV_X1 U10472 ( .A(n8271), .ZN(n8269) );
  NAND2_X1 U10473 ( .A1(n8269), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8297) );
  INV_X1 U10474 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8270) );
  NAND2_X1 U10475 ( .A1(n8271), .A2(n8270), .ZN(n8272) );
  NAND2_X1 U10476 ( .A1(n8297), .A2(n8272), .ZN(n11554) );
  OR2_X1 U10477 ( .A1(n11554), .A2(n8585), .ZN(n8274) );
  AOI22_X1 U10478 ( .A1(n8564), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n6571), .B2(
        P2_REG0_REG_15__SCAN_IN), .ZN(n8273) );
  OAI211_X1 U10479 ( .C1(n8614), .C2(n8275), .A(n8274), .B(n8273), .ZN(n12979)
         );
  NAND2_X1 U10480 ( .A1(n12979), .A2(n8616), .ZN(n8276) );
  NAND2_X1 U10481 ( .A1(n8277), .A2(n8276), .ZN(n8279) );
  AOI22_X1 U10482 ( .A1(n13369), .A2(n8617), .B1(n8615), .B2(n12979), .ZN(
        n8278) );
  INV_X1 U10483 ( .A(n8285), .ZN(n8281) );
  NAND2_X1 U10484 ( .A1(n8281), .A2(SI_15_), .ZN(n8286) );
  NAND2_X1 U10485 ( .A1(n8284), .A2(SI_14_), .ZN(n8282) );
  NOR2_X1 U10486 ( .A1(n8284), .A2(SI_14_), .ZN(n8287) );
  AOI22_X1 U10487 ( .A1(n8287), .A2(n8286), .B1(n12360), .B2(n8285), .ZN(n8288) );
  MUX2_X1 U10488 ( .A(n10340), .B(n10331), .S(n8510), .Z(n8310) );
  XNOR2_X1 U10489 ( .A(n8310), .B(SI_16_), .ZN(n8307) );
  XNOR2_X1 U10490 ( .A(n8308), .B(n8307), .ZN(n13495) );
  NAND2_X1 U10491 ( .A1(n13495), .A2(n8400), .ZN(n8294) );
  NAND2_X1 U10492 ( .A1(n8290), .A2(n8289), .ZN(n8291) );
  NAND2_X1 U10493 ( .A1(n8291), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8292) );
  XNOR2_X1 U10494 ( .A(n8292), .B(P2_IR_REG_16__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U10495 ( .A1(n10803), .A2(n8334), .B1(n8361), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U10496 ( .A1(n13364), .A2(n8617), .ZN(n8302) );
  INV_X1 U10497 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11586) );
  INV_X1 U10498 ( .A(n8297), .ZN(n8295) );
  NAND2_X1 U10499 ( .A1(n8295), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8317) );
  INV_X1 U10500 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U10501 ( .A1(n8297), .A2(n8296), .ZN(n8298) );
  NAND2_X1 U10502 ( .A1(n8317), .A2(n8298), .ZN(n12898) );
  OR2_X1 U10503 ( .A1(n12898), .A2(n8585), .ZN(n8300) );
  AOI22_X1 U10504 ( .A1(n8564), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n6571), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n8299) );
  OAI211_X1 U10505 ( .C1(n8614), .C2(n11586), .A(n8300), .B(n8299), .ZN(n12978) );
  NAND2_X1 U10506 ( .A1(n12978), .A2(n8615), .ZN(n8301) );
  INV_X1 U10507 ( .A(n12978), .ZN(n12908) );
  NAND2_X1 U10508 ( .A1(n13364), .A2(n8615), .ZN(n8303) );
  OAI21_X1 U10509 ( .B1(n12908), .B2(n8592), .A(n8303), .ZN(n8304) );
  MUX2_X1 U10510 ( .A(n12347), .B(n10466), .S(n13436), .Z(n8329) );
  XNOR2_X1 U10511 ( .A(n8329), .B(SI_17_), .ZN(n8311) );
  XNOR2_X1 U10512 ( .A(n8331), .B(n8311), .ZN(n13507) );
  NAND2_X1 U10513 ( .A1(n13507), .A2(n8400), .ZN(n8316) );
  OR2_X1 U10514 ( .A1(n8313), .A2(n8312), .ZN(n8332) );
  NAND2_X1 U10515 ( .A1(n8332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8314) );
  XNOR2_X1 U10516 ( .A(n8314), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U10517 ( .A1(n8361), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n15304), 
        .B2(n9476), .ZN(n8315) );
  NAND2_X1 U10518 ( .A1(n13069), .A2(n8615), .ZN(n8325) );
  NAND2_X1 U10519 ( .A1(n8317), .A2(n12902), .ZN(n8318) );
  AND2_X1 U10520 ( .A1(n8338), .A2(n8318), .ZN(n12906) );
  NAND2_X1 U10521 ( .A1(n12906), .A2(n8160), .ZN(n8323) );
  INV_X1 U10522 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11343) );
  NAND2_X1 U10523 ( .A1(n8586), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8320) );
  NAND2_X1 U10524 ( .A1(n6571), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8319) );
  OAI211_X1 U10525 ( .C1(n7997), .C2(n11343), .A(n8320), .B(n8319), .ZN(n8321)
         );
  INV_X1 U10526 ( .A(n8321), .ZN(n8322) );
  NAND2_X1 U10527 ( .A1(n8323), .A2(n8322), .ZN(n13065) );
  NAND2_X1 U10528 ( .A1(n13065), .A2(n8617), .ZN(n8324) );
  NAND2_X1 U10529 ( .A1(n8325), .A2(n8324), .ZN(n8327) );
  AOI22_X1 U10530 ( .A1(n13069), .A2(n8617), .B1(n8615), .B2(n13065), .ZN(
        n8326) );
  MUX2_X1 U10531 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n8510), .Z(n8354) );
  XNOR2_X1 U10532 ( .A(n8353), .B(n8354), .ZN(n13522) );
  NAND2_X1 U10533 ( .A1(n13522), .A2(n8400), .ZN(n8336) );
  OAI21_X1 U10534 ( .B1(n8332), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8333) );
  XNOR2_X1 U10535 ( .A(n8333), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U10536 ( .A1(n8361), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n13014), 
        .B2(n8334), .ZN(n8335) );
  NAND2_X1 U10537 ( .A1(n13353), .A2(n8617), .ZN(n8347) );
  INV_X1 U10538 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n12953) );
  NAND2_X1 U10539 ( .A1(n8338), .A2(n12953), .ZN(n8339) );
  NAND2_X1 U10540 ( .A1(n8365), .A2(n8339), .ZN(n12952) );
  OR2_X1 U10541 ( .A1(n12952), .A2(n8585), .ZN(n8345) );
  INV_X1 U10542 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U10543 ( .A1(n8564), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U10544 ( .A1(n6571), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8340) );
  OAI211_X1 U10545 ( .C1(n8342), .C2(n8614), .A(n8341), .B(n8340), .ZN(n8343)
         );
  INV_X1 U10546 ( .A(n8343), .ZN(n8344) );
  NAND2_X1 U10547 ( .A1(n8345), .A2(n8344), .ZN(n13042) );
  NAND2_X1 U10548 ( .A1(n13042), .A2(n8615), .ZN(n8346) );
  NAND2_X1 U10549 ( .A1(n8347), .A2(n8346), .ZN(n8350) );
  INV_X1 U10550 ( .A(n13042), .ZN(n13071) );
  NAND2_X1 U10551 ( .A1(n13353), .A2(n8615), .ZN(n8348) );
  OAI21_X1 U10552 ( .B1(n13071), .B2(n8592), .A(n8348), .ZN(n8349) );
  NAND2_X1 U10553 ( .A1(n8355), .A2(SI_18_), .ZN(n8356) );
  MUX2_X1 U10554 ( .A(n10944), .B(n10947), .S(n13436), .Z(n8358) );
  NAND2_X1 U10555 ( .A1(n8358), .A2(n10139), .ZN(n8377) );
  INV_X1 U10556 ( .A(n8358), .ZN(n8359) );
  NAND2_X1 U10557 ( .A1(n8359), .A2(SI_19_), .ZN(n8360) );
  NAND2_X1 U10558 ( .A1(n8377), .A2(n8360), .ZN(n8378) );
  XNOR2_X1 U10559 ( .A(n8379), .B(n8378), .ZN(n13461) );
  NAND2_X1 U10560 ( .A1(n13461), .A2(n8400), .ZN(n8363) );
  INV_X1 U10561 ( .A(n10945), .ZN(n13024) );
  AOI22_X1 U10562 ( .A1(n8361), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n13024), 
        .B2(n8334), .ZN(n8362) );
  NAND2_X1 U10563 ( .A1(n13348), .A2(n8615), .ZN(n8373) );
  NAND2_X1 U10564 ( .A1(n8365), .A2(n8364), .ZN(n8366) );
  AND2_X1 U10565 ( .A1(n8384), .A2(n8366), .ZN(n13249) );
  NAND2_X1 U10566 ( .A1(n13249), .A2(n8160), .ZN(n8371) );
  INV_X1 U10567 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13253) );
  NAND2_X1 U10568 ( .A1(n6571), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8368) );
  INV_X1 U10569 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13017) );
  OR2_X1 U10570 ( .A1(n7997), .A2(n13017), .ZN(n8367) );
  OAI211_X1 U10571 ( .C1(n13253), .C2(n8614), .A(n8368), .B(n8367), .ZN(n8369)
         );
  INV_X1 U10572 ( .A(n8369), .ZN(n8370) );
  NAND2_X1 U10573 ( .A1(n8371), .A2(n8370), .ZN(n13043) );
  NAND2_X1 U10574 ( .A1(n13043), .A2(n8616), .ZN(n8372) );
  NAND2_X1 U10575 ( .A1(n8373), .A2(n8372), .ZN(n8375) );
  AOI22_X1 U10576 ( .A1(n13348), .A2(n8616), .B1(n8615), .B2(n13043), .ZN(
        n8374) );
  XNOR2_X1 U10577 ( .A(n8420), .B(SI_20_), .ZN(n8395) );
  INV_X1 U10578 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11331) );
  MUX2_X1 U10579 ( .A(n13542), .B(n11331), .S(n13436), .Z(n8421) );
  XNOR2_X1 U10580 ( .A(n8395), .B(n8421), .ZN(n13541) );
  NAND2_X1 U10581 ( .A1(n13541), .A2(n8400), .ZN(n8381) );
  NAND2_X1 U10582 ( .A1(n8561), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8380) );
  NAND2_X1 U10583 ( .A1(n13343), .A2(n8616), .ZN(n8392) );
  INV_X1 U10584 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U10585 ( .A1(n8384), .A2(n8383), .ZN(n8385) );
  NAND2_X1 U10586 ( .A1(n8404), .A2(n8385), .ZN(n13237) );
  OR2_X1 U10587 ( .A1(n13237), .A2(n8585), .ZN(n8390) );
  INV_X1 U10588 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13238) );
  NAND2_X1 U10589 ( .A1(n8564), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10590 ( .A1(n6571), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8386) );
  OAI211_X1 U10591 ( .C1(n13238), .C2(n8614), .A(n8387), .B(n8386), .ZN(n8388)
         );
  INV_X1 U10592 ( .A(n8388), .ZN(n8389) );
  NAND2_X1 U10593 ( .A1(n8390), .A2(n8389), .ZN(n13047) );
  NAND2_X1 U10594 ( .A1(n13047), .A2(n8615), .ZN(n8391) );
  NAND2_X1 U10595 ( .A1(n8392), .A2(n8391), .ZN(n8394) );
  AOI22_X1 U10596 ( .A1(n13343), .A2(n8615), .B1(n13047), .B2(n8617), .ZN(
        n8393) );
  INV_X1 U10597 ( .A(n8421), .ZN(n8419) );
  NAND2_X1 U10598 ( .A1(n8395), .A2(n8419), .ZN(n8397) );
  INV_X1 U10599 ( .A(SI_20_), .ZN(n10404) );
  OR2_X1 U10600 ( .A1(n8420), .A2(n10404), .ZN(n8396) );
  NAND2_X1 U10601 ( .A1(n8397), .A2(n8396), .ZN(n8399) );
  MUX2_X1 U10602 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n13436), .Z(n8422) );
  XNOR2_X1 U10603 ( .A(n8422), .B(SI_21_), .ZN(n8398) );
  NAND2_X1 U10604 ( .A1(n13450), .A2(n8400), .ZN(n8402) );
  NAND2_X1 U10605 ( .A1(n8361), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U10606 ( .A1(n13337), .A2(n8615), .ZN(n8413) );
  NAND2_X1 U10607 ( .A1(n8404), .A2(n8403), .ZN(n8405) );
  NAND2_X1 U10608 ( .A1(n8427), .A2(n8405), .ZN(n13219) );
  OR2_X1 U10609 ( .A1(n13219), .A2(n8585), .ZN(n8411) );
  INV_X1 U10610 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U10611 ( .A1(n8564), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U10612 ( .A1(n6571), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8406) );
  OAI211_X1 U10613 ( .C1(n8408), .C2(n8614), .A(n8407), .B(n8406), .ZN(n8409)
         );
  INV_X1 U10614 ( .A(n8409), .ZN(n8410) );
  NAND2_X1 U10615 ( .A1(n8411), .A2(n8410), .ZN(n13048) );
  NAND2_X1 U10616 ( .A1(n13048), .A2(n8616), .ZN(n8412) );
  NAND2_X1 U10617 ( .A1(n8413), .A2(n8412), .ZN(n8418) );
  NAND2_X1 U10618 ( .A1(n13337), .A2(n8617), .ZN(n8415) );
  NAND2_X1 U10619 ( .A1(n13048), .A2(n8615), .ZN(n8414) );
  NAND2_X1 U10620 ( .A1(n8415), .A2(n8414), .ZN(n8416) );
  NOR2_X1 U10621 ( .A1(n8421), .A2(n10404), .ZN(n8423) );
  AOI22_X1 U10622 ( .A1(n8423), .A2(n6598), .B1(n8422), .B2(SI_21_), .ZN(n8424) );
  MUX2_X1 U10623 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n13436), .Z(n8439) );
  XNOR2_X1 U10624 ( .A(n13437), .B(n8439), .ZN(n11404) );
  NAND2_X1 U10625 ( .A1(n11404), .A2(n8532), .ZN(n8426) );
  NAND2_X1 U10626 ( .A1(n8561), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U10627 ( .A1(n13330), .A2(n8616), .ZN(n8436) );
  INV_X1 U10628 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12942) );
  NAND2_X1 U10629 ( .A1(n8427), .A2(n12942), .ZN(n8428) );
  AND2_X1 U10630 ( .A1(n8447), .A2(n8428), .ZN(n13203) );
  NAND2_X1 U10631 ( .A1(n13203), .A2(n8160), .ZN(n8434) );
  INV_X1 U10632 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U10633 ( .A1(n8564), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8430) );
  NAND2_X1 U10634 ( .A1(n6571), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8429) );
  OAI211_X1 U10635 ( .C1(n8431), .C2(n8614), .A(n8430), .B(n8429), .ZN(n8432)
         );
  INV_X1 U10636 ( .A(n8432), .ZN(n8433) );
  NAND2_X1 U10637 ( .A1(n8434), .A2(n8433), .ZN(n12977) );
  NAND2_X1 U10638 ( .A1(n12977), .A2(n8615), .ZN(n8435) );
  NAND2_X1 U10639 ( .A1(n8436), .A2(n8435), .ZN(n8438) );
  AOI22_X1 U10640 ( .A1(n13330), .A2(n8615), .B1(n12977), .B2(n8617), .ZN(
        n8437) );
  INV_X1 U10641 ( .A(n8439), .ZN(n8440) );
  NAND2_X1 U10642 ( .A1(n8441), .A2(SI_22_), .ZN(n8442) );
  MUX2_X1 U10643 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n6568), .Z(n8463) );
  XNOR2_X1 U10644 ( .A(n8463), .B(SI_23_), .ZN(n8443) );
  XNOR2_X1 U10645 ( .A(n8462), .B(n8443), .ZN(n13564) );
  NAND2_X1 U10646 ( .A1(n13564), .A2(n8400), .ZN(n8445) );
  NAND2_X1 U10647 ( .A1(n8361), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8444) );
  NAND2_X2 U10648 ( .A1(n8445), .A2(n8444), .ZN(n13325) );
  NAND2_X1 U10649 ( .A1(n13325), .A2(n8615), .ZN(n8455) );
  INV_X1 U10650 ( .A(n8447), .ZN(n8446) );
  NAND2_X1 U10651 ( .A1(n8446), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8470) );
  INV_X1 U10652 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12853) );
  NAND2_X1 U10653 ( .A1(n8447), .A2(n12853), .ZN(n8448) );
  NAND2_X1 U10654 ( .A1(n8470), .A2(n8448), .ZN(n13188) );
  OR2_X1 U10655 ( .A1(n13188), .A2(n8585), .ZN(n8453) );
  INV_X1 U10656 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n12345) );
  NAND2_X1 U10657 ( .A1(n8586), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U10658 ( .A1(n6571), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8449) );
  OAI211_X1 U10659 ( .C1(n7997), .C2(n12345), .A(n8450), .B(n8449), .ZN(n8451)
         );
  INV_X1 U10660 ( .A(n8451), .ZN(n8452) );
  NAND2_X1 U10661 ( .A1(n13051), .A2(n8616), .ZN(n8454) );
  NAND2_X1 U10662 ( .A1(n13325), .A2(n8617), .ZN(n8457) );
  NAND2_X1 U10663 ( .A1(n13051), .A2(n8615), .ZN(n8456) );
  NAND2_X1 U10664 ( .A1(n8457), .A2(n8456), .ZN(n8458) );
  INV_X1 U10665 ( .A(n8463), .ZN(n8460) );
  INV_X1 U10666 ( .A(SI_23_), .ZN(n10795) );
  NAND2_X1 U10667 ( .A1(n8460), .A2(n10795), .ZN(n8461) );
  NAND2_X1 U10668 ( .A1(n8463), .A2(SI_23_), .ZN(n8464) );
  MUX2_X1 U10669 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n8510), .Z(n8486) );
  NAND2_X1 U10670 ( .A1(n13582), .A2(n8400), .ZN(n8467) );
  NAND2_X1 U10671 ( .A1(n8361), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8466) );
  NAND2_X2 U10672 ( .A1(n8467), .A2(n8466), .ZN(n13318) );
  NAND2_X1 U10673 ( .A1(n13318), .A2(n8616), .ZN(n8478) );
  INV_X1 U10674 ( .A(n8470), .ZN(n8468) );
  NAND2_X1 U10675 ( .A1(n8468), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8495) );
  INV_X1 U10676 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8469) );
  NAND2_X1 U10677 ( .A1(n8470), .A2(n8469), .ZN(n8471) );
  NAND2_X1 U10678 ( .A1(n8495), .A2(n8471), .ZN(n13177) );
  OR2_X1 U10679 ( .A1(n13177), .A2(n8585), .ZN(n8476) );
  INV_X1 U10680 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13176) );
  NAND2_X1 U10681 ( .A1(n8564), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U10682 ( .A1(n6571), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8472) );
  OAI211_X1 U10683 ( .C1(n13176), .C2(n8614), .A(n8473), .B(n8472), .ZN(n8474)
         );
  INV_X1 U10684 ( .A(n8474), .ZN(n8475) );
  NAND2_X1 U10685 ( .A1(n8476), .A2(n8475), .ZN(n13052) );
  NAND2_X1 U10686 ( .A1(n13052), .A2(n8615), .ZN(n8477) );
  NAND2_X1 U10687 ( .A1(n8478), .A2(n8477), .ZN(n8482) );
  INV_X1 U10688 ( .A(n13052), .ZN(n12886) );
  NAND2_X1 U10689 ( .A1(n13318), .A2(n8615), .ZN(n8479) );
  OAI21_X1 U10690 ( .B1(n12886), .B2(n8592), .A(n8479), .ZN(n8480) );
  NAND2_X1 U10691 ( .A1(n8481), .A2(n8480), .ZN(n8485) );
  INV_X1 U10692 ( .A(n8482), .ZN(n8483) );
  NAND2_X1 U10693 ( .A1(n8487), .A2(SI_24_), .ZN(n8488) );
  NAND2_X1 U10694 ( .A1(n8489), .A2(n8488), .ZN(n8509) );
  INV_X1 U10695 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14568) );
  MUX2_X1 U10696 ( .A(n14568), .B(n13413), .S(n8510), .Z(n8490) );
  INV_X1 U10697 ( .A(SI_25_), .ZN(n11295) );
  NAND2_X1 U10698 ( .A1(n8490), .A2(n11295), .ZN(n8507) );
  INV_X1 U10699 ( .A(n8490), .ZN(n8491) );
  NAND2_X1 U10700 ( .A1(n8491), .A2(SI_25_), .ZN(n8492) );
  NAND2_X1 U10701 ( .A1(n8507), .A2(n8492), .ZN(n8508) );
  XNOR2_X1 U10702 ( .A(n8509), .B(n8508), .ZN(n13598) );
  NAND2_X1 U10703 ( .A1(n13598), .A2(n8400), .ZN(n8494) );
  NAND2_X1 U10704 ( .A1(n8361), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8493) );
  NAND2_X1 U10705 ( .A1(n13313), .A2(n8615), .ZN(n8503) );
  NAND2_X1 U10706 ( .A1(n8495), .A2(n12887), .ZN(n8496) );
  NAND2_X1 U10707 ( .A1(n13162), .A2(n8160), .ZN(n8501) );
  INV_X1 U10708 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13164) );
  NAND2_X1 U10709 ( .A1(n8564), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8498) );
  NAND2_X1 U10710 ( .A1(n6571), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8497) );
  OAI211_X1 U10711 ( .C1(n13164), .C2(n8614), .A(n8498), .B(n8497), .ZN(n8499)
         );
  INV_X1 U10712 ( .A(n8499), .ZN(n8500) );
  NAND2_X1 U10713 ( .A1(n8501), .A2(n8500), .ZN(n13053) );
  NAND2_X1 U10714 ( .A1(n13053), .A2(n8616), .ZN(n8502) );
  NAND2_X1 U10715 ( .A1(n8503), .A2(n8502), .ZN(n8506) );
  NAND2_X1 U10716 ( .A1(n13313), .A2(n8616), .ZN(n8504) );
  OAI21_X1 U10717 ( .B1(n13086), .B2(n8635), .A(n8504), .ZN(n8505) );
  MUX2_X1 U10718 ( .A(n14565), .B(n13410), .S(n8510), .Z(n8529) );
  XNOR2_X1 U10719 ( .A(n8529), .B(SI_26_), .ZN(n8511) );
  XNOR2_X1 U10720 ( .A(n8530), .B(n8511), .ZN(n13614) );
  NAND2_X1 U10721 ( .A1(n13614), .A2(n8400), .ZN(n8513) );
  NAND2_X1 U10722 ( .A1(n8361), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8512) );
  NAND2_X1 U10723 ( .A1(n13307), .A2(n8616), .ZN(n8524) );
  INV_X1 U10724 ( .A(n8516), .ZN(n8514) );
  NAND2_X1 U10725 ( .A1(n8514), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8535) );
  INV_X1 U10726 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U10727 ( .A1(n8516), .A2(n8515), .ZN(n8517) );
  NAND2_X1 U10728 ( .A1(n8535), .A2(n8517), .ZN(n12964) );
  OR2_X1 U10729 ( .A1(n12964), .A2(n8585), .ZN(n8522) );
  INV_X1 U10730 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n12174) );
  NAND2_X1 U10731 ( .A1(n8564), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U10732 ( .A1(n8586), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8518) );
  OAI211_X1 U10733 ( .C1(n8092), .C2(n12174), .A(n8519), .B(n8518), .ZN(n8520)
         );
  INV_X1 U10734 ( .A(n8520), .ZN(n8521) );
  NAND2_X1 U10735 ( .A1(n13087), .A2(n8615), .ZN(n8523) );
  NAND2_X1 U10736 ( .A1(n8524), .A2(n8523), .ZN(n8527) );
  NAND2_X1 U10737 ( .A1(n13307), .A2(n8615), .ZN(n8525) );
  OAI21_X1 U10738 ( .B1(n13088), .B2(n8592), .A(n8525), .ZN(n8526) );
  INV_X1 U10739 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14562) );
  INV_X1 U10740 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13408) );
  MUX2_X1 U10741 ( .A(n14562), .B(n13408), .S(n13436), .Z(n8544) );
  XNOR2_X1 U10742 ( .A(n8544), .B(SI_27_), .ZN(n8531) );
  XNOR2_X1 U10743 ( .A(n8547), .B(n8531), .ZN(n13420) );
  NAND2_X1 U10744 ( .A1(n13420), .A2(n8532), .ZN(n8534) );
  NAND2_X1 U10745 ( .A1(n8561), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U10746 ( .A1(n13301), .A2(n8615), .ZN(n8543) );
  INV_X1 U10747 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12843) );
  NAND2_X1 U10748 ( .A1(n8535), .A2(n12843), .ZN(n8536) );
  NAND2_X1 U10749 ( .A1(n13129), .A2(n8160), .ZN(n8541) );
  INV_X1 U10750 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13131) );
  NAND2_X1 U10751 ( .A1(n8564), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U10752 ( .A1(n6571), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8537) );
  OAI211_X1 U10753 ( .C1(n13131), .C2(n8614), .A(n8538), .B(n8537), .ZN(n8539)
         );
  INV_X1 U10754 ( .A(n8539), .ZN(n8540) );
  NAND2_X1 U10755 ( .A1(n13089), .A2(n8616), .ZN(n8542) );
  NAND2_X1 U10756 ( .A1(n8543), .A2(n8542), .ZN(n8599) );
  INV_X1 U10757 ( .A(SI_27_), .ZN(n11495) );
  INV_X1 U10758 ( .A(n8544), .ZN(n8545) );
  NAND2_X1 U10759 ( .A1(n8546), .A2(n8545), .ZN(n8550) );
  INV_X1 U10760 ( .A(n8547), .ZN(n8548) );
  MUX2_X1 U10761 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6568), .Z(n8551) );
  XNOR2_X1 U10762 ( .A(n8551), .B(SI_28_), .ZN(n8568) );
  INV_X1 U10763 ( .A(n8551), .ZN(n8552) );
  INV_X1 U10764 ( .A(SI_28_), .ZN(n11697) );
  NAND2_X1 U10765 ( .A1(n8552), .A2(n11697), .ZN(n8553) );
  INV_X1 U10766 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13849) );
  INV_X1 U10767 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13401) );
  MUX2_X1 U10768 ( .A(n13849), .B(n13401), .S(n6568), .Z(n8554) );
  XNOR2_X1 U10769 ( .A(n8554), .B(SI_29_), .ZN(n8581) );
  INV_X1 U10770 ( .A(SI_29_), .ZN(n12783) );
  NAND2_X1 U10771 ( .A1(n8554), .A2(n12783), .ZN(n8555) );
  MUX2_X1 U10772 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8510), .Z(n8556) );
  XNOR2_X1 U10773 ( .A(n8556), .B(SI_30_), .ZN(n8608) );
  NAND2_X1 U10774 ( .A1(n8556), .A2(SI_30_), .ZN(n8557) );
  OAI21_X1 U10775 ( .B1(n8609), .B2(n8608), .A(n8557), .ZN(n8560) );
  MUX2_X1 U10776 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6568), .Z(n8558) );
  XNOR2_X1 U10777 ( .A(n8558), .B(SI_31_), .ZN(n8559) );
  NAND2_X1 U10778 ( .A1(n14560), .A2(n8400), .ZN(n8563) );
  NAND2_X1 U10779 ( .A1(n8561), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8562) );
  NAND2_X1 U10780 ( .A1(n8563), .A2(n8562), .ZN(n8631) );
  INV_X1 U10781 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U10782 ( .A1(n8564), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U10783 ( .A1(n6571), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8565) );
  OAI211_X1 U10784 ( .C1(n8614), .C2(n8567), .A(n8566), .B(n8565), .ZN(n13033)
         );
  NOR2_X1 U10785 ( .A1(n8631), .A2(n13033), .ZN(n8607) );
  AOI21_X1 U10786 ( .B1(n8631), .B2(n13033), .A(n8607), .ZN(n8661) );
  INV_X1 U10787 ( .A(n8661), .ZN(n8596) );
  NAND2_X1 U10788 ( .A1(n13676), .A2(n8400), .ZN(n8571) );
  NAND2_X1 U10789 ( .A1(n8361), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8570) );
  INV_X1 U10790 ( .A(n8574), .ZN(n8572) );
  NAND2_X1 U10791 ( .A1(n8572), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13060) );
  INV_X1 U10792 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U10793 ( .A1(n8574), .A2(n8573), .ZN(n8575) );
  NAND2_X1 U10794 ( .A1(n13060), .A2(n8575), .ZN(n12871) );
  OR2_X1 U10795 ( .A1(n12871), .A2(n8585), .ZN(n8580) );
  INV_X1 U10796 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n12176) );
  NAND2_X1 U10797 ( .A1(n8586), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8577) );
  INV_X1 U10798 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n12223) );
  OR2_X1 U10799 ( .A1(n8092), .A2(n12223), .ZN(n8576) );
  OAI211_X1 U10800 ( .C1(n7997), .C2(n12176), .A(n8577), .B(n8576), .ZN(n8578)
         );
  INV_X1 U10801 ( .A(n8578), .ZN(n8579) );
  AOI22_X1 U10802 ( .A1(n13107), .A2(n8616), .B1(n8615), .B2(n13096), .ZN(
        n8603) );
  OAI22_X1 U10803 ( .A1(n13292), .A2(n8635), .B1(n13058), .B2(n8592), .ZN(
        n8602) );
  XNOR2_X1 U10804 ( .A(n8582), .B(n8581), .ZN(n13848) );
  NAND2_X1 U10805 ( .A1(n13848), .A2(n8400), .ZN(n8584) );
  NAND2_X1 U10806 ( .A1(n8361), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8583) );
  OR2_X1 U10807 ( .A1(n13060), .A2(n8585), .ZN(n8591) );
  INV_X1 U10808 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n12257) );
  NAND2_X1 U10809 ( .A1(n8586), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U10810 ( .A1(n8564), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8587) );
  OAI211_X1 U10811 ( .C1(n8092), .C2(n12257), .A(n8588), .B(n8587), .ZN(n8589)
         );
  INV_X1 U10812 ( .A(n8589), .ZN(n8590) );
  OAI22_X1 U10813 ( .A1(n13063), .A2(n8592), .B1(n8593), .B2(n8635), .ZN(n8621) );
  AOI22_X1 U10814 ( .A1(n13289), .A2(n8615), .B1(n12976), .B2(n8616), .ZN(
        n8622) );
  NAND2_X1 U10815 ( .A1(n8621), .A2(n8622), .ZN(n8601) );
  OAI21_X1 U10816 ( .B1(n8603), .B2(n8602), .A(n8601), .ZN(n8594) );
  NAND2_X1 U10817 ( .A1(n8596), .A2(n8595), .ZN(n8597) );
  AOI22_X1 U10818 ( .A1(n13301), .A2(n8616), .B1(n8615), .B2(n13089), .ZN(
        n8598) );
  INV_X1 U10819 ( .A(n8601), .ZN(n8606) );
  INV_X1 U10820 ( .A(n8602), .ZN(n8605) );
  INV_X1 U10821 ( .A(n8603), .ZN(n8604) );
  NOR4_X1 U10822 ( .A1(n8661), .A2(n8606), .A3(n8605), .A4(n8604), .ZN(n8628)
         );
  AOI22_X1 U10823 ( .A1(n8631), .A2(n8617), .B1(n8615), .B2(n13033), .ZN(n8626) );
  INV_X1 U10824 ( .A(n8607), .ZN(n8633) );
  INV_X1 U10825 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11726) );
  OAI22_X1 U10826 ( .A1(n13837), .A2(n8611), .B1(n8610), .B2(n11726), .ZN(
        n13040) );
  INV_X1 U10827 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13037) );
  NAND2_X1 U10828 ( .A1(n8564), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U10829 ( .A1(n6571), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8612) );
  OAI211_X1 U10830 ( .C1(n8614), .C2(n13037), .A(n8613), .B(n8612), .ZN(n13097) );
  AOI22_X1 U10831 ( .A1(n13040), .A2(n8616), .B1(n8615), .B2(n13097), .ZN(
        n8630) );
  AND2_X1 U10832 ( .A1(n13033), .A2(n8617), .ZN(n8632) );
  INV_X1 U10833 ( .A(n10147), .ZN(n9696) );
  NAND2_X1 U10834 ( .A1(n10945), .A2(n7288), .ZN(n9707) );
  OAI211_X1 U10835 ( .C1(n9696), .C2(n10146), .A(n9939), .B(n9707), .ZN(n8619)
         );
  OAI21_X1 U10836 ( .B1(n8632), .B2(n8619), .A(n13097), .ZN(n8620) );
  OAI21_X1 U10837 ( .B1(n13287), .B2(n8635), .A(n8620), .ZN(n8629) );
  INV_X1 U10838 ( .A(n8621), .ZN(n8624) );
  INV_X1 U10839 ( .A(n8622), .ZN(n8623) );
  AOI22_X1 U10840 ( .A1(n8630), .A2(n8629), .B1(n8624), .B2(n8623), .ZN(n8625)
         );
  AOI21_X1 U10841 ( .B1(n8626), .B2(n8633), .A(n8625), .ZN(n8627) );
  NOR2_X1 U10842 ( .A1(n8630), .A2(n8629), .ZN(n8637) );
  INV_X1 U10843 ( .A(n8632), .ZN(n8634) );
  OAI211_X1 U10844 ( .C1(n13284), .C2(n8635), .A(n8634), .B(n8633), .ZN(n8636)
         );
  XNOR2_X1 U10845 ( .A(n13287), .B(n13097), .ZN(n8660) );
  XOR2_X1 U10846 ( .A(n12976), .B(n13289), .Z(n13092) );
  NOR2_X1 U10847 ( .A1(n13107), .A2(n13058), .ZN(n13091) );
  AOI21_X1 U10848 ( .B1(n13058), .B2(n13107), .A(n13091), .ZN(n13057) );
  XNOR2_X1 U10849 ( .A(n13313), .B(n13086), .ZN(n13154) );
  NAND2_X1 U10850 ( .A1(n13318), .A2(n12886), .ZN(n13085) );
  OR2_X1 U10851 ( .A1(n13318), .A2(n12886), .ZN(n8638) );
  NAND2_X1 U10852 ( .A1(n13085), .A2(n8638), .ZN(n13084) );
  XNOR2_X1 U10853 ( .A(n13325), .B(n13051), .ZN(n13184) );
  INV_X1 U10854 ( .A(n13047), .ZN(n13044) );
  OR2_X1 U10855 ( .A1(n13343), .A2(n13044), .ZN(n13077) );
  NAND2_X1 U10856 ( .A1(n13343), .A2(n13044), .ZN(n13213) );
  NAND2_X1 U10857 ( .A1(n13077), .A2(n13213), .ZN(n13231) );
  XOR2_X1 U10858 ( .A(n13042), .B(n13353), .Z(n13267) );
  INV_X1 U10859 ( .A(n13043), .ZN(n13075) );
  XNOR2_X1 U10860 ( .A(n13348), .B(n13075), .ZN(n13255) );
  XNOR2_X1 U10861 ( .A(n13369), .B(n12979), .ZN(n11575) );
  XNOR2_X1 U10862 ( .A(n13069), .B(n13065), .ZN(n11595) );
  XNOR2_X1 U10863 ( .A(n13364), .B(n12908), .ZN(n11572) );
  INV_X1 U10864 ( .A(n12981), .ZN(n11300) );
  XNOR2_X1 U10865 ( .A(n13374), .B(n11300), .ZN(n11198) );
  INV_X1 U10866 ( .A(n12982), .ZN(n11196) );
  XNOR2_X1 U10867 ( .A(n11195), .B(n11196), .ZN(n11068) );
  INV_X1 U10868 ( .A(n12984), .ZN(n8639) );
  NAND2_X1 U10869 ( .A1(n11003), .A2(n8639), .ZN(n10988) );
  OR2_X1 U10870 ( .A1(n11003), .A2(n8639), .ZN(n8640) );
  XNOR2_X1 U10871 ( .A(n10745), .B(n12985), .ZN(n10537) );
  INV_X1 U10872 ( .A(n12986), .ZN(n10527) );
  XNOR2_X1 U10873 ( .A(n10647), .B(n10527), .ZN(n10538) );
  INV_X1 U10874 ( .A(n12987), .ZN(n10455) );
  INV_X1 U10875 ( .A(n10300), .ZN(n10135) );
  NAND2_X1 U10876 ( .A1(n10135), .A2(n12989), .ZN(n8641) );
  INV_X1 U10877 ( .A(n12989), .ZN(n10307) );
  NAND2_X1 U10878 ( .A1(n10300), .A2(n10307), .ZN(n10304) );
  NAND2_X1 U10879 ( .A1(n10115), .A2(n8021), .ZN(n10122) );
  OR2_X1 U10880 ( .A1(n15348), .A2(n9920), .ZN(n8642) );
  NAND2_X1 U10881 ( .A1(n15348), .A2(n9920), .ZN(n10121) );
  INV_X1 U10882 ( .A(n7166), .ZN(n15342) );
  NAND2_X1 U10883 ( .A1(n15342), .A2(n12992), .ZN(n8644) );
  INV_X1 U10884 ( .A(n12992), .ZN(n8643) );
  NAND2_X1 U10885 ( .A1(n7166), .A2(n8643), .ZN(n10120) );
  NAND2_X1 U10886 ( .A1(n8644), .A2(n10120), .ZN(n10119) );
  NAND2_X1 U10887 ( .A1(n10130), .A2(n12994), .ZN(n8647) );
  INV_X1 U10888 ( .A(n12994), .ZN(n8646) );
  NAND2_X1 U10889 ( .A1(n8646), .A2(n6574), .ZN(n10118) );
  INV_X1 U10890 ( .A(n8648), .ZN(n9881) );
  NAND2_X1 U10891 ( .A1(n9881), .A2(n10260), .ZN(n10253) );
  NAND2_X1 U10892 ( .A1(n10253), .A2(n8649), .ZN(n15331) );
  NOR4_X1 U10893 ( .A1(n10119), .A2(n7288), .A3(n10252), .A4(n15331), .ZN(
        n8650) );
  NAND4_X1 U10894 ( .A1(n10124), .A2(n10435), .A3(n10204), .A4(n8650), .ZN(
        n8651) );
  NOR4_X1 U10895 ( .A1(n10538), .A2(n10344), .A3(n10446), .A4(n8651), .ZN(
        n8652) );
  XNOR2_X1 U10896 ( .A(n11066), .B(n12983), .ZN(n10990) );
  NAND4_X1 U10897 ( .A1(n10746), .A2(n10537), .A3(n8652), .A4(n10990), .ZN(
        n8653) );
  NOR4_X1 U10898 ( .A1(n11572), .A2(n11198), .A3(n11068), .A4(n8653), .ZN(
        n8654) );
  XNOR2_X1 U10899 ( .A(n11505), .B(n12980), .ZN(n11307) );
  NAND4_X1 U10900 ( .A1(n11575), .A2(n11595), .A3(n8654), .A4(n11307), .ZN(
        n8655) );
  NOR4_X1 U10901 ( .A1(n13231), .A2(n13267), .A3(n13255), .A4(n8655), .ZN(
        n8656) );
  XNOR2_X1 U10902 ( .A(n13330), .B(n12977), .ZN(n13196) );
  XNOR2_X1 U10903 ( .A(n13337), .B(n13048), .ZN(n13222) );
  NAND4_X1 U10904 ( .A1(n13184), .A2(n8656), .A3(n13196), .A4(n13222), .ZN(
        n8657) );
  NOR3_X1 U10905 ( .A1(n13154), .A2(n13084), .A3(n8657), .ZN(n8658) );
  XNOR2_X1 U10906 ( .A(n13307), .B(n13087), .ZN(n13148) );
  XNOR2_X1 U10907 ( .A(n13301), .B(n13089), .ZN(n13055) );
  NAND4_X1 U10908 ( .A1(n13057), .A2(n8658), .A3(n13148), .A4(n13055), .ZN(
        n8659) );
  NOR4_X1 U10909 ( .A1(n8661), .A2(n8660), .A3(n13092), .A4(n8659), .ZN(n8662)
         );
  XOR2_X1 U10910 ( .A(n10945), .B(n8662), .Z(n8663) );
  INV_X1 U10911 ( .A(n9707), .ZN(n8664) );
  AOI21_X1 U10912 ( .B1(n9939), .B2(n10945), .A(n8664), .ZN(n8665) );
  OAI21_X1 U10913 ( .B1(n9712), .B2(n11403), .A(n8665), .ZN(n8666) );
  INV_X1 U10914 ( .A(n9939), .ZN(n11387) );
  MUX2_X1 U10915 ( .A(n11387), .B(n10146), .S(n7288), .Z(n8667) );
  NOR2_X1 U10916 ( .A1(n8667), .A2(n10945), .ZN(n8668) );
  OAI21_X1 U10917 ( .B1(n8671), .B2(n8670), .A(n8669), .ZN(n8680) );
  NAND3_X1 U10918 ( .A1(n8675), .A2(n8674), .A3(n8673), .ZN(n8676) );
  NAND2_X1 U10919 ( .A1(n8676), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8678) );
  OR2_X1 U10920 ( .A1(n8678), .A2(n8677), .ZN(n8679) );
  NOR2_X1 U10921 ( .A1(n9475), .A2(P2_U3088), .ZN(n11491) );
  NAND2_X1 U10922 ( .A1(n8684), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8685) );
  MUX2_X1 U10923 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8685), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8686) );
  NAND2_X1 U10924 ( .A1(n8687), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8688) );
  MUX2_X1 U10925 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8688), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8689) );
  AND2_X1 U10926 ( .A1(n9697), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15327) );
  INV_X1 U10927 ( .A(n15327), .ZN(n15324) );
  NAND2_X1 U10928 ( .A1(n8683), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U10929 ( .A1(n8694), .A2(n8693), .ZN(n8691) );
  NAND2_X1 U10930 ( .A1(n8691), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8692) );
  XNOR2_X1 U10931 ( .A(n8694), .B(n8693), .ZN(n13409) );
  NOR4_X1 U10932 ( .A1(n15324), .A2(n9707), .A3(n12916), .A4(n13409), .ZN(
        n8697) );
  INV_X1 U10933 ( .A(n11491), .ZN(n8695) );
  OAI21_X1 U10934 ( .B1(n8695), .B2(n11403), .A(P2_B_REG_SCAN_IN), .ZN(n8696)
         );
  OR2_X1 U10935 ( .A1(n8697), .A2(n8696), .ZN(n8698) );
  NAND2_X1 U10936 ( .A1(n8699), .A2(n8698), .ZN(P2_U3328) );
  INV_X1 U10937 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8710) );
  XNOR2_X1 U10938 ( .A(n8726), .B(P3_B_REG_SCAN_IN), .ZN(n8721) );
  NAND2_X1 U10939 ( .A1(n6651), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8719) );
  MUX2_X1 U10940 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8719), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8720) );
  NAND2_X1 U10941 ( .A1(n8721), .A2(n11297), .ZN(n8725) );
  NAND2_X1 U10942 ( .A1(n6604), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8722) );
  MUX2_X1 U10943 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8722), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8723) );
  NAND2_X1 U10944 ( .A1(n8726), .A2(n11402), .ZN(n8727) );
  NOR2_X1 U10945 ( .A1(n8718), .A2(n8709), .ZN(n8729) );
  MUX2_X1 U10946 ( .A(n8709), .B(n8729), .S(P3_IR_REG_20__SCAN_IN), .Z(n8730)
         );
  INV_X1 U10947 ( .A(n11932), .ZN(n10582) );
  NOR2_X1 U10948 ( .A1(n8731), .A2(n8709), .ZN(n8732) );
  MUX2_X1 U10949 ( .A(n8709), .B(n8732), .S(P3_IR_REG_19__SCAN_IN), .Z(n8733)
         );
  INV_X1 U10950 ( .A(n8733), .ZN(n8735) );
  INV_X1 U10951 ( .A(n8718), .ZN(n8734) );
  AOI21_X1 U10952 ( .B1(n10582), .B2(n10403), .A(n9382), .ZN(n8736) );
  OR2_X1 U10953 ( .A1(n6570), .A2(SI_4_), .ZN(n8756) );
  XNOR2_X1 U10954 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8798) );
  INV_X1 U10955 ( .A(n8797), .ZN(n8743) );
  NAND2_X1 U10956 ( .A1(n8798), .A2(n8743), .ZN(n8745) );
  INV_X1 U10957 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U10958 ( .A1(n9422), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U10959 ( .A1(n8745), .A2(n8744), .ZN(n8772) );
  XNOR2_X1 U10960 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8771) );
  NAND2_X1 U10961 ( .A1(n8772), .A2(n8771), .ZN(n8747) );
  INV_X1 U10962 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U10963 ( .A1(n9426), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8746) );
  NAND2_X1 U10964 ( .A1(n8747), .A2(n8746), .ZN(n8815) );
  XNOR2_X1 U10965 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8814) );
  NAND2_X1 U10966 ( .A1(n8815), .A2(n8814), .ZN(n8749) );
  NAND2_X1 U10967 ( .A1(n9447), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U10968 ( .A1(n8749), .A2(n8748), .ZN(n8829) );
  XNOR2_X1 U10969 ( .A(n8829), .B(n8828), .ZN(n9439) );
  OR2_X1 U10970 ( .A1(n8799), .A2(n9439), .ZN(n8755) );
  AND2_X1 U10971 ( .A1(n8750), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8751) );
  NAND2_X1 U10972 ( .A1(n8751), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8753) );
  INV_X1 U10973 ( .A(n8751), .ZN(n8752) );
  NAND2_X1 U10974 ( .A1(n8752), .A2(n8844), .ZN(n8832) );
  OR2_X1 U10975 ( .A1(n10163), .A2(n10375), .ZN(n8754) );
  XNOR2_X1 U10976 ( .A(n10473), .B(n10831), .ZN(n8827) );
  INV_X1 U10977 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12774) );
  NAND2_X1 U10978 ( .A1(n8788), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8770) );
  AND2_X2 U10979 ( .A1(n8764), .A2(n12781), .ZN(n8790) );
  NAND2_X1 U10980 ( .A1(n8790), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8769) );
  AND2_X1 U10981 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8765) );
  NOR2_X1 U10982 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8837) );
  OR2_X1 U10983 ( .A1(n8765), .A2(n8837), .ZN(n10957) );
  NAND2_X1 U10984 ( .A1(n8789), .A2(n10957), .ZN(n8768) );
  NAND2_X1 U10985 ( .A1(n9354), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8767) );
  OR2_X1 U10986 ( .A1(n8795), .A2(SI_2_), .ZN(n8777) );
  XNOR2_X1 U10987 ( .A(n8772), .B(n8771), .ZN(n9437) );
  OR2_X1 U10988 ( .A1(n8799), .A2(n9437), .ZN(n8776) );
  OR2_X1 U10989 ( .A1(n10163), .A2(n10371), .ZN(n8775) );
  XNOR2_X1 U10990 ( .A(n8804), .B(n10704), .ZN(n8813) );
  NAND2_X1 U10991 ( .A1(n9354), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8779) );
  NAND2_X1 U10992 ( .A1(n8790), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8778) );
  INV_X1 U10993 ( .A(n8812), .ZN(n12106) );
  INV_X1 U10994 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n15402) );
  OR2_X1 U10995 ( .A1(n6570), .A2(n9962), .ZN(n8783) );
  NAND2_X1 U10996 ( .A1(n8780), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8781) );
  AND2_X1 U10997 ( .A1(n8797), .A2(n8781), .ZN(n9425) );
  OR2_X1 U10998 ( .A1(n8799), .A2(n9425), .ZN(n8782) );
  NAND2_X1 U10999 ( .A1(n8789), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U11000 ( .A1(n8788), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8786) );
  NAND2_X1 U11001 ( .A1(n8790), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U11002 ( .A1(n9354), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8784) );
  NAND2_X1 U11003 ( .A1(n9354), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8793) );
  NAND2_X1 U11004 ( .A1(n8788), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8792) );
  NAND2_X1 U11005 ( .A1(n8790), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8791) );
  INV_X1 U11006 ( .A(SI_1_), .ZN(n9427) );
  NAND2_X1 U11007 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8794) );
  XNOR2_X1 U11008 ( .A(n8798), .B(n8797), .ZN(n9428) );
  INV_X1 U11009 ( .A(n8802), .ZN(n9302) );
  NAND2_X1 U11010 ( .A1(n9267), .A2(n8804), .ZN(n8809) );
  NAND2_X1 U11011 ( .A1(n10708), .A2(n8802), .ZN(n11936) );
  NAND2_X1 U11012 ( .A1(n10708), .A2(n8803), .ZN(n8805) );
  NOR2_X1 U11013 ( .A1(n8804), .A2(n9302), .ZN(n8807) );
  NAND2_X1 U11014 ( .A1(n12108), .A2(n10317), .ZN(n10586) );
  INV_X1 U11015 ( .A(n8810), .ZN(n8811) );
  OR2_X1 U11016 ( .A1(n6569), .A2(SI_3_), .ZN(n8819) );
  XNOR2_X1 U11017 ( .A(n8815), .B(n8814), .ZN(n9435) );
  OR2_X1 U11018 ( .A1(n8799), .A2(n9435), .ZN(n8818) );
  NAND2_X1 U11019 ( .A1(n8774), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8816) );
  XNOR2_X1 U11020 ( .A(n8816), .B(P3_IR_REG_3__SCAN_IN), .ZN(n15418) );
  OR2_X1 U11021 ( .A1(n10163), .A2(n15418), .ZN(n8817) );
  XNOR2_X1 U11022 ( .A(n8804), .B(n9311), .ZN(n8825) );
  INV_X1 U11023 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10784) );
  NAND2_X1 U11024 ( .A1(n8789), .A2(n10784), .ZN(n8824) );
  NAND2_X1 U11025 ( .A1(n8788), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8823) );
  INV_X1 U11026 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n8820) );
  OR2_X1 U11027 ( .A1(n8962), .A2(n8820), .ZN(n8822) );
  NAND2_X1 U11028 ( .A1(n9354), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8821) );
  XNOR2_X1 U11029 ( .A(n8825), .B(n9268), .ZN(n10783) );
  INV_X1 U11030 ( .A(n8825), .ZN(n8826) );
  XNOR2_X1 U11031 ( .A(n8827), .B(n12105), .ZN(n10960) );
  OR2_X1 U11032 ( .A1(n6570), .A2(SI_5_), .ZN(n8836) );
  NAND2_X1 U11033 ( .A1(n8829), .A2(n8828), .ZN(n8831) );
  NAND2_X1 U11034 ( .A1(n9467), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8830) );
  XNOR2_X1 U11035 ( .A(n8848), .B(n8847), .ZN(n9441) );
  OR2_X1 U11036 ( .A1(n8799), .A2(n9441), .ZN(n8835) );
  NAND2_X1 U11037 ( .A1(n8832), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8833) );
  XNOR2_X1 U11038 ( .A(n8833), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10378) );
  OR2_X1 U11039 ( .A1(n10163), .A2(n10378), .ZN(n8834) );
  XNOR2_X1 U11040 ( .A(n10473), .B(n11112), .ZN(n8843) );
  NAND2_X1 U11041 ( .A1(n8788), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U11042 ( .A1(n9354), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8841) );
  NAND2_X1 U11043 ( .A1(n8837), .A2(n11099), .ZN(n8854) );
  OR2_X1 U11044 ( .A1(n8837), .A2(n11099), .ZN(n8838) );
  NAND2_X1 U11045 ( .A1(n8854), .A2(n8838), .ZN(n11113) );
  NAND2_X1 U11046 ( .A1(n8789), .A2(n11113), .ZN(n8840) );
  NAND2_X1 U11047 ( .A1(n8790), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8839) );
  INV_X1 U11048 ( .A(n11206), .ZN(n12104) );
  XNOR2_X1 U11049 ( .A(n8843), .B(n12104), .ZN(n11097) );
  NAND2_X1 U11050 ( .A1(n8844), .A2(n6818), .ZN(n8845) );
  NOR2_X1 U11051 ( .A1(n8750), .A2(n8845), .ZN(n8868) );
  OR2_X1 U11052 ( .A1(n8868), .A2(n8709), .ZN(n8846) );
  XNOR2_X1 U11053 ( .A(n8846), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10555) );
  INV_X1 U11054 ( .A(SI_6_), .ZN(n9429) );
  OR2_X1 U11055 ( .A1(n6569), .A2(n9429), .ZN(n8853) );
  INV_X1 U11056 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8849) );
  NAND2_X1 U11057 ( .A1(n8849), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8850) );
  XNOR2_X1 U11058 ( .A(n9549), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8851) );
  XNOR2_X1 U11059 ( .A(n8872), .B(n8851), .ZN(n9430) );
  OR2_X1 U11060 ( .A1(n8799), .A2(n9430), .ZN(n8852) );
  OAI211_X1 U11061 ( .C1(n10163), .C2(n10547), .A(n8853), .B(n8852), .ZN(n9315) );
  INV_X1 U11062 ( .A(n9315), .ZN(n11205) );
  XNOR2_X1 U11063 ( .A(n10473), .B(n11205), .ZN(n8860) );
  NAND2_X1 U11064 ( .A1(n8788), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8859) );
  NAND2_X1 U11065 ( .A1(n9354), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U11066 ( .A1(n8854), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8855) );
  NAND2_X1 U11067 ( .A1(n8861), .A2(n8855), .ZN(n11185) );
  NAND2_X1 U11068 ( .A1(n8789), .A2(n11185), .ZN(n8857) );
  NAND2_X1 U11069 ( .A1(n8790), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8856) );
  XNOR2_X1 U11070 ( .A(n8860), .B(n11288), .ZN(n11204) );
  NAND2_X1 U11071 ( .A1(n9354), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8866) );
  NAND2_X1 U11072 ( .A1(n8788), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8865) );
  AND2_X1 U11073 ( .A1(n8861), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8862) );
  OR2_X1 U11074 ( .A1(n8862), .A2(n8888), .ZN(n11284) );
  NAND2_X1 U11075 ( .A1(n8789), .A2(n11284), .ZN(n8864) );
  NAND2_X1 U11076 ( .A1(n8790), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8863) );
  NAND4_X1 U11077 ( .A1(n8866), .A2(n8865), .A3(n8864), .A4(n8863), .ZN(n12102) );
  INV_X1 U11078 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8867) );
  NAND2_X1 U11079 ( .A1(n8868), .A2(n8867), .ZN(n8882) );
  NAND2_X1 U11080 ( .A1(n8882), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8870) );
  INV_X1 U11081 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8869) );
  XNOR2_X1 U11082 ( .A(n8870), .B(n8869), .ZN(n12393) );
  AND2_X1 U11083 ( .A1(n9549), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8871) );
  XNOR2_X1 U11084 ( .A(n9553), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8877) );
  XNOR2_X1 U11085 ( .A(n8879), .B(n8877), .ZN(n9431) );
  OR2_X1 U11086 ( .A1(n8799), .A2(n9431), .ZN(n8874) );
  OR2_X1 U11087 ( .A1(n6570), .A2(SI_7_), .ZN(n8873) );
  OAI211_X1 U11088 ( .C1(n12381), .C2(n10163), .A(n8874), .B(n8873), .ZN(
        n11965) );
  XNOR2_X1 U11089 ( .A(n12102), .B(n11965), .ZN(n11912) );
  XNOR2_X1 U11090 ( .A(n11912), .B(n8803), .ZN(n11286) );
  NAND2_X1 U11091 ( .A1(n11287), .A2(n11286), .ZN(n11285) );
  INV_X1 U11092 ( .A(n11286), .ZN(n8875) );
  NAND2_X1 U11093 ( .A1(n8875), .A2(n12102), .ZN(n8876) );
  NAND2_X1 U11094 ( .A1(n11285), .A2(n8876), .ZN(n11393) );
  INV_X1 U11095 ( .A(SI_8_), .ZN(n9423) );
  OR2_X1 U11096 ( .A1(n6570), .A2(n9423), .ZN(n8886) );
  INV_X1 U11097 ( .A(n8877), .ZN(n8878) );
  NAND2_X1 U11098 ( .A1(n9553), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U11099 ( .A1(n8881), .A2(n8880), .ZN(n8900) );
  XNOR2_X1 U11100 ( .A(n8900), .B(n8899), .ZN(n9424) );
  OR2_X1 U11101 ( .A1(n8799), .A2(n9424), .ZN(n8885) );
  NAND2_X1 U11102 ( .A1(n8896), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8883) );
  XNOR2_X1 U11103 ( .A(n8883), .B(P3_IR_REG_8__SCAN_IN), .ZN(n14640) );
  OR2_X1 U11104 ( .A1(n10163), .A2(n14601), .ZN(n8884) );
  XNOR2_X1 U11105 ( .A(n8804), .B(n11971), .ZN(n8894) );
  NAND2_X1 U11106 ( .A1(n8788), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8893) );
  NAND2_X1 U11107 ( .A1(n8790), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8892) );
  NOR2_X1 U11108 ( .A1(n8888), .A2(n8887), .ZN(n8889) );
  OR2_X1 U11109 ( .A1(n8906), .A2(n8889), .ZN(n11390) );
  NAND2_X1 U11110 ( .A1(n8789), .A2(n11390), .ZN(n8891) );
  NAND2_X1 U11111 ( .A1(n9354), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8890) );
  XNOR2_X1 U11112 ( .A(n8894), .B(n11564), .ZN(n11392) );
  NAND2_X1 U11113 ( .A1(n8894), .A2(n12101), .ZN(n8895) );
  NAND2_X1 U11114 ( .A1(n11391), .A2(n8895), .ZN(n11561) );
  OAI21_X1 U11115 ( .B1(n8896), .B2(P3_IR_REG_8__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8898) );
  INV_X1 U11116 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8897) );
  XNOR2_X1 U11117 ( .A(n8898), .B(n8897), .ZN(n15467) );
  OR2_X1 U11118 ( .A1(n6569), .A2(SI_9_), .ZN(n8905) );
  NAND2_X1 U11119 ( .A1(n8900), .A2(n8899), .ZN(n8903) );
  NAND2_X1 U11120 ( .A1(n8901), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8902) );
  XNOR2_X1 U11121 ( .A(n8917), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n8914) );
  XNOR2_X1 U11122 ( .A(n8916), .B(n8914), .ZN(n9433) );
  OR2_X1 U11123 ( .A1(n8799), .A2(n9433), .ZN(n8904) );
  OAI211_X1 U11124 ( .C1(n14642), .C2(n10163), .A(n8905), .B(n8904), .ZN(
        n11979) );
  INV_X1 U11125 ( .A(n11979), .ZN(n11977) );
  XNOR2_X1 U11126 ( .A(n10473), .B(n11977), .ZN(n8912) );
  NAND2_X1 U11127 ( .A1(n8788), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U11128 ( .A1(n9354), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U11129 ( .A1(n8906), .A2(n11563), .ZN(n8925) );
  OR2_X1 U11130 ( .A1(n8906), .A2(n11563), .ZN(n8907) );
  NAND2_X1 U11131 ( .A1(n8925), .A2(n8907), .ZN(n11566) );
  NAND2_X1 U11132 ( .A1(n8789), .A2(n11566), .ZN(n8909) );
  NAND2_X1 U11133 ( .A1(n8790), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8908) );
  NAND4_X1 U11134 ( .A1(n8911), .A2(n8910), .A3(n8909), .A4(n8908), .ZN(n12100) );
  INV_X1 U11135 ( .A(n12100), .ZN(n11609) );
  XNOR2_X1 U11136 ( .A(n8912), .B(n11609), .ZN(n11562) );
  NAND2_X1 U11137 ( .A1(n8912), .A2(n11609), .ZN(n8913) );
  INV_X1 U11138 ( .A(n8914), .ZN(n8915) );
  NAND2_X1 U11139 ( .A1(n8917), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8918) );
  XNOR2_X1 U11140 ( .A(n12307), .B(P1_DATAO_REG_10__SCAN_IN), .ZN(n8934) );
  XNOR2_X1 U11141 ( .A(n8936), .B(n8934), .ZN(n9445) );
  OR2_X1 U11142 ( .A1(n8799), .A2(n9445), .ZN(n8924) );
  OR2_X1 U11143 ( .A1(n6570), .A2(SI_10_), .ZN(n8923) );
  OR2_X1 U11144 ( .A1(n8919), .A2(n8709), .ZN(n8921) );
  XNOR2_X1 U11145 ( .A(n8921), .B(n8920), .ZN(n15485) );
  OR2_X1 U11146 ( .A1(n10163), .A2(n14644), .ZN(n8922) );
  XNOR2_X1 U11147 ( .A(n10473), .B(n11472), .ZN(n8932) );
  NAND2_X1 U11148 ( .A1(n9354), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8930) );
  NAND2_X1 U11149 ( .A1(n8788), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8929) );
  NAND2_X1 U11150 ( .A1(n8925), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8926) );
  NAND2_X1 U11151 ( .A1(n8946), .A2(n8926), .ZN(n11473) );
  NAND2_X1 U11152 ( .A1(n8789), .A2(n11473), .ZN(n8928) );
  NAND2_X1 U11153 ( .A1(n8790), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8927) );
  XNOR2_X1 U11154 ( .A(n8932), .B(n11836), .ZN(n11604) );
  INV_X1 U11155 ( .A(n8932), .ZN(n8933) );
  INV_X1 U11156 ( .A(n8934), .ZN(n8935) );
  NAND2_X1 U11157 ( .A1(n12307), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U11158 ( .A1(n8938), .A2(n8937), .ZN(n8954) );
  XNOR2_X1 U11159 ( .A(n9811), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8939) );
  XNOR2_X1 U11160 ( .A(n8954), .B(n8939), .ZN(n9458) );
  OR2_X1 U11161 ( .A1(n8799), .A2(n9458), .ZN(n8945) );
  OR2_X1 U11162 ( .A1(n6570), .A2(SI_11_), .ZN(n8944) );
  NAND2_X1 U11163 ( .A1(n8940), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8941) );
  MUX2_X1 U11164 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8941), .S(
        P3_IR_REG_11__SCAN_IN), .Z(n8942) );
  NAND2_X1 U11165 ( .A1(n8942), .A2(n6584), .ZN(n15501) );
  OR2_X1 U11166 ( .A1(n10163), .A2(n14646), .ZN(n8943) );
  XNOR2_X1 U11167 ( .A(n8804), .B(n11414), .ZN(n8970) );
  NAND2_X1 U11168 ( .A1(n8788), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U11169 ( .A1(n9354), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U11170 ( .A1(n8946), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U11171 ( .A1(n8963), .A2(n8947), .ZN(n11838) );
  NAND2_X1 U11172 ( .A1(n8789), .A2(n11838), .ZN(n8949) );
  NAND2_X1 U11173 ( .A1(n8790), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8948) );
  NAND2_X1 U11174 ( .A1(n6584), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8952) );
  XNOR2_X1 U11175 ( .A(n8952), .B(P3_IR_REG_12__SCAN_IN), .ZN(n14648) );
  NAND2_X1 U11176 ( .A1(n9811), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U11177 ( .A1(n9933), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8976) );
  NAND2_X1 U11178 ( .A1(n9927), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8956) );
  NAND2_X1 U11179 ( .A1(n8976), .A2(n8956), .ZN(n8957) );
  NAND2_X1 U11180 ( .A1(n8958), .A2(n8957), .ZN(n8959) );
  NAND2_X1 U11181 ( .A1(n8977), .A2(n8959), .ZN(n9473) );
  OR2_X1 U11182 ( .A1(n8799), .A2(n9473), .ZN(n8961) );
  OR2_X1 U11183 ( .A1(n6569), .A2(n9474), .ZN(n8960) );
  OAI211_X1 U11184 ( .C1(n10163), .C2(n15519), .A(n8961), .B(n8960), .ZN(
        n12637) );
  INV_X1 U11185 ( .A(n12637), .ZN(n11765) );
  XNOR2_X1 U11186 ( .A(n10473), .B(n11765), .ZN(n11762) );
  NAND2_X1 U11187 ( .A1(n8788), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8968) );
  NAND2_X1 U11188 ( .A1(n8790), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8967) );
  AND2_X1 U11189 ( .A1(n8963), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8964) );
  OR2_X1 U11190 ( .A1(n8964), .A2(n8984), .ZN(n12638) );
  NAND2_X1 U11191 ( .A1(n8789), .A2(n12638), .ZN(n8966) );
  NAND2_X1 U11192 ( .A1(n9354), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U11193 ( .A1(n11762), .A2(n12616), .ZN(n8969) );
  OAI21_X1 U11194 ( .B1(n8970), .B2(n11832), .A(n8969), .ZN(n8975) );
  INV_X1 U11195 ( .A(n11762), .ZN(n8973) );
  INV_X1 U11196 ( .A(n8969), .ZN(n8971) );
  INV_X1 U11197 ( .A(n8970), .ZN(n11761) );
  NOR3_X1 U11198 ( .A1(n8971), .A2(n12632), .A3(n11761), .ZN(n8972) );
  AOI21_X1 U11199 ( .B1(n11820), .B2(n8973), .A(n8972), .ZN(n8974) );
  NAND2_X1 U11200 ( .A1(n8978), .A2(n10048), .ZN(n8992) );
  INV_X1 U11201 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10046) );
  NAND2_X1 U11202 ( .A1(n6690), .A2(n10046), .ZN(n8979) );
  NAND2_X1 U11203 ( .A1(n8993), .A2(n8979), .ZN(n9613) );
  NAND2_X1 U11204 ( .A1(n9613), .A2(n11887), .ZN(n8983) );
  INV_X1 U11205 ( .A(n10163), .ZN(n9077) );
  OR2_X1 U11206 ( .A1(n6584), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8995) );
  NAND2_X1 U11207 ( .A1(n8995), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8981) );
  INV_X1 U11208 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8980) );
  XNOR2_X1 U11209 ( .A(n8981), .B(n8980), .ZN(n15537) );
  AOI22_X1 U11210 ( .A1(n9063), .A2(n9614), .B1(n9077), .B2(n15537), .ZN(n8982) );
  NAND2_X1 U11211 ( .A1(n8983), .A2(n8982), .ZN(n12622) );
  XNOR2_X1 U11212 ( .A(n12622), .B(n10473), .ZN(n11815) );
  NAND2_X1 U11213 ( .A1(n9354), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U11214 ( .A1(n8788), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U11215 ( .A1(n8984), .A2(n11818), .ZN(n9003) );
  OR2_X1 U11216 ( .A1(n8984), .A2(n11818), .ZN(n8985) );
  NAND2_X1 U11217 ( .A1(n9003), .A2(n8985), .ZN(n12623) );
  NAND2_X1 U11218 ( .A1(n8789), .A2(n12623), .ZN(n8987) );
  NAND2_X1 U11219 ( .A1(n8790), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8986) );
  NOR2_X1 U11220 ( .A1(n11815), .A2(n12634), .ZN(n8991) );
  INV_X1 U11221 ( .A(n11815), .ZN(n8990) );
  XNOR2_X1 U11222 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8994) );
  XNOR2_X1 U11223 ( .A(n9010), .B(n8994), .ZN(n9675) );
  NAND2_X1 U11224 ( .A1(n9675), .A2(n11887), .ZN(n9002) );
  INV_X1 U11225 ( .A(SI_14_), .ZN(n9676) );
  NOR2_X1 U11226 ( .A1(n8995), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8999) );
  NOR2_X1 U11227 ( .A1(n8999), .A2(n8709), .ZN(n8996) );
  MUX2_X1 U11228 ( .A(n8709), .B(n8996), .S(P3_IR_REG_14__SCAN_IN), .Z(n8997)
         );
  INV_X1 U11229 ( .A(n8997), .ZN(n9000) );
  INV_X1 U11230 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U11231 ( .A1(n8999), .A2(n8998), .ZN(n9013) );
  NAND2_X1 U11232 ( .A1(n9000), .A2(n9013), .ZN(n15554) );
  AOI22_X1 U11233 ( .A1(n9063), .A2(n9676), .B1(n9077), .B2(n15554), .ZN(n9001) );
  XOR2_X1 U11234 ( .A(n8804), .B(n12769), .Z(n11729) );
  NAND2_X1 U11235 ( .A1(n9354), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U11236 ( .A1(n8788), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U11237 ( .A1(n9003), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U11238 ( .A1(n9017), .A2(n9004), .ZN(n12606) );
  NAND2_X1 U11239 ( .A1(n8789), .A2(n12606), .ZN(n9006) );
  NAND2_X1 U11240 ( .A1(n8790), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9005) );
  NAND4_X1 U11241 ( .A1(n9008), .A2(n9007), .A3(n9006), .A4(n9005), .ZN(n12617) );
  INV_X1 U11242 ( .A(n12617), .ZN(n12586) );
  NAND2_X1 U11243 ( .A1(n12254), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U11244 ( .A1(n10342), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9011) );
  XNOR2_X1 U11245 ( .A(n10572), .B(P2_DATAO_REG_15__SCAN_IN), .ZN(n9026) );
  XNOR2_X1 U11246 ( .A(n9028), .B(n9026), .ZN(n9807) );
  NAND2_X1 U11247 ( .A1(n9807), .A2(n11887), .ZN(n9016) );
  NAND2_X1 U11248 ( .A1(n9013), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9012) );
  MUX2_X1 U11249 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9012), .S(
        P3_IR_REG_15__SCAN_IN), .Z(n9014) );
  NAND2_X1 U11250 ( .A1(n9014), .A2(n9047), .ZN(n14827) );
  INV_X1 U11251 ( .A(n14827), .ZN(n14623) );
  AOI22_X1 U11252 ( .A1(n9063), .A2(SI_15_), .B1(n9077), .B2(n14623), .ZN(
        n9015) );
  NAND2_X1 U11253 ( .A1(n9016), .A2(n9015), .ZN(n11862) );
  XNOR2_X1 U11254 ( .A(n11862), .B(n10473), .ZN(n9023) );
  NAND2_X1 U11255 ( .A1(n9354), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U11256 ( .A1(n8788), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9021) );
  AND2_X1 U11257 ( .A1(n9017), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9018) );
  OR2_X1 U11258 ( .A1(n9018), .A2(n9034), .ZN(n12593) );
  NAND2_X1 U11259 ( .A1(n8789), .A2(n12593), .ZN(n9020) );
  NAND2_X1 U11260 ( .A1(n8790), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9019) );
  NAND4_X1 U11261 ( .A1(n9022), .A2(n9021), .A3(n9020), .A4(n9019), .ZN(n12603) );
  XNOR2_X1 U11262 ( .A(n9023), .B(n12603), .ZN(n11865) );
  INV_X1 U11263 ( .A(n9023), .ZN(n9024) );
  NAND2_X1 U11264 ( .A1(n9024), .A2(n12603), .ZN(n9025) );
  INV_X1 U11265 ( .A(n9026), .ZN(n9027) );
  NAND2_X1 U11266 ( .A1(n10573), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9029) );
  XNOR2_X1 U11267 ( .A(n10331), .B(P2_DATAO_REG_16__SCAN_IN), .ZN(n9040) );
  XNOR2_X1 U11268 ( .A(n9042), .B(n9040), .ZN(n9867) );
  NAND2_X1 U11269 ( .A1(n9867), .A2(n11887), .ZN(n9032) );
  NAND2_X1 U11270 ( .A1(n9047), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9030) );
  XNOR2_X1 U11271 ( .A(n9030), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14655) );
  AOI22_X1 U11272 ( .A1(n9063), .A2(SI_16_), .B1(n9077), .B2(n14655), .ZN(
        n9031) );
  NAND2_X1 U11273 ( .A1(n9032), .A2(n9031), .ZN(n12701) );
  XOR2_X1 U11274 ( .A(n8804), .B(n12701), .Z(n11782) );
  NAND2_X1 U11275 ( .A1(n9354), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U11276 ( .A1(n8788), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9038) );
  NOR2_X1 U11277 ( .A1(n9034), .A2(n9033), .ZN(n9035) );
  OR2_X1 U11278 ( .A1(n9051), .A2(n9035), .ZN(n12577) );
  NAND2_X1 U11279 ( .A1(n8789), .A2(n12577), .ZN(n9037) );
  NAND2_X1 U11280 ( .A1(n8790), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9036) );
  INV_X1 U11281 ( .A(n12588), .ZN(n12557) );
  INV_X1 U11282 ( .A(n9040), .ZN(n9041) );
  NAND2_X1 U11283 ( .A1(n10340), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9043) );
  AOI22_X1 U11284 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10466), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n12347), .ZN(n9045) );
  INV_X1 U11285 ( .A(n9045), .ZN(n9046) );
  XNOR2_X1 U11286 ( .A(n9058), .B(n9046), .ZN(n9886) );
  NAND2_X1 U11287 ( .A1(n9886), .A2(n11887), .ZN(n9050) );
  OAI21_X1 U11288 ( .B1(n9047), .B2(P3_IR_REG_16__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9048) );
  XNOR2_X1 U11289 ( .A(n9048), .B(P3_IR_REG_17__SCAN_IN), .ZN(n14628) );
  AOI22_X1 U11290 ( .A1(n9063), .A2(SI_17_), .B1(n9077), .B2(n14628), .ZN(
        n9049) );
  NAND2_X1 U11291 ( .A1(n9050), .A2(n9049), .ZN(n12697) );
  XNOR2_X1 U11292 ( .A(n12697), .B(n10473), .ZN(n11790) );
  NAND2_X1 U11293 ( .A1(n8788), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U11294 ( .A1(n8790), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9055) );
  OR2_X1 U11295 ( .A1(n9051), .A2(n12256), .ZN(n9052) );
  NAND2_X1 U11296 ( .A1(n9066), .A2(n9052), .ZN(n12563) );
  NAND2_X1 U11297 ( .A1(n8789), .A2(n12563), .ZN(n9054) );
  NAND2_X1 U11298 ( .A1(n9354), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U11299 ( .A1(n10466), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U11300 ( .A1(n12269), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U11301 ( .A1(n10792), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9060) );
  XNOR2_X1 U11302 ( .A(n9074), .B(n9072), .ZN(n14781) );
  NAND2_X1 U11303 ( .A1(n14781), .A2(n11887), .ZN(n9065) );
  NAND2_X1 U11304 ( .A1(n9061), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9062) );
  XNOR2_X1 U11305 ( .A(n9062), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14660) );
  AOI22_X1 U11306 ( .A1(n9063), .A2(SI_18_), .B1(n9077), .B2(n14660), .ZN(
        n9064) );
  NAND2_X1 U11307 ( .A1(n9065), .A2(n9064), .ZN(n12550) );
  XOR2_X1 U11308 ( .A(n10473), .B(n12550), .Z(n11842) );
  NAND2_X1 U11309 ( .A1(n9354), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U11310 ( .A1(n8788), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U11311 ( .A1(n9066), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9067) );
  NAND2_X1 U11312 ( .A1(n9080), .A2(n9067), .ZN(n12551) );
  NAND2_X1 U11313 ( .A1(n8789), .A2(n12551), .ZN(n9069) );
  NAND2_X1 U11314 ( .A1(n8790), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9068) );
  INV_X1 U11315 ( .A(n9072), .ZN(n9073) );
  NAND2_X1 U11316 ( .A1(n10944), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9089) );
  NAND2_X1 U11317 ( .A1(n10947), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9076) );
  XNOR2_X1 U11318 ( .A(n9088), .B(n9087), .ZN(n10140) );
  NAND2_X1 U11319 ( .A1(n10140), .A2(n11887), .ZN(n9079) );
  AOI22_X1 U11320 ( .A1(n9063), .A2(n10139), .B1(n9077), .B2(n14638), .ZN(
        n9078) );
  XNOR2_X1 U11321 ( .A(n12755), .B(n10473), .ZN(n9086) );
  NAND2_X1 U11322 ( .A1(n9354), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9085) );
  NAND2_X1 U11323 ( .A1(n8788), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9084) );
  AND2_X1 U11324 ( .A1(n9080), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9081) );
  OR2_X1 U11325 ( .A1(n9081), .A2(n9093), .ZN(n12537) );
  NAND2_X1 U11326 ( .A1(n8789), .A2(n12537), .ZN(n9083) );
  NAND2_X1 U11327 ( .A1(n8790), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9082) );
  NAND4_X1 U11328 ( .A1(n9085), .A2(n9084), .A3(n9083), .A4(n9082), .ZN(n12098) );
  INV_X1 U11329 ( .A(n12098), .ZN(n12549) );
  XNOR2_X1 U11330 ( .A(n9086), .B(n12549), .ZN(n11746) );
  XNOR2_X1 U11331 ( .A(n9106), .B(n13542), .ZN(n10402) );
  NAND2_X1 U11332 ( .A1(n10402), .A2(n11887), .ZN(n9092) );
  OR2_X1 U11333 ( .A1(n6569), .A2(n10404), .ZN(n9091) );
  XNOR2_X1 U11334 ( .A(n12524), .B(n10473), .ZN(n9099) );
  NAND2_X1 U11335 ( .A1(n9354), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9098) );
  NOR2_X1 U11336 ( .A1(n9093), .A2(n11809), .ZN(n9094) );
  OR2_X1 U11337 ( .A1(n9102), .A2(n9094), .ZN(n12525) );
  NAND2_X1 U11338 ( .A1(n8789), .A2(n12525), .ZN(n9097) );
  NAND2_X1 U11339 ( .A1(n8788), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9096) );
  NAND2_X1 U11340 ( .A1(n8790), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9095) );
  XNOR2_X1 U11341 ( .A(n9099), .B(n12509), .ZN(n11807) );
  INV_X1 U11342 ( .A(n9099), .ZN(n9100) );
  NAND2_X1 U11343 ( .A1(n9100), .A2(n12534), .ZN(n9101) );
  OR2_X1 U11344 ( .A1(n9102), .A2(n12199), .ZN(n9103) );
  NAND2_X1 U11345 ( .A1(n9122), .A2(n9103), .ZN(n12512) );
  AOI22_X1 U11346 ( .A1(n12512), .A2(n8789), .B1(n8790), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n9105) );
  AOI22_X1 U11347 ( .A1(n9354), .A2(P3_REG0_REG_21__SCAN_IN), .B1(n8788), .B2(
        P3_REG1_REG_21__SCAN_IN), .ZN(n9104) );
  INV_X1 U11348 ( .A(n9107), .ZN(n9108) );
  NAND2_X1 U11349 ( .A1(n9108), .A2(n11331), .ZN(n9109) );
  XNOR2_X1 U11350 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .ZN(n9114) );
  XNOR2_X1 U11351 ( .A(n9115), .B(n9114), .ZN(n10630) );
  NAND2_X1 U11352 ( .A1(n10630), .A2(n11887), .ZN(n9111) );
  INV_X1 U11353 ( .A(SI_21_), .ZN(n10631) );
  OR2_X1 U11354 ( .A1(n6570), .A2(n10631), .ZN(n9110) );
  XNOR2_X1 U11355 ( .A(n12516), .B(n10473), .ZN(n9112) );
  XOR2_X1 U11356 ( .A(n12522), .B(n9112), .Z(n11752) );
  NOR2_X1 U11357 ( .A1(n9112), .A2(n12522), .ZN(n9113) );
  INV_X1 U11358 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11388) );
  NAND2_X1 U11359 ( .A1(n11388), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9116) );
  XNOR2_X1 U11360 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .ZN(n9127) );
  XNOR2_X1 U11361 ( .A(n9128), .B(n9127), .ZN(n14788) );
  NAND2_X1 U11362 ( .A1(n14788), .A2(n11887), .ZN(n9119) );
  INV_X1 U11363 ( .A(SI_22_), .ZN(n9117) );
  OR2_X1 U11364 ( .A1(n6569), .A2(n9117), .ZN(n9118) );
  XNOR2_X1 U11365 ( .A(n11829), .B(n10473), .ZN(n9121) );
  INV_X1 U11366 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U11367 ( .A1(n9122), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9123) );
  NAND2_X1 U11368 ( .A1(n9137), .A2(n9123), .ZN(n12498) );
  NAND2_X1 U11369 ( .A1(n12498), .A2(n8789), .ZN(n9125) );
  AOI22_X1 U11370 ( .A1(n9354), .A2(P3_REG0_REG_22__SCAN_IN), .B1(n8788), .B2(
        P3_REG1_REG_22__SCAN_IN), .ZN(n9124) );
  INV_X1 U11371 ( .A(n9135), .ZN(n9133) );
  INV_X1 U11372 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n9129) );
  XNOR2_X1 U11373 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9142) );
  XNOR2_X1 U11374 ( .A(n9143), .B(n9142), .ZN(n10793) );
  NAND2_X1 U11375 ( .A1(n10793), .A2(n11887), .ZN(n9131) );
  OR2_X1 U11376 ( .A1(n6570), .A2(n10795), .ZN(n9130) );
  XNOR2_X1 U11377 ( .A(n11742), .B(n10473), .ZN(n9134) );
  INV_X1 U11378 ( .A(n9134), .ZN(n9132) );
  NAND2_X1 U11379 ( .A1(n9133), .A2(n9132), .ZN(n9136) );
  NAND2_X1 U11380 ( .A1(n9136), .A2(n11798), .ZN(n11738) );
  NAND2_X1 U11381 ( .A1(n9137), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9138) );
  NAND2_X1 U11382 ( .A1(n9151), .A2(n9138), .ZN(n12488) );
  NAND2_X1 U11383 ( .A1(n12488), .A2(n8789), .ZN(n9141) );
  AOI22_X1 U11384 ( .A1(n9354), .A2(P3_REG0_REG_23__SCAN_IN), .B1(n8788), .B2(
        P3_REG1_REG_23__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U11385 ( .A1(n8790), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9139) );
  NAND2_X1 U11386 ( .A1(n9143), .A2(n9142), .ZN(n9146) );
  INV_X1 U11387 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9144) );
  NAND2_X1 U11388 ( .A1(n9144), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U11389 ( .A1(n9147), .A2(n13416), .ZN(n9148) );
  INV_X1 U11390 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n14572) );
  XNOR2_X1 U11391 ( .A(n9159), .B(n14572), .ZN(n11700) );
  NAND2_X1 U11392 ( .A1(n11700), .A2(n11887), .ZN(n9150) );
  OR2_X1 U11393 ( .A1(n6569), .A2(n7624), .ZN(n9149) );
  XNOR2_X1 U11394 ( .A(n12478), .B(n10473), .ZN(n9156) );
  AND2_X1 U11395 ( .A1(n9151), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9152) );
  OR2_X1 U11396 ( .A1(n9152), .A2(n9165), .ZN(n12474) );
  INV_X1 U11397 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12476) );
  NAND2_X1 U11398 ( .A1(n9354), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9154) );
  NAND2_X1 U11399 ( .A1(n8788), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9153) );
  OAI211_X1 U11400 ( .C1(n12476), .C2(n8962), .A(n9154), .B(n9153), .ZN(n9155)
         );
  NAND2_X1 U11401 ( .A1(n9156), .A2(n12487), .ZN(n11771) );
  INV_X1 U11402 ( .A(n9156), .ZN(n9157) );
  INV_X1 U11403 ( .A(n12487), .ZN(n12453) );
  NAND2_X1 U11404 ( .A1(n9157), .A2(n12453), .ZN(n9158) );
  AND2_X1 U11405 ( .A1(n11771), .A2(n9158), .ZN(n11799) );
  AOI22_X1 U11406 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n14568), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n13413), .ZN(n9161) );
  INV_X1 U11407 ( .A(n9161), .ZN(n9162) );
  XNOR2_X1 U11408 ( .A(n9176), .B(n9162), .ZN(n11294) );
  NAND2_X1 U11409 ( .A1(n11294), .A2(n11887), .ZN(n9164) );
  OR2_X1 U11410 ( .A1(n6570), .A2(n11295), .ZN(n9163) );
  XNOR2_X1 U11411 ( .A(n9301), .B(n10473), .ZN(n9170) );
  NAND2_X1 U11412 ( .A1(n9165), .A2(n11777), .ZN(n9180) );
  OR2_X1 U11413 ( .A1(n9165), .A2(n11777), .ZN(n9166) );
  NAND2_X1 U11414 ( .A1(n9180), .A2(n9166), .ZN(n12461) );
  INV_X1 U11415 ( .A(n9354), .ZN(n9252) );
  INV_X1 U11416 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U11417 ( .A1(n8790), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U11418 ( .A1(n8788), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9167) );
  OAI211_X1 U11419 ( .C1(n9252), .C2(n12729), .A(n9168), .B(n9167), .ZN(n9169)
         );
  NAND2_X1 U11420 ( .A1(n9170), .A2(n12473), .ZN(n9174) );
  INV_X1 U11421 ( .A(n9170), .ZN(n9171) );
  INV_X1 U11422 ( .A(n12473), .ZN(n12096) );
  NAND2_X1 U11423 ( .A1(n9171), .A2(n12096), .ZN(n9172) );
  AND2_X1 U11424 ( .A1(n9174), .A2(n9172), .ZN(n11772) );
  NAND2_X1 U11425 ( .A1(n13413), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U11426 ( .A1(n14568), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9177) );
  AOI22_X1 U11427 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(
        P2_DATAO_REG_26__SCAN_IN), .B1(n14565), .B2(n13410), .ZN(n9178) );
  OR2_X1 U11428 ( .A1(n6570), .A2(n11401), .ZN(n9179) );
  XNOR2_X1 U11429 ( .A(n12727), .B(n10473), .ZN(n9187) );
  NAND2_X1 U11430 ( .A1(n9180), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9181) );
  NAND2_X1 U11431 ( .A1(n9196), .A2(n9181), .ZN(n12446) );
  NAND2_X1 U11432 ( .A1(n12446), .A2(n8789), .ZN(n9186) );
  INV_X1 U11433 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12725) );
  NAND2_X1 U11434 ( .A1(n8790), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9183) );
  NAND2_X1 U11435 ( .A1(n8788), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9182) );
  OAI211_X1 U11436 ( .C1(n9252), .C2(n12725), .A(n9183), .B(n9182), .ZN(n9184)
         );
  INV_X1 U11437 ( .A(n9184), .ZN(n9185) );
  NOR2_X1 U11438 ( .A1(n9187), .A2(n12095), .ZN(n9188) );
  AOI21_X1 U11439 ( .B1(n9187), .B2(n12095), .A(n9188), .ZN(n11856) );
  INV_X1 U11440 ( .A(n9207), .ZN(n9205) );
  AND2_X1 U11441 ( .A1(n14565), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9189) );
  NAND2_X1 U11442 ( .A1(n13410), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9191) );
  AOI22_X1 U11443 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(
        P2_DATAO_REG_27__SCAN_IN), .B1(n14562), .B2(n13408), .ZN(n9192) );
  INV_X1 U11444 ( .A(n9192), .ZN(n9193) );
  XNOR2_X1 U11445 ( .A(n9279), .B(n9193), .ZN(n11494) );
  NAND2_X1 U11446 ( .A1(n11494), .A2(n11887), .ZN(n9195) );
  OR2_X1 U11447 ( .A1(n6570), .A2(n11495), .ZN(n9194) );
  XNOR2_X1 U11448 ( .A(n9349), .B(n8803), .ZN(n11707) );
  INV_X1 U11449 ( .A(n9247), .ZN(n9198) );
  NAND2_X1 U11450 ( .A1(n9196), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9197) );
  NAND2_X1 U11451 ( .A1(n9198), .A2(n9197), .ZN(n12435) );
  NAND2_X1 U11452 ( .A1(n12435), .A2(n8789), .ZN(n9203) );
  INV_X1 U11453 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12722) );
  NAND2_X1 U11454 ( .A1(n8788), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9200) );
  NAND2_X1 U11455 ( .A1(n8790), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9199) );
  OAI211_X1 U11456 ( .C1(n12722), .C2(n9252), .A(n9200), .B(n9199), .ZN(n9201)
         );
  INV_X1 U11457 ( .A(n9201), .ZN(n9202) );
  NOR2_X1 U11458 ( .A1(n11707), .A2(n12094), .ZN(n11703) );
  AOI21_X1 U11459 ( .B1(n11707), .B2(n12094), .A(n11703), .ZN(n9206) );
  NAND2_X1 U11460 ( .A1(n9205), .A2(n9204), .ZN(n9208) );
  NAND2_X1 U11461 ( .A1(n9208), .A2(n11713), .ZN(n9234) );
  INV_X1 U11462 ( .A(n9376), .ZN(n12773) );
  NAND2_X1 U11463 ( .A1(n11402), .A2(n11297), .ZN(n9210) );
  NOR4_X1 U11464 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9220) );
  NOR4_X1 U11465 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9215) );
  NOR4_X1 U11466 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9214) );
  NOR4_X1 U11467 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9213) );
  NOR4_X1 U11468 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9212) );
  NAND4_X1 U11469 ( .A1(n9215), .A2(n9214), .A3(n9213), .A4(n9212), .ZN(n9216)
         );
  NOR4_X1 U11470 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        n9217), .A4(n9216), .ZN(n9219) );
  NOR4_X1 U11471 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n9218) );
  AND3_X1 U11472 ( .A1(n9220), .A2(n9219), .A3(n9218), .ZN(n9221) );
  OR2_X1 U11473 ( .A1(n9209), .A2(n9221), .ZN(n9377) );
  NAND2_X1 U11474 ( .A1(n11932), .A2(n10403), .ZN(n9381) );
  INV_X1 U11475 ( .A(n14790), .ZN(n12086) );
  XNOR2_X1 U11476 ( .A(n9381), .B(n12086), .ZN(n9226) );
  NAND2_X1 U11477 ( .A1(n11932), .A2(n14638), .ZN(n9225) );
  NAND2_X1 U11478 ( .A1(n9226), .A2(n9225), .ZN(n9362) );
  NAND2_X1 U11479 ( .A1(n9362), .A2(n12621), .ZN(n10467) );
  NAND2_X1 U11480 ( .A1(n9376), .A2(n9377), .ZN(n9227) );
  OR2_X1 U11481 ( .A1(n14790), .A2(n14638), .ZN(n9383) );
  INV_X1 U11482 ( .A(n9383), .ZN(n9229) );
  NAND2_X1 U11483 ( .A1(n9229), .A2(n9228), .ZN(n9365) );
  OAI22_X1 U11484 ( .A1(n9367), .A2(n10467), .B1(n9364), .B2(n9365), .ZN(n9233) );
  INV_X1 U11485 ( .A(n8726), .ZN(n9231) );
  NOR2_X1 U11486 ( .A1(n11402), .A2(n11297), .ZN(n9230) );
  NAND2_X1 U11487 ( .A1(n9234), .A2(n11863), .ZN(n9266) );
  NAND2_X1 U11488 ( .A1(n10160), .A2(n14898), .ZN(n9235) );
  OR2_X1 U11489 ( .A1(n9367), .A2(n9235), .ZN(n9237) );
  INV_X1 U11490 ( .A(n10705), .ZN(n12076) );
  NOR2_X1 U11491 ( .A1(n12621), .A2(n12076), .ZN(n9236) );
  NAND2_X1 U11492 ( .A1(n9367), .A2(n9362), .ZN(n9242) );
  OAI211_X1 U11493 ( .C1(n9382), .C2(n12044), .A(n9420), .B(n10161), .ZN(n9238) );
  INV_X1 U11494 ( .A(n9238), .ZN(n9241) );
  INV_X1 U11495 ( .A(n9365), .ZN(n9239) );
  NAND2_X1 U11496 ( .A1(n9364), .A2(n9239), .ZN(n9240) );
  NAND3_X1 U11497 ( .A1(n9242), .A2(n9241), .A3(n9240), .ZN(n9243) );
  NAND2_X1 U11498 ( .A1(n9243), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9245) );
  NAND2_X1 U11499 ( .A1(n10160), .A2(n9382), .ZN(n9259) );
  NAND2_X1 U11500 ( .A1(n9364), .A2(n9368), .ZN(n9244) );
  INV_X1 U11501 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9246) );
  NOR2_X1 U11502 ( .A1(n9247), .A2(n9246), .ZN(n9248) );
  INV_X1 U11503 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U11504 ( .A1(n8790), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9250) );
  NAND2_X1 U11505 ( .A1(n8788), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9249) );
  OAI211_X1 U11506 ( .C1(n9252), .C2(n9251), .A(n9250), .B(n9249), .ZN(n9253)
         );
  INV_X1 U11507 ( .A(n9364), .ZN(n9257) );
  INV_X1 U11508 ( .A(n9254), .ZN(n12083) );
  NAND2_X1 U11509 ( .A1(n12083), .A2(n10182), .ZN(n10164) );
  NAND2_X1 U11510 ( .A1(n10163), .A2(n10164), .ZN(n9258) );
  NOR2_X1 U11511 ( .A1(n12589), .A2(n9259), .ZN(n9256) );
  NAND2_X1 U11512 ( .A1(n9257), .A2(n9256), .ZN(n11870) );
  INV_X1 U11513 ( .A(n9259), .ZN(n12084) );
  NAND2_X1 U11514 ( .A1(n12631), .A2(n12084), .ZN(n9260) );
  INV_X2 U11515 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  AOI22_X1 U11516 ( .A1(n12095), .A2(n11868), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9261) );
  OAI21_X1 U11517 ( .B1(n6575), .B2(n11870), .A(n9261), .ZN(n9262) );
  AOI21_X1 U11518 ( .B1(n12435), .B2(n11872), .A(n9262), .ZN(n9263) );
  INV_X1 U11519 ( .A(n9264), .ZN(n9265) );
  NAND2_X1 U11520 ( .A1(n9266), .A2(n9265), .ZN(P3_U3154) );
  INV_X1 U11521 ( .A(n10704), .ZN(n9306) );
  NAND2_X1 U11522 ( .A1(n12106), .A2(n9306), .ZN(n11941) );
  NAND2_X1 U11523 ( .A1(n11942), .A2(n11941), .ZN(n9305) );
  NAND2_X1 U11524 ( .A1(n9268), .A2(n10934), .ZN(n11946) );
  NAND2_X1 U11525 ( .A1(n10964), .A2(n9311), .ZN(n11945) );
  NAND2_X1 U11526 ( .A1(n10663), .A2(n9309), .ZN(n10662) );
  NAND2_X1 U11527 ( .A1(n10662), .A2(n11945), .ZN(n10824) );
  NAND2_X1 U11528 ( .A1(n11106), .A2(n10831), .ZN(n11951) );
  INV_X1 U11529 ( .A(n10831), .ZN(n10963) );
  NAND2_X1 U11530 ( .A1(n12105), .A2(n10963), .ZN(n11952) );
  NAND2_X1 U11531 ( .A1(n11951), .A2(n11952), .ZN(n11911) );
  NAND2_X1 U11532 ( .A1(n11206), .A2(n11112), .ZN(n11956) );
  INV_X1 U11533 ( .A(n11112), .ZN(n11100) );
  NAND2_X1 U11534 ( .A1(n12104), .A2(n11100), .ZN(n11955) );
  NAND2_X1 U11535 ( .A1(n11288), .A2(n9315), .ZN(n11959) );
  NAND2_X1 U11536 ( .A1(n12103), .A2(n11205), .ZN(n11960) );
  INV_X1 U11537 ( .A(n11912), .ZN(n11962) );
  INV_X1 U11538 ( .A(n12102), .ZN(n11394) );
  INV_X1 U11539 ( .A(n11965), .ZN(n9319) );
  NAND2_X1 U11540 ( .A1(n11394), .A2(n9319), .ZN(n11966) );
  NAND2_X1 U11541 ( .A1(n11278), .A2(n11966), .ZN(n11366) );
  XNOR2_X1 U11542 ( .A(n12101), .B(n9320), .ZN(n11969) );
  NAND2_X1 U11543 ( .A1(n11366), .A2(n11969), .ZN(n11368) );
  NAND2_X1 U11544 ( .A1(n11564), .A2(n9320), .ZN(n11973) );
  NAND2_X1 U11545 ( .A1(n11350), .A2(n11977), .ZN(n9269) );
  NAND2_X1 U11546 ( .A1(n11836), .A2(n11472), .ZN(n11987) );
  INV_X1 U11547 ( .A(n11472), .ZN(n11608) );
  NAND2_X1 U11548 ( .A1(n12099), .A2(n11608), .ZN(n11410) );
  INV_X1 U11549 ( .A(n11980), .ZN(n9271) );
  NAND2_X1 U11550 ( .A1(n11832), .A2(n11414), .ZN(n11984) );
  INV_X1 U11551 ( .A(n11414), .ZN(n11835) );
  NAND2_X1 U11552 ( .A1(n12632), .A2(n11835), .ZN(n11990) );
  INV_X1 U11553 ( .A(n11410), .ZN(n9272) );
  NOR2_X1 U11554 ( .A1(n11917), .A2(n9272), .ZN(n11983) );
  NAND2_X1 U11555 ( .A1(n11412), .A2(n11984), .ZN(n12643) );
  NAND2_X1 U11556 ( .A1(n11820), .A2(n12637), .ZN(n11993) );
  NAND2_X1 U11557 ( .A1(n12616), .A2(n11765), .ZN(n11989) );
  NAND2_X1 U11558 ( .A1(n11993), .A2(n11989), .ZN(n12642) );
  INV_X1 U11559 ( .A(n12642), .ZN(n12630) );
  NOR2_X1 U11560 ( .A1(n12622), .A2(n12634), .ZN(n11998) );
  NAND2_X1 U11561 ( .A1(n12622), .A2(n12634), .ZN(n11916) );
  OR2_X1 U11562 ( .A1(n12769), .A2(n12617), .ZN(n12001) );
  NAND2_X1 U11563 ( .A1(n12769), .A2(n12617), .ZN(n12002) );
  INV_X1 U11564 ( .A(n12603), .ZN(n11733) );
  OR2_X1 U11565 ( .A1(n11862), .A2(n11733), .ZN(n12005) );
  NAND2_X1 U11566 ( .A1(n11862), .A2(n11733), .ZN(n12004) );
  OR2_X1 U11567 ( .A1(n12701), .A2(n12588), .ZN(n12011) );
  NAND2_X1 U11568 ( .A1(n12701), .A2(n12588), .ZN(n12012) );
  NAND2_X1 U11569 ( .A1(n12011), .A2(n12012), .ZN(n9335) );
  NAND2_X1 U11570 ( .A1(n12574), .A2(n12573), .ZN(n12576) );
  NAND2_X1 U11571 ( .A1(n12576), .A2(n12012), .ZN(n12562) );
  OR2_X1 U11572 ( .A1(n12697), .A2(n12548), .ZN(n12016) );
  NAND2_X1 U11573 ( .A1(n12697), .A2(n12548), .ZN(n12020) );
  NAND2_X1 U11574 ( .A1(n12016), .A2(n12020), .ZN(n12013) );
  NAND2_X1 U11575 ( .A1(n12562), .A2(n12561), .ZN(n12560) );
  NAND2_X1 U11576 ( .A1(n12550), .A2(n9274), .ZN(n12019) );
  NAND2_X1 U11577 ( .A1(n12755), .A2(n12098), .ZN(n12025) );
  OR2_X1 U11578 ( .A1(n12755), .A2(n12098), .ZN(n12024) );
  NAND2_X1 U11579 ( .A1(n12524), .A2(n12509), .ZN(n12030) );
  NAND2_X1 U11580 ( .A1(n12029), .A2(n12030), .ZN(n12519) );
  NAND2_X1 U11581 ( .A1(n12516), .A2(n12522), .ZN(n12034) );
  INV_X1 U11582 ( .A(n12507), .ZN(n11756) );
  NAND2_X1 U11583 ( .A1(n11829), .A2(n11756), .ZN(n11908) );
  NOR2_X1 U11584 ( .A1(n11829), .A2(n11756), .ZN(n12039) );
  NAND2_X1 U11585 ( .A1(n11742), .A2(n12495), .ZN(n9276) );
  NAND2_X1 U11586 ( .A1(n12042), .A2(n9276), .ZN(n12483) );
  OR2_X1 U11587 ( .A1(n12478), .A2(n12487), .ZN(n12043) );
  NAND2_X1 U11588 ( .A1(n12478), .A2(n12487), .ZN(n9277) );
  NAND2_X1 U11589 ( .A1(n12043), .A2(n9277), .ZN(n12469) );
  NOR2_X1 U11590 ( .A1(n12467), .A2(n12469), .ZN(n12466) );
  INV_X1 U11591 ( .A(n9277), .ZN(n12046) );
  OR2_X1 U11592 ( .A1(n9301), .A2(n12473), .ZN(n12050) );
  NAND2_X1 U11593 ( .A1(n9301), .A2(n12473), .ZN(n9278) );
  NAND2_X1 U11594 ( .A1(n12050), .A2(n9278), .ZN(n12458) );
  INV_X1 U11595 ( .A(n9278), .ZN(n12052) );
  NOR2_X1 U11596 ( .A1(n9348), .A2(n12456), .ZN(n12057) );
  NAND2_X1 U11597 ( .A1(n9348), .A2(n12456), .ZN(n12055) );
  XNOR2_X1 U11598 ( .A(n9349), .B(n12443), .ZN(n12428) );
  INV_X1 U11599 ( .A(n12428), .ZN(n11907) );
  AND2_X1 U11600 ( .A1(n9349), .A2(n12443), .ZN(n12064) );
  INV_X1 U11601 ( .A(n9279), .ZN(n9281) );
  NAND2_X1 U11602 ( .A1(n13408), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9280) );
  NAND2_X1 U11603 ( .A1(n9281), .A2(n9280), .ZN(n9283) );
  NAND2_X1 U11604 ( .A1(n14562), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9282) );
  INV_X1 U11605 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13407) );
  INV_X1 U11606 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13677) );
  AOI22_X1 U11607 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(
        P1_DATAO_REG_28__SCAN_IN), .B1(n13407), .B2(n13677), .ZN(n9284) );
  XNOR2_X1 U11608 ( .A(n9288), .B(n9284), .ZN(n11695) );
  NAND2_X1 U11609 ( .A1(n11695), .A2(n11887), .ZN(n9286) );
  OR2_X1 U11610 ( .A1(n6569), .A2(n11697), .ZN(n9285) );
  NAND2_X1 U11611 ( .A1(n12652), .A2(n6575), .ZN(n12061) );
  NOR2_X1 U11612 ( .A1(n13407), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9287) );
  NAND2_X1 U11613 ( .A1(n13407), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9289) );
  XNOR2_X1 U11614 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n11722) );
  XNOR2_X1 U11615 ( .A(n11723), .B(n11722), .ZN(n12780) );
  NOR2_X1 U11616 ( .A1(n6569), .A2(n12783), .ZN(n9290) );
  NAND2_X1 U11617 ( .A1(n12408), .A2(n8789), .ZN(n11894) );
  INV_X1 U11618 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11619 ( .A1(n9354), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U11620 ( .A1(n8790), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9291) );
  OAI211_X1 U11621 ( .C1(n9293), .C2(n7009), .A(n9292), .B(n9291), .ZN(n9294)
         );
  INV_X1 U11622 ( .A(n9294), .ZN(n9295) );
  NAND2_X1 U11623 ( .A1(n11894), .A2(n9295), .ZN(n12092) );
  NOR2_X1 U11624 ( .A1(n11718), .A2(n12092), .ZN(n11895) );
  INV_X1 U11625 ( .A(n11718), .ZN(n9296) );
  INV_X1 U11626 ( .A(n12092), .ZN(n12413) );
  NOR2_X1 U11627 ( .A1(n9296), .A2(n12413), .ZN(n11876) );
  NOR2_X1 U11628 ( .A1(n11895), .A2(n11876), .ZN(n9351) );
  INV_X1 U11629 ( .A(n9351), .ZN(n9297) );
  AND2_X1 U11630 ( .A1(n12621), .A2(n9382), .ZN(n9298) );
  NAND2_X1 U11631 ( .A1(n9362), .A2(n9298), .ZN(n9300) );
  NAND2_X1 U11632 ( .A1(n9353), .A2(n14638), .ZN(n9299) );
  OR2_X1 U11633 ( .A1(n14790), .A2(n9299), .ZN(n9380) );
  NAND2_X1 U11634 ( .A1(n10705), .A2(n14790), .ZN(n12656) );
  NAND2_X1 U11635 ( .A1(n10708), .A2(n9302), .ZN(n9303) );
  NAND2_X1 U11636 ( .A1(n9304), .A2(n9303), .ZN(n10706) );
  NAND2_X1 U11637 ( .A1(n8812), .A2(n9306), .ZN(n9307) );
  NAND2_X1 U11638 ( .A1(n9268), .A2(n9311), .ZN(n9312) );
  NAND2_X1 U11639 ( .A1(n10664), .A2(n9312), .ZN(n10826) );
  NAND2_X1 U11640 ( .A1(n12105), .A2(n10831), .ZN(n9313) );
  NAND2_X1 U11641 ( .A1(n11206), .A2(n11100), .ZN(n9314) );
  NAND2_X1 U11642 ( .A1(n12103), .A2(n9315), .ZN(n9316) );
  NAND2_X1 U11643 ( .A1(n11564), .A2(n11971), .ZN(n9318) );
  AND2_X1 U11644 ( .A1(n11912), .A2(n9318), .ZN(n9317) );
  INV_X1 U11645 ( .A(n9318), .ZN(n9323) );
  NAND2_X1 U11646 ( .A1(n12102), .A2(n9319), .ZN(n11363) );
  NAND2_X1 U11647 ( .A1(n12101), .A2(n9320), .ZN(n9321) );
  AND2_X1 U11648 ( .A1(n11363), .A2(n9321), .ZN(n9322) );
  OR2_X1 U11649 ( .A1(n9323), .A2(n9322), .ZN(n9324) );
  XNOR2_X1 U11650 ( .A(n12100), .B(n11979), .ZN(n11352) );
  NAND2_X1 U11651 ( .A1(n12099), .A2(n11472), .ZN(n9325) );
  NAND2_X1 U11652 ( .A1(n12629), .A2(n12642), .ZN(n9327) );
  NAND2_X1 U11653 ( .A1(n12616), .A2(n12637), .ZN(n9326) );
  NOR2_X1 U11654 ( .A1(n9329), .A2(n12622), .ZN(n9328) );
  NAND2_X1 U11655 ( .A1(n9329), .A2(n12622), .ZN(n9330) );
  OR2_X1 U11656 ( .A1(n12769), .A2(n12586), .ZN(n9331) );
  OR2_X1 U11657 ( .A1(n11862), .A2(n12603), .ZN(n9332) );
  NAND2_X1 U11658 ( .A1(n12583), .A2(n9332), .ZN(n9334) );
  NAND2_X1 U11659 ( .A1(n11862), .A2(n12603), .ZN(n9333) );
  NAND2_X1 U11660 ( .A1(n9334), .A2(n9333), .ZN(n12568) );
  NAND2_X1 U11661 ( .A1(n12568), .A2(n9335), .ZN(n9337) );
  NAND2_X1 U11662 ( .A1(n12701), .A2(n12557), .ZN(n9336) );
  NAND2_X1 U11663 ( .A1(n9337), .A2(n9336), .ZN(n12556) );
  NAND2_X1 U11664 ( .A1(n12697), .A2(n12570), .ZN(n9338) );
  OR2_X1 U11665 ( .A1(n12550), .A2(n12558), .ZN(n9341) );
  OR2_X1 U11666 ( .A1(n12755), .A2(n12549), .ZN(n9343) );
  NAND2_X1 U11667 ( .A1(n12033), .A2(n12034), .ZN(n12503) );
  INV_X1 U11668 ( .A(n12516), .ZN(n12747) );
  NAND2_X1 U11669 ( .A1(n11829), .A2(n12507), .ZN(n9345) );
  NAND2_X1 U11670 ( .A1(n11742), .A2(n9346), .ZN(n9347) );
  NAND2_X1 U11671 ( .A1(n12482), .A2(n9347), .ZN(n12470) );
  NAND2_X1 U11672 ( .A1(n12468), .A2(n7886), .ZN(n12452) );
  INV_X1 U11673 ( .A(n6575), .ZN(n12093) );
  XNOR2_X1 U11674 ( .A(n9352), .B(n9351), .ZN(n9361) );
  NAND2_X1 U11675 ( .A1(n10582), .A2(n9353), .ZN(n11905) );
  INV_X1 U11676 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n14896) );
  NAND2_X1 U11677 ( .A1(n9354), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U11678 ( .A1(n8788), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9355) );
  OAI211_X1 U11679 ( .C1(n14896), .C2(n8962), .A(n9356), .B(n9355), .ZN(n9357)
         );
  INV_X1 U11680 ( .A(n9357), .ZN(n9358) );
  AND2_X1 U11681 ( .A1(n11894), .A2(n9358), .ZN(n11898) );
  AND2_X1 U11682 ( .A1(n12083), .A2(P3_B_REG_SCAN_IN), .ZN(n9359) );
  OR2_X1 U11683 ( .A1(n12589), .A2(n9359), .ZN(n12406) );
  OAI22_X1 U11684 ( .A1(n6575), .A2(n12587), .B1(n11898), .B2(n12406), .ZN(
        n9360) );
  INV_X1 U11685 ( .A(n9362), .ZN(n9363) );
  OAI22_X1 U11686 ( .A1(n9367), .A2(n9365), .B1(n9364), .B2(n9363), .ZN(n9366)
         );
  NAND2_X1 U11687 ( .A1(n9366), .A2(n10160), .ZN(n9371) );
  INV_X1 U11688 ( .A(n9367), .ZN(n9369) );
  NAND2_X1 U11689 ( .A1(n9369), .A2(n9368), .ZN(n9370) );
  INV_X1 U11690 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9372) );
  NAND2_X1 U11691 ( .A1(n15601), .A2(n9372), .ZN(n9373) );
  NAND2_X1 U11692 ( .A1(n9374), .A2(n9373), .ZN(n9375) );
  NAND2_X1 U11693 ( .A1(n9375), .A2(n7877), .ZN(P3_U3456) );
  XNOR2_X1 U11694 ( .A(n9376), .B(n12771), .ZN(n9379) );
  INV_X1 U11695 ( .A(n9380), .ZN(n10576) );
  MUX2_X1 U11696 ( .A(n9382), .B(n10576), .S(n12044), .Z(n10578) );
  NAND2_X1 U11697 ( .A1(n9381), .A2(n14790), .ZN(n9384) );
  INV_X1 U11698 ( .A(n9382), .ZN(n12075) );
  NAND3_X1 U11699 ( .A1(n9384), .A2(n12075), .A3(n9383), .ZN(n9385) );
  AND2_X1 U11700 ( .A1(n9385), .A2(n12044), .ZN(n9387) );
  INV_X1 U11701 ( .A(n12771), .ZN(n9386) );
  MUX2_X1 U11702 ( .A(n10578), .B(n9387), .S(n9386), .Z(n9388) );
  NAND2_X1 U11703 ( .A1(n9391), .A2(n7883), .ZN(P3_U3488) );
  NOR2_X1 U11704 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9395) );
  NAND2_X1 U11705 ( .A1(n9414), .A2(n9416), .ZN(n9401) );
  XNOR2_X1 U11706 ( .A(n9400), .B(n9399), .ZN(n14570) );
  NAND2_X1 U11707 ( .A1(n9401), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9403) );
  NOR2_X1 U11708 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9406) );
  NOR2_X1 U11709 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9405) );
  NOR2_X1 U11710 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n9404) );
  NOR2_X1 U11711 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n9407) );
  INV_X1 U11712 ( .A(n9410), .ZN(n9411) );
  OAI21_X1 U11713 ( .B1(n9409), .B2(n9411), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9412) );
  MUX2_X1 U11714 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9412), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9413) );
  INV_X1 U11715 ( .A(n9414), .ZN(n9415) );
  NAND2_X1 U11716 ( .A1(n9415), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9417) );
  NAND3_X1 U11717 ( .A1(n13414), .A2(n9419), .A3(n9475), .ZN(n9479) );
  INV_X4 U11718 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U11719 ( .A(n9420), .ZN(n9421) );
  INV_X2 U11720 ( .A(n13397), .ZN(n13417) );
  INV_X2 U11721 ( .A(n13404), .ZN(n13399) );
  INV_X1 U11722 ( .A(n9515), .ZN(n9524) );
  OAI222_X1 U11723 ( .A1(n13417), .A2(n9422), .B1(n13399), .B2(n10021), .C1(
        n9524), .C2(P2_U3088), .ZN(P2_U3326) );
  INV_X1 U11724 ( .A(n14780), .ZN(n14787) );
  OAI222_X1 U11725 ( .A1(n14787), .A2(n9424), .B1(n12784), .B2(n9423), .C1(
        P3_U3151), .C2(n14601), .ZN(P3_U3287) );
  OAI222_X1 U11726 ( .A1(P3_U3151), .A2(n15402), .B1(n14787), .B2(n9425), .C1(
        n9962), .C2(n12784), .ZN(P3_U3295) );
  INV_X1 U11727 ( .A(n10071), .ZN(n9450) );
  INV_X1 U11728 ( .A(n9531), .ZN(n9542) );
  OAI222_X1 U11729 ( .A1(n13417), .A2(n9426), .B1(n13399), .B2(n9450), .C1(
        n9542), .C2(P2_U3088), .ZN(P2_U3325) );
  OAI222_X1 U11730 ( .A1(n14787), .A2(n9428), .B1(n12784), .B2(n9427), .C1(
        P3_U3151), .C2(n10279), .ZN(P3_U3294) );
  OAI222_X1 U11731 ( .A1(P3_U3151), .A2(n10547), .B1(n14787), .B2(n9430), .C1(
        n9429), .C2(n12784), .ZN(P3_U3289) );
  INV_X1 U11732 ( .A(n12784), .ZN(n14779) );
  AOI222_X1 U11733 ( .A1(n9431), .A2(n14780), .B1(SI_7_), .B2(n14779), .C1(
        n12381), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9432) );
  INV_X1 U11734 ( .A(n9432), .ZN(P3_U3288) );
  AOI222_X1 U11735 ( .A1(n9433), .A2(n14780), .B1(SI_9_), .B2(n14779), .C1(
        n14642), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9434) );
  INV_X1 U11736 ( .A(n9434), .ZN(P3_U3286) );
  AOI222_X1 U11737 ( .A1(n9435), .A2(n14780), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15418), .C1(SI_3_), .C2(n14779), .ZN(n9436) );
  INV_X1 U11738 ( .A(n9436), .ZN(P3_U3292) );
  AOI222_X1 U11739 ( .A1(n9437), .A2(n14780), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10371), .C1(SI_2_), .C2(n14779), .ZN(n9438) );
  INV_X1 U11740 ( .A(n9438), .ZN(P3_U3293) );
  AOI222_X1 U11741 ( .A1(n9439), .A2(n14780), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10375), .C1(SI_4_), .C2(n14779), .ZN(n9440) );
  INV_X1 U11742 ( .A(n9440), .ZN(P3_U3291) );
  AOI222_X1 U11743 ( .A1(n9441), .A2(n14780), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10378), .C1(SI_5_), .C2(n14779), .ZN(n9442) );
  INV_X1 U11744 ( .A(n9442), .ZN(P3_U3290) );
  NAND2_X2 U11745 ( .A1(n6568), .A2(P1_U3086), .ZN(n14571) );
  INV_X1 U11746 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9444) );
  NAND2_X1 U11747 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9443) );
  XNOR2_X1 U11748 ( .A(n9444), .B(n9443), .ZN(n14069) );
  OAI222_X1 U11749 ( .A1(n14571), .A2(n7606), .B1(n11699), .B2(n10021), .C1(
        P1_U3086), .C2(n14069), .ZN(P1_U3354) );
  AOI222_X1 U11750 ( .A1(n9445), .A2(n14780), .B1(SI_10_), .B2(n14779), .C1(
        n14644), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9446) );
  INV_X1 U11751 ( .A(n9446), .ZN(P3_U3285) );
  INV_X1 U11752 ( .A(n10215), .ZN(n9456) );
  INV_X1 U11753 ( .A(n9562), .ZN(n9511) );
  OAI222_X1 U11754 ( .A1(n13417), .A2(n9447), .B1(n13399), .B2(n9456), .C1(
        P2_U3088), .C2(n9511), .ZN(P2_U3324) );
  OR2_X1 U11755 ( .A1(n9448), .A2(n10335), .ZN(n9449) );
  XNOR2_X1 U11756 ( .A(n9449), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14088) );
  INV_X1 U11757 ( .A(n14088), .ZN(n9451) );
  OAI222_X1 U11758 ( .A1(P1_U3086), .A2(n9451), .B1(n11699), .B2(n9450), .C1(
        n7591), .C2(n14571), .ZN(P1_U3353) );
  NAND2_X1 U11759 ( .A1(n9452), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9453) );
  MUX2_X1 U11760 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9453), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9454) );
  OR2_X1 U11761 ( .A1(n9452), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9468) );
  INV_X1 U11762 ( .A(n14102), .ZN(n9457) );
  INV_X1 U11763 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9455) );
  OAI222_X1 U11764 ( .A1(n9457), .A2(P1_U3086), .B1(n11699), .B2(n9456), .C1(
        n9455), .C2(n14571), .ZN(P1_U3352) );
  INV_X1 U11765 ( .A(n9458), .ZN(n9459) );
  OAI222_X1 U11766 ( .A1(P3_U3151), .A2(n15501), .B1(n12784), .B2(n9460), .C1(
        n14787), .C2(n9459), .ZN(P3_U3284) );
  AOI22_X1 U11767 ( .A1(n9583), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n13397), .ZN(n9462) );
  OAI21_X1 U11768 ( .B1(n9461), .B2(n13399), .A(n9462), .ZN(P2_U3322) );
  NAND2_X1 U11769 ( .A1(n9468), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9463) );
  XNOR2_X1 U11770 ( .A(n9463), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14994) );
  INV_X1 U11771 ( .A(n14994), .ZN(n9465) );
  INV_X1 U11772 ( .A(n10216), .ZN(n9466) );
  INV_X1 U11773 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9464) );
  OAI222_X1 U11774 ( .A1(n9465), .A2(P1_U3086), .B1(n11699), .B2(n9466), .C1(
        n9464), .C2(n14571), .ZN(P1_U3351) );
  INV_X1 U11775 ( .A(n9599), .ZN(n9609) );
  OAI222_X1 U11776 ( .A1(n13417), .A2(n9467), .B1(n13399), .B2(n9466), .C1(
        P2_U3088), .C2(n9609), .ZN(P2_U3323) );
  INV_X1 U11777 ( .A(n9468), .ZN(n9470) );
  NAND2_X1 U11778 ( .A1(n9470), .A2(n9469), .ZN(n9543) );
  NAND2_X1 U11779 ( .A1(n9543), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9471) );
  XNOR2_X1 U11780 ( .A(n9471), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10408) );
  INV_X1 U11781 ( .A(n10408), .ZN(n9806) );
  INV_X1 U11782 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9472) );
  OAI222_X1 U11783 ( .A1(P1_U3086), .A2(n9806), .B1(n11699), .B2(n9461), .C1(
        n9472), .C2(n14571), .ZN(P1_U3350) );
  OAI222_X1 U11784 ( .A1(n12784), .A2(n9474), .B1(n14787), .B2(n9473), .C1(
        n15519), .C2(P3_U3151), .ZN(P3_U3283) );
  NAND2_X1 U11785 ( .A1(n9475), .A2(n9703), .ZN(n9477) );
  NAND2_X1 U11786 ( .A1(n9477), .A2(n7923), .ZN(n9478) );
  NAND2_X1 U11787 ( .A1(n9479), .A2(n9478), .ZN(n9493) );
  INV_X1 U11788 ( .A(n9704), .ZN(n9480) );
  AND2_X1 U11789 ( .A1(n9493), .A2(n9480), .ZN(n15277) );
  NAND2_X1 U11790 ( .A1(n9704), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13405) );
  NOR2_X1 U11791 ( .A1(n13405), .A2(n13409), .ZN(n9481) );
  NAND2_X1 U11792 ( .A1(n9493), .A2(n9481), .ZN(n15270) );
  INV_X1 U11793 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10207) );
  MUX2_X1 U11794 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10207), .S(n9562), .Z(n9487) );
  INV_X1 U11795 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9532) );
  MUX2_X1 U11796 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9532), .S(n9531), .Z(n9485)
         );
  INV_X1 U11797 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9516) );
  MUX2_X1 U11798 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9516), .S(n9515), .Z(n9483)
         );
  AND2_X1 U11799 ( .A1(n15229), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U11800 ( .A1(n9483), .A2(n9482), .ZN(n9534) );
  NAND2_X1 U11801 ( .A1(n9515), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9533) );
  NAND2_X1 U11802 ( .A1(n9534), .A2(n9533), .ZN(n9484) );
  NAND2_X1 U11803 ( .A1(n9485), .A2(n9484), .ZN(n9536) );
  NAND2_X1 U11804 ( .A1(n9531), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U11805 ( .A1(n9536), .A2(n9488), .ZN(n9486) );
  NAND2_X1 U11806 ( .A1(n9487), .A2(n9486), .ZN(n9602) );
  MUX2_X1 U11807 ( .A(n10207), .B(P2_REG2_REG_3__SCAN_IN), .S(n9562), .Z(n9489) );
  NAND3_X1 U11808 ( .A1(n9489), .A2(n9536), .A3(n9488), .ZN(n9490) );
  NAND2_X1 U11809 ( .A1(n9602), .A2(n9490), .ZN(n9491) );
  NOR2_X1 U11810 ( .A1(n15270), .A2(n9491), .ZN(n9509) );
  INV_X1 U11811 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9507) );
  INV_X1 U11812 ( .A(n13409), .ZN(n13032) );
  NOR2_X1 U11813 ( .A1(n13405), .A2(n13032), .ZN(n9492) );
  NAND2_X1 U11814 ( .A1(n9493), .A2(n9492), .ZN(n15265) );
  INV_X1 U11815 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9494) );
  MUX2_X1 U11816 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9494), .S(n9562), .Z(n9502)
         );
  INV_X1 U11817 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9495) );
  MUX2_X1 U11818 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9495), .S(n9531), .Z(n9500)
         );
  INV_X1 U11819 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9496) );
  MUX2_X1 U11820 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9496), .S(n9515), .Z(n9498)
         );
  AND2_X1 U11821 ( .A1(n15229), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U11822 ( .A1(n9498), .A2(n9497), .ZN(n9526) );
  NAND2_X1 U11823 ( .A1(n9515), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9525) );
  NAND2_X1 U11824 ( .A1(n9526), .A2(n9525), .ZN(n9499) );
  NAND2_X1 U11825 ( .A1(n9500), .A2(n9499), .ZN(n9528) );
  NAND2_X1 U11826 ( .A1(n9531), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U11827 ( .A1(n9528), .A2(n9503), .ZN(n9501) );
  NAND2_X1 U11828 ( .A1(n9502), .A2(n9501), .ZN(n9595) );
  MUX2_X1 U11829 ( .A(n9494), .B(P2_REG1_REG_3__SCAN_IN), .S(n9562), .Z(n9504)
         );
  NAND3_X1 U11830 ( .A1(n9504), .A2(n9528), .A3(n9503), .ZN(n9505) );
  NAND2_X1 U11831 ( .A1(n9595), .A2(n9505), .ZN(n9506) );
  OAI22_X1 U11832 ( .A1(n15260), .A2(n9507), .B1(n15265), .B2(n9506), .ZN(
        n9508) );
  AOI211_X1 U11833 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(P2_U3088), .A(n9509), 
        .B(n9508), .ZN(n9510) );
  OAI21_X1 U11834 ( .B1(n9511), .B2(n15262), .A(n9510), .ZN(P2_U3217) );
  INV_X1 U11835 ( .A(n15260), .ZN(n15299) );
  MUX2_X1 U11836 ( .A(n9496), .B(P2_REG1_REG_1__SCAN_IN), .S(n9515), .Z(n9512)
         );
  OAI21_X1 U11837 ( .B1(n7908), .B2(n9518), .A(n9512), .ZN(n9513) );
  NAND2_X1 U11838 ( .A1(n9513), .A2(n9526), .ZN(n9514) );
  NOR2_X1 U11839 ( .A1(n15265), .A2(n9514), .ZN(n9522) );
  INV_X1 U11840 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9949) );
  MUX2_X1 U11841 ( .A(n9516), .B(P2_REG2_REG_1__SCAN_IN), .S(n9515), .Z(n9517)
         );
  OAI21_X1 U11842 ( .B1(n9949), .B2(n9518), .A(n9517), .ZN(n9519) );
  NAND2_X1 U11843 ( .A1(n9519), .A2(n9534), .ZN(n9520) );
  INV_X1 U11844 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10257) );
  OAI22_X1 U11845 ( .A1(n15270), .A2(n9520), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10257), .ZN(n9521) );
  AOI211_X1 U11846 ( .C1(n15299), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n9522), .B(
        n9521), .ZN(n9523) );
  OAI21_X1 U11847 ( .B1(n9524), .B2(n15262), .A(n9523), .ZN(P2_U3215) );
  MUX2_X1 U11848 ( .A(n9495), .B(P2_REG1_REG_2__SCAN_IN), .S(n9531), .Z(n9527)
         );
  NAND3_X1 U11849 ( .A1(n9527), .A2(n9526), .A3(n9525), .ZN(n9529) );
  NAND2_X1 U11850 ( .A1(n9529), .A2(n9528), .ZN(n9530) );
  NOR2_X1 U11851 ( .A1(n15265), .A2(n9530), .ZN(n9540) );
  MUX2_X1 U11852 ( .A(n9532), .B(P2_REG2_REG_2__SCAN_IN), .S(n9531), .Z(n9535)
         );
  NAND3_X1 U11853 ( .A1(n9535), .A2(n9534), .A3(n9533), .ZN(n9537) );
  NAND2_X1 U11854 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  INV_X1 U11855 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10395) );
  OAI22_X1 U11856 ( .A1(n15270), .A2(n9538), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10395), .ZN(n9539) );
  AOI211_X1 U11857 ( .C1(n15299), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n9540), .B(
        n9539), .ZN(n9541) );
  OAI21_X1 U11858 ( .B1(n9542), .B2(n15262), .A(n9541), .ZN(P2_U3216) );
  OAI21_X1 U11859 ( .B1(n9543), .B2(P1_IR_REG_5__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9544) );
  MUX2_X1 U11860 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9544), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n9546) );
  AND2_X1 U11861 ( .A1(n9546), .A2(n9545), .ZN(n10853) );
  INV_X1 U11862 ( .A(n10853), .ZN(n9761) );
  INV_X1 U11863 ( .A(n10852), .ZN(n9548) );
  OAI222_X1 U11864 ( .A1(n9761), .A2(P1_U3086), .B1(n11699), .B2(n9548), .C1(
        n9547), .C2(n14571), .ZN(P1_U3349) );
  INV_X1 U11865 ( .A(n9634), .ZN(n9592) );
  OAI222_X1 U11866 ( .A1(n13417), .A2(n9549), .B1(n13399), .B2(n9548), .C1(
        P2_U3088), .C2(n9592), .ZN(P2_U3321) );
  INV_X1 U11867 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9551) );
  INV_X1 U11868 ( .A(n15232), .ZN(n9550) );
  OAI222_X1 U11869 ( .A1(n13417), .A2(n9551), .B1(n13399), .B2(n10857), .C1(
        n9550), .C2(P2_U3088), .ZN(P2_U3320) );
  NAND2_X1 U11870 ( .A1(n9545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9552) );
  XNOR2_X1 U11871 ( .A(n9552), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10858) );
  INV_X1 U11872 ( .A(n10858), .ZN(n9866) );
  OAI222_X1 U11873 ( .A1(P1_U3086), .A2(n9866), .B1(n11699), .B2(n10857), .C1(
        n9553), .C2(n14571), .ZN(P1_U3348) );
  INV_X1 U11874 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15616) );
  NAND2_X1 U11875 ( .A1(n9562), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U11876 ( .A1(n9602), .A2(n9601), .ZN(n9555) );
  INV_X1 U11877 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10438) );
  MUX2_X1 U11878 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10438), .S(n9599), .Z(n9554) );
  NAND2_X1 U11879 ( .A1(n9555), .A2(n9554), .ZN(n9604) );
  NAND2_X1 U11880 ( .A1(n9599), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9559) );
  NAND2_X1 U11881 ( .A1(n9604), .A2(n9559), .ZN(n9557) );
  INV_X1 U11882 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10128) );
  MUX2_X1 U11883 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10128), .S(n9583), .Z(n9556) );
  NAND2_X1 U11884 ( .A1(n9557), .A2(n9556), .ZN(n9588) );
  MUX2_X1 U11885 ( .A(n10128), .B(P2_REG2_REG_5__SCAN_IN), .S(n9583), .Z(n9558) );
  NAND3_X1 U11886 ( .A1(n9604), .A2(n9559), .A3(n9558), .ZN(n9560) );
  NAND2_X1 U11887 ( .A1(n9588), .A2(n9560), .ZN(n9561) );
  OAI22_X1 U11888 ( .A1(n15616), .A2(n15260), .B1(n15270), .B2(n9561), .ZN(
        n9574) );
  INV_X1 U11889 ( .A(n15265), .ZN(n15300) );
  NAND2_X1 U11890 ( .A1(n9562), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9594) );
  NAND2_X1 U11891 ( .A1(n9595), .A2(n9594), .ZN(n9565) );
  INV_X1 U11892 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9563) );
  MUX2_X1 U11893 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9563), .S(n9599), .Z(n9564)
         );
  NAND2_X1 U11894 ( .A1(n9565), .A2(n9564), .ZN(n9597) );
  NAND2_X1 U11895 ( .A1(n9599), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9570) );
  NAND2_X1 U11896 ( .A1(n9597), .A2(n9570), .ZN(n9568) );
  INV_X1 U11897 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9566) );
  MUX2_X1 U11898 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9566), .S(n9583), .Z(n9567)
         );
  NAND2_X1 U11899 ( .A1(n9568), .A2(n9567), .ZN(n9577) );
  MUX2_X1 U11900 ( .A(n9566), .B(P2_REG1_REG_5__SCAN_IN), .S(n9583), .Z(n9569)
         );
  NAND3_X1 U11901 ( .A1(n9597), .A2(n9570), .A3(n9569), .ZN(n9571) );
  NAND3_X1 U11902 ( .A1(n15300), .A2(n9577), .A3(n9571), .ZN(n9572) );
  NAND2_X1 U11903 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10098) );
  NAND2_X1 U11904 ( .A1(n9572), .A2(n10098), .ZN(n9573) );
  AOI211_X1 U11905 ( .C1(n9583), .C2(n15305), .A(n9574), .B(n9573), .ZN(n9575)
         );
  INV_X1 U11906 ( .A(n9575), .ZN(P2_U3219) );
  NAND2_X1 U11907 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10322) );
  NAND2_X1 U11908 ( .A1(n9583), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U11909 ( .A1(n9577), .A2(n9576), .ZN(n9580) );
  INV_X1 U11910 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9578) );
  MUX2_X1 U11911 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9578), .S(n9634), .Z(n9579)
         );
  NAND2_X1 U11912 ( .A1(n9580), .A2(n9579), .ZN(n9628) );
  OAI211_X1 U11913 ( .C1(n9580), .C2(n9579), .A(n15300), .B(n9628), .ZN(n9581)
         );
  NAND2_X1 U11914 ( .A1(n10322), .A2(n9581), .ZN(n9582) );
  AOI21_X1 U11915 ( .B1(n15299), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9582), .ZN(
        n9591) );
  NAND2_X1 U11916 ( .A1(n9583), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U11917 ( .A1(n9588), .A2(n9587), .ZN(n9585) );
  INV_X1 U11918 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10310) );
  MUX2_X1 U11919 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10310), .S(n9634), .Z(n9584) );
  NAND2_X1 U11920 ( .A1(n9585), .A2(n9584), .ZN(n9636) );
  MUX2_X1 U11921 ( .A(n10310), .B(P2_REG2_REG_6__SCAN_IN), .S(n9634), .Z(n9586) );
  NAND3_X1 U11922 ( .A1(n9588), .A2(n9587), .A3(n9586), .ZN(n9589) );
  NAND3_X1 U11923 ( .A1(n15306), .A2(n9636), .A3(n9589), .ZN(n9590) );
  OAI211_X1 U11924 ( .C1(n15262), .C2(n9592), .A(n9591), .B(n9590), .ZN(
        P2_U3220) );
  MUX2_X1 U11925 ( .A(n9563), .B(P2_REG1_REG_4__SCAN_IN), .S(n9599), .Z(n9593)
         );
  NAND3_X1 U11926 ( .A1(n9595), .A2(n9594), .A3(n9593), .ZN(n9596) );
  NAND2_X1 U11927 ( .A1(n9597), .A2(n9596), .ZN(n9598) );
  NOR2_X1 U11928 ( .A1(n15265), .A2(n9598), .ZN(n9607) );
  MUX2_X1 U11929 ( .A(n10438), .B(P2_REG2_REG_4__SCAN_IN), .S(n9599), .Z(n9600) );
  NAND3_X1 U11930 ( .A1(n9602), .A2(n9601), .A3(n9600), .ZN(n9603) );
  NAND3_X1 U11931 ( .A1(n15306), .A2(n9604), .A3(n9603), .ZN(n9605) );
  NAND2_X1 U11932 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U11933 ( .A1(n9605), .A2(n9917), .ZN(n9606) );
  AOI211_X1 U11934 ( .C1(n15299), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n9607), .B(
        n9606), .ZN(n9608) );
  OAI21_X1 U11935 ( .B1(n9609), .B2(n15262), .A(n9608), .ZN(P2_U3218) );
  NOR2_X1 U11936 ( .A1(n9545), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9750) );
  OR2_X1 U11937 ( .A1(n9750), .A2(n10335), .ZN(n9624) );
  XNOR2_X1 U11938 ( .A(n9624), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10871) );
  INV_X1 U11939 ( .A(n14571), .ZN(n9722) );
  AOI22_X1 U11940 ( .A1(n10871), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9722), .ZN(n9610) );
  OAI21_X1 U11941 ( .B1(n10870), .B2(n11699), .A(n9610), .ZN(P1_U3347) );
  INV_X1 U11942 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9611) );
  OAI222_X1 U11943 ( .A1(n13417), .A2(n9611), .B1(n13399), .B2(n10870), .C1(
        n13001), .C2(P2_U3088), .ZN(P2_U3319) );
  NAND2_X1 U11944 ( .A1(n8648), .A2(n12993), .ZN(n9612) );
  OAI21_X1 U11945 ( .B1(n12993), .B2(n8780), .A(n9612), .ZN(P2_U3531) );
  OAI222_X1 U11946 ( .A1(P3_U3151), .A2(n15537), .B1(n12784), .B2(n9614), .C1(
        n14787), .C2(n9613), .ZN(P3_U3282) );
  NAND2_X1 U11947 ( .A1(n14570), .A2(P1_B_REG_SCAN_IN), .ZN(n9615) );
  MUX2_X1 U11948 ( .A(P1_B_REG_SCAN_IN), .B(n9615), .S(n14574), .Z(n9617) );
  INV_X1 U11949 ( .A(n14567), .ZN(n9616) );
  INV_X1 U11950 ( .A(n14570), .ZN(n9619) );
  NAND2_X1 U11951 ( .A1(n9618), .A2(n14567), .ZN(n9621) );
  OAI22_X1 U11952 ( .A1(n15136), .A2(P1_D_REG_1__SCAN_IN), .B1(n9619), .B2(
        n9621), .ZN(n9620) );
  INV_X1 U11953 ( .A(n9620), .ZN(P1_U3446) );
  INV_X1 U11954 ( .A(n14574), .ZN(n9622) );
  OAI22_X1 U11955 ( .A1(n15136), .A2(P1_D_REG_0__SCAN_IN), .B1(n9622), .B2(
        n9621), .ZN(n9623) );
  INV_X1 U11956 ( .A(n9623), .ZN(P1_U3445) );
  INV_X1 U11957 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U11958 ( .A1(n9624), .A2(n9748), .ZN(n9625) );
  NAND2_X1 U11959 ( .A1(n9625), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9719) );
  XNOR2_X1 U11960 ( .A(n9719), .B(P1_IR_REG_9__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U11961 ( .A1(n14122), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9722), .ZN(n9626) );
  OAI21_X1 U11962 ( .B1(n11035), .B2(n11699), .A(n9626), .ZN(P1_U3346) );
  INV_X1 U11963 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10654) );
  NOR2_X1 U11964 ( .A1(n15265), .A2(n10654), .ZN(n9644) );
  NAND2_X1 U11965 ( .A1(n9634), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9627) );
  NAND2_X1 U11966 ( .A1(n9628), .A2(n9627), .ZN(n15235) );
  INV_X1 U11967 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9629) );
  MUX2_X1 U11968 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9629), .S(n15232), .Z(
        n15234) );
  NAND2_X1 U11969 ( .A1(n15235), .A2(n15234), .ZN(n15233) );
  NAND2_X1 U11970 ( .A1(n15232), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n12998) );
  NAND2_X1 U11971 ( .A1(n15233), .A2(n12998), .ZN(n9632) );
  INV_X1 U11972 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9630) );
  MUX2_X1 U11973 ( .A(n9630), .B(P2_REG1_REG_8__SCAN_IN), .S(n13001), .Z(n9631) );
  NAND2_X1 U11974 ( .A1(n9632), .A2(n9631), .ZN(n13000) );
  NAND2_X1 U11975 ( .A1(n9640), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9633) );
  NAND2_X1 U11976 ( .A1(n13000), .A2(n9633), .ZN(n9652) );
  NAND2_X1 U11977 ( .A1(n9634), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U11978 ( .A1(n9636), .A2(n9635), .ZN(n15238) );
  INV_X1 U11979 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9637) );
  MUX2_X1 U11980 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9637), .S(n15232), .Z(
        n15237) );
  NAND2_X1 U11981 ( .A1(n15238), .A2(n15237), .ZN(n15236) );
  NAND2_X1 U11982 ( .A1(n15232), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n13003) );
  NAND2_X1 U11983 ( .A1(n15236), .A2(n13003), .ZN(n9639) );
  INV_X1 U11984 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10484) );
  MUX2_X1 U11985 ( .A(n10484), .B(P2_REG2_REG_8__SCAN_IN), .S(n13001), .Z(
        n9638) );
  NAND2_X1 U11986 ( .A1(n9639), .A2(n9638), .ZN(n13005) );
  NAND2_X1 U11987 ( .A1(n9640), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9641) );
  NAND2_X1 U11988 ( .A1(n13005), .A2(n9641), .ZN(n9646) );
  INV_X1 U11989 ( .A(n9646), .ZN(n9642) );
  INV_X1 U11990 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9732) );
  NOR3_X1 U11991 ( .A1(n9642), .A2(n9732), .A3(n15270), .ZN(n9643) );
  AOI211_X1 U11992 ( .C1(n9644), .C2(n9652), .A(n15305), .B(n9643), .ZN(n9657)
         );
  INV_X1 U11993 ( .A(n9650), .ZN(n9733) );
  AND2_X1 U11994 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10625) );
  MUX2_X1 U11995 ( .A(n9732), .B(P2_REG2_REG_9__SCAN_IN), .S(n9650), .Z(n9645)
         );
  OR2_X1 U11996 ( .A1(n9646), .A2(n9645), .ZN(n9735) );
  NAND3_X1 U11997 ( .A1(n9646), .A2(n9733), .A3(n9732), .ZN(n9647) );
  AOI21_X1 U11998 ( .B1(n9735), .B2(n9647), .A(n15270), .ZN(n9648) );
  AOI211_X1 U11999 ( .C1(n15299), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n10625), .B(
        n9648), .ZN(n9656) );
  INV_X1 U12000 ( .A(n9652), .ZN(n9649) );
  NOR3_X1 U12001 ( .A1(n9649), .A2(n9650), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n9654) );
  MUX2_X1 U12002 ( .A(n10654), .B(P2_REG1_REG_9__SCAN_IN), .S(n9650), .Z(n9651) );
  OR2_X1 U12003 ( .A1(n9652), .A2(n9651), .ZN(n9728) );
  INV_X1 U12004 ( .A(n9728), .ZN(n9653) );
  OAI21_X1 U12005 ( .B1(n9654), .B2(n9653), .A(n15300), .ZN(n9655) );
  OAI211_X1 U12006 ( .C1(n9657), .C2(n9733), .A(n9656), .B(n9655), .ZN(
        P2_U3223) );
  INV_X1 U12007 ( .A(n14052), .ZN(n9659) );
  INV_X1 U12008 ( .A(n9663), .ZN(n9658) );
  NAND2_X1 U12009 ( .A1(n9658), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14055) );
  NAND2_X1 U12010 ( .A1(n9659), .A2(n14055), .ZN(n9669) );
  NAND2_X1 U12011 ( .A1(n6643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9662) );
  INV_X1 U12012 ( .A(n14023), .ZN(n10036) );
  NAND2_X1 U12013 ( .A1(n10036), .A2(n9663), .ZN(n9666) );
  NAND2_X1 U12014 ( .A1(n9666), .A2(n10020), .ZN(n9667) );
  AND2_X1 U12015 ( .A1(n9669), .A2(n9667), .ZN(n15018) );
  INV_X1 U12016 ( .A(n9667), .ZN(n9668) );
  INV_X1 U12017 ( .A(n6573), .ZN(n14051) );
  NOR2_X1 U12018 ( .A1(n6573), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9670) );
  OAI21_X1 U12019 ( .B1(n14051), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6761), .ZN(
        n9671) );
  XNOR2_X1 U12020 ( .A(n9671), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9672) );
  AOI22_X1 U12021 ( .A1(n9767), .A2(n9672), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9673) );
  OAI21_X1 U12022 ( .B1(n15047), .B2(n6910), .A(n9673), .ZN(P1_U3243) );
  INV_X1 U12023 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9674) );
  OAI222_X1 U12024 ( .A1(n13417), .A2(n9674), .B1(n13399), .B2(n11035), .C1(
        n9733), .C2(P2_U3088), .ZN(P2_U3318) );
  OAI222_X1 U12025 ( .A1(P3_U3151), .A2(n15554), .B1(n12784), .B2(n9676), .C1(
        n14787), .C2(n9675), .ZN(P3_U3281) );
  AND2_X1 U12026 ( .A1(n9724), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12027 ( .A1(n9724), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12028 ( .A1(n9724), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12029 ( .A1(n9724), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12030 ( .A1(n9724), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12031 ( .A1(n9724), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12032 ( .A1(n9724), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12033 ( .A1(n9724), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12034 ( .A1(n9724), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12035 ( .A1(n9724), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12036 ( .A1(n9724), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12037 ( .A1(n9724), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12038 ( .A1(n9724), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12039 ( .A1(n9724), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12040 ( .A1(n9724), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  INV_X1 U12041 ( .A(P2_B_REG_SCAN_IN), .ZN(n9677) );
  XNOR2_X1 U12042 ( .A(n13414), .B(n9677), .ZN(n9678) );
  NAND2_X1 U12043 ( .A1(n9678), .A2(n13412), .ZN(n9679) );
  INV_X1 U12044 ( .A(n13411), .ZN(n9693) );
  INV_X1 U12045 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15325) );
  NAND2_X1 U12046 ( .A1(n15314), .A2(n15325), .ZN(n9681) );
  NAND2_X1 U12047 ( .A1(n13411), .A2(n13412), .ZN(n9680) );
  NOR4_X1 U12048 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9685) );
  NOR4_X1 U12049 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9684) );
  NOR4_X1 U12050 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9683) );
  NOR4_X1 U12051 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9682) );
  AND4_X1 U12052 ( .A1(n9685), .A2(n9684), .A3(n9683), .A4(n9682), .ZN(n9691)
         );
  NOR2_X1 U12053 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .ZN(
        n9689) );
  NOR4_X1 U12054 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9688) );
  NOR4_X1 U12055 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9687) );
  NOR4_X1 U12056 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n9686) );
  AND4_X1 U12057 ( .A1(n9689), .A2(n9688), .A3(n9687), .A4(n9686), .ZN(n9690)
         );
  NAND2_X1 U12058 ( .A1(n9691), .A2(n9690), .ZN(n9692) );
  AND2_X1 U12059 ( .A1(n15314), .A2(n9692), .ZN(n10144) );
  INV_X1 U12060 ( .A(n9935), .ZN(n9710) );
  INV_X1 U12061 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15323) );
  NAND2_X1 U12062 ( .A1(n15314), .A2(n15323), .ZN(n9695) );
  OR2_X1 U12063 ( .A1(n9693), .A2(n13414), .ZN(n9694) );
  NAND2_X1 U12064 ( .A1(n9695), .A2(n9694), .ZN(n10153) );
  INV_X1 U12065 ( .A(n9701), .ZN(n10142) );
  OAI21_X1 U12066 ( .B1(n9710), .B2(n10153), .A(n10142), .ZN(n9699) );
  NAND2_X1 U12067 ( .A1(n9703), .A2(n9707), .ZN(n10141) );
  AND2_X1 U12068 ( .A1(n9697), .A2(n10141), .ZN(n9698) );
  NAND2_X1 U12069 ( .A1(n9699), .A2(n9698), .ZN(n9890) );
  NOR2_X1 U12070 ( .A1(n9890), .A2(P2_U3088), .ZN(n9956) );
  OR2_X1 U12071 ( .A1(n10153), .A2(n15324), .ZN(n15322) );
  INV_X1 U12072 ( .A(n15322), .ZN(n9700) );
  NOR2_X1 U12073 ( .A1(n9711), .A2(n7288), .ZN(n10133) );
  NAND3_X1 U12074 ( .A1(n9700), .A2(n9935), .A3(n10133), .ZN(n9702) );
  OR3_X1 U12075 ( .A1(n9710), .A2(n15322), .A3(n9707), .ZN(n12967) );
  INV_X1 U12076 ( .A(n12967), .ZN(n12925) );
  INV_X1 U12077 ( .A(n9703), .ZN(n9708) );
  INV_X1 U12078 ( .A(n13031), .ZN(n12963) );
  NAND2_X1 U12079 ( .A1(n12963), .A2(n12992), .ZN(n9706) );
  NAND2_X1 U12080 ( .A1(n13095), .A2(n8648), .ZN(n9705) );
  NAND2_X1 U12081 ( .A1(n9706), .A2(n9705), .ZN(n10255) );
  AOI22_X1 U12082 ( .A1(n12972), .A2(n6574), .B1(n12925), .B2(n10255), .ZN(
        n9718) );
  INV_X1 U12083 ( .A(n9711), .ZN(n9945) );
  NAND2_X1 U12084 ( .A1(n15376), .A2(n9708), .ZN(n9709) );
  OR3_X2 U12085 ( .A1(n9710), .A2(n15322), .A3(n9709), .ZN(n12968) );
  AND2_X1 U12086 ( .A1(n8648), .A2(n10260), .ZN(n10251) );
  NOR2_X2 U12087 ( .A1(n9711), .A2(n9938), .ZN(n13294) );
  NAND2_X1 U12088 ( .A1(n13294), .A2(n10945), .ZN(n10289) );
  NAND2_X1 U12089 ( .A1(n10251), .A2(n10289), .ZN(n9882) );
  NAND2_X1 U12090 ( .A1(n12806), .A2(n10129), .ZN(n9713) );
  AND2_X1 U12091 ( .A1(n9882), .A2(n9713), .ZN(n9715) );
  XNOR2_X1 U12092 ( .A(n11315), .B(n6574), .ZN(n9950) );
  NAND2_X1 U12093 ( .A1(n10289), .A2(n12994), .ZN(n9891) );
  XNOR2_X1 U12094 ( .A(n9950), .B(n9891), .ZN(n9714) );
  NAND2_X1 U12095 ( .A1(n9714), .A2(n9715), .ZN(n9958) );
  OAI21_X1 U12096 ( .B1(n9715), .B2(n9714), .A(n9958), .ZN(n9716) );
  NAND2_X1 U12097 ( .A1(n12961), .A2(n9716), .ZN(n9717) );
  OAI211_X1 U12098 ( .C1(n9956), .C2(n10257), .A(n9718), .B(n9717), .ZN(
        P2_U3194) );
  CLKBUF_X2 U12099 ( .A(P1_U4016), .Z(n14081) );
  NOR2_X1 U12100 ( .A1(n15018), .A2(n14081), .ZN(P1_U3085) );
  INV_X1 U12101 ( .A(n11141), .ZN(n9725) );
  INV_X1 U12102 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9747) );
  NAND2_X1 U12103 ( .A1(n9719), .A2(n9747), .ZN(n9720) );
  NAND2_X1 U12104 ( .A1(n9720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9721) );
  XNOR2_X1 U12105 ( .A(n9721), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11142) );
  AOI22_X1 U12106 ( .A1(n11142), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9722), .ZN(n9723) );
  OAI21_X1 U12107 ( .B1(n9725), .B2(n11699), .A(n9723), .ZN(P1_U3345) );
  INV_X1 U12108 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n12292) );
  NOR2_X1 U12109 ( .A1(n9889), .A2(n12292), .ZN(P3_U3243) );
  INV_X1 U12110 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n12190) );
  NOR2_X1 U12111 ( .A1(n9889), .A2(n12190), .ZN(P3_U3253) );
  INV_X1 U12112 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n12322) );
  NOR2_X1 U12113 ( .A1(n9889), .A2(n12322), .ZN(P3_U3251) );
  INV_X1 U12114 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9726) );
  INV_X1 U12115 ( .A(n9817), .ZN(n9742) );
  OAI222_X1 U12116 ( .A1(n13417), .A2(n9726), .B1(n13399), .B2(n9725), .C1(
        P2_U3088), .C2(n9742), .ZN(P2_U3317) );
  NAND2_X1 U12117 ( .A1(n9733), .A2(n10654), .ZN(n9727) );
  NAND2_X1 U12118 ( .A1(n9728), .A2(n9727), .ZN(n9731) );
  INV_X1 U12119 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11008) );
  MUX2_X1 U12120 ( .A(n11008), .B(P2_REG1_REG_10__SCAN_IN), .S(n9817), .Z(
        n9730) );
  OR2_X1 U12121 ( .A1(n9731), .A2(n9730), .ZN(n9823) );
  INV_X1 U12122 ( .A(n9823), .ZN(n9729) );
  AOI211_X1 U12123 ( .C1(n9731), .C2(n9730), .A(n15265), .B(n9729), .ZN(n9745)
         );
  NAND2_X1 U12124 ( .A1(n9733), .A2(n9732), .ZN(n9734) );
  NAND2_X1 U12125 ( .A1(n9735), .A2(n9734), .ZN(n9739) );
  INV_X1 U12126 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9736) );
  MUX2_X1 U12127 ( .A(n9736), .B(P2_REG2_REG_10__SCAN_IN), .S(n9817), .Z(n9738) );
  OR2_X1 U12128 ( .A1(n9739), .A2(n9738), .ZN(n9813) );
  INV_X1 U12129 ( .A(n9813), .ZN(n9737) );
  AOI211_X1 U12130 ( .C1(n9739), .C2(n9738), .A(n15270), .B(n9737), .ZN(n9744)
         );
  NOR2_X1 U12131 ( .A1(n9740), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10683) );
  AOI21_X1 U12132 ( .B1(n15299), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10683), 
        .ZN(n9741) );
  OAI21_X1 U12133 ( .B1(n15262), .B2(n9742), .A(n9741), .ZN(n9743) );
  OR3_X1 U12134 ( .A1(n9745), .A2(n9744), .A3(n9743), .ZN(P2_U3224) );
  INV_X1 U12135 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14955) );
  INV_X1 U12136 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10335) );
  INV_X1 U12137 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9746) );
  AND3_X1 U12138 ( .A1(n9748), .A2(n9747), .A3(n9746), .ZN(n9749) );
  AND2_X1 U12139 ( .A1(n9750), .A2(n9749), .ZN(n9752) );
  NOR2_X1 U12140 ( .A1(n9752), .A2(n10335), .ZN(n9751) );
  MUX2_X1 U12141 ( .A(n10335), .B(n9751), .S(P1_IR_REG_11__SCAN_IN), .Z(n9753)
         );
  NOR2_X1 U12142 ( .A1(n9753), .A2(n9931), .ZN(n11149) );
  MUX2_X1 U12143 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n14955), .S(n11149), .Z(
        n9764) );
  INV_X1 U12144 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15216) );
  INV_X1 U12145 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10079) );
  MUX2_X1 U12146 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10079), .S(n14102), .Z(
        n9760) );
  INV_X1 U12147 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9754) );
  MUX2_X1 U12148 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9754), .S(n14088), .Z(n9758) );
  INV_X1 U12149 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10015) );
  MUX2_X1 U12150 ( .A(n10015), .B(P1_REG1_REG_1__SCAN_IN), .S(n14069), .Z(
        n9756) );
  AND2_X1 U12151 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9755) );
  NAND2_X1 U12152 ( .A1(n9756), .A2(n9755), .ZN(n14090) );
  OR2_X1 U12153 ( .A1(n14069), .A2(n10015), .ZN(n14089) );
  NAND2_X1 U12154 ( .A1(n14090), .A2(n14089), .ZN(n9757) );
  NAND2_X1 U12155 ( .A1(n9758), .A2(n9757), .ZN(n14099) );
  NAND2_X1 U12156 ( .A1(n14088), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14098) );
  NAND2_X1 U12157 ( .A1(n14099), .A2(n14098), .ZN(n9759) );
  NAND2_X1 U12158 ( .A1(n9760), .A2(n9759), .ZN(n14991) );
  NAND2_X1 U12159 ( .A1(n14102), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14990) );
  INV_X1 U12160 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10246) );
  MUX2_X1 U12161 ( .A(n10246), .B(P1_REG1_REG_4__SCAN_IN), .S(n14994), .Z(
        n14989) );
  AOI21_X1 U12162 ( .B1(n14991), .B2(n14990), .A(n14989), .ZN(n14988) );
  AOI21_X1 U12163 ( .B1(n14994), .B2(P1_REG1_REG_4__SCAN_IN), .A(n14988), .ZN(
        n9796) );
  INV_X1 U12164 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10429) );
  MUX2_X1 U12165 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10429), .S(n10408), .Z(
        n9797) );
  NAND2_X1 U12166 ( .A1(n9796), .A2(n9797), .ZN(n9795) );
  OAI21_X1 U12167 ( .B1(n10408), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9795), .ZN(
        n9877) );
  INV_X1 U12168 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n15214) );
  MUX2_X1 U12169 ( .A(n15214), .B(P1_REG1_REG_6__SCAN_IN), .S(n10853), .Z(
        n9876) );
  NOR2_X1 U12170 ( .A1(n9877), .A2(n9876), .ZN(n9875) );
  NOR2_X1 U12171 ( .A1(n9761), .A2(n15214), .ZN(n9854) );
  MUX2_X1 U12172 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n15216), .S(n10858), .Z(
        n9762) );
  OAI21_X1 U12173 ( .B1(n9875), .B2(n9854), .A(n9762), .ZN(n9857) );
  OAI21_X1 U12174 ( .B1(n15216), .B2(n9866), .A(n9857), .ZN(n9844) );
  INV_X1 U12175 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10874) );
  MUX2_X1 U12176 ( .A(n10874), .B(P1_REG1_REG_8__SCAN_IN), .S(n10871), .Z(
        n9845) );
  NOR2_X1 U12177 ( .A1(n9844), .A2(n9845), .ZN(n14113) );
  NOR2_X1 U12178 ( .A1(n10871), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n14111) );
  INV_X1 U12179 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15219) );
  MUX2_X1 U12180 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15219), .S(n14122), .Z(
        n14112) );
  OAI21_X1 U12181 ( .B1(n14113), .B2(n14111), .A(n14112), .ZN(n14110) );
  OAI21_X1 U12182 ( .B1(n14122), .B2(P1_REG1_REG_9__SCAN_IN), .A(n14110), .ZN(
        n9834) );
  INV_X1 U12183 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n15222) );
  MUX2_X1 U12184 ( .A(n15222), .B(P1_REG1_REG_10__SCAN_IN), .S(n11142), .Z(
        n9833) );
  NOR2_X1 U12185 ( .A1(n9834), .A2(n9833), .ZN(n9832) );
  AOI21_X1 U12186 ( .B1(n11142), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9832), .ZN(
        n9763) );
  NAND2_X1 U12187 ( .A1(n9763), .A2(n9764), .ZN(n15008) );
  OAI21_X1 U12188 ( .B1(n9764), .B2(n9763), .A(n15008), .ZN(n9793) );
  OR2_X1 U12189 ( .A1(n9765), .A2(n14051), .ZN(n15041) );
  INV_X1 U12190 ( .A(n15041), .ZN(n15028) );
  INV_X1 U12191 ( .A(n11694), .ZN(n14079) );
  INV_X1 U12192 ( .A(n11149), .ZN(n10052) );
  NOR2_X1 U12193 ( .A1(n11694), .A2(n6573), .ZN(n9766) );
  AND2_X1 U12194 ( .A1(n9767), .A2(n9766), .ZN(n15024) );
  INV_X1 U12195 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10080) );
  MUX2_X1 U12196 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10080), .S(n14102), .Z(
        n9771) );
  INV_X1 U12197 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10039) );
  MUX2_X1 U12198 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10039), .S(n14088), .Z(
        n9769) );
  INV_X1 U12199 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n14435) );
  MUX2_X1 U12200 ( .A(n14435), .B(P1_REG2_REG_1__SCAN_IN), .S(n14069), .Z(
        n14073) );
  AND2_X1 U12201 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n14078) );
  NAND2_X1 U12202 ( .A1(n14073), .A2(n14078), .ZN(n14084) );
  OR2_X1 U12203 ( .A1(n14069), .A2(n14435), .ZN(n14083) );
  NAND2_X1 U12204 ( .A1(n14084), .A2(n14083), .ZN(n9768) );
  NAND2_X1 U12205 ( .A1(n9769), .A2(n9768), .ZN(n14104) );
  NAND2_X1 U12206 ( .A1(n14088), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14103) );
  NAND2_X1 U12207 ( .A1(n14104), .A2(n14103), .ZN(n9770) );
  NAND2_X1 U12208 ( .A1(n9771), .A2(n9770), .ZN(n14985) );
  NAND2_X1 U12209 ( .A1(n14102), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14984) );
  NAND2_X1 U12210 ( .A1(n14985), .A2(n14984), .ZN(n9773) );
  INV_X1 U12211 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10219) );
  MUX2_X1 U12212 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10219), .S(n14994), .Z(
        n9772) );
  NAND2_X1 U12213 ( .A1(n9773), .A2(n9772), .ZN(n14987) );
  NAND2_X1 U12214 ( .A1(n14994), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9799) );
  NAND2_X1 U12215 ( .A1(n14987), .A2(n9799), .ZN(n9775) );
  INV_X1 U12216 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10234) );
  MUX2_X1 U12217 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10234), .S(n10408), .Z(
        n9774) );
  NAND2_X1 U12218 ( .A1(n9775), .A2(n9774), .ZN(n9872) );
  NAND2_X1 U12219 ( .A1(n10408), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9871) );
  NAND2_X1 U12220 ( .A1(n9872), .A2(n9871), .ZN(n9777) );
  INV_X1 U12221 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n15082) );
  MUX2_X1 U12222 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n15082), .S(n10853), .Z(
        n9776) );
  NAND2_X1 U12223 ( .A1(n9777), .A2(n9776), .ZN(n9874) );
  NAND2_X1 U12224 ( .A1(n10853), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U12225 ( .A1(n9874), .A2(n9778), .ZN(n9861) );
  INV_X1 U12226 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11028) );
  MUX2_X1 U12227 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11028), .S(n10858), .Z(
        n9860) );
  NAND2_X1 U12228 ( .A1(n9861), .A2(n9860), .ZN(n9859) );
  NAND2_X1 U12229 ( .A1(n10858), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9849) );
  NAND2_X1 U12230 ( .A1(n9859), .A2(n9849), .ZN(n9780) );
  INV_X1 U12231 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10877) );
  MUX2_X1 U12232 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10877), .S(n10871), .Z(
        n9779) );
  NAND2_X1 U12233 ( .A1(n9780), .A2(n9779), .ZN(n14119) );
  NAND2_X1 U12234 ( .A1(n10871), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n14118) );
  NAND2_X1 U12235 ( .A1(n14119), .A2(n14118), .ZN(n9782) );
  INV_X1 U12236 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11051) );
  MUX2_X1 U12237 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11051), .S(n14122), .Z(
        n9781) );
  NAND2_X1 U12238 ( .A1(n9782), .A2(n9781), .ZN(n14121) );
  NAND2_X1 U12239 ( .A1(n14122), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9836) );
  NAND2_X1 U12240 ( .A1(n14121), .A2(n9836), .ZN(n9784) );
  INV_X1 U12241 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11043) );
  MUX2_X1 U12242 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11043), .S(n11142), .Z(
        n9783) );
  NAND2_X1 U12243 ( .A1(n9784), .A2(n9783), .ZN(n9838) );
  NAND2_X1 U12244 ( .A1(n11142), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9788) );
  NAND2_X1 U12245 ( .A1(n9838), .A2(n9788), .ZN(n9786) );
  INV_X1 U12246 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11164) );
  MUX2_X1 U12247 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11164), .S(n11149), .Z(
        n9785) );
  NAND2_X1 U12248 ( .A1(n9786), .A2(n9785), .ZN(n10061) );
  MUX2_X1 U12249 ( .A(n11164), .B(P1_REG2_REG_11__SCAN_IN), .S(n11149), .Z(
        n9787) );
  NAND3_X1 U12250 ( .A1(n9838), .A2(n9788), .A3(n9787), .ZN(n9789) );
  NAND3_X1 U12251 ( .A1(n15024), .A2(n10061), .A3(n9789), .ZN(n9791) );
  AND2_X1 U12252 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11656) );
  AOI21_X1 U12253 ( .B1(n15018), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n11656), 
        .ZN(n9790) );
  OAI211_X1 U12254 ( .C1(n15043), .C2(n10052), .A(n9791), .B(n9790), .ZN(n9792) );
  AOI21_X1 U12255 ( .B1(n9793), .B2(n15028), .A(n9792), .ZN(n9794) );
  INV_X1 U12256 ( .A(n9794), .ZN(P1_U3254) );
  OAI21_X1 U12257 ( .B1(n9797), .B2(n9796), .A(n9795), .ZN(n9802) );
  MUX2_X1 U12258 ( .A(n10234), .B(P1_REG2_REG_5__SCAN_IN), .S(n10408), .Z(
        n9798) );
  NAND3_X1 U12259 ( .A1(n14987), .A2(n9799), .A3(n9798), .ZN(n9800) );
  AND3_X1 U12260 ( .A1(n15024), .A2(n9872), .A3(n9800), .ZN(n9801) );
  AOI21_X1 U12261 ( .B1(n15028), .B2(n9802), .A(n9801), .ZN(n9805) );
  NAND2_X1 U12262 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10733) );
  INV_X1 U12263 ( .A(n10733), .ZN(n9803) );
  AOI21_X1 U12264 ( .B1(n15018), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9803), .ZN(
        n9804) );
  OAI211_X1 U12265 ( .C1(n9806), .C2(n15043), .A(n9805), .B(n9804), .ZN(
        P1_U3248) );
  INV_X1 U12266 ( .A(n9807), .ZN(n9808) );
  OAI222_X1 U12267 ( .A1(P3_U3151), .A2(n14827), .B1(n12784), .B2(n12360), 
        .C1(n14787), .C2(n9808), .ZN(P3_U3280) );
  INV_X1 U12268 ( .A(n11148), .ZN(n9810) );
  OAI222_X1 U12269 ( .A1(n10052), .A2(P1_U3086), .B1(n11699), .B2(n9810), .C1(
        n9809), .C2(n14571), .ZN(P1_U3344) );
  INV_X1 U12270 ( .A(n10806), .ZN(n9828) );
  OAI222_X1 U12271 ( .A1(n13417), .A2(n9811), .B1(n13399), .B2(n9810), .C1(
        P2_U3088), .C2(n9828), .ZN(P2_U3316) );
  NAND2_X1 U12272 ( .A1(n9817), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9812) );
  AND2_X1 U12273 ( .A1(n9813), .A2(n9812), .ZN(n9816) );
  INV_X1 U12274 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9814) );
  MUX2_X1 U12275 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n9814), .S(n10806), .Z(
        n9815) );
  NAND2_X1 U12276 ( .A1(n9816), .A2(n9815), .ZN(n15245) );
  OAI21_X1 U12277 ( .B1(n9816), .B2(n9815), .A(n15245), .ZN(n9830) );
  NAND2_X1 U12278 ( .A1(n9817), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9822) );
  NAND2_X1 U12279 ( .A1(n9823), .A2(n9822), .ZN(n9820) );
  INV_X1 U12280 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9818) );
  MUX2_X1 U12281 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9818), .S(n10806), .Z(
        n9819) );
  NAND2_X1 U12282 ( .A1(n9820), .A2(n9819), .ZN(n10808) );
  MUX2_X1 U12283 ( .A(n9818), .B(P2_REG1_REG_11__SCAN_IN), .S(n10806), .Z(
        n9821) );
  NAND3_X1 U12284 ( .A1(n9823), .A2(n9822), .A3(n9821), .ZN(n9824) );
  NAND3_X1 U12285 ( .A1(n10808), .A2(n15300), .A3(n9824), .ZN(n9827) );
  NAND2_X1 U12286 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n10979)
         );
  INV_X1 U12287 ( .A(n10979), .ZN(n9825) );
  AOI21_X1 U12288 ( .B1(n15299), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9825), .ZN(
        n9826) );
  OAI211_X1 U12289 ( .C1(n15262), .C2(n9828), .A(n9827), .B(n9826), .ZN(n9829)
         );
  AOI21_X1 U12290 ( .B1(n15306), .B2(n9830), .A(n9829), .ZN(n9831) );
  INV_X1 U12291 ( .A(n9831), .ZN(P2_U3225) );
  AOI211_X1 U12292 ( .C1(n9834), .C2(n9833), .A(n15041), .B(n9832), .ZN(n9843)
         );
  INV_X1 U12293 ( .A(n11142), .ZN(n9841) );
  MUX2_X1 U12294 ( .A(n11043), .B(P1_REG2_REG_10__SCAN_IN), .S(n11142), .Z(
        n9835) );
  NAND3_X1 U12295 ( .A1(n14121), .A2(n9836), .A3(n9835), .ZN(n9837) );
  NAND3_X1 U12296 ( .A1(n15024), .A2(n9838), .A3(n9837), .ZN(n9840) );
  NOR2_X1 U12297 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12362), .ZN(n11464) );
  AOI21_X1 U12298 ( .B1(n15018), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11464), 
        .ZN(n9839) );
  OAI211_X1 U12299 ( .C1(n15043), .C2(n9841), .A(n9840), .B(n9839), .ZN(n9842)
         );
  OR2_X1 U12300 ( .A1(n9843), .A2(n9842), .ZN(P1_U3253) );
  AOI21_X1 U12301 ( .B1(n9845), .B2(n9844), .A(n14113), .ZN(n9853) );
  NAND2_X1 U12302 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9846) );
  OAI21_X1 U12303 ( .B1(n15047), .B2(n14685), .A(n9846), .ZN(n9847) );
  AOI21_X1 U12304 ( .B1(n10871), .B2(n15012), .A(n9847), .ZN(n9852) );
  MUX2_X1 U12305 ( .A(n10877), .B(P1_REG2_REG_8__SCAN_IN), .S(n10871), .Z(
        n9848) );
  NAND3_X1 U12306 ( .A1(n9859), .A2(n9849), .A3(n9848), .ZN(n9850) );
  NAND3_X1 U12307 ( .A1(n15024), .A2(n14119), .A3(n9850), .ZN(n9851) );
  OAI211_X1 U12308 ( .C1(n9853), .C2(n15041), .A(n9852), .B(n9851), .ZN(
        P1_U3251) );
  INV_X1 U12309 ( .A(n9854), .ZN(n9856) );
  MUX2_X1 U12310 ( .A(n15216), .B(P1_REG1_REG_7__SCAN_IN), .S(n10858), .Z(
        n9855) );
  NAND2_X1 U12311 ( .A1(n9856), .A2(n9855), .ZN(n9858) );
  OAI211_X1 U12312 ( .C1(n9875), .C2(n9858), .A(n15028), .B(n9857), .ZN(n9865)
         );
  NAND2_X1 U12313 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11089) );
  OAI211_X1 U12314 ( .C1(n9861), .C2(n9860), .A(n15024), .B(n9859), .ZN(n9862)
         );
  NAND2_X1 U12315 ( .A1(n11089), .A2(n9862), .ZN(n9863) );
  AOI21_X1 U12316 ( .B1(n15018), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9863), .ZN(
        n9864) );
  OAI211_X1 U12317 ( .C1(n15043), .C2(n9866), .A(n9865), .B(n9864), .ZN(
        P1_U3250) );
  AOI222_X1 U12318 ( .A1(n9867), .A2(n14780), .B1(n14655), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_16_), .C2(n14779), .ZN(n9868) );
  INV_X1 U12319 ( .A(n9868), .ZN(P3_U3279) );
  NAND2_X1 U12320 ( .A1(n15012), .A2(n10853), .ZN(n9869) );
  NAND2_X1 U12321 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10924) );
  OAI211_X1 U12322 ( .C1(n14731), .C2(n15047), .A(n9869), .B(n10924), .ZN(
        n9880) );
  MUX2_X1 U12323 ( .A(n15082), .B(P1_REG2_REG_6__SCAN_IN), .S(n10853), .Z(
        n9870) );
  NAND3_X1 U12324 ( .A1(n9872), .A2(n9871), .A3(n9870), .ZN(n9873) );
  AND3_X1 U12325 ( .A1(n15024), .A2(n9874), .A3(n9873), .ZN(n9879) );
  AOI211_X1 U12326 ( .C1(n9877), .C2(n9876), .A(n9875), .B(n15041), .ZN(n9878)
         );
  OR3_X1 U12327 ( .A1(n9880), .A2(n9879), .A3(n9878), .ZN(P1_U3249) );
  INV_X1 U12328 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n12234) );
  NAND2_X1 U12329 ( .A1(n12961), .A2(n12824), .ZN(n12958) );
  OAI22_X1 U12330 ( .A1(n12958), .A2(n9881), .B1(n10129), .B2(n12968), .ZN(
        n9883) );
  NAND2_X1 U12331 ( .A1(n9883), .A2(n9882), .ZN(n9885) );
  AND2_X1 U12332 ( .A1(n12963), .A2(n12994), .ZN(n9942) );
  AOI22_X1 U12333 ( .A1(n12972), .A2(n10260), .B1(n12925), .B2(n9942), .ZN(
        n9884) );
  OAI211_X1 U12334 ( .C1(n9956), .C2(n12234), .A(n9885), .B(n9884), .ZN(
        P2_U3204) );
  INV_X1 U12335 ( .A(n14628), .ZN(n14868) );
  INV_X1 U12336 ( .A(n9886), .ZN(n9888) );
  INV_X1 U12337 ( .A(SI_17_), .ZN(n9887) );
  OAI222_X1 U12338 ( .A1(n14868), .A2(P3_U3151), .B1(n14787), .B2(n9888), .C1(
        n9887), .C2(n12784), .ZN(P3_U3278) );
  AND2_X1 U12339 ( .A1(n9724), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12340 ( .A1(n9724), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12341 ( .A1(n9724), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12342 ( .A1(n9724), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12343 ( .A1(n9724), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12344 ( .A1(n9724), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12345 ( .A1(n9724), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12346 ( .A1(n9724), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12347 ( .A1(n9724), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12348 ( .A1(n9724), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12349 ( .A1(n9724), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12350 ( .A1(n9724), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  INV_X1 U12351 ( .A(n9891), .ZN(n9892) );
  OR2_X1 U12352 ( .A1(n9950), .A2(n9892), .ZN(n9893) );
  NAND2_X1 U12353 ( .A1(n9958), .A2(n9893), .ZN(n9894) );
  XNOR2_X1 U12354 ( .A(n7166), .B(n11315), .ZN(n9895) );
  NAND2_X1 U12355 ( .A1(n10289), .A2(n12992), .ZN(n9896) );
  XNOR2_X1 U12356 ( .A(n9895), .B(n9896), .ZN(n9951) );
  NAND2_X1 U12357 ( .A1(n9894), .A2(n9951), .ZN(n9961) );
  INV_X1 U12358 ( .A(n9895), .ZN(n9897) );
  NAND2_X1 U12359 ( .A1(n9897), .A2(n9896), .ZN(n9898) );
  NAND2_X1 U12360 ( .A1(n9961), .A2(n9898), .ZN(n9904) );
  AND2_X1 U12361 ( .A1(n12824), .A2(n12991), .ZN(n9900) );
  NAND2_X1 U12362 ( .A1(n9899), .A2(n9900), .ZN(n9913) );
  INV_X1 U12363 ( .A(n9900), .ZN(n9901) );
  NAND2_X1 U12364 ( .A1(n9913), .A2(n9902), .ZN(n9903) );
  INV_X1 U12365 ( .A(n9914), .ZN(n9916) );
  AOI211_X1 U12366 ( .C1(n9904), .C2(n9903), .A(n12968), .B(n9916), .ZN(n9905)
         );
  INV_X1 U12367 ( .A(n9905), .ZN(n9912) );
  NAND2_X1 U12368 ( .A1(n12963), .A2(n12990), .ZN(n9907) );
  NAND2_X1 U12369 ( .A1(n13095), .A2(n12992), .ZN(n9906) );
  NAND2_X1 U12370 ( .A1(n9907), .A2(n9906), .ZN(n10205) );
  INV_X1 U12371 ( .A(n10205), .ZN(n9909) );
  INV_X1 U12372 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9908) );
  OAI22_X1 U12373 ( .A1(n12967), .A2(n9909), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9908), .ZN(n9910) );
  AOI21_X1 U12374 ( .B1(n15348), .B2(n12972), .A(n9910), .ZN(n9911) );
  OAI211_X1 U12375 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n12928), .A(n9912), .B(
        n9911), .ZN(P2_U3190) );
  XNOR2_X1 U12376 ( .A(n10115), .B(n12869), .ZN(n10099) );
  NAND2_X1 U12377 ( .A1(n12824), .A2(n12990), .ZN(n10090) );
  XNOR2_X1 U12378 ( .A(n10099), .B(n10090), .ZN(n9921) );
  INV_X1 U12379 ( .A(n9921), .ZN(n9915) );
  NAND3_X1 U12380 ( .A1(n9914), .A2(n9921), .A3(n9913), .ZN(n10093) );
  INV_X1 U12381 ( .A(n10093), .ZN(n10102) );
  AOI21_X1 U12382 ( .B1(n9916), .B2(n9915), .A(n10102), .ZN(n9926) );
  INV_X1 U12383 ( .A(n10441), .ZN(n9924) );
  INV_X1 U12384 ( .A(n10115), .ZN(n15358) );
  OAI22_X1 U12385 ( .A1(n9920), .A2(n12916), .B1(n10307), .B2(n13031), .ZN(
        n10436) );
  NAND2_X1 U12386 ( .A1(n12925), .A2(n10436), .ZN(n9918) );
  OAI211_X1 U12387 ( .C1(n12957), .C2(n15358), .A(n9918), .B(n9917), .ZN(n9923) );
  NOR4_X1 U12388 ( .A1(n9921), .A2(n12958), .A3(n9920), .A4(n9919), .ZN(n9922)
         );
  AOI211_X1 U12389 ( .C1(n12965), .C2(n9924), .A(n9923), .B(n9922), .ZN(n9925)
         );
  OAI21_X1 U12390 ( .B1(n9926), .B2(n12968), .A(n9925), .ZN(P2_U3202) );
  INV_X1 U12391 ( .A(n10810), .ZN(n15256) );
  INV_X1 U12392 ( .A(n11232), .ZN(n9934) );
  OAI222_X1 U12393 ( .A1(P2_U3088), .A2(n15256), .B1(n13399), .B2(n9934), .C1(
        n9927), .C2(n13417), .ZN(P2_U3315) );
  NOR2_X1 U12394 ( .A1(n9931), .A2(n10335), .ZN(n9928) );
  MUX2_X1 U12395 ( .A(n10335), .B(n9928), .S(P1_IR_REG_12__SCAN_IN), .Z(n9929)
         );
  INV_X1 U12396 ( .A(n9929), .ZN(n9932) );
  INV_X1 U12397 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9930) );
  NAND2_X1 U12398 ( .A1(n9931), .A2(n9930), .ZN(n10050) );
  INV_X1 U12399 ( .A(n15013), .ZN(n10053) );
  OAI222_X1 U12400 ( .A1(P1_U3086), .A2(n10053), .B1(n11699), .B2(n9934), .C1(
        n9933), .C2(n14571), .ZN(P1_U3343) );
  NAND4_X1 U12401 ( .A1(n9935), .A2(n15327), .A3(n10153), .A4(n10141), .ZN(
        n9936) );
  NAND2_X1 U12402 ( .A1(n13252), .A2(n10197), .ZN(n10756) );
  INV_X1 U12403 ( .A(n10756), .ZN(n9937) );
  NAND2_X1 U12404 ( .A1(n9937), .A2(n15331), .ZN(n9948) );
  NAND2_X1 U12405 ( .A1(n9939), .A2(n9938), .ZN(n9941) );
  NAND2_X1 U12406 ( .A1(n11403), .A2(n13024), .ZN(n9940) );
  OAI21_X1 U12407 ( .B1(n15362), .B2(n13264), .A(n15331), .ZN(n9944) );
  INV_X1 U12408 ( .A(n9942), .ZN(n9943) );
  NAND2_X1 U12409 ( .A1(n9944), .A2(n9943), .ZN(n15329) );
  NAND2_X1 U12410 ( .A1(n10260), .A2(n9945), .ZN(n15328) );
  OAI22_X1 U12411 ( .A1(n13236), .A2(n12234), .B1(n10147), .B2(n15328), .ZN(
        n9946) );
  OAI21_X1 U12412 ( .B1(n15329), .B2(n9946), .A(n13252), .ZN(n9947) );
  OAI211_X1 U12413 ( .C1(n9949), .C2(n13252), .A(n9948), .B(n9947), .ZN(
        P2_U3265) );
  INV_X1 U12414 ( .A(n12958), .ZN(n12940) );
  AOI22_X1 U12415 ( .A1(n12940), .A2(n12994), .B1(n12961), .B2(n9950), .ZN(
        n9952) );
  NOR2_X1 U12416 ( .A1(n9952), .A2(n9951), .ZN(n9959) );
  NAND2_X1 U12417 ( .A1(n12963), .A2(n12991), .ZN(n9954) );
  NAND2_X1 U12418 ( .A1(n13095), .A2(n12994), .ZN(n9953) );
  NAND2_X1 U12419 ( .A1(n9954), .A2(n9953), .ZN(n10393) );
  AOI22_X1 U12420 ( .A1(n12972), .A2(n7166), .B1(n12925), .B2(n10393), .ZN(
        n9955) );
  OAI21_X1 U12421 ( .B1(n9956), .B2(n10395), .A(n9955), .ZN(n9957) );
  AOI21_X1 U12422 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(n9960) );
  OAI21_X1 U12423 ( .B1(n9961), .B2(n12968), .A(n9960), .ZN(P2_U3209) );
  INV_X1 U12424 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14071) );
  NOR2_X1 U12425 ( .A1(n6568), .A2(n9962), .ZN(n9963) );
  XNOR2_X1 U12426 ( .A(n9963), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14576) );
  MUX2_X1 U12427 ( .A(n14071), .B(n14576), .S(n10020), .Z(n15140) );
  OR2_X1 U12428 ( .A1(n9979), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U12429 ( .A1(n14570), .A2(n14567), .ZN(n9964) );
  NAND2_X1 U12430 ( .A1(n9965), .A2(n9964), .ZN(n10764) );
  OR2_X1 U12431 ( .A1(n9979), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U12432 ( .A1(n14574), .A2(n14567), .ZN(n9966) );
  NAND2_X1 U12433 ( .A1(n9967), .A2(n9966), .ZN(n10765) );
  NOR4_X1 U12434 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9971) );
  NOR4_X1 U12435 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9970) );
  NOR4_X1 U12436 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9969) );
  NOR4_X1 U12437 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n9968) );
  NAND4_X1 U12438 ( .A1(n9971), .A2(n9970), .A3(n9969), .A4(n9968), .ZN(n9977)
         );
  NOR2_X1 U12439 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .ZN(
        n9975) );
  NOR4_X1 U12440 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9974) );
  NOR4_X1 U12441 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n9973) );
  NOR4_X1 U12442 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9972) );
  NAND4_X1 U12443 ( .A1(n9975), .A2(n9974), .A3(n9973), .A4(n9972), .ZN(n9976)
         );
  NOR2_X1 U12444 ( .A1(n9977), .A2(n9976), .ZN(n9978) );
  OR2_X1 U12445 ( .A1(n9979), .A2(n9978), .ZN(n10007) );
  INV_X1 U12446 ( .A(n10007), .ZN(n9984) );
  INV_X1 U12447 ( .A(n13861), .ZN(n9981) );
  NAND2_X1 U12448 ( .A1(n9409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9980) );
  NAND2_X1 U12449 ( .A1(n6679), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9982) );
  MUX2_X1 U12450 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9982), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9983) );
  OAI21_X1 U12451 ( .B1(n10013), .B2(n9984), .A(n10769), .ZN(n10494) );
  INV_X1 U12452 ( .A(n15139), .ZN(n13862) );
  INV_X1 U12453 ( .A(n11298), .ZN(n13864) );
  NAND2_X1 U12454 ( .A1(n13862), .A2(n13864), .ZN(n14032) );
  INV_X1 U12455 ( .A(n13782), .ZN(n13801) );
  INV_X1 U12456 ( .A(n14265), .ZN(n13462) );
  NAND2_X1 U12457 ( .A1(n13861), .A2(n13462), .ZN(n9985) );
  NAND2_X1 U12458 ( .A1(n15139), .A2(n13864), .ZN(n13863) );
  NAND2_X1 U12459 ( .A1(n13772), .A2(n14050), .ZN(n10087) );
  NAND2_X1 U12460 ( .A1(n15139), .A2(n11298), .ZN(n13856) );
  INV_X1 U12461 ( .A(n15140), .ZN(n10928) );
  NAND2_X1 U12462 ( .A1(n13627), .A2(n10928), .ZN(n10002) );
  INV_X1 U12463 ( .A(n13856), .ZN(n10229) );
  NAND2_X1 U12464 ( .A1(n13832), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9998) );
  INV_X1 U12465 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10929) );
  OR2_X1 U12466 ( .A1(n13692), .A2(n10929), .ZN(n9997) );
  INV_X1 U12467 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9992) );
  OR2_X1 U12468 ( .A1(n10037), .A2(n9992), .ZN(n9996) );
  INV_X1 U12469 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9994) );
  OR2_X1 U12470 ( .A1(n13842), .A2(n9994), .ZN(n9995) );
  NAND2_X1 U12471 ( .A1(n10717), .A2(n10212), .ZN(n10001) );
  INV_X1 U12472 ( .A(n9986), .ZN(n9999) );
  NAND2_X1 U12473 ( .A1(n9999), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10000) );
  INV_X1 U12474 ( .A(n10212), .ZN(n14426) );
  OAI22_X1 U12475 ( .A1(n13681), .A2(n15140), .B1(n9986), .B2(n14071), .ZN(
        n10003) );
  INV_X1 U12476 ( .A(n10003), .ZN(n10004) );
  OAI21_X1 U12477 ( .B1(n13680), .B2(n14426), .A(n10004), .ZN(n10006) );
  INV_X1 U12478 ( .A(n10032), .ZN(n10005) );
  AOI21_X1 U12479 ( .B1(n10030), .B2(n10006), .A(n10005), .ZN(n14077) );
  INV_X1 U12480 ( .A(n10013), .ZN(n10010) );
  NAND2_X1 U12481 ( .A1(n10007), .A2(n14052), .ZN(n10012) );
  NAND2_X1 U12482 ( .A1(n15191), .A2(n14023), .ZN(n10008) );
  NOR2_X1 U12483 ( .A1(n10012), .A2(n10008), .ZN(n10009) );
  INV_X1 U12484 ( .A(n14050), .ZN(n10011) );
  INV_X1 U12485 ( .A(n13650), .ZN(n13795) );
  INV_X1 U12486 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10014) );
  OR2_X1 U12487 ( .A1(n10037), .A2(n10015), .ZN(n10016) );
  OR2_X1 U12488 ( .A1(n14023), .A2(n14079), .ZN(n14156) );
  INV_X2 U12489 ( .A(n14156), .ZN(n15059) );
  NAND2_X1 U12490 ( .A1(n14066), .A2(n15059), .ZN(n15138) );
  OAI22_X1 U12491 ( .A1(n14077), .A2(n13784), .B1(n13795), .B2(n15138), .ZN(
        n10017) );
  AOI21_X1 U12492 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n10087), .A(n10017), .ZN(
        n10018) );
  OAI21_X1 U12493 ( .B1(n15140), .B2(n13801), .A(n10018), .ZN(P1_U3232) );
  INV_X1 U12494 ( .A(n13772), .ZN(n13766) );
  OR2_X1 U12495 ( .A1(n13850), .A2(n7606), .ZN(n10024) );
  OR2_X1 U12496 ( .A1(n13836), .A2(n10021), .ZN(n10023) );
  OR2_X1 U12497 ( .A1(n10020), .A2(n14069), .ZN(n10022) );
  INV_X1 U12498 ( .A(n14423), .ZN(n14421) );
  NAND2_X1 U12499 ( .A1(n15200), .A2(n14421), .ZN(n15146) );
  NOR2_X1 U12500 ( .A1(n13681), .A2(n14423), .ZN(n10025) );
  NAND2_X1 U12501 ( .A1(n13861), .A2(n14265), .ZN(n10026) );
  OAI21_X1 U12502 ( .B1(n10028), .B2(n10027), .A(n10074), .ZN(n10029) );
  INV_X1 U12503 ( .A(n10029), .ZN(n10034) );
  NAND2_X1 U12504 ( .A1(n10032), .A2(n10031), .ZN(n10033) );
  OAI21_X1 U12505 ( .B1(n10034), .B2(n10033), .A(n10075), .ZN(n10035) );
  AOI22_X1 U12506 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n10087), .B1(n10035), 
        .B2(n13790), .ZN(n10045) );
  AND2_X2 U12507 ( .A1(n10036), .A2(n14079), .ZN(n15049) );
  INV_X1 U12508 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10950) );
  OR2_X1 U12509 ( .A1(n13692), .A2(n10950), .ZN(n10042) );
  INV_X1 U12510 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10038) );
  OR2_X1 U12511 ( .A1(n13844), .A2(n10038), .ZN(n10041) );
  OR2_X1 U12512 ( .A1(n13842), .A2(n10039), .ZN(n10040) );
  AOI22_X1 U12513 ( .A1(n13777), .A2(n10212), .B1(n13776), .B2(n14434), .ZN(
        n10044) );
  OAI211_X1 U12514 ( .C1(n13766), .C2(n15146), .A(n10045), .B(n10044), .ZN(
        P1_U3222) );
  INV_X1 U12515 ( .A(n11422), .ZN(n10049) );
  OAI222_X1 U12516 ( .A1(P2_U3088), .A2(n15261), .B1(n13399), .B2(n10049), 
        .C1(n10046), .C2(n13417), .ZN(P2_U3314) );
  NAND2_X1 U12517 ( .A1(n10050), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10047) );
  XNOR2_X1 U12518 ( .A(n10047), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11423) );
  INV_X1 U12519 ( .A(n11423), .ZN(n15021) );
  OAI222_X1 U12520 ( .A1(P1_U3086), .A2(n15021), .B1(n11699), .B2(n10049), 
        .C1(n10048), .C2(n14571), .ZN(P1_U3342) );
  OAI21_X1 U12521 ( .B1(n10050), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10051) );
  XNOR2_X1 U12522 ( .A(n10051), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11515) );
  INV_X1 U12523 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14942) );
  INV_X1 U12524 ( .A(n11515), .ZN(n10516) );
  AOI22_X1 U12525 ( .A1(n11515), .A2(n14942), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n10516), .ZN(n10055) );
  INV_X1 U12526 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n14949) );
  INV_X1 U12527 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14803) );
  NAND2_X1 U12528 ( .A1(n10052), .A2(n14955), .ZN(n15006) );
  MUX2_X1 U12529 ( .A(n14803), .B(P1_REG1_REG_12__SCAN_IN), .S(n15013), .Z(
        n15007) );
  AOI21_X1 U12530 ( .B1(n15008), .B2(n15006), .A(n15007), .ZN(n15005) );
  AOI21_X1 U12531 ( .B1(n14803), .B2(n10053), .A(n15005), .ZN(n15030) );
  MUX2_X1 U12532 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n14949), .S(n11423), .Z(
        n15029) );
  NAND2_X1 U12533 ( .A1(n15030), .A2(n15029), .ZN(n15027) );
  OAI21_X1 U12534 ( .B1(n15021), .B2(n14949), .A(n15027), .ZN(n10054) );
  NOR2_X1 U12535 ( .A1(n10055), .A2(n10054), .ZN(n10512) );
  AOI21_X1 U12536 ( .B1(n10055), .B2(n10054), .A(n10512), .ZN(n10070) );
  NAND2_X1 U12537 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n13652)
         );
  NAND2_X1 U12538 ( .A1(n15018), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n10056) );
  OAI211_X1 U12539 ( .C1(n15043), .C2(n10516), .A(n13652), .B(n10056), .ZN(
        n10057) );
  INV_X1 U12540 ( .A(n10057), .ZN(n10069) );
  NAND2_X1 U12541 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n11423), .ZN(n10065) );
  INV_X1 U12542 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10058) );
  MUX2_X1 U12543 ( .A(n10058), .B(P1_REG2_REG_13__SCAN_IN), .S(n11423), .Z(
        n10059) );
  INV_X1 U12544 ( .A(n10059), .ZN(n15025) );
  NAND2_X1 U12545 ( .A1(n11149), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10060) );
  AND2_X1 U12546 ( .A1(n10061), .A2(n10060), .ZN(n15003) );
  INV_X1 U12547 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10062) );
  MUX2_X1 U12548 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10062), .S(n15013), .Z(
        n15004) );
  NAND2_X1 U12549 ( .A1(n15003), .A2(n15004), .ZN(n15002) );
  INV_X1 U12550 ( .A(n15002), .ZN(n10064) );
  NOR2_X1 U12551 ( .A1(n15013), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U12552 ( .A1(n10064), .A2(n10063), .ZN(n15026) );
  NAND2_X1 U12553 ( .A1(n15025), .A2(n15026), .ZN(n15023) );
  NAND2_X1 U12554 ( .A1(n10065), .A2(n15023), .ZN(n10067) );
  INV_X1 U12555 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11525) );
  MUX2_X1 U12556 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11525), .S(n11515), .Z(
        n10066) );
  NAND2_X1 U12557 ( .A1(n10066), .A2(n10067), .ZN(n10515) );
  OAI211_X1 U12558 ( .C1(n10067), .C2(n10066), .A(n15024), .B(n10515), .ZN(
        n10068) );
  OAI211_X1 U12559 ( .C1(n10070), .C2(n15041), .A(n10069), .B(n10068), .ZN(
        P1_U3257) );
  XNOR2_X1 U12560 ( .A(n10073), .B(n13517), .ZN(n10503) );
  OAI22_X1 U12561 ( .A1(n13680), .A2(n13876), .B1(n15156), .B2(n13681), .ZN(
        n10501) );
  XNOR2_X1 U12562 ( .A(n10503), .B(n10501), .ZN(n10077) );
  NAND2_X1 U12563 ( .A1(n10075), .A2(n10074), .ZN(n10076) );
  NAND2_X1 U12564 ( .A1(n10078), .A2(n13790), .ZN(n10089) );
  NAND2_X1 U12565 ( .A1(n13832), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n10084) );
  OR2_X1 U12566 ( .A1(n10037), .A2(n10079), .ZN(n10083) );
  OR2_X1 U12567 ( .A1(n13842), .A2(n10080), .ZN(n10082) );
  OR2_X1 U12568 ( .A1(n13692), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10081) );
  NAND2_X1 U12569 ( .A1(n14065), .A2(n15059), .ZN(n10086) );
  NAND2_X1 U12570 ( .A1(n14066), .A2(n15049), .ZN(n10085) );
  NAND2_X1 U12571 ( .A1(n10086), .A2(n10085), .ZN(n15153) );
  AOI22_X1 U12572 ( .A1(n10087), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n13650), 
        .B2(n15153), .ZN(n10088) );
  OAI211_X1 U12573 ( .C1(n15156), .C2(n13801), .A(n10089), .B(n10088), .ZN(
        P1_U3237) );
  INV_X1 U12574 ( .A(n10099), .ZN(n10091) );
  NAND2_X1 U12575 ( .A1(n10091), .A2(n10090), .ZN(n10092) );
  NAND2_X1 U12576 ( .A1(n10093), .A2(n10092), .ZN(n10094) );
  XNOR2_X1 U12577 ( .A(n10300), .B(n12869), .ZN(n10280) );
  NAND2_X1 U12578 ( .A1(n12824), .A2(n12989), .ZN(n10281) );
  INV_X1 U12579 ( .A(n10134), .ZN(n10105) );
  NAND2_X1 U12580 ( .A1(n12963), .A2(n12988), .ZN(n10096) );
  NAND2_X1 U12581 ( .A1(n13095), .A2(n12990), .ZN(n10095) );
  NAND2_X1 U12582 ( .A1(n10096), .A2(n10095), .ZN(n10126) );
  NAND2_X1 U12583 ( .A1(n12925), .A2(n10126), .ZN(n10097) );
  OAI211_X1 U12584 ( .C1(n12957), .C2(n10135), .A(n10098), .B(n10097), .ZN(
        n10104) );
  AOI22_X1 U12585 ( .A1(n12940), .A2(n12990), .B1(n12961), .B2(n10099), .ZN(
        n10101) );
  NOR3_X1 U12586 ( .A1(n10102), .A2(n10101), .A3(n10100), .ZN(n10103) );
  AOI211_X1 U12587 ( .C1(n12965), .C2(n10105), .A(n10104), .B(n10103), .ZN(
        n10106) );
  OAI21_X1 U12588 ( .B1(n10284), .B2(n12968), .A(n10106), .ZN(P2_U3199) );
  INV_X1 U12589 ( .A(n10251), .ZN(n10107) );
  NAND2_X1 U12590 ( .A1(n10252), .A2(n10107), .ZN(n10109) );
  OR2_X1 U12591 ( .A1(n12994), .A2(n6574), .ZN(n10108) );
  NAND2_X1 U12592 ( .A1(n10109), .A2(n10108), .ZN(n10389) );
  NAND2_X1 U12593 ( .A1(n10389), .A2(n10119), .ZN(n10111) );
  OR2_X1 U12594 ( .A1(n7166), .A2(n12992), .ZN(n10110) );
  NAND2_X1 U12595 ( .A1(n10111), .A2(n10110), .ZN(n10196) );
  NAND2_X1 U12596 ( .A1(n10112), .A2(n10196), .ZN(n10114) );
  OR2_X1 U12597 ( .A1(n15348), .A2(n12991), .ZN(n10113) );
  NAND2_X1 U12598 ( .A1(n10114), .A2(n10113), .ZN(n10432) );
  NAND2_X1 U12599 ( .A1(n10432), .A2(n7331), .ZN(n10117) );
  OR2_X1 U12600 ( .A1(n10115), .A2(n12990), .ZN(n10116) );
  XNOR2_X1 U12601 ( .A(n10303), .B(n10124), .ZN(n10151) );
  NAND2_X1 U12602 ( .A1(n10254), .A2(n10118), .ZN(n10391) );
  INV_X1 U12603 ( .A(n10119), .ZN(n10392) );
  NAND2_X1 U12604 ( .A1(n10391), .A2(n10392), .ZN(n10390) );
  NAND2_X1 U12605 ( .A1(n10123), .A2(n10124), .ZN(n10305) );
  OAI21_X1 U12606 ( .B1(n10124), .B2(n10123), .A(n10305), .ZN(n10127) );
  AOI211_X1 U12607 ( .C1(n13264), .C2(n10127), .A(n10126), .B(n10125), .ZN(
        n10150) );
  MUX2_X1 U12608 ( .A(n10128), .B(n10150), .S(n13252), .Z(n10138) );
  NAND2_X1 U12609 ( .A1(n10130), .A2(n10129), .ZN(n10396) );
  INV_X1 U12610 ( .A(n10131), .ZN(n10439) );
  INV_X1 U12611 ( .A(n10311), .ZN(n10132) );
  AOI211_X1 U12612 ( .C1(n10300), .C2(n10439), .A(n13270), .B(n10132), .ZN(
        n10148) );
  OAI22_X1 U12613 ( .A1(n13277), .A2(n10135), .B1(n13236), .B2(n10134), .ZN(
        n10136) );
  AOI21_X1 U12614 ( .B1(n10148), .B2(n13272), .A(n10136), .ZN(n10137) );
  OAI211_X1 U12615 ( .C1(n10151), .C2(n10756), .A(n10138), .B(n10137), .ZN(
        P2_U3260) );
  OAI222_X1 U12616 ( .A1(P3_U3151), .A2(n14638), .B1(n14787), .B2(n10140), 
        .C1(n10139), .C2(n12784), .ZN(P3_U3276) );
  NAND3_X1 U12617 ( .A1(n15327), .A2(n10142), .A3(n10141), .ZN(n10143) );
  NOR2_X1 U12618 ( .A1(n10144), .A2(n10143), .ZN(n10145) );
  AND2_X2 U12619 ( .A1(n10155), .A2(n10153), .ZN(n15383) );
  INV_X1 U12620 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n12206) );
  AOI21_X1 U12621 ( .B1(n15366), .B2(n10300), .A(n10148), .ZN(n10149) );
  OAI211_X1 U12622 ( .C1(n10151), .C2(n15369), .A(n10150), .B(n10149), .ZN(
        n10156) );
  NAND2_X1 U12623 ( .A1(n10156), .A2(n15383), .ZN(n10152) );
  OAI21_X1 U12624 ( .B1(n15383), .B2(n12206), .A(n10152), .ZN(P2_U3445) );
  INV_X1 U12625 ( .A(n10153), .ZN(n10154) );
  AND2_X2 U12626 ( .A1(n10155), .A2(n10154), .ZN(n15392) );
  NAND2_X1 U12627 ( .A1(n10156), .A2(n15392), .ZN(n10157) );
  OAI21_X1 U12628 ( .B1(n15392), .B2(n9566), .A(n10157), .ZN(P2_U3504) );
  INV_X1 U12629 ( .A(n10161), .ZN(n10158) );
  NAND2_X1 U12630 ( .A1(n10158), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12088) );
  INV_X1 U12631 ( .A(n12088), .ZN(n10159) );
  OR2_X1 U12632 ( .A1(n10160), .A2(n10159), .ZN(n10171) );
  NAND2_X1 U12633 ( .A1(n12070), .A2(n10161), .ZN(n10162) );
  AND2_X1 U12634 ( .A1(n10163), .A2(n10162), .ZN(n10169) );
  NAND2_X1 U12635 ( .A1(n10171), .A2(n10169), .ZN(n10178) );
  INV_X1 U12636 ( .A(n10178), .ZN(n10166) );
  INV_X1 U12637 ( .A(n10164), .ZN(n10165) );
  INV_X1 U12638 ( .A(n15571), .ZN(n15398) );
  XNOR2_X1 U12639 ( .A(n10371), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10168) );
  INV_X1 U12640 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10184) );
  NOR2_X1 U12641 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10184), .ZN(n15396) );
  INV_X1 U12642 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U12643 ( .A1(n10268), .A2(n6606), .ZN(n10167) );
  NAND2_X1 U12644 ( .A1(n10168), .A2(n10167), .ZN(n10370) );
  OAI21_X1 U12645 ( .B1(n10168), .B2(n10167), .A(n10370), .ZN(n10181) );
  INV_X1 U12646 ( .A(n10169), .ZN(n10170) );
  AOI22_X1 U12647 ( .A1(n15535), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10177) );
  NOR2_X2 U12648 ( .A1(n10178), .A2(n10182), .ZN(n15562) );
  INV_X1 U12649 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10186) );
  NAND2_X1 U12650 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n15402), .ZN(n10172) );
  INV_X1 U12651 ( .A(n10172), .ZN(n15399) );
  OAI21_X1 U12652 ( .B1(n10279), .B2(n15399), .A(n7882), .ZN(n10269) );
  INV_X1 U12653 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10605) );
  OR2_X1 U12654 ( .A1(n10269), .A2(n10605), .ZN(n10271) );
  NAND2_X1 U12655 ( .A1(n10271), .A2(n7882), .ZN(n10173) );
  OAI21_X1 U12656 ( .B1(n10174), .B2(n10173), .A(n10365), .ZN(n10175) );
  NAND2_X1 U12657 ( .A1(n15562), .A2(n10175), .ZN(n10176) );
  NAND2_X1 U12658 ( .A1(n10177), .A2(n10176), .ZN(n10180) );
  INV_X1 U12659 ( .A(P3_U3897), .ZN(n12107) );
  INV_X1 U12660 ( .A(n10371), .ZN(n10188) );
  NOR2_X1 U12661 ( .A1(n15555), .A2(n10188), .ZN(n10179) );
  AOI211_X1 U12662 ( .C1(n15398), .C2(n10181), .A(n10180), .B(n10179), .ZN(
        n10195) );
  INV_X1 U12663 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10183) );
  MUX2_X1 U12664 ( .A(n10184), .B(n10183), .S(n14633), .Z(n15394) );
  AND2_X1 U12665 ( .A1(n15394), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15397) );
  NAND2_X1 U12666 ( .A1(n10264), .A2(n15397), .ZN(n10263) );
  INV_X1 U12667 ( .A(n10185), .ZN(n10192) );
  INV_X1 U12668 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10714) );
  MUX2_X1 U12669 ( .A(n10714), .B(n10186), .S(n14633), .Z(n10187) );
  NAND2_X1 U12670 ( .A1(n10187), .A2(n10371), .ZN(n10357) );
  INV_X1 U12671 ( .A(n10187), .ZN(n10189) );
  NAND2_X1 U12672 ( .A1(n10189), .A2(n10188), .ZN(n10190) );
  NAND2_X1 U12673 ( .A1(n10357), .A2(n10190), .ZN(n10191) );
  AND3_X1 U12674 ( .A1(n10263), .A2(n10192), .A3(n10191), .ZN(n10193) );
  OAI21_X1 U12675 ( .B1(n15413), .B2(n10193), .A(n15543), .ZN(n10194) );
  NAND2_X1 U12676 ( .A1(n10195), .A2(n10194), .ZN(P3_U3184) );
  XNOR2_X1 U12677 ( .A(n10196), .B(n10204), .ZN(n15351) );
  INV_X1 U12678 ( .A(n10197), .ZN(n10198) );
  AOI211_X1 U12679 ( .C1(n15348), .C2(n10397), .A(n13270), .B(n10440), .ZN(
        n15347) );
  INV_X1 U12680 ( .A(n15348), .ZN(n10200) );
  OAI22_X1 U12681 ( .A1(n13277), .A2(n10200), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13236), .ZN(n10201) );
  AOI21_X1 U12682 ( .B1(n13272), .B2(n15347), .A(n10201), .ZN(n10209) );
  OAI21_X1 U12683 ( .B1(n10204), .B2(n10203), .A(n10202), .ZN(n10206) );
  AOI21_X1 U12684 ( .B1(n10206), .B2(n13264), .A(n10205), .ZN(n15349) );
  MUX2_X1 U12685 ( .A(n10207), .B(n15349), .S(n13252), .Z(n10208) );
  OAI211_X1 U12686 ( .C1(n15351), .C2(n13256), .A(n10209), .B(n10208), .ZN(
        P2_U3262) );
  INV_X1 U12687 ( .A(n10765), .ZN(n10210) );
  AND3_X1 U12688 ( .A1(n10210), .A2(n10769), .A3(n10764), .ZN(n10211) );
  NAND2_X1 U12689 ( .A1(n14428), .A2(n14421), .ZN(n13872) );
  NAND2_X1 U12690 ( .A1(n13857), .A2(n13872), .ZN(n13868) );
  NAND2_X1 U12691 ( .A1(n14066), .A2(n14423), .ZN(n13871) );
  NAND2_X1 U12692 ( .A1(n10948), .A2(n13809), .ZN(n10214) );
  NAND2_X1 U12693 ( .A1(n13876), .A2(n13880), .ZN(n10213) );
  NAND2_X1 U12694 ( .A1(n10214), .A2(n10213), .ZN(n10771) );
  NAND2_X1 U12695 ( .A1(n10216), .A2(n11615), .ZN(n10218) );
  AOI22_X1 U12696 ( .A1(n13524), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n13523), 
        .B2(n14994), .ZN(n10217) );
  NAND2_X1 U12697 ( .A1(n13832), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10223) );
  OR2_X1 U12698 ( .A1(n13842), .A2(n10219), .ZN(n10222) );
  OR2_X1 U12699 ( .A1(n10037), .A2(n10246), .ZN(n10221) );
  XNOR2_X1 U12700 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10839) );
  OR2_X1 U12701 ( .A1(n13692), .A2(n10839), .ZN(n10220) );
  XNOR2_X1 U12702 ( .A(n7261), .B(n13891), .ZN(n13812) );
  XNOR2_X1 U12703 ( .A(n10412), .B(n13812), .ZN(n10849) );
  NAND2_X1 U12704 ( .A1(n10212), .A2(n10928), .ZN(n14420) );
  OR2_X1 U12705 ( .A1(n14066), .A2(n14421), .ZN(n10224) );
  INV_X1 U12706 ( .A(n13809), .ZN(n10953) );
  NAND2_X1 U12707 ( .A1(n10954), .A2(n10953), .ZN(n10226) );
  NAND2_X1 U12708 ( .A1(n13876), .A2(n15156), .ZN(n10225) );
  NAND2_X1 U12709 ( .A1(n10226), .A2(n10225), .ZN(n10763) );
  OR2_X1 U12710 ( .A1(n14065), .A2(n10777), .ZN(n10228) );
  XNOR2_X1 U12711 ( .A(n10407), .B(n13812), .ZN(n10846) );
  NAND2_X1 U12712 ( .A1(n10229), .A2(n13861), .ZN(n10230) );
  NAND2_X1 U12713 ( .A1(n10230), .A2(n14265), .ZN(n10231) );
  AND2_X1 U12714 ( .A1(n14423), .A2(n15140), .ZN(n14425) );
  INV_X1 U12715 ( .A(n10424), .ZN(n10232) );
  OAI211_X1 U12716 ( .C1(n13892), .C2(n6756), .A(n10232), .B(n15076), .ZN(
        n10840) );
  AOI21_X1 U12717 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10233) );
  NOR2_X1 U12718 ( .A1(n10233), .A2(n10415), .ZN(n15092) );
  NAND2_X1 U12719 ( .A1(n13553), .A2(n15092), .ZN(n10239) );
  OR2_X1 U12720 ( .A1(n13842), .A2(n10234), .ZN(n10238) );
  OR2_X1 U12721 ( .A1(n10037), .A2(n10429), .ZN(n10237) );
  INV_X1 U12722 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10235) );
  OR2_X1 U12723 ( .A1(n13844), .A2(n10235), .ZN(n10236) );
  NAND4_X1 U12724 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n14063) );
  NAND2_X1 U12725 ( .A1(n14063), .A2(n15059), .ZN(n10241) );
  NAND2_X1 U12726 ( .A1(n14065), .A2(n15049), .ZN(n10240) );
  NAND2_X1 U12727 ( .A1(n10241), .A2(n10240), .ZN(n10841) );
  INV_X1 U12728 ( .A(n10841), .ZN(n10242) );
  OAI211_X1 U12729 ( .C1(n13892), .C2(n15191), .A(n10840), .B(n10242), .ZN(
        n10243) );
  AOI21_X1 U12730 ( .B1(n10846), .B2(n15207), .A(n10243), .ZN(n10244) );
  OAI21_X1 U12731 ( .B1(n15178), .B2(n10849), .A(n10244), .ZN(n10249) );
  NAND2_X1 U12732 ( .A1(n10249), .A2(n15224), .ZN(n10245) );
  OAI21_X1 U12733 ( .B1(n15224), .B2(n10246), .A(n10245), .ZN(P1_U3532) );
  NAND3_X1 U12734 ( .A1(n10764), .A2(n10765), .A3(n10769), .ZN(n10247) );
  INV_X1 U12735 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n12243) );
  NAND2_X1 U12736 ( .A1(n10249), .A2(n15209), .ZN(n10250) );
  OAI21_X1 U12737 ( .B1(n15209), .B2(n12243), .A(n10250), .ZN(P1_U3471) );
  XNOR2_X1 U12738 ( .A(n10252), .B(n10251), .ZN(n15336) );
  INV_X2 U12739 ( .A(n13252), .ZN(n13282) );
  OAI21_X1 U12740 ( .B1(n6572), .B2(n6762), .A(n10254), .ZN(n10256) );
  AOI21_X1 U12741 ( .B1(n10256), .B2(n13264), .A(n10255), .ZN(n15334) );
  OAI22_X1 U12742 ( .A1(n13282), .A2(n15334), .B1(n10257), .B2(n13236), .ZN(
        n10258) );
  AOI21_X1 U12743 ( .B1(n13282), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10258), .ZN(
        n10262) );
  INV_X1 U12744 ( .A(n10396), .ZN(n10259) );
  AOI211_X1 U12745 ( .C1(n10260), .C2(n6574), .A(n13270), .B(n10259), .ZN(
        n15333) );
  AOI22_X1 U12746 ( .A1(n13240), .A2(n6574), .B1(n13272), .B2(n15333), .ZN(
        n10261) );
  OAI211_X1 U12747 ( .C1(n15336), .C2(n13256), .A(n10262), .B(n10261), .ZN(
        P2_U3264) );
  OAI21_X1 U12748 ( .B1(n15397), .B2(n10264), .A(n10263), .ZN(n10277) );
  NAND2_X1 U12749 ( .A1(n10266), .A2(n10265), .ZN(n10267) );
  AND2_X1 U12750 ( .A1(n10268), .A2(n10267), .ZN(n10275) );
  AOI22_X1 U12751 ( .A1(n15535), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10274) );
  NAND2_X1 U12752 ( .A1(n10269), .A2(n10605), .ZN(n10270) );
  NAND2_X1 U12753 ( .A1(n10271), .A2(n10270), .ZN(n10272) );
  NAND2_X1 U12754 ( .A1(n15562), .A2(n10272), .ZN(n10273) );
  OAI211_X1 U12755 ( .C1(n15571), .C2(n10275), .A(n10274), .B(n10273), .ZN(
        n10276) );
  AOI21_X1 U12756 ( .B1(n10277), .B2(n15543), .A(n10276), .ZN(n10278) );
  OAI21_X1 U12757 ( .B1(n10279), .B2(n15555), .A(n10278), .ZN(P3_U3183) );
  INV_X1 U12758 ( .A(n10564), .ZN(n10349) );
  INV_X1 U12759 ( .A(n10280), .ZN(n10282) );
  NAND2_X1 U12760 ( .A1(n10282), .A2(n10281), .ZN(n10283) );
  XNOR2_X1 U12761 ( .A(n15365), .B(n11315), .ZN(n10285) );
  AND2_X1 U12762 ( .A1(n12824), .A2(n12988), .ZN(n10286) );
  NAND2_X1 U12763 ( .A1(n10285), .A2(n10286), .ZN(n10291) );
  INV_X1 U12764 ( .A(n10285), .ZN(n10290) );
  INV_X1 U12765 ( .A(n10286), .ZN(n10287) );
  NAND2_X1 U12766 ( .A1(n10290), .A2(n10287), .ZN(n10288) );
  NAND2_X1 U12767 ( .A1(n10291), .A2(n10288), .ZN(n10327) );
  NAND2_X1 U12768 ( .A1(n12824), .A2(n12987), .ZN(n10612) );
  XNOR2_X1 U12769 ( .A(n10614), .B(n10612), .ZN(n10292) );
  AOI21_X1 U12770 ( .B1(n10324), .B2(n7306), .A(n12968), .ZN(n10295) );
  NOR3_X1 U12771 ( .A1(n10290), .A2(n10350), .A3(n12958), .ZN(n10294) );
  OAI21_X1 U12772 ( .B1(n10295), .B2(n10294), .A(n10616), .ZN(n10299) );
  INV_X1 U12773 ( .A(n10296), .ZN(n10563) );
  AOI22_X1 U12774 ( .A1(n12963), .A2(n12986), .B1(n13095), .B2(n12988), .ZN(
        n10353) );
  NAND2_X1 U12775 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n15230) );
  OAI21_X1 U12776 ( .B1(n12967), .B2(n10353), .A(n15230), .ZN(n10297) );
  AOI21_X1 U12777 ( .B1(n12965), .B2(n10563), .A(n10297), .ZN(n10298) );
  OAI211_X1 U12778 ( .C1(n10349), .C2(n12957), .A(n10299), .B(n10298), .ZN(
        P2_U3185) );
  NOR2_X1 U12779 ( .A1(n10300), .A2(n12989), .ZN(n10302) );
  NAND2_X1 U12780 ( .A1(n10300), .A2(n12989), .ZN(n10301) );
  XNOR2_X1 U12781 ( .A(n10345), .B(n10344), .ZN(n15370) );
  NAND2_X1 U12782 ( .A1(n10305), .A2(n10304), .ZN(n10306) );
  NAND2_X1 U12783 ( .A1(n10306), .A2(n7774), .ZN(n10352) );
  OAI21_X1 U12784 ( .B1(n10306), .B2(n7774), .A(n10352), .ZN(n10309) );
  OAI22_X1 U12785 ( .A1(n10455), .A2(n13031), .B1(n10307), .B2(n12916), .ZN(
        n10320) );
  AOI211_X1 U12786 ( .C1(n13264), .C2(n10309), .A(n10320), .B(n10308), .ZN(
        n15368) );
  MUX2_X1 U12787 ( .A(n10310), .B(n15368), .S(n13252), .Z(n10314) );
  INV_X1 U12788 ( .A(n10347), .ZN(n10346) );
  AOI211_X1 U12789 ( .C1(n15365), .C2(n10311), .A(n13270), .B(n10346), .ZN(
        n15364) );
  OAI22_X1 U12790 ( .A1(n13277), .A2(n7527), .B1(n13236), .B2(n10323), .ZN(
        n10312) );
  AOI21_X1 U12791 ( .B1(n15364), .B2(n13272), .A(n10312), .ZN(n10313) );
  OAI211_X1 U12792 ( .C1(n15370), .C2(n10756), .A(n10314), .B(n10313), .ZN(
        P2_U3259) );
  NAND2_X1 U12793 ( .A1(n12108), .A2(n10316), .ZN(n11929) );
  INV_X1 U12794 ( .A(n11929), .ZN(n11931) );
  NOR2_X1 U12795 ( .A1(n10315), .A2(n11931), .ZN(n11910) );
  NAND2_X1 U12796 ( .A1(n11613), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10598) );
  NAND2_X1 U12797 ( .A1(n10598), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10319) );
  INV_X1 U12798 ( .A(n11870), .ZN(n11845) );
  AOI22_X1 U12799 ( .A1(n11850), .A2(n10317), .B1(n11845), .B2(n8806), .ZN(
        n10318) );
  OAI211_X1 U12800 ( .C1(n11910), .C2(n11852), .A(n10319), .B(n10318), .ZN(
        P3_U3172) );
  NAND2_X1 U12801 ( .A1(n12925), .A2(n10320), .ZN(n10321) );
  OAI211_X1 U12802 ( .C1(n12928), .C2(n10323), .A(n10322), .B(n10321), .ZN(
        n10329) );
  INV_X1 U12803 ( .A(n10324), .ZN(n10325) );
  AOI211_X1 U12804 ( .C1(n10327), .C2(n10326), .A(n12968), .B(n10325), .ZN(
        n10328) );
  AOI211_X1 U12805 ( .C1(n15365), .C2(n12972), .A(n10329), .B(n10328), .ZN(
        n10330) );
  INV_X1 U12806 ( .A(n10330), .ZN(P2_U3211) );
  INV_X1 U12807 ( .A(n10803), .ZN(n11341) );
  INV_X1 U12808 ( .A(n13495), .ZN(n10341) );
  OAI222_X1 U12809 ( .A1(P2_U3088), .A2(n11341), .B1(n13399), .B2(n10341), 
        .C1(n10331), .C2(n13417), .ZN(P2_U3311) );
  INV_X1 U12810 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10333) );
  NOR2_X1 U12811 ( .A1(n10337), .A2(n10335), .ZN(n10334) );
  MUX2_X1 U12812 ( .A(n10335), .B(n10334), .S(P1_IR_REG_16__SCAN_IN), .Z(
        n10339) );
  INV_X1 U12813 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10336) );
  NAND2_X1 U12814 ( .A1(n10337), .A2(n10336), .ZN(n10463) );
  INV_X1 U12815 ( .A(n10463), .ZN(n10338) );
  NOR2_X1 U12816 ( .A1(n10339), .A2(n10338), .ZN(n13496) );
  INV_X1 U12817 ( .A(n13496), .ZN(n11173) );
  OAI222_X1 U12818 ( .A1(P1_U3086), .A2(n11173), .B1(n11699), .B2(n10341), 
        .C1(n10340), .C2(n14571), .ZN(P1_U3339) );
  INV_X1 U12819 ( .A(n10812), .ZN(n15278) );
  INV_X1 U12820 ( .A(n11514), .ZN(n10343) );
  OAI222_X1 U12821 ( .A1(P2_U3088), .A2(n15278), .B1(n13399), .B2(n10343), 
        .C1(n12254), .C2(n13417), .ZN(P2_U3313) );
  OAI222_X1 U12822 ( .A1(P1_U3086), .A2(n10516), .B1(n11699), .B2(n10343), 
        .C1(n10342), .C2(n14571), .ZN(P1_U3341) );
  XOR2_X1 U12823 ( .A(n10446), .B(n10447), .Z(n10570) );
  NAND2_X1 U12824 ( .A1(n10349), .A2(n10346), .ZN(n10450) );
  AOI21_X1 U12825 ( .B1(n10564), .B2(n10347), .A(n13270), .ZN(n10348) );
  NAND2_X1 U12826 ( .A1(n10450), .A2(n10348), .ZN(n10566) );
  OAI21_X1 U12827 ( .B1(n10349), .B2(n15376), .A(n10566), .ZN(n10355) );
  NAND2_X1 U12828 ( .A1(n15365), .A2(n10350), .ZN(n10351) );
  XNOR2_X1 U12829 ( .A(n10452), .B(n10446), .ZN(n10354) );
  OAI21_X1 U12830 ( .B1(n10354), .B2(n13247), .A(n10353), .ZN(n10567) );
  AOI211_X1 U12831 ( .C1(n15373), .C2(n10570), .A(n10355), .B(n10567), .ZN(
        n10491) );
  NAND2_X1 U12832 ( .A1(n15390), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10356) );
  OAI21_X1 U12833 ( .B1(n10491), .B2(n15390), .A(n10356), .ZN(P2_U3506) );
  MUX2_X1 U12834 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n14633), .Z(n10548) );
  XNOR2_X1 U12835 ( .A(n10548), .B(n10547), .ZN(n10549) );
  MUX2_X1 U12836 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n14633), .Z(n10363) );
  INV_X1 U12837 ( .A(n10375), .ZN(n15433) );
  INV_X1 U12838 ( .A(n10357), .ZN(n15412) );
  INV_X1 U12839 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10358) );
  MUX2_X1 U12840 ( .A(n8820), .B(n10358), .S(n14633), .Z(n10359) );
  NAND2_X1 U12841 ( .A1(n10359), .A2(n15418), .ZN(n10362) );
  INV_X1 U12842 ( .A(n10359), .ZN(n10360) );
  INV_X1 U12843 ( .A(n15418), .ZN(n10372) );
  NAND2_X1 U12844 ( .A1(n10360), .A2(n10372), .ZN(n10361) );
  AND2_X1 U12845 ( .A1(n10362), .A2(n10361), .ZN(n15411) );
  XNOR2_X1 U12846 ( .A(n10363), .B(n10375), .ZN(n15429) );
  OAI21_X1 U12847 ( .B1(n10363), .B2(n15433), .A(n15428), .ZN(n15450) );
  MUX2_X1 U12848 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n14633), .Z(n10364) );
  INV_X1 U12849 ( .A(n10378), .ZN(n15453) );
  NAND2_X1 U12850 ( .A1(n10364), .A2(n15453), .ZN(n15446) );
  NOR2_X1 U12851 ( .A1(n10364), .A2(n15453), .ZN(n15448) );
  AOI21_X1 U12852 ( .B1(n15450), .B2(n15446), .A(n15448), .ZN(n10550) );
  XOR2_X1 U12853 ( .A(n10549), .B(n10550), .Z(n10388) );
  OAI21_X1 U12854 ( .B1(n10371), .B2(n10186), .A(n10365), .ZN(n10366) );
  XNOR2_X1 U12855 ( .A(n10366), .B(n15418), .ZN(n15420) );
  AOI22_X1 U12856 ( .A1(n15420), .A2(P3_REG1_REG_3__SCAN_IN), .B1(n10372), 
        .B2(n10366), .ZN(n15437) );
  INV_X1 U12857 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10940) );
  MUX2_X1 U12858 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10940), .S(n10375), .Z(
        n15436) );
  NOR2_X1 U12859 ( .A1(n15437), .A2(n15436), .ZN(n15439) );
  INV_X1 U12860 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10367) );
  INV_X1 U12861 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U12862 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n10547), .B1(n10555), 
        .B2(n11128), .ZN(n10368) );
  NAND2_X1 U12863 ( .A1(n10368), .A2(n10369), .ZN(n10554) );
  OAI21_X1 U12864 ( .B1(n10369), .B2(n10368), .A(n10554), .ZN(n10386) );
  OAI21_X1 U12865 ( .B1(n10371), .B2(n10714), .A(n10370), .ZN(n10373) );
  XNOR2_X1 U12866 ( .A(n10373), .B(n10372), .ZN(n15408) );
  INV_X1 U12867 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10376) );
  MUX2_X1 U12868 ( .A(n10376), .B(P3_REG2_REG_4__SCAN_IN), .S(n10375), .Z(
        n10377) );
  INV_X1 U12869 ( .A(n10377), .ZN(n15426) );
  INV_X1 U12870 ( .A(n10379), .ZN(n10380) );
  INV_X1 U12871 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15445) );
  INV_X1 U12872 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U12873 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n10555), .B1(n10547), 
        .B2(n12279), .ZN(n10381) );
  AOI21_X1 U12874 ( .B1(n6758), .B2(n10381), .A(n10544), .ZN(n10383) );
  AND2_X1 U12875 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11208) );
  AOI21_X1 U12876 ( .B1(n15535), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11208), .ZN(
        n10382) );
  OAI21_X1 U12877 ( .B1(n15571), .B2(n10383), .A(n10382), .ZN(n10385) );
  NOR2_X1 U12878 ( .A1(n15555), .A2(n10547), .ZN(n10384) );
  AOI211_X1 U12879 ( .C1(n15562), .C2(n10386), .A(n10385), .B(n10384), .ZN(
        n10387) );
  OAI21_X1 U12880 ( .B1(n10388), .B2(n15564), .A(n10387), .ZN(P3_U3188) );
  XNOR2_X1 U12881 ( .A(n10392), .B(n10389), .ZN(n15339) );
  OAI21_X1 U12882 ( .B1(n10392), .B2(n10391), .A(n10390), .ZN(n10394) );
  AOI21_X1 U12883 ( .B1(n10394), .B2(n13264), .A(n10393), .ZN(n15341) );
  OAI22_X1 U12884 ( .A1(n13282), .A2(n15341), .B1(n10395), .B2(n13236), .ZN(
        n10400) );
  AOI21_X1 U12885 ( .B1(n10396), .B2(n7166), .A(n13270), .ZN(n10398) );
  NAND2_X1 U12886 ( .A1(n10398), .A2(n10397), .ZN(n15340) );
  OAI22_X1 U12887 ( .A1(n13206), .A2(n15340), .B1(n15342), .B2(n13277), .ZN(
        n10399) );
  AOI211_X1 U12888 ( .C1(n13282), .C2(P2_REG2_REG_2__SCAN_IN), .A(n10400), .B(
        n10399), .ZN(n10401) );
  OAI21_X1 U12889 ( .B1(n13256), .B2(n15339), .A(n10401), .ZN(P2_U3263) );
  INV_X1 U12890 ( .A(n10402), .ZN(n10405) );
  OAI222_X1 U12891 ( .A1(n14787), .A2(n10405), .B1(n12784), .B2(n10404), .C1(
        P3_U3151), .C2(n10403), .ZN(P3_U3275) );
  AND2_X1 U12892 ( .A1(n13892), .A2(n13891), .ZN(n10406) );
  OR2_X1 U12893 ( .A1(n9461), .A2(n13836), .ZN(n10410) );
  AOI22_X1 U12894 ( .A1(n13524), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n13523), 
        .B2(n10408), .ZN(n10409) );
  NAND2_X1 U12895 ( .A1(n10410), .A2(n10409), .ZN(n13899) );
  XNOR2_X1 U12896 ( .A(n13899), .B(n14063), .ZN(n13895) );
  OAI21_X1 U12897 ( .B1(n6750), .B2(n7821), .A(n10851), .ZN(n15101) );
  INV_X1 U12898 ( .A(n15101), .ZN(n10427) );
  INV_X1 U12899 ( .A(n13891), .ZN(n14064) );
  NOR2_X1 U12900 ( .A1(n13892), .A2(n14064), .ZN(n10411) );
  NAND2_X1 U12901 ( .A1(n13892), .A2(n14064), .ZN(n10413) );
  XNOR2_X1 U12902 ( .A(n10891), .B(n13895), .ZN(n10414) );
  NOR2_X1 U12903 ( .A1(n10414), .A2(n15178), .ZN(n10423) );
  INV_X1 U12904 ( .A(n15049), .ZN(n14432) );
  OR2_X1 U12905 ( .A1(n13891), .A2(n14432), .ZN(n10422) );
  NAND2_X1 U12906 ( .A1(n13688), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10420) );
  OR2_X1 U12907 ( .A1(n13842), .A2(n15082), .ZN(n10419) );
  NAND2_X1 U12908 ( .A1(n10415), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10862) );
  OAI21_X1 U12909 ( .B1(n10415), .B2(P1_REG3_REG_6__SCAN_IN), .A(n10862), .ZN(
        n15081) );
  OR2_X1 U12910 ( .A1(n13692), .A2(n15081), .ZN(n10418) );
  INV_X1 U12911 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10416) );
  OR2_X1 U12912 ( .A1(n13844), .A2(n10416), .ZN(n10417) );
  NAND4_X1 U12913 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n10417), .ZN(
        n14062) );
  NAND2_X1 U12914 ( .A1(n14062), .A2(n15059), .ZN(n10421) );
  NAND2_X1 U12915 ( .A1(n10422), .A2(n10421), .ZN(n10732) );
  AOI211_X1 U12916 ( .C1(n15101), .C2(n15074), .A(n10423), .B(n10732), .ZN(
        n15104) );
  OR2_X1 U12917 ( .A1(n15095), .A2(n10424), .ZN(n10425) );
  AND2_X1 U12918 ( .A1(n10425), .A2(n15075), .ZN(n15098) );
  AOI22_X1 U12919 ( .A1(n15098), .A2(n15076), .B1(n13899), .B2(n15200), .ZN(
        n10426) );
  OAI211_X1 U12920 ( .C1(n10427), .C2(n14795), .A(n15104), .B(n10426), .ZN(
        n10430) );
  NAND2_X1 U12921 ( .A1(n10430), .A2(n15224), .ZN(n10428) );
  OAI21_X1 U12922 ( .B1(n15224), .B2(n10429), .A(n10428), .ZN(P1_U3533) );
  NAND2_X1 U12923 ( .A1(n10430), .A2(n15209), .ZN(n10431) );
  OAI21_X1 U12924 ( .B1(n15209), .B2(n10235), .A(n10431), .ZN(P1_U3474) );
  XNOR2_X1 U12925 ( .A(n10432), .B(n10435), .ZN(n15355) );
  OAI21_X1 U12926 ( .B1(n10435), .B2(n10434), .A(n10433), .ZN(n10437) );
  AOI21_X1 U12927 ( .B1(n10437), .B2(n13264), .A(n10436), .ZN(n15357) );
  MUX2_X1 U12928 ( .A(n10438), .B(n15357), .S(n13252), .Z(n10445) );
  OAI211_X1 U12929 ( .C1(n15358), .C2(n10440), .A(n10439), .B(n13294), .ZN(
        n15356) );
  INV_X1 U12930 ( .A(n15356), .ZN(n10443) );
  OAI22_X1 U12931 ( .A1(n13277), .A2(n15358), .B1(n10441), .B2(n13236), .ZN(
        n10442) );
  AOI21_X1 U12932 ( .B1(n13272), .B2(n10443), .A(n10442), .ZN(n10444) );
  OAI211_X1 U12933 ( .C1(n13256), .C2(n15355), .A(n10445), .B(n10444), .ZN(
        P2_U3261) );
  NAND2_X1 U12934 ( .A1(n10447), .A2(n10446), .ZN(n10449) );
  NAND2_X1 U12935 ( .A1(n10564), .A2(n12987), .ZN(n10448) );
  XNOR2_X1 U12936 ( .A(n10539), .B(n10538), .ZN(n10490) );
  AOI211_X1 U12937 ( .C1(n10647), .C2(n10450), .A(n13270), .B(n10532), .ZN(
        n10487) );
  AOI21_X1 U12938 ( .B1(n15366), .B2(n10647), .A(n10487), .ZN(n10457) );
  OR2_X1 U12939 ( .A1(n10564), .A2(n10455), .ZN(n10451) );
  NAND2_X1 U12940 ( .A1(n10452), .A2(n10451), .ZN(n10454) );
  NAND2_X1 U12941 ( .A1(n10564), .A2(n10455), .ZN(n10453) );
  NAND2_X1 U12942 ( .A1(n10454), .A2(n10453), .ZN(n10526) );
  INV_X1 U12943 ( .A(n10538), .ZN(n10525) );
  XNOR2_X1 U12944 ( .A(n10526), .B(n10525), .ZN(n10456) );
  INV_X1 U12945 ( .A(n12985), .ZN(n10744) );
  OAI22_X1 U12946 ( .A1(n10455), .A2(n12916), .B1(n10744), .B2(n13031), .ZN(
        n10634) );
  AOI21_X1 U12947 ( .B1(n10456), .B2(n13264), .A(n10634), .ZN(n10483) );
  OAI211_X1 U12948 ( .C1(n15352), .C2(n10490), .A(n10457), .B(n10483), .ZN(
        n10459) );
  NAND2_X1 U12949 ( .A1(n10459), .A2(n15392), .ZN(n10458) );
  OAI21_X1 U12950 ( .B1(n15392), .B2(n9630), .A(n10458), .ZN(P2_U3507) );
  INV_X1 U12951 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U12952 ( .A1(n10459), .A2(n15383), .ZN(n10460) );
  OAI21_X1 U12953 ( .B1(n15383), .B2(n10461), .A(n10460), .ZN(P2_U3454) );
  NAND2_X1 U12954 ( .A1(n10463), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10462) );
  MUX2_X1 U12955 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10462), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n10464) );
  AND2_X1 U12956 ( .A1(n10464), .A2(n10788), .ZN(n13508) );
  INV_X1 U12957 ( .A(n13508), .ZN(n14128) );
  INV_X1 U12958 ( .A(n13507), .ZN(n10465) );
  OAI222_X1 U12959 ( .A1(P1_U3086), .A2(n14128), .B1(n11699), .B2(n10465), 
        .C1(n12347), .C2(n14571), .ZN(P1_U3338) );
  INV_X1 U12960 ( .A(n15304), .ZN(n11342) );
  OAI222_X1 U12961 ( .A1(n13417), .A2(n10466), .B1(n13399), .B2(n10465), .C1(
        n11342), .C2(P2_U3088), .ZN(P2_U3310) );
  AND2_X1 U12962 ( .A1(n10467), .A2(n12584), .ZN(n10468) );
  OR2_X1 U12963 ( .A1(n11910), .A2(n10468), .ZN(n10470) );
  OR2_X1 U12964 ( .A1(n10708), .A2(n12589), .ZN(n10469) );
  NAND2_X1 U12965 ( .A1(n10470), .A2(n10469), .ZN(n10761) );
  INV_X1 U12966 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n12339) );
  NOR2_X1 U12967 ( .A1(n15599), .A2(n12339), .ZN(n10471) );
  AOI21_X1 U12968 ( .B1(n15599), .B2(n10761), .A(n10471), .ZN(n10472) );
  OAI21_X1 U12969 ( .B1(n10316), .B2(n12770), .A(n10472), .ZN(P3_U3390) );
  INV_X1 U12970 ( .A(n10598), .ZN(n10482) );
  INV_X1 U12971 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10481) );
  INV_X1 U12972 ( .A(n10315), .ZN(n10585) );
  OAI211_X1 U12973 ( .C1(n10476), .C2(n10586), .A(n10475), .B(n10474), .ZN(
        n10477) );
  NAND2_X1 U12974 ( .A1(n10477), .A2(n11863), .ZN(n10480) );
  INV_X1 U12975 ( .A(n11868), .ZN(n11848) );
  OAI22_X1 U12976 ( .A1(n11848), .A2(n7415), .B1(n8812), .B2(n11870), .ZN(
        n10478) );
  AOI21_X1 U12977 ( .B1(n8802), .B2(n11850), .A(n10478), .ZN(n10479) );
  OAI211_X1 U12978 ( .C1(n10482), .C2(n10481), .A(n10480), .B(n10479), .ZN(
        P3_U3162) );
  MUX2_X1 U12979 ( .A(n10484), .B(n10483), .S(n13252), .Z(n10489) );
  INV_X1 U12980 ( .A(n10647), .ZN(n10485) );
  OAI22_X1 U12981 ( .A1(n10485), .A2(n13277), .B1(n13236), .B2(n10636), .ZN(
        n10486) );
  AOI21_X1 U12982 ( .B1(n10487), .B2(n13272), .A(n10486), .ZN(n10488) );
  OAI211_X1 U12983 ( .C1(n10490), .C2(n13256), .A(n10489), .B(n10488), .ZN(
        P2_U3257) );
  INV_X1 U12984 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10493) );
  OR2_X1 U12985 ( .A1(n10491), .A2(n15381), .ZN(n10492) );
  OAI21_X1 U12986 ( .B1(n15383), .B2(n10493), .A(n10492), .ZN(P2_U3451) );
  INV_X1 U12987 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14096) );
  NAND3_X1 U12988 ( .A1(n10494), .A2(n9986), .A3(n14050), .ZN(n10495) );
  NAND2_X1 U12989 ( .A1(n10495), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10496) );
  INV_X1 U12990 ( .A(n13780), .ZN(n13798) );
  INV_X1 U12991 ( .A(n13776), .ZN(n13762) );
  NAND2_X1 U12992 ( .A1(n13782), .A2(n10777), .ZN(n10498) );
  AOI22_X1 U12993 ( .A1(n13777), .A2(n14434), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10497) );
  OAI211_X1 U12994 ( .C1(n13891), .C2(n13762), .A(n10498), .B(n10497), .ZN(
        n10510) );
  INV_X1 U12995 ( .A(n14065), .ZN(n10500) );
  OAI22_X1 U12996 ( .A1(n10500), .A2(n13681), .B1(n10072), .B2(n15163), .ZN(
        n10499) );
  INV_X2 U12997 ( .A(n13517), .ZN(n13682) );
  XNOR2_X1 U12998 ( .A(n10499), .B(n13682), .ZN(n10671) );
  OAI22_X1 U12999 ( .A1(n13680), .A2(n10500), .B1(n15163), .B2(n13681), .ZN(
        n10670) );
  XNOR2_X1 U13000 ( .A(n10671), .B(n10670), .ZN(n10508) );
  INV_X1 U13001 ( .A(n10501), .ZN(n10502) );
  NAND2_X1 U13002 ( .A1(n10503), .A2(n10502), .ZN(n10504) );
  INV_X1 U13003 ( .A(n10673), .ZN(n10506) );
  AOI211_X1 U13004 ( .C1(n10508), .C2(n10507), .A(n13784), .B(n10506), .ZN(
        n10509) );
  AOI211_X1 U13005 ( .C1(n14096), .C2(n13798), .A(n10510), .B(n10509), .ZN(
        n10511) );
  INV_X1 U13006 ( .A(n10511), .ZN(P1_U3218) );
  AOI21_X1 U13007 ( .B1(n10516), .B2(n14942), .A(n10512), .ZN(n10689) );
  XNOR2_X1 U13008 ( .A(n10513), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11617) );
  XNOR2_X1 U13009 ( .A(n10689), .B(n11617), .ZN(n10514) );
  NOR2_X1 U13010 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10514), .ZN(n10690) );
  AOI21_X1 U13011 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n10514), .A(n10690), 
        .ZN(n10524) );
  OAI21_X1 U13012 ( .B1(n11525), .B2(n10516), .A(n10515), .ZN(n10693) );
  INV_X1 U13013 ( .A(n11617), .ZN(n10575) );
  XOR2_X1 U13014 ( .A(n10693), .B(n10575), .Z(n10517) );
  NOR2_X1 U13015 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n10517), .ZN(n10694) );
  AOI21_X1 U13016 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n10517), .A(n10694), 
        .ZN(n10518) );
  INV_X1 U13017 ( .A(n15024), .ZN(n15039) );
  NOR2_X1 U13018 ( .A1(n10518), .A2(n15039), .ZN(n10522) );
  INV_X1 U13019 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n13793) );
  NOR2_X1 U13020 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13793), .ZN(n10519) );
  AOI21_X1 U13021 ( .B1(n15018), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n10519), 
        .ZN(n10520) );
  OAI21_X1 U13022 ( .B1(n10575), .B2(n15043), .A(n10520), .ZN(n10521) );
  NOR2_X1 U13023 ( .A1(n10522), .A2(n10521), .ZN(n10523) );
  OAI21_X1 U13024 ( .B1(n10524), .B2(n15041), .A(n10523), .ZN(P1_U3258) );
  NAND2_X1 U13025 ( .A1(n10647), .A2(n10527), .ZN(n10528) );
  XNOR2_X1 U13026 ( .A(n10743), .B(n10537), .ZN(n10531) );
  NAND2_X1 U13027 ( .A1(n12963), .A2(n12984), .ZN(n10530) );
  NAND2_X1 U13028 ( .A1(n13095), .A2(n12986), .ZN(n10529) );
  NAND2_X1 U13029 ( .A1(n10530), .A2(n10529), .ZN(n10626) );
  AOI21_X1 U13030 ( .B1(n10531), .B2(n13264), .A(n10626), .ZN(n10650) );
  INV_X1 U13031 ( .A(n10745), .ZN(n10629) );
  INV_X1 U13032 ( .A(n10751), .ZN(n10533) );
  AOI211_X1 U13033 ( .C1(n10745), .C2(n10534), .A(n13270), .B(n10533), .ZN(
        n10649) );
  INV_X1 U13034 ( .A(n10623), .ZN(n10535) );
  INV_X1 U13035 ( .A(n13236), .ZN(n13273) );
  AOI22_X1 U13036 ( .A1(n13282), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10535), 
        .B2(n13273), .ZN(n10536) );
  OAI21_X1 U13037 ( .B1(n10629), .B2(n13277), .A(n10536), .ZN(n10542) );
  INV_X1 U13038 ( .A(n10537), .ZN(n10739) );
  NAND2_X1 U13039 ( .A1(n10647), .A2(n12986), .ZN(n10540) );
  XNOR2_X1 U13040 ( .A(n10739), .B(n10738), .ZN(n10652) );
  NOR2_X1 U13041 ( .A1(n10652), .A2(n13256), .ZN(n10541) );
  AOI211_X1 U13042 ( .C1(n10649), .C2(n13272), .A(n10542), .B(n10541), .ZN(
        n10543) );
  OAI21_X1 U13043 ( .B1(n13282), .B2(n10650), .A(n10543), .ZN(P2_U3256) );
  XNOR2_X1 U13044 ( .A(n12380), .B(n12381), .ZN(n10546) );
  INV_X1 U13045 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10545) );
  NOR2_X1 U13046 ( .A1(n10545), .A2(n10546), .ZN(n12382) );
  AOI21_X1 U13047 ( .B1(n10546), .B2(n10545), .A(n12382), .ZN(n10562) );
  OAI22_X1 U13048 ( .A1(n10550), .A2(n10549), .B1(n10548), .B2(n10547), .ZN(
        n10552) );
  MUX2_X1 U13049 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n14633), .Z(n12386) );
  XNOR2_X1 U13050 ( .A(n12386), .B(n12381), .ZN(n10551) );
  NAND2_X1 U13051 ( .A1(n10552), .A2(n10551), .ZN(n12387) );
  OAI21_X1 U13052 ( .B1(n10552), .B2(n10551), .A(n12387), .ZN(n10553) );
  NAND2_X1 U13053 ( .A1(n10553), .A2(n15543), .ZN(n10561) );
  OAI21_X1 U13054 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10556), .A(n12394), .ZN(
        n10559) );
  INV_X1 U13055 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n12173) );
  NOR2_X1 U13056 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12173), .ZN(n11290) );
  AOI21_X1 U13057 ( .B1(n15535), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11290), .ZN(
        n10557) );
  OAI21_X1 U13058 ( .B1(n15555), .B2(n12393), .A(n10557), .ZN(n10558) );
  AOI21_X1 U13059 ( .B1(n10559), .B2(n15562), .A(n10558), .ZN(n10560) );
  OAI211_X1 U13060 ( .C1(n10562), .C2(n15571), .A(n10561), .B(n10560), .ZN(
        P3_U3189) );
  AOI22_X1 U13061 ( .A1(n13240), .A2(n10564), .B1(n10563), .B2(n13273), .ZN(
        n10565) );
  OAI21_X1 U13062 ( .B1(n10566), .B2(n13206), .A(n10565), .ZN(n10569) );
  MUX2_X1 U13063 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10567), .S(n13252), .Z(
        n10568) );
  AOI211_X1 U13064 ( .C1(n13280), .C2(n10570), .A(n10569), .B(n10568), .ZN(
        n10571) );
  INV_X1 U13065 ( .A(n10571), .ZN(P2_U3258) );
  INV_X1 U13066 ( .A(n11616), .ZN(n10574) );
  INV_X1 U13067 ( .A(n15290), .ZN(n10814) );
  OAI222_X1 U13068 ( .A1(n13417), .A2(n10572), .B1(n13399), .B2(n10574), .C1(
        n10814), .C2(P2_U3088), .ZN(P2_U3312) );
  OAI222_X1 U13069 ( .A1(P1_U3086), .A2(n10575), .B1(n11699), .B2(n10574), 
        .C1(n10573), .C2(n14571), .ZN(P1_U3340) );
  OAI21_X1 U13070 ( .B1(n10576), .B2(n12070), .A(n12771), .ZN(n10577) );
  OAI21_X1 U13071 ( .B1(n12771), .B2(n10578), .A(n10577), .ZN(n10579) );
  INV_X1 U13072 ( .A(n10579), .ZN(n10580) );
  AND2_X1 U13073 ( .A1(n10582), .A2(n10705), .ZN(n10583) );
  NAND2_X1 U13074 ( .A1(n14895), .A2(n10583), .ZN(n11357) );
  INV_X1 U13075 ( .A(n12433), .ZN(n11370) );
  NAND2_X1 U13076 ( .A1(n14895), .A2(n11370), .ZN(n10584) );
  NAND2_X1 U13077 ( .A1(n12108), .A2(n12631), .ZN(n10587) );
  OAI21_X1 U13078 ( .B1(n8812), .B2(n12589), .A(n10587), .ZN(n10588) );
  AOI21_X1 U13079 ( .B1(n10589), .B2(n12636), .A(n10588), .ZN(n10603) );
  AND2_X1 U13080 ( .A1(n8802), .A2(n14898), .ZN(n10601) );
  AOI22_X1 U13081 ( .A1(n10601), .A2(n12076), .B1(n12624), .B2(
        P3_REG3_REG_1__SCAN_IN), .ZN(n10590) );
  NAND2_X1 U13082 ( .A1(n10603), .A2(n10590), .ZN(n10591) );
  MUX2_X1 U13083 ( .A(P3_REG2_REG_1__SCAN_IN), .B(n10591), .S(n14895), .Z(
        n10592) );
  AOI21_X1 U13084 ( .B1(n12627), .B2(n10602), .A(n10592), .ZN(n10593) );
  INV_X1 U13085 ( .A(n10593), .ZN(P3_U3232) );
  XOR2_X1 U13086 ( .A(n10595), .B(n10594), .Z(n10600) );
  AOI22_X1 U13087 ( .A1(n11845), .A2(n9268), .B1(n11868), .B2(n8806), .ZN(
        n10596) );
  OAI21_X1 U13088 ( .B1(n11875), .B2(n9306), .A(n10596), .ZN(n10597) );
  AOI21_X1 U13089 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10598), .A(n10597), .ZN(
        n10599) );
  OAI21_X1 U13090 ( .B1(n10600), .B2(n11852), .A(n10599), .ZN(P3_U3177) );
  AOI21_X1 U13091 ( .B1(n10602), .B2(n15595), .A(n10601), .ZN(n10604) );
  AND2_X1 U13092 ( .A1(n10604), .A2(n10603), .ZN(n15573) );
  MUX2_X1 U13093 ( .A(n10605), .B(n15573), .S(n15611), .Z(n10606) );
  INV_X1 U13094 ( .A(n10606), .ZN(P3_U3460) );
  XNOR2_X1 U13095 ( .A(n10745), .B(n12806), .ZN(n10607) );
  NAND2_X1 U13096 ( .A1(n12824), .A2(n12985), .ZN(n10608) );
  NAND2_X1 U13097 ( .A1(n10607), .A2(n10608), .ZN(n10681) );
  INV_X1 U13098 ( .A(n10607), .ZN(n10610) );
  INV_X1 U13099 ( .A(n10608), .ZN(n10609) );
  NAND2_X1 U13100 ( .A1(n10610), .A2(n10609), .ZN(n10611) );
  AND2_X1 U13101 ( .A1(n10681), .A2(n10611), .ZN(n10621) );
  INV_X1 U13102 ( .A(n10612), .ZN(n10613) );
  NAND2_X1 U13103 ( .A1(n10614), .A2(n10613), .ZN(n10615) );
  XNOR2_X1 U13104 ( .A(n10647), .B(n11315), .ZN(n10639) );
  AND2_X1 U13105 ( .A1(n12824), .A2(n12986), .ZN(n10617) );
  AND2_X1 U13106 ( .A1(n10639), .A2(n10617), .ZN(n10637) );
  INV_X1 U13107 ( .A(n10639), .ZN(n10619) );
  INV_X1 U13108 ( .A(n10617), .ZN(n10618) );
  NAND2_X1 U13109 ( .A1(n10619), .A2(n10618), .ZN(n10641) );
  OAI21_X1 U13110 ( .B1(n10621), .B2(n10620), .A(n10682), .ZN(n10622) );
  NAND2_X1 U13111 ( .A1(n10622), .A2(n12961), .ZN(n10628) );
  NOR2_X1 U13112 ( .A1(n12928), .A2(n10623), .ZN(n10624) );
  AOI211_X1 U13113 ( .C1(n12925), .C2(n10626), .A(n10625), .B(n10624), .ZN(
        n10627) );
  OAI211_X1 U13114 ( .C1(n10629), .C2(n12957), .A(n10628), .B(n10627), .ZN(
        P2_U3203) );
  INV_X1 U13115 ( .A(n10630), .ZN(n10632) );
  OAI222_X1 U13116 ( .A1(P3_U3151), .A2(n11932), .B1(n14787), .B2(n10632), 
        .C1(n10631), .C2(n12784), .ZN(P3_U3274) );
  NOR2_X1 U13117 ( .A1(n10633), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12996) );
  AOI21_X1 U13118 ( .B1(n12925), .B2(n10634), .A(n12996), .ZN(n10635) );
  OAI21_X1 U13119 ( .B1(n12928), .B2(n10636), .A(n10635), .ZN(n10646) );
  INV_X1 U13120 ( .A(n10641), .ZN(n10638) );
  NOR3_X1 U13121 ( .A1(n10638), .A2(n10637), .A3(n12968), .ZN(n10644) );
  NAND3_X1 U13122 ( .A1(n10639), .A2(n12940), .A3(n12986), .ZN(n10640) );
  OAI21_X1 U13123 ( .B1(n10641), .B2(n12968), .A(n10640), .ZN(n10643) );
  MUX2_X1 U13124 ( .A(n10644), .B(n10643), .S(n10642), .Z(n10645) );
  AOI211_X1 U13125 ( .C1(n10647), .C2(n12972), .A(n10646), .B(n10645), .ZN(
        n10648) );
  INV_X1 U13126 ( .A(n10648), .ZN(P2_U3193) );
  AOI21_X1 U13127 ( .B1(n15366), .B2(n10745), .A(n10649), .ZN(n10651) );
  OAI211_X1 U13128 ( .C1(n15352), .C2(n10652), .A(n10651), .B(n10650), .ZN(
        n10655) );
  NAND2_X1 U13129 ( .A1(n10655), .A2(n15392), .ZN(n10653) );
  OAI21_X1 U13130 ( .B1(n15392), .B2(n10654), .A(n10653), .ZN(P2_U3508) );
  INV_X1 U13131 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10657) );
  NAND2_X1 U13132 ( .A1(n10655), .A2(n15383), .ZN(n10656) );
  OAI21_X1 U13133 ( .B1(n15383), .B2(n10657), .A(n10656), .ZN(P2_U3457) );
  MUX2_X1 U13134 ( .A(n10761), .B(P3_REG2_REG_0__SCAN_IN), .S(n12648), .Z(
        n10661) );
  INV_X1 U13135 ( .A(n12641), .ZN(n11415) );
  INV_X1 U13136 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10659) );
  OAI22_X1 U13137 ( .A1(n12595), .A2(n10316), .B1(n12639), .B2(n10659), .ZN(
        n10660) );
  OR2_X1 U13138 ( .A1(n10661), .A2(n10660), .ZN(P3_U3233) );
  OAI21_X1 U13139 ( .B1(n10663), .B2(n9309), .A(n10662), .ZN(n10938) );
  AOI22_X1 U13140 ( .A1(n12631), .A2(n12106), .B1(n12105), .B2(n12633), .ZN(
        n10665) );
  NAND2_X1 U13141 ( .A1(n10666), .A2(n10665), .ZN(n10935) );
  AOI21_X1 U13142 ( .B1(n15595), .B2(n10938), .A(n10935), .ZN(n10910) );
  INV_X1 U13143 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n10667) );
  OAI22_X1 U13144 ( .A1(n10934), .A2(n12770), .B1(n15599), .B2(n10667), .ZN(
        n10668) );
  INV_X1 U13145 ( .A(n10668), .ZN(n10669) );
  OAI21_X1 U13146 ( .B1(n10910), .B2(n15601), .A(n10669), .ZN(P3_U3399) );
  NAND2_X1 U13147 ( .A1(n10671), .A2(n10670), .ZN(n10672) );
  OAI22_X1 U13148 ( .A1(n13680), .A2(n13891), .B1(n13892), .B2(n13681), .ZN(
        n10728) );
  INV_X1 U13149 ( .A(n10728), .ZN(n10674) );
  OAI22_X1 U13150 ( .A1(n13892), .A2(n10072), .B1(n13681), .B2(n13891), .ZN(
        n10675) );
  XNOR2_X1 U13151 ( .A(n10675), .B(n13682), .ZN(n10726) );
  XOR2_X1 U13152 ( .A(n10727), .B(n10726), .Z(n10679) );
  NAND2_X1 U13153 ( .A1(n13782), .A2(n7261), .ZN(n10677) );
  AND2_X1 U13154 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14995) );
  AOI21_X1 U13155 ( .B1(n13650), .B2(n10841), .A(n14995), .ZN(n10676) );
  OAI211_X1 U13156 ( .C1(n13780), .C2(n10839), .A(n10677), .B(n10676), .ZN(
        n10678) );
  AOI21_X1 U13157 ( .B1(n10679), .B2(n13790), .A(n10678), .ZN(n10680) );
  INV_X1 U13158 ( .A(n10680), .ZN(P1_U3230) );
  XNOR2_X1 U13159 ( .A(n11003), .B(n12806), .ZN(n10971) );
  NAND2_X1 U13160 ( .A1(n12824), .A2(n12984), .ZN(n10972) );
  XNOR2_X1 U13161 ( .A(n10971), .B(n10972), .ZN(n10969) );
  XNOR2_X1 U13162 ( .A(n10970), .B(n10969), .ZN(n10688) );
  INV_X1 U13163 ( .A(n10752), .ZN(n10685) );
  INV_X1 U13164 ( .A(n12983), .ZN(n11059) );
  OAI22_X1 U13165 ( .A1(n11059), .A2(n13031), .B1(n10744), .B2(n12916), .ZN(
        n10750) );
  AOI21_X1 U13166 ( .B1(n12925), .B2(n10750), .A(n10683), .ZN(n10684) );
  OAI21_X1 U13167 ( .B1(n12928), .B2(n10685), .A(n10684), .ZN(n10686) );
  AOI21_X1 U13168 ( .B1(n11003), .B2(n12972), .A(n10686), .ZN(n10687) );
  OAI21_X1 U13169 ( .B1(n10688), .B2(n12968), .A(n10687), .ZN(P2_U3189) );
  XNOR2_X1 U13170 ( .A(n13496), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11174) );
  NOR2_X1 U13171 ( .A1(n11617), .A2(n10689), .ZN(n10691) );
  NOR2_X1 U13172 ( .A1(n10691), .A2(n10690), .ZN(n11171) );
  XOR2_X1 U13173 ( .A(n11174), .B(n11171), .Z(n10702) );
  NAND2_X1 U13174 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13725)
         );
  INV_X1 U13175 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11170) );
  NOR2_X1 U13176 ( .A1(n11173), .A2(n11170), .ZN(n10692) );
  AOI21_X1 U13177 ( .B1(n11170), .B2(n11173), .A(n10692), .ZN(n10697) );
  NOR2_X1 U13178 ( .A1(n11617), .A2(n10693), .ZN(n10695) );
  NOR2_X1 U13179 ( .A1(n10695), .A2(n10694), .ZN(n10696) );
  NAND2_X1 U13180 ( .A1(n10696), .A2(n10697), .ZN(n11169) );
  OAI211_X1 U13181 ( .C1(n10697), .C2(n10696), .A(n15024), .B(n11169), .ZN(
        n10698) );
  NAND2_X1 U13182 ( .A1(n13725), .A2(n10698), .ZN(n10700) );
  NOR2_X1 U13183 ( .A1(n15043), .A2(n11173), .ZN(n10699) );
  AOI211_X1 U13184 ( .C1(n15018), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n10700), 
        .B(n10699), .ZN(n10701) );
  OAI21_X1 U13185 ( .B1(n10702), .B2(n15041), .A(n10701), .ZN(P1_U3259) );
  INV_X1 U13186 ( .A(n15578), .ZN(n10716) );
  NAND2_X1 U13187 ( .A1(n10704), .A2(n14898), .ZN(n15575) );
  NOR2_X1 U13188 ( .A1(n15575), .A2(n10705), .ZN(n10712) );
  XNOR2_X1 U13189 ( .A(n10707), .B(n10706), .ZN(n10711) );
  OAI22_X1 U13190 ( .A1(n10708), .A2(n12587), .B1(n10964), .B2(n12589), .ZN(
        n10709) );
  AOI21_X1 U13191 ( .B1(n15578), .B2(n11370), .A(n10709), .ZN(n10710) );
  OAI21_X1 U13192 ( .B1(n12584), .B2(n10711), .A(n10710), .ZN(n15576) );
  AOI211_X1 U13193 ( .C1(n12624), .C2(P3_REG3_REG_2__SCAN_IN), .A(n10712), .B(
        n15576), .ZN(n10713) );
  MUX2_X1 U13194 ( .A(n10714), .B(n10713), .S(n14895), .Z(n10715) );
  OAI21_X1 U13195 ( .B1(n10716), .B2(n11357), .A(n10715), .ZN(P3_U3231) );
  NAND2_X1 U13196 ( .A1(n13899), .A2(n13627), .ZN(n10719) );
  NAND2_X1 U13197 ( .A1(n13607), .A2(n14063), .ZN(n10718) );
  NAND2_X1 U13198 ( .A1(n10719), .A2(n10718), .ZN(n10720) );
  XNOR2_X1 U13199 ( .A(n10720), .B(n13517), .ZN(n10722) );
  AOI22_X1 U13200 ( .A1(n13626), .A2(n14063), .B1(n13607), .B2(n13899), .ZN(
        n10723) );
  NAND2_X1 U13201 ( .A1(n10722), .A2(n10723), .ZN(n10911) );
  INV_X1 U13202 ( .A(n10722), .ZN(n10725) );
  INV_X1 U13203 ( .A(n10723), .ZN(n10724) );
  NAND2_X1 U13204 ( .A1(n10725), .A2(n10724), .ZN(n10913) );
  NAND2_X1 U13205 ( .A1(n10911), .A2(n10913), .ZN(n10731) );
  NAND2_X1 U13206 ( .A1(n10729), .A2(n10728), .ZN(n10730) );
  XOR2_X1 U13207 ( .A(n10731), .B(n10912), .Z(n10737) );
  NAND2_X1 U13208 ( .A1(n13650), .A2(n10732), .ZN(n10734) );
  OAI211_X1 U13209 ( .C1(n13801), .C2(n15095), .A(n10734), .B(n10733), .ZN(
        n10735) );
  AOI21_X1 U13210 ( .B1(n15092), .B2(n13798), .A(n10735), .ZN(n10736) );
  OAI21_X1 U13211 ( .B1(n10737), .B2(n13784), .A(n10736), .ZN(P1_U3227) );
  NAND2_X1 U13212 ( .A1(n10745), .A2(n12985), .ZN(n10740) );
  XNOR2_X1 U13213 ( .A(n10985), .B(n10746), .ZN(n10755) );
  AND2_X1 U13214 ( .A1(n10745), .A2(n10744), .ZN(n10742) );
  INV_X1 U13215 ( .A(n10746), .ZN(n10984) );
  NAND2_X1 U13216 ( .A1(n10747), .A2(n10984), .ZN(n10748) );
  AOI21_X1 U13217 ( .B1(n10989), .B2(n10748), .A(n13247), .ZN(n10749) );
  AOI211_X1 U13218 ( .C1(n15362), .C2(n10755), .A(n10750), .B(n10749), .ZN(
        n11005) );
  AOI211_X1 U13219 ( .C1(n11003), .C2(n10751), .A(n13270), .B(n10995), .ZN(
        n11002) );
  INV_X1 U13220 ( .A(n11003), .ZN(n10754) );
  AOI22_X1 U13221 ( .A1(n13282), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10752), 
        .B2(n13273), .ZN(n10753) );
  OAI21_X1 U13222 ( .B1(n10754), .B2(n13277), .A(n10753), .ZN(n10758) );
  INV_X1 U13223 ( .A(n10755), .ZN(n11006) );
  NOR2_X1 U13224 ( .A1(n11006), .A2(n10756), .ZN(n10757) );
  AOI211_X1 U13225 ( .C1(n11002), .C2(n13272), .A(n10758), .B(n10757), .ZN(
        n10759) );
  OAI21_X1 U13226 ( .B1(n11005), .B2(n13282), .A(n10759), .ZN(P2_U3255) );
  NOR2_X1 U13227 ( .A1(n15611), .A2(n10183), .ZN(n10760) );
  AOI21_X1 U13228 ( .B1(n10761), .B2(n15611), .A(n10760), .ZN(n10762) );
  OAI21_X1 U13229 ( .B1(n10316), .B2(n12715), .A(n10762), .ZN(P3_U3459) );
  XNOR2_X1 U13230 ( .A(n10763), .B(n13885), .ZN(n10775) );
  INV_X1 U13231 ( .A(n10775), .ZN(n15166) );
  INV_X1 U13232 ( .A(n10764), .ZN(n10766) );
  INV_X1 U13233 ( .A(n10769), .ZN(n10770) );
  OR2_X1 U13234 ( .A1(n13856), .A2(n14265), .ZN(n14024) );
  XNOR2_X1 U13235 ( .A(n10771), .B(n13885), .ZN(n10773) );
  OAI22_X1 U13236 ( .A1(n13891), .A2(n14156), .B1(n13876), .B2(n14432), .ZN(
        n10772) );
  AOI21_X1 U13237 ( .B1(n10773), .B2(n15196), .A(n10772), .ZN(n10774) );
  OAI21_X1 U13238 ( .B1(n10775), .B2(n10844), .A(n10774), .ZN(n15164) );
  MUX2_X1 U13239 ( .A(n15164), .B(P1_REG2_REG_3__SCAN_IN), .S(n15105), .Z(
        n10780) );
  AOI211_X1 U13240 ( .C1(n10777), .C2(n10949), .A(n15147), .B(n6756), .ZN(
        n15161) );
  INV_X1 U13241 ( .A(n15080), .ZN(n15091) );
  AOI22_X1 U13242 ( .A1(n15063), .A2(n15161), .B1(n15091), .B2(n14096), .ZN(
        n10778) );
  OAI21_X1 U13243 ( .B1(n15163), .B2(n15096), .A(n10778), .ZN(n10779) );
  AOI211_X1 U13244 ( .C1(n15166), .C2(n15100), .A(n10780), .B(n10779), .ZN(
        n10781) );
  INV_X1 U13245 ( .A(n10781), .ZN(P1_U3290) );
  OAI211_X1 U13246 ( .C1(n10783), .C2(n10782), .A(n6759), .B(n11863), .ZN(
        n10787) );
  NOR2_X1 U13247 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10784), .ZN(n15409) );
  OAI22_X1 U13248 ( .A1(n8812), .A2(n11848), .B1(n11875), .B2(n10934), .ZN(
        n10785) );
  AOI211_X1 U13249 ( .C1(n11845), .C2(n12105), .A(n15409), .B(n10785), .ZN(
        n10786) );
  OAI211_X1 U13250 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11613), .A(n10787), .B(
        n10786), .ZN(P3_U3158) );
  NAND2_X1 U13251 ( .A1(n10788), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10789) );
  XNOR2_X1 U13252 ( .A(n10789), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14139) );
  INV_X1 U13253 ( .A(n14139), .ZN(n15042) );
  INV_X1 U13254 ( .A(n13522), .ZN(n10791) );
  OAI222_X1 U13255 ( .A1(n15042), .A2(P1_U3086), .B1(n11699), .B2(n10791), 
        .C1(n12269), .C2(n14571), .ZN(P1_U3337) );
  INV_X1 U13256 ( .A(n13014), .ZN(n10790) );
  OAI222_X1 U13257 ( .A1(n13417), .A2(n10792), .B1(n13399), .B2(n10791), .C1(
        P2_U3088), .C2(n10790), .ZN(P2_U3309) );
  NAND2_X1 U13258 ( .A1(n10793), .A2(n14780), .ZN(n10794) );
  OAI211_X1 U13259 ( .C1(n10795), .C2(n12784), .A(n10794), .B(n12088), .ZN(
        P3_U3272) );
  OR2_X1 U13260 ( .A1(n10806), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n15243) );
  NAND2_X1 U13261 ( .A1(n15245), .A2(n15243), .ZN(n10797) );
  INV_X1 U13262 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10796) );
  MUX2_X1 U13263 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n10796), .S(n10810), .Z(
        n15242) );
  NAND2_X1 U13264 ( .A1(n10797), .A2(n15242), .ZN(n15247) );
  OAI21_X1 U13265 ( .B1(n10810), .B2(P2_REG2_REG_12__SCAN_IN), .A(n15247), 
        .ZN(n15271) );
  INV_X1 U13266 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10798) );
  MUX2_X1 U13267 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n10798), .S(n15261), .Z(
        n15272) );
  NOR2_X1 U13268 ( .A1(n15271), .A2(n15272), .ZN(n15269) );
  AOI21_X1 U13269 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n10811), .A(n15269), 
        .ZN(n10799) );
  OR2_X1 U13270 ( .A1(n10799), .A2(n15278), .ZN(n10800) );
  XNOR2_X1 U13271 ( .A(n10799), .B(n10812), .ZN(n15282) );
  NAND2_X1 U13272 ( .A1(n15282), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n15281) );
  NAND2_X1 U13273 ( .A1(n10800), .A2(n15281), .ZN(n10801) );
  NAND2_X1 U13274 ( .A1(n15290), .A2(n10801), .ZN(n10802) );
  XNOR2_X1 U13275 ( .A(n10814), .B(n10801), .ZN(n15292) );
  NAND2_X1 U13276 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15292), .ZN(n15291) );
  NAND2_X1 U13277 ( .A1(n10802), .A2(n15291), .ZN(n10805) );
  XNOR2_X1 U13278 ( .A(n10803), .B(n11586), .ZN(n10804) );
  NAND2_X1 U13279 ( .A1(n10804), .A2(n10805), .ZN(n11334) );
  OAI211_X1 U13280 ( .C1(n10805), .C2(n10804), .A(n15306), .B(n11334), .ZN(
        n10822) );
  NAND2_X1 U13281 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n12897)
         );
  NAND2_X1 U13282 ( .A1(n10806), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10807) );
  NAND2_X1 U13283 ( .A1(n10808), .A2(n10807), .ZN(n15250) );
  INV_X1 U13284 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10809) );
  MUX2_X1 U13285 ( .A(n10809), .B(P2_REG1_REG_12__SCAN_IN), .S(n10810), .Z(
        n15249) );
  OAI21_X1 U13286 ( .B1(n10810), .B2(P2_REG1_REG_12__SCAN_IN), .A(n15252), 
        .ZN(n15266) );
  XNOR2_X1 U13287 ( .A(n10811), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n15267) );
  NOR2_X1 U13288 ( .A1(n15266), .A2(n15267), .ZN(n15264) );
  AOI21_X1 U13289 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n10811), .A(n15264), 
        .ZN(n15283) );
  XNOR2_X1 U13290 ( .A(n10812), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n15284) );
  INV_X1 U13291 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10813) );
  OAI22_X1 U13292 ( .A1(n15283), .A2(n15284), .B1(n15278), .B2(n10813), .ZN(
        n10815) );
  NAND2_X1 U13293 ( .A1(n15290), .A2(n10815), .ZN(n10816) );
  XNOR2_X1 U13294 ( .A(n10815), .B(n10814), .ZN(n15294) );
  NAND2_X1 U13295 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15294), .ZN(n15293) );
  NAND2_X1 U13296 ( .A1(n10816), .A2(n15293), .ZN(n10818) );
  XNOR2_X1 U13297 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n11341), .ZN(n10817) );
  NAND2_X1 U13298 ( .A1(n10817), .A2(n10818), .ZN(n11339) );
  OAI211_X1 U13299 ( .C1(n10818), .C2(n10817), .A(n15300), .B(n11339), .ZN(
        n10819) );
  NAND2_X1 U13300 ( .A1(n12897), .A2(n10819), .ZN(n10820) );
  AOI21_X1 U13301 ( .B1(n15299), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n10820), 
        .ZN(n10821) );
  OAI211_X1 U13302 ( .C1(n15262), .C2(n11341), .A(n10822), .B(n10821), .ZN(
        P2_U3230) );
  OAI21_X1 U13303 ( .B1(n10824), .B2(n11948), .A(n10823), .ZN(n10825) );
  INV_X1 U13304 ( .A(n10825), .ZN(n10835) );
  INV_X1 U13305 ( .A(n10826), .ZN(n10827) );
  AOI21_X1 U13306 ( .B1(n10827), .B2(n11948), .A(n12584), .ZN(n10830) );
  OAI22_X1 U13307 ( .A1(n10964), .A2(n12587), .B1(n11206), .B2(n12589), .ZN(
        n10828) );
  AOI21_X1 U13308 ( .B1(n10830), .B2(n10829), .A(n10828), .ZN(n10834) );
  MUX2_X1 U13309 ( .A(n10376), .B(n10834), .S(n14895), .Z(n10833) );
  INV_X1 U13310 ( .A(n12595), .ZN(n14893) );
  AOI22_X1 U13311 ( .A1(n14893), .A2(n10831), .B1(n12624), .B2(n10957), .ZN(
        n10832) );
  OAI211_X1 U13312 ( .C1(n12644), .C2(n10835), .A(n10833), .B(n10832), .ZN(
        P3_U3229) );
  OAI21_X1 U13313 ( .B1(n14910), .B2(n10835), .A(n10834), .ZN(n10942) );
  INV_X1 U13314 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n10836) );
  OAI22_X1 U13315 ( .A1(n10963), .A2(n12770), .B1(n15599), .B2(n10836), .ZN(
        n10837) );
  AOI21_X1 U13316 ( .B1(n10942), .B2(n15599), .A(n10837), .ZN(n10838) );
  INV_X1 U13317 ( .A(n10838), .ZN(P3_U3402) );
  OR2_X1 U13318 ( .A1(n15105), .A2(n15178), .ZN(n14273) );
  OAI22_X1 U13319 ( .A1(n15087), .A2(n10840), .B1(n10839), .B2(n15080), .ZN(
        n10843) );
  MUX2_X1 U13320 ( .A(n10841), .B(P1_REG2_REG_4__SCAN_IN), .S(n15105), .Z(
        n10842) );
  AOI211_X1 U13321 ( .C1(n15085), .C2(n7261), .A(n10843), .B(n10842), .ZN(
        n10848) );
  AND2_X1 U13322 ( .A1(n10844), .A2(n14024), .ZN(n10845) );
  NAND2_X1 U13323 ( .A1(n15065), .A2(n10846), .ZN(n10847) );
  OAI211_X1 U13324 ( .C1(n10849), .C2(n14273), .A(n10848), .B(n10847), .ZN(
        P1_U3289) );
  INV_X1 U13325 ( .A(n14063), .ZN(n10889) );
  NAND2_X1 U13326 ( .A1(n15095), .A2(n10889), .ZN(n10850) );
  NAND2_X1 U13327 ( .A1(n10852), .A2(n11615), .ZN(n10855) );
  AOI22_X1 U13328 ( .A1(n13524), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n13523), 
        .B2(n10853), .ZN(n10854) );
  NAND2_X1 U13329 ( .A1(n10855), .A2(n10854), .ZN(n15084) );
  XNOR2_X1 U13330 ( .A(n15084), .B(n14062), .ZN(n13814) );
  OR2_X1 U13331 ( .A1(n15084), .A2(n14062), .ZN(n10856) );
  NAND2_X1 U13332 ( .A1(n15069), .A2(n10856), .ZN(n11025) );
  OR2_X1 U13333 ( .A1(n10857), .A2(n13836), .ZN(n10860) );
  AOI22_X1 U13334 ( .A1(n13524), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n13523), 
        .B2(n10858), .ZN(n10859) );
  NAND2_X1 U13335 ( .A1(n10860), .A2(n10859), .ZN(n13906) );
  NAND2_X1 U13336 ( .A1(n13688), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10868) );
  OR2_X1 U13337 ( .A1(n13842), .A2(n11028), .ZN(n10867) );
  INV_X1 U13338 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10861) );
  AND2_X1 U13339 ( .A1(n10862), .A2(n10861), .ZN(n10863) );
  NOR2_X1 U13340 ( .A1(n10862), .A2(n10861), .ZN(n10875) );
  OR2_X1 U13341 ( .A1(n10863), .A2(n10875), .ZN(n11096) );
  OR2_X1 U13342 ( .A1(n13692), .A2(n11096), .ZN(n10866) );
  INV_X1 U13343 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10864) );
  OR2_X1 U13344 ( .A1(n13844), .A2(n10864), .ZN(n10865) );
  NAND4_X1 U13345 ( .A1(n10868), .A2(n10867), .A3(n10866), .A4(n10865), .ZN(
        n14061) );
  INV_X1 U13346 ( .A(n14061), .ZN(n11085) );
  XNOR2_X1 U13347 ( .A(n13906), .B(n11085), .ZN(n13813) );
  NAND2_X1 U13348 ( .A1(n11025), .A2(n13813), .ZN(n11024) );
  OR2_X1 U13349 ( .A1(n13906), .A2(n14061), .ZN(n10869) );
  NAND2_X1 U13350 ( .A1(n11024), .A2(n10869), .ZN(n10883) );
  OR2_X1 U13351 ( .A1(n10870), .A2(n13836), .ZN(n10873) );
  AOI22_X1 U13352 ( .A1(n13524), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n13523), 
        .B2(n10871), .ZN(n10872) );
  NAND2_X1 U13353 ( .A1(n10873), .A2(n10872), .ZN(n13913) );
  NAND2_X1 U13354 ( .A1(n13832), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10881) );
  OR2_X1 U13355 ( .A1(n10037), .A2(n10874), .ZN(n10880) );
  NAND2_X1 U13356 ( .A1(n10875), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10897) );
  OR2_X1 U13357 ( .A1(n10875), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10876) );
  NAND2_X1 U13358 ( .A1(n10897), .A2(n10876), .ZN(n11271) );
  OR2_X1 U13359 ( .A1(n13692), .A2(n11271), .ZN(n10879) );
  OR2_X1 U13360 ( .A1(n13842), .A2(n10877), .ZN(n10878) );
  NAND4_X1 U13361 ( .A1(n10881), .A2(n10880), .A3(n10879), .A4(n10878), .ZN(
        n14060) );
  XNOR2_X1 U13362 ( .A(n13913), .B(n14060), .ZN(n13815) );
  INV_X1 U13363 ( .A(n13815), .ZN(n10882) );
  NAND2_X1 U13364 ( .A1(n10883), .A2(n10882), .ZN(n11034) );
  OAI21_X1 U13365 ( .B1(n10883), .B2(n10882), .A(n11034), .ZN(n15188) );
  INV_X1 U13366 ( .A(n13906), .ZN(n15177) );
  AOI21_X1 U13367 ( .B1(n11026), .B2(n13913), .A(n15147), .ZN(n10884) );
  AND2_X1 U13368 ( .A1(n10884), .A2(n11052), .ZN(n15185) );
  NAND2_X1 U13369 ( .A1(n15185), .A2(n15063), .ZN(n10887) );
  NOR2_X1 U13370 ( .A1(n15080), .A2(n11271), .ZN(n10885) );
  AOI21_X1 U13371 ( .B1(n15105), .B2(P1_REG2_REG_8__SCAN_IN), .A(n10885), .ZN(
        n10886) );
  OAI211_X1 U13372 ( .C1(n7592), .C2(n15096), .A(n10887), .B(n10886), .ZN(
        n10888) );
  AOI21_X1 U13373 ( .B1(n15188), .B2(n15065), .A(n10888), .ZN(n10907) );
  NOR2_X1 U13374 ( .A1(n13899), .A2(n10889), .ZN(n10890) );
  INV_X1 U13375 ( .A(n14062), .ZN(n10917) );
  NAND2_X1 U13376 ( .A1(n15084), .A2(n10917), .ZN(n10892) );
  OR2_X1 U13377 ( .A1(n13906), .A2(n11085), .ZN(n10894) );
  XNOR2_X1 U13378 ( .A(n11039), .B(n13815), .ZN(n10895) );
  NOR2_X1 U13379 ( .A1(n10895), .A2(n15178), .ZN(n15186) );
  NAND2_X1 U13380 ( .A1(n14061), .A2(n15049), .ZN(n10905) );
  NAND2_X1 U13381 ( .A1(n13831), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10903) );
  OR2_X1 U13382 ( .A1(n10037), .A2(n15219), .ZN(n10902) );
  INV_X1 U13383 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10896) );
  NAND2_X1 U13384 ( .A1(n10897), .A2(n10896), .ZN(n10898) );
  NAND2_X1 U13385 ( .A1(n11040), .A2(n10898), .ZN(n11487) );
  OR2_X1 U13386 ( .A1(n13692), .A2(n11487), .ZN(n10901) );
  INV_X1 U13387 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10899) );
  OR2_X1 U13388 ( .A1(n13844), .A2(n10899), .ZN(n10900) );
  NAND4_X1 U13389 ( .A1(n10903), .A2(n10902), .A3(n10901), .A4(n10900), .ZN(
        n15050) );
  NAND2_X1 U13390 ( .A1(n15050), .A2(n15059), .ZN(n10904) );
  NAND2_X1 U13391 ( .A1(n10905), .A2(n10904), .ZN(n15183) );
  OAI21_X1 U13392 ( .B1(n15186), .B2(n15183), .A(n14379), .ZN(n10906) );
  NAND2_X1 U13393 ( .A1(n10907), .A2(n10906), .ZN(P1_U3285) );
  OAI22_X1 U13394 ( .A1(n12715), .A2(n10934), .B1(n15611), .B2(n10358), .ZN(
        n10908) );
  INV_X1 U13395 ( .A(n10908), .ZN(n10909) );
  OAI21_X1 U13396 ( .B1(n10910), .B2(n15608), .A(n10909), .ZN(P3_U3462) );
  NAND2_X1 U13397 ( .A1(n15084), .A2(n13627), .ZN(n10915) );
  NAND2_X1 U13398 ( .A1(n13607), .A2(n14062), .ZN(n10914) );
  NAND2_X1 U13399 ( .A1(n10915), .A2(n10914), .ZN(n10916) );
  XNOR2_X1 U13400 ( .A(n10916), .B(n13682), .ZN(n11079) );
  NOR2_X1 U13401 ( .A1(n13680), .A2(n10917), .ZN(n10918) );
  AOI21_X1 U13402 ( .B1(n15084), .B2(n13607), .A(n10918), .ZN(n11077) );
  XNOR2_X1 U13403 ( .A(n11079), .B(n11077), .ZN(n10919) );
  OAI211_X1 U13404 ( .C1(n10920), .C2(n10919), .A(n11081), .B(n13790), .ZN(
        n10927) );
  INV_X1 U13405 ( .A(n15084), .ZN(n10921) );
  NOR2_X1 U13406 ( .A1(n10921), .A2(n15191), .ZN(n15168) );
  NAND2_X1 U13407 ( .A1(n14061), .A2(n15059), .ZN(n10923) );
  NAND2_X1 U13408 ( .A1(n14063), .A2(n15049), .ZN(n10922) );
  AND2_X1 U13409 ( .A1(n10923), .A2(n10922), .ZN(n15170) );
  OAI21_X1 U13410 ( .B1(n13795), .B2(n15170), .A(n10924), .ZN(n10925) );
  AOI21_X1 U13411 ( .B1(n13772), .B2(n15168), .A(n10925), .ZN(n10926) );
  OAI211_X1 U13412 ( .C1(n13780), .C2(n15081), .A(n10927), .B(n10926), .ZN(
        P1_U3239) );
  XNOR2_X1 U13413 ( .A(n10212), .B(n10928), .ZN(n15137) );
  INV_X1 U13414 ( .A(n14273), .ZN(n15064) );
  NOR2_X1 U13415 ( .A1(n15064), .A2(n15065), .ZN(n10933) );
  OAI22_X1 U13416 ( .A1(n15105), .A2(n15138), .B1(n10929), .B2(n15080), .ZN(
        n10931) );
  NAND2_X1 U13417 ( .A1(n15063), .A2(n15076), .ZN(n14422) );
  AOI21_X1 U13418 ( .B1(n14422), .B2(n15096), .A(n15140), .ZN(n10930) );
  AOI211_X1 U13419 ( .C1(n15105), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10931), .B(
        n10930), .ZN(n10932) );
  OAI21_X1 U13420 ( .B1(n15137), .B2(n10933), .A(n10932), .ZN(P1_U3293) );
  OAI22_X1 U13421 ( .A1(n12595), .A2(n10934), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n12639), .ZN(n10937) );
  MUX2_X1 U13422 ( .A(n10935), .B(P3_REG2_REG_3__SCAN_IN), .S(n12648), .Z(
        n10936) );
  AOI211_X1 U13423 ( .C1(n12627), .C2(n10938), .A(n10937), .B(n10936), .ZN(
        n10939) );
  INV_X1 U13424 ( .A(n10939), .ZN(P3_U3230) );
  OAI22_X1 U13425 ( .A1(n12715), .A2(n10963), .B1(n15611), .B2(n10940), .ZN(
        n10941) );
  AOI21_X1 U13426 ( .B1(n10942), .B2(n15611), .A(n10941), .ZN(n10943) );
  INV_X1 U13427 ( .A(n10943), .ZN(P3_U3463) );
  INV_X1 U13428 ( .A(n13461), .ZN(n10946) );
  OAI222_X1 U13429 ( .A1(n14265), .A2(P1_U3086), .B1(n11699), .B2(n10946), 
        .C1(n10944), .C2(n14571), .ZN(P1_U3336) );
  OAI222_X1 U13430 ( .A1(n13417), .A2(n10947), .B1(n13399), .B2(n10946), .C1(
        n10945), .C2(P2_U3088), .ZN(P2_U3308) );
  XNOR2_X1 U13431 ( .A(n10948), .B(n10953), .ZN(n15157) );
  OAI211_X1 U13432 ( .C1(n14425), .C2(n15156), .A(n15076), .B(n10949), .ZN(
        n15154) );
  OAI22_X1 U13433 ( .A1(n15087), .A2(n15154), .B1(n10950), .B2(n15080), .ZN(
        n10952) );
  NOR2_X1 U13434 ( .A1(n14379), .A2(n10039), .ZN(n10951) );
  AOI211_X1 U13435 ( .C1(n14379), .C2(n15153), .A(n10952), .B(n10951), .ZN(
        n10956) );
  XNOR2_X1 U13436 ( .A(n10954), .B(n10953), .ZN(n15160) );
  AOI22_X1 U13437 ( .A1(n15160), .A2(n15065), .B1(n15085), .B2(n13880), .ZN(
        n10955) );
  OAI211_X1 U13438 ( .C1(n14273), .C2(n15157), .A(n10956), .B(n10955), .ZN(
        P1_U3291) );
  INV_X1 U13439 ( .A(n10957), .ZN(n10968) );
  OAI21_X1 U13440 ( .B1(n10960), .B2(n10959), .A(n10958), .ZN(n10961) );
  NAND2_X1 U13441 ( .A1(n10961), .A2(n11863), .ZN(n10967) );
  INV_X1 U13442 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10962) );
  NOR2_X1 U13443 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10962), .ZN(n15431) );
  OAI22_X1 U13444 ( .A1(n10964), .A2(n11848), .B1(n11875), .B2(n10963), .ZN(
        n10965) );
  AOI211_X1 U13445 ( .C1(n11845), .C2(n12104), .A(n15431), .B(n10965), .ZN(
        n10966) );
  OAI211_X1 U13446 ( .C1(n10968), .C2(n11613), .A(n10967), .B(n10966), .ZN(
        P3_U3170) );
  AND2_X1 U13447 ( .A1(n12824), .A2(n12983), .ZN(n11012) );
  XNOR2_X1 U13448 ( .A(n11066), .B(n11315), .ZN(n11011) );
  OAI21_X1 U13449 ( .B1(n11012), .B2(n11011), .A(n6749), .ZN(n10976) );
  INV_X1 U13450 ( .A(n10971), .ZN(n10974) );
  INV_X1 U13451 ( .A(n10972), .ZN(n10973) );
  NAND2_X1 U13452 ( .A1(n10974), .A2(n10973), .ZN(n10975) );
  XOR2_X1 U13453 ( .A(n10976), .B(n11013), .Z(n10983) );
  NOR2_X1 U13454 ( .A1(n12928), .A2(n10996), .ZN(n10981) );
  NAND2_X1 U13455 ( .A1(n12963), .A2(n12982), .ZN(n10978) );
  NAND2_X1 U13456 ( .A1(n13095), .A2(n12984), .ZN(n10977) );
  AND2_X1 U13457 ( .A1(n10978), .A2(n10977), .ZN(n10993) );
  OAI21_X1 U13458 ( .B1(n12967), .B2(n10993), .A(n10979), .ZN(n10980) );
  AOI211_X1 U13459 ( .C1(n11066), .C2(n12972), .A(n10981), .B(n10980), .ZN(
        n10982) );
  OAI21_X1 U13460 ( .B1(n10983), .B2(n12968), .A(n10982), .ZN(P2_U3208) );
  NAND2_X1 U13461 ( .A1(n10985), .A2(n10984), .ZN(n10987) );
  NAND2_X1 U13462 ( .A1(n11003), .A2(n12984), .ZN(n10986) );
  XNOR2_X1 U13463 ( .A(n11065), .B(n10990), .ZN(n15374) );
  INV_X1 U13464 ( .A(n15374), .ZN(n11001) );
  NAND2_X1 U13465 ( .A1(n10989), .A2(n10988), .ZN(n10991) );
  NAND2_X1 U13466 ( .A1(n10991), .A2(n10990), .ZN(n11061) );
  OAI21_X1 U13467 ( .B1(n10991), .B2(n10990), .A(n11061), .ZN(n10992) );
  NAND2_X1 U13468 ( .A1(n10992), .A2(n13264), .ZN(n10994) );
  NAND2_X1 U13469 ( .A1(n10994), .A2(n10993), .ZN(n15380) );
  INV_X1 U13470 ( .A(n11066), .ZN(n15377) );
  NAND2_X1 U13471 ( .A1(n15377), .A2(n10995), .ZN(n11069) );
  OAI211_X1 U13472 ( .C1(n15377), .C2(n10995), .A(n13294), .B(n11069), .ZN(
        n15375) );
  OAI22_X1 U13473 ( .A1(n13252), .A2(n9814), .B1(n10996), .B2(n13236), .ZN(
        n10997) );
  AOI21_X1 U13474 ( .B1(n11066), .B2(n13240), .A(n10997), .ZN(n10998) );
  OAI21_X1 U13475 ( .B1(n15375), .B2(n13206), .A(n10998), .ZN(n10999) );
  AOI21_X1 U13476 ( .B1(n15380), .B2(n13252), .A(n10999), .ZN(n11000) );
  OAI21_X1 U13477 ( .B1(n11001), .B2(n13256), .A(n11000), .ZN(P2_U3254) );
  AOI21_X1 U13478 ( .B1(n15366), .B2(n11003), .A(n11002), .ZN(n11004) );
  OAI211_X1 U13479 ( .C1(n15369), .C2(n11006), .A(n11005), .B(n11004), .ZN(
        n11009) );
  NAND2_X1 U13480 ( .A1(n11009), .A2(n15392), .ZN(n11007) );
  OAI21_X1 U13481 ( .B1(n15392), .B2(n11008), .A(n11007), .ZN(P2_U3509) );
  INV_X1 U13482 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U13483 ( .A1(n11009), .A2(n15383), .ZN(n11010) );
  OAI21_X1 U13484 ( .B1(n15383), .B2(n12340), .A(n11010), .ZN(P2_U3460) );
  XNOR2_X1 U13485 ( .A(n11195), .B(n12869), .ZN(n11212) );
  NAND2_X1 U13486 ( .A1(n12824), .A2(n12982), .ZN(n11213) );
  NAND3_X1 U13487 ( .A1(n11013), .A2(n12940), .A3(n12983), .ZN(n11014) );
  OAI21_X1 U13488 ( .B1(n11015), .B2(n12968), .A(n11014), .ZN(n11016) );
  NAND2_X1 U13489 ( .A1(n11016), .A2(n6747), .ZN(n11022) );
  NOR2_X1 U13490 ( .A1(n12928), .A2(n11071), .ZN(n11020) );
  NAND2_X1 U13491 ( .A1(n12963), .A2(n12981), .ZN(n11018) );
  NAND2_X1 U13492 ( .A1(n13095), .A2(n12983), .ZN(n11017) );
  AND2_X1 U13493 ( .A1(n11018), .A2(n11017), .ZN(n11062) );
  NAND2_X1 U13494 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15258)
         );
  OAI21_X1 U13495 ( .B1(n12967), .B2(n11062), .A(n15258), .ZN(n11019) );
  AOI211_X1 U13496 ( .C1(n11195), .C2(n12972), .A(n11020), .B(n11019), .ZN(
        n11021) );
  OAI211_X1 U13497 ( .C1(n12968), .C2(n11216), .A(n11022), .B(n11021), .ZN(
        P2_U3196) );
  XNOR2_X1 U13498 ( .A(n11023), .B(n13813), .ZN(n15179) );
  OAI21_X1 U13499 ( .B1(n11025), .B2(n13813), .A(n11024), .ZN(n15182) );
  OAI211_X1 U13500 ( .C1(n15079), .C2(n15177), .A(n15076), .B(n11026), .ZN(
        n15176) );
  INV_X1 U13501 ( .A(n11096), .ZN(n11027) );
  AOI22_X1 U13502 ( .A1(n15085), .A2(n13906), .B1(n15091), .B2(n11027), .ZN(
        n11030) );
  AOI22_X1 U13503 ( .A1(n15049), .A2(n14062), .B1(n14060), .B2(n15059), .ZN(
        n15175) );
  MUX2_X1 U13504 ( .A(n15175), .B(n11028), .S(n15105), .Z(n11029) );
  OAI211_X1 U13505 ( .C1(n15176), .C2(n15087), .A(n11030), .B(n11029), .ZN(
        n11031) );
  AOI21_X1 U13506 ( .B1(n15182), .B2(n15065), .A(n11031), .ZN(n11032) );
  OAI21_X1 U13507 ( .B1(n15179), .B2(n14273), .A(n11032), .ZN(P1_U3286) );
  OR2_X1 U13508 ( .A1(n13913), .A2(n14060), .ZN(n11033) );
  NAND2_X1 U13509 ( .A1(n11034), .A2(n11033), .ZN(n11038) );
  OR2_X1 U13510 ( .A1(n11035), .A2(n13836), .ZN(n11037) );
  AOI22_X1 U13511 ( .A1(n13524), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n13523), 
        .B2(n14122), .ZN(n11036) );
  XNOR2_X1 U13512 ( .A(n13917), .B(n15050), .ZN(n13817) );
  NAND2_X1 U13513 ( .A1(n11038), .A2(n6857), .ZN(n11161) );
  OAI21_X1 U13514 ( .B1(n11038), .B2(n6857), .A(n11161), .ZN(n15194) );
  INV_X1 U13515 ( .A(n15194), .ZN(n11058) );
  INV_X1 U13516 ( .A(n15100), .ZN(n14384) );
  INV_X1 U13517 ( .A(n14060), .ZN(n11260) );
  XNOR2_X1 U13518 ( .A(n11139), .B(n6857), .ZN(n11050) );
  NAND2_X1 U13519 ( .A1(n13688), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11047) );
  NAND2_X1 U13520 ( .A1(n11040), .A2(n12362), .ZN(n11041) );
  NAND2_X1 U13521 ( .A1(n11153), .A2(n11041), .ZN(n15068) );
  OR2_X1 U13522 ( .A1(n13692), .A2(n15068), .ZN(n11046) );
  INV_X1 U13523 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11042) );
  OR2_X1 U13524 ( .A1(n13844), .A2(n11042), .ZN(n11045) );
  OR2_X1 U13525 ( .A1(n13842), .A2(n11043), .ZN(n11044) );
  NAND4_X1 U13526 ( .A1(n11047), .A2(n11046), .A3(n11045), .A4(n11044), .ZN(
        n14059) );
  OAI22_X1 U13527 ( .A1(n11654), .A2(n14156), .B1(n11260), .B2(n14432), .ZN(
        n11048) );
  AOI21_X1 U13528 ( .B1(n15194), .B2(n15074), .A(n11048), .ZN(n11049) );
  OAI21_X1 U13529 ( .B1(n15178), .B2(n11050), .A(n11049), .ZN(n15192) );
  NAND2_X1 U13530 ( .A1(n15192), .A2(n14379), .ZN(n11057) );
  OAI22_X1 U13531 ( .A1(n14379), .A2(n11051), .B1(n11487), .B2(n15080), .ZN(
        n11055) );
  INV_X1 U13532 ( .A(n11052), .ZN(n11053) );
  OAI211_X1 U13533 ( .C1(n7265), .C2(n11053), .A(n7266), .B(n15076), .ZN(
        n15190) );
  NOR2_X1 U13534 ( .A1(n15190), .A2(n15087), .ZN(n11054) );
  AOI211_X1 U13535 ( .C1(n15085), .C2(n13917), .A(n11055), .B(n11054), .ZN(
        n11056) );
  OAI211_X1 U13536 ( .C1(n11058), .C2(n14384), .A(n11057), .B(n11056), .ZN(
        P1_U3284) );
  NAND2_X1 U13537 ( .A1(n11066), .A2(n11059), .ZN(n11060) );
  XNOR2_X1 U13538 ( .A(n11190), .B(n11068), .ZN(n11063) );
  OAI21_X1 U13539 ( .B1(n11063), .B2(n13247), .A(n11062), .ZN(n14928) );
  INV_X1 U13540 ( .A(n14928), .ZN(n11076) );
  AND2_X1 U13541 ( .A1(n11066), .A2(n12983), .ZN(n11064) );
  OR2_X1 U13542 ( .A1(n11066), .A2(n12983), .ZN(n11067) );
  XNOR2_X1 U13543 ( .A(n11197), .B(n11068), .ZN(n14930) );
  INV_X1 U13544 ( .A(n11069), .ZN(n11070) );
  INV_X1 U13545 ( .A(n11195), .ZN(n14927) );
  OAI211_X1 U13546 ( .C1(n11070), .C2(n14927), .A(n13294), .B(n11193), .ZN(
        n14926) );
  OAI22_X1 U13547 ( .A1(n13252), .A2(n10796), .B1(n11071), .B2(n13236), .ZN(
        n11072) );
  AOI21_X1 U13548 ( .B1(n11195), .B2(n13240), .A(n11072), .ZN(n11073) );
  OAI21_X1 U13549 ( .B1(n14926), .B2(n13206), .A(n11073), .ZN(n11074) );
  AOI21_X1 U13550 ( .B1(n14930), .B2(n13280), .A(n11074), .ZN(n11075) );
  OAI21_X1 U13551 ( .B1(n11076), .B2(n13282), .A(n11075), .ZN(P2_U3253) );
  INV_X1 U13552 ( .A(n11077), .ZN(n11078) );
  NAND2_X1 U13553 ( .A1(n11079), .A2(n11078), .ZN(n11080) );
  NAND2_X1 U13554 ( .A1(n11081), .A2(n11080), .ZN(n11088) );
  NAND2_X1 U13555 ( .A1(n13906), .A2(n13627), .ZN(n11083) );
  NAND2_X1 U13556 ( .A1(n13607), .A2(n14061), .ZN(n11082) );
  NAND2_X1 U13557 ( .A1(n11083), .A2(n11082), .ZN(n11084) );
  XNOR2_X1 U13558 ( .A(n11084), .B(n13682), .ZN(n11264) );
  NOR2_X1 U13559 ( .A1(n13680), .A2(n11085), .ZN(n11086) );
  AOI21_X1 U13560 ( .B1(n13906), .B2(n13607), .A(n11086), .ZN(n11262) );
  XNOR2_X1 U13561 ( .A(n11264), .B(n11262), .ZN(n11087) );
  OAI211_X1 U13562 ( .C1(n11088), .C2(n11087), .A(n11266), .B(n13790), .ZN(
        n11095) );
  NAND2_X1 U13563 ( .A1(n13782), .A2(n13906), .ZN(n11092) );
  INV_X1 U13564 ( .A(n11089), .ZN(n11090) );
  AOI21_X1 U13565 ( .B1(n13777), .B2(n14062), .A(n11090), .ZN(n11091) );
  OAI211_X1 U13566 ( .C1(n11260), .C2(n13762), .A(n11092), .B(n11091), .ZN(
        n11093) );
  INV_X1 U13567 ( .A(n11093), .ZN(n11094) );
  OAI211_X1 U13568 ( .C1(n13780), .C2(n11096), .A(n11095), .B(n11094), .ZN(
        P1_U3213) );
  XOR2_X1 U13569 ( .A(n11098), .B(n11097), .Z(n11104) );
  NOR2_X1 U13570 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11099), .ZN(n15451) );
  OAI22_X1 U13571 ( .A1(n11106), .A2(n11848), .B1(n11875), .B2(n11100), .ZN(
        n11101) );
  AOI211_X1 U13572 ( .C1(n11845), .C2(n12103), .A(n15451), .B(n11101), .ZN(
        n11103) );
  NAND2_X1 U13573 ( .A1(n11872), .A2(n11113), .ZN(n11102) );
  OAI211_X1 U13574 ( .C1(n11104), .C2(n11852), .A(n11103), .B(n11102), .ZN(
        P3_U3167) );
  XNOR2_X1 U13575 ( .A(n11105), .B(n7430), .ZN(n15583) );
  INV_X1 U13576 ( .A(n15583), .ZN(n11116) );
  OAI22_X1 U13577 ( .A1(n11106), .A2(n12587), .B1(n11288), .B2(n12589), .ZN(
        n11111) );
  NAND2_X1 U13578 ( .A1(n11107), .A2(n7430), .ZN(n11108) );
  AOI21_X1 U13579 ( .B1(n11109), .B2(n11108), .A(n12584), .ZN(n11110) );
  AOI211_X1 U13580 ( .C1(n15583), .C2(n11370), .A(n11111), .B(n11110), .ZN(
        n15580) );
  MUX2_X1 U13581 ( .A(n15445), .B(n15580), .S(n14895), .Z(n11115) );
  AND2_X1 U13582 ( .A1(n11112), .A2(n14898), .ZN(n15582) );
  AOI22_X1 U13583 ( .A1(n11415), .A2(n15582), .B1(n12624), .B2(n11113), .ZN(
        n11114) );
  OAI211_X1 U13584 ( .C1(n11116), .C2(n11357), .A(n11115), .B(n11114), .ZN(
        P3_U3228) );
  OR2_X1 U13585 ( .A1(n11117), .A2(n11909), .ZN(n11118) );
  NAND2_X1 U13586 ( .A1(n11119), .A2(n11118), .ZN(n11187) );
  OR2_X1 U13587 ( .A1(n11120), .A2(n11909), .ZN(n11122) );
  NAND2_X1 U13588 ( .A1(n11120), .A2(n11909), .ZN(n11121) );
  NAND3_X1 U13589 ( .A1(n11122), .A2(n12636), .A3(n11121), .ZN(n11124) );
  AOI22_X1 U13590 ( .A1(n12104), .A2(n12631), .B1(n12633), .B2(n12102), .ZN(
        n11123) );
  NAND2_X1 U13591 ( .A1(n11124), .A2(n11123), .ZN(n11183) );
  AOI21_X1 U13592 ( .B1(n15595), .B2(n11187), .A(n11183), .ZN(n11131) );
  INV_X1 U13593 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11125) );
  OAI22_X1 U13594 ( .A1(n11205), .A2(n12770), .B1(n15599), .B2(n11125), .ZN(
        n11126) );
  INV_X1 U13595 ( .A(n11126), .ZN(n11127) );
  OAI21_X1 U13596 ( .B1(n11131), .B2(n15601), .A(n11127), .ZN(P3_U3408) );
  OAI22_X1 U13597 ( .A1(n12715), .A2(n11205), .B1(n15611), .B2(n11128), .ZN(
        n11129) );
  INV_X1 U13598 ( .A(n11129), .ZN(n11130) );
  OAI21_X1 U13599 ( .B1(n11131), .B2(n15608), .A(n11130), .ZN(P3_U3465) );
  NAND2_X1 U13600 ( .A1(n13832), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11138) );
  OR2_X1 U13601 ( .A1(n13842), .A2(n10062), .ZN(n11137) );
  OR2_X1 U13602 ( .A1(n10037), .A2(n14803), .ZN(n11136) );
  INV_X1 U13603 ( .A(n11153), .ZN(n11132) );
  AOI21_X1 U13604 ( .B1(n11132), .B2(P1_REG3_REG_11__SCAN_IN), .A(
        P1_REG3_REG_12__SCAN_IN), .ZN(n11134) );
  NAND2_X1 U13605 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n11133) );
  NOR2_X1 U13606 ( .A1(n11153), .A2(n11133), .ZN(n11240) );
  OR2_X1 U13607 ( .A1(n11134), .A2(n11240), .ZN(n11672) );
  OR2_X1 U13608 ( .A1(n13692), .A2(n11672), .ZN(n11135) );
  INV_X1 U13609 ( .A(n15050), .ZN(n11452) );
  NAND2_X1 U13610 ( .A1(n13917), .A2(n11452), .ZN(n11140) );
  INV_X1 U13611 ( .A(n15055), .ZN(n11146) );
  NAND2_X1 U13612 ( .A1(n11141), .A2(n11615), .ZN(n11144) );
  AOI22_X1 U13613 ( .A1(n13524), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n13523), 
        .B2(n11142), .ZN(n11143) );
  XNOR2_X1 U13614 ( .A(n15201), .B(n11654), .ZN(n15054) );
  INV_X1 U13615 ( .A(n15054), .ZN(n11145) );
  OR2_X1 U13616 ( .A1(n15201), .A2(n11654), .ZN(n11147) );
  NAND2_X1 U13617 ( .A1(n11148), .A2(n11615), .ZN(n11151) );
  AOI22_X1 U13618 ( .A1(n13524), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n13523), 
        .B2(n11149), .ZN(n11150) );
  NAND2_X1 U13619 ( .A1(n13831), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11158) );
  OR2_X1 U13620 ( .A1(n10037), .A2(n14955), .ZN(n11157) );
  INV_X1 U13621 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11152) );
  XNOR2_X1 U13622 ( .A(n11153), .B(n11152), .ZN(n11658) );
  OR2_X1 U13623 ( .A1(n13692), .A2(n11658), .ZN(n11156) );
  INV_X1 U13624 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11154) );
  OR2_X1 U13625 ( .A1(n13844), .A2(n11154), .ZN(n11155) );
  NAND4_X1 U13626 ( .A1(n11158), .A2(n11157), .A3(n11156), .A4(n11155), .ZN(
        n15060) );
  XNOR2_X1 U13627 ( .A(n13924), .B(n13925), .ZN(n13819) );
  XNOR2_X1 U13628 ( .A(n11235), .B(n13819), .ZN(n11159) );
  AOI222_X1 U13629 ( .A1(n14058), .A2(n15059), .B1(n14059), .B2(n15049), .C1(
        n15196), .C2(n11159), .ZN(n14951) );
  OR2_X1 U13630 ( .A1(n13917), .A2(n15050), .ZN(n11160) );
  NAND2_X1 U13631 ( .A1(n11161), .A2(n11160), .ZN(n15053) );
  OR2_X1 U13632 ( .A1(n15201), .A2(n14059), .ZN(n11162) );
  XNOR2_X1 U13633 ( .A(n11231), .B(n13819), .ZN(n14954) );
  INV_X1 U13634 ( .A(n15201), .ZN(n11163) );
  INV_X1 U13635 ( .A(n13924), .ZN(n14952) );
  OAI211_X1 U13636 ( .C1(n6601), .C2(n14952), .A(n15076), .B(n11251), .ZN(
        n14950) );
  OAI22_X1 U13637 ( .A1(n14379), .A2(n11164), .B1(n11658), .B2(n15080), .ZN(
        n11165) );
  AOI21_X1 U13638 ( .B1(n13924), .B2(n15085), .A(n11165), .ZN(n11166) );
  OAI21_X1 U13639 ( .B1(n14950), .B2(n15087), .A(n11166), .ZN(n11167) );
  AOI21_X1 U13640 ( .B1(n14954), .B2(n15065), .A(n11167), .ZN(n11168) );
  OAI21_X1 U13641 ( .B1(n14951), .B2(n15093), .A(n11168), .ZN(P1_U3282) );
  NAND2_X1 U13642 ( .A1(n13508), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14137) );
  OAI21_X1 U13643 ( .B1(n13508), .B2(P1_REG2_REG_17__SCAN_IN), .A(n14137), 
        .ZN(n14133) );
  OAI21_X1 U13644 ( .B1(n11170), .B2(n11173), .A(n11169), .ZN(n14135) );
  XOR2_X1 U13645 ( .A(n14133), .B(n14135), .Z(n11182) );
  NAND2_X1 U13646 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13734)
         );
  XNOR2_X1 U13647 ( .A(n14128), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11177) );
  INV_X1 U13648 ( .A(n11171), .ZN(n11175) );
  INV_X1 U13649 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11172) );
  OAI22_X1 U13650 ( .A1(n11175), .A2(n11174), .B1(n11173), .B2(n11172), .ZN(
        n11176) );
  NAND2_X1 U13651 ( .A1(n11176), .A2(n11177), .ZN(n14127) );
  OAI211_X1 U13652 ( .C1(n11177), .C2(n11176), .A(n15028), .B(n14127), .ZN(
        n11178) );
  NAND2_X1 U13653 ( .A1(n13734), .A2(n11178), .ZN(n11180) );
  NOR2_X1 U13654 ( .A1(n15043), .A2(n14128), .ZN(n11179) );
  AOI211_X1 U13655 ( .C1(n15018), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n11180), 
        .B(n11179), .ZN(n11181) );
  OAI21_X1 U13656 ( .B1(n11182), .B2(n15039), .A(n11181), .ZN(P1_U3260) );
  MUX2_X1 U13657 ( .A(n11183), .B(P3_REG2_REG_6__SCAN_IN), .S(n12648), .Z(
        n11184) );
  INV_X1 U13658 ( .A(n11184), .ZN(n11189) );
  INV_X1 U13659 ( .A(n11185), .ZN(n11211) );
  OAI22_X1 U13660 ( .A1(n12595), .A2(n11205), .B1(n11211), .B2(n12639), .ZN(
        n11186) );
  AOI21_X1 U13661 ( .B1(n11187), .B2(n12627), .A(n11186), .ZN(n11188) );
  NAND2_X1 U13662 ( .A1(n11189), .A2(n11188), .ZN(P3_U3227) );
  NAND2_X1 U13663 ( .A1(n11190), .A2(n11195), .ZN(n11191) );
  XOR2_X1 U13664 ( .A(n11198), .B(n11299), .Z(n11192) );
  OAI22_X1 U13665 ( .A1(n11499), .A2(n13031), .B1(n11196), .B2(n12916), .ZN(
        n11224) );
  AOI21_X1 U13666 ( .B1(n11192), .B2(n13264), .A(n11224), .ZN(n13376) );
  AOI211_X1 U13667 ( .C1(n13374), .C2(n11193), .A(n13270), .B(n11309), .ZN(
        n13373) );
  AOI22_X1 U13668 ( .A1(n13282), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11228), 
        .B2(n13273), .ZN(n11194) );
  OAI21_X1 U13669 ( .B1(n7537), .B2(n13277), .A(n11194), .ZN(n11200) );
  XNOR2_X1 U13670 ( .A(n11304), .B(n11198), .ZN(n13377) );
  NOR2_X1 U13671 ( .A1(n13377), .A2(n13256), .ZN(n11199) );
  AOI211_X1 U13672 ( .C1(n13373), .C2(n13272), .A(n11200), .B(n11199), .ZN(
        n11201) );
  OAI21_X1 U13673 ( .B1(n13282), .B2(n13376), .A(n11201), .ZN(P2_U3252) );
  OAI211_X1 U13674 ( .C1(n11202), .C2(n11204), .A(n11203), .B(n11863), .ZN(
        n11210) );
  OAI22_X1 U13675 ( .A1(n11206), .A2(n11848), .B1(n11875), .B2(n11205), .ZN(
        n11207) );
  AOI211_X1 U13676 ( .C1(n11845), .C2(n12102), .A(n11208), .B(n11207), .ZN(
        n11209) );
  OAI211_X1 U13677 ( .C1(n11211), .C2(n11613), .A(n11210), .B(n11209), .ZN(
        P3_U3179) );
  INV_X1 U13678 ( .A(n11212), .ZN(n11214) );
  NAND2_X1 U13679 ( .A1(n11214), .A2(n11213), .ZN(n11215) );
  XNOR2_X1 U13680 ( .A(n13374), .B(n11315), .ZN(n11317) );
  AND2_X1 U13681 ( .A1(n12981), .A2(n12824), .ZN(n11217) );
  NAND2_X1 U13682 ( .A1(n11317), .A2(n11217), .ZN(n11316) );
  INV_X1 U13683 ( .A(n11317), .ZN(n11219) );
  INV_X1 U13684 ( .A(n11217), .ZN(n11218) );
  NAND2_X1 U13685 ( .A1(n11219), .A2(n11218), .ZN(n11220) );
  NAND2_X1 U13686 ( .A1(n11316), .A2(n11220), .ZN(n11221) );
  AOI21_X1 U13687 ( .B1(n11222), .B2(n11221), .A(n12968), .ZN(n11223) );
  NAND2_X1 U13688 ( .A1(n11223), .A2(n11319), .ZN(n11230) );
  INV_X1 U13689 ( .A(n11224), .ZN(n11226) );
  OAI22_X1 U13690 ( .A1(n12967), .A2(n11226), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11225), .ZN(n11227) );
  AOI21_X1 U13691 ( .B1(n12965), .B2(n11228), .A(n11227), .ZN(n11229) );
  OAI211_X1 U13692 ( .C1(n7537), .C2(n12957), .A(n11230), .B(n11229), .ZN(
        P2_U3206) );
  NAND2_X1 U13693 ( .A1(n11232), .A2(n11615), .ZN(n11234) );
  AOI22_X1 U13694 ( .A1(n13524), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n15013), 
        .B2(n13523), .ZN(n11233) );
  XNOR2_X1 U13695 ( .A(n13930), .B(n13929), .ZN(n13820) );
  XNOR2_X1 U13696 ( .A(n11420), .B(n13820), .ZN(n14799) );
  NAND2_X1 U13697 ( .A1(n13924), .A2(n13925), .ZN(n11236) );
  NAND2_X1 U13698 ( .A1(n11237), .A2(n11236), .ZN(n11238) );
  NAND2_X1 U13699 ( .A1(n11238), .A2(n13820), .ZN(n11239) );
  NAND2_X1 U13700 ( .A1(n11239), .A2(n15196), .ZN(n11249) );
  NAND2_X1 U13701 ( .A1(n13832), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11245) );
  OR2_X1 U13702 ( .A1(n10037), .A2(n14949), .ZN(n11244) );
  OR2_X1 U13703 ( .A1(n13842), .A2(n10058), .ZN(n11243) );
  NAND2_X1 U13704 ( .A1(n11240), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11530) );
  OR2_X1 U13705 ( .A1(n11240), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11241) );
  NAND2_X1 U13706 ( .A1(n11530), .A2(n11241), .ZN(n11689) );
  OR2_X1 U13707 ( .A1(n13692), .A2(n11689), .ZN(n11242) );
  NAND4_X1 U13708 ( .A1(n11245), .A2(n11244), .A3(n11243), .A4(n11242), .ZN(
        n14057) );
  NAND2_X1 U13709 ( .A1(n14057), .A2(n15059), .ZN(n11247) );
  NAND2_X1 U13710 ( .A1(n15060), .A2(n15049), .ZN(n11246) );
  NAND2_X1 U13711 ( .A1(n11247), .A2(n11246), .ZN(n11675) );
  INV_X1 U13712 ( .A(n11675), .ZN(n11248) );
  OAI21_X1 U13713 ( .B1(n11426), .B2(n11249), .A(n11248), .ZN(n11250) );
  AOI21_X1 U13714 ( .B1(n14799), .B2(n15074), .A(n11250), .ZN(n14801) );
  INV_X1 U13715 ( .A(n11251), .ZN(n11252) );
  NAND2_X1 U13716 ( .A1(n14797), .A2(n11252), .ZN(n11434) );
  OAI211_X1 U13717 ( .C1(n14797), .C2(n11252), .A(n15076), .B(n11434), .ZN(
        n14796) );
  OAI22_X1 U13718 ( .A1(n14379), .A2(n10062), .B1(n11672), .B2(n15080), .ZN(
        n11253) );
  AOI21_X1 U13719 ( .B1(n13930), .B2(n15085), .A(n11253), .ZN(n11254) );
  OAI21_X1 U13720 ( .B1(n14796), .B2(n15087), .A(n11254), .ZN(n11255) );
  AOI21_X1 U13721 ( .B1(n14799), .B2(n15100), .A(n11255), .ZN(n11256) );
  OAI21_X1 U13722 ( .B1(n14801), .B2(n15093), .A(n11256), .ZN(P1_U3281) );
  NAND2_X1 U13723 ( .A1(n13913), .A2(n13627), .ZN(n11258) );
  NAND2_X1 U13724 ( .A1(n13607), .A2(n14060), .ZN(n11257) );
  NAND2_X1 U13725 ( .A1(n11258), .A2(n11257), .ZN(n11259) );
  XNOR2_X1 U13726 ( .A(n11259), .B(n13517), .ZN(n11449) );
  NOR2_X1 U13727 ( .A1(n13680), .A2(n11260), .ZN(n11261) );
  AOI21_X1 U13728 ( .B1(n13913), .B2(n13607), .A(n11261), .ZN(n11448) );
  XNOR2_X1 U13729 ( .A(n11449), .B(n11448), .ZN(n11269) );
  INV_X1 U13730 ( .A(n11262), .ZN(n11263) );
  NAND2_X1 U13731 ( .A1(n11264), .A2(n11263), .ZN(n11265) );
  INV_X1 U13732 ( .A(n11451), .ZN(n11267) );
  AOI21_X1 U13733 ( .B1(n11269), .B2(n11268), .A(n11267), .ZN(n11274) );
  NOR2_X1 U13734 ( .A1(n7592), .A2(n15191), .ZN(n15184) );
  AOI22_X1 U13735 ( .A1(n13650), .A2(n15183), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11270) );
  OAI21_X1 U13736 ( .B1(n13780), .B2(n11271), .A(n11270), .ZN(n11272) );
  AOI21_X1 U13737 ( .B1(n13772), .B2(n15184), .A(n11272), .ZN(n11273) );
  OAI21_X1 U13738 ( .B1(n11274), .B2(n13784), .A(n11273), .ZN(P1_U3221) );
  NAND2_X1 U13739 ( .A1(n11275), .A2(n11912), .ZN(n11364) );
  OAI211_X1 U13740 ( .C1(n11275), .C2(n11912), .A(n11364), .B(n12636), .ZN(
        n11277) );
  OR2_X1 U13741 ( .A1(n11288), .A2(n12587), .ZN(n11276) );
  OAI211_X1 U13742 ( .C1(n11564), .C2(n12589), .A(n11277), .B(n11276), .ZN(
        n11378) );
  INV_X1 U13743 ( .A(n11378), .ZN(n11283) );
  OAI21_X1 U13744 ( .B1(n11279), .B2(n11962), .A(n11278), .ZN(n11379) );
  AOI22_X1 U13745 ( .A1(n12648), .A2(P3_REG2_REG_7__SCAN_IN), .B1(n12624), 
        .B2(n11284), .ZN(n11280) );
  OAI21_X1 U13746 ( .B1(n12595), .B2(n11965), .A(n11280), .ZN(n11281) );
  AOI21_X1 U13747 ( .B1(n11379), .B2(n12627), .A(n11281), .ZN(n11282) );
  OAI21_X1 U13748 ( .B1(n11283), .B2(n12648), .A(n11282), .ZN(P3_U3226) );
  INV_X1 U13749 ( .A(n11284), .ZN(n11293) );
  OAI211_X1 U13750 ( .C1(n11287), .C2(n11286), .A(n11285), .B(n11863), .ZN(
        n11292) );
  OAI22_X1 U13751 ( .A1(n11288), .A2(n11848), .B1(n11875), .B2(n11965), .ZN(
        n11289) );
  AOI211_X1 U13752 ( .C1(n11845), .C2(n12101), .A(n11290), .B(n11289), .ZN(
        n11291) );
  OAI211_X1 U13753 ( .C1(n11293), .C2(n11613), .A(n11292), .B(n11291), .ZN(
        P3_U3153) );
  INV_X1 U13754 ( .A(n11294), .ZN(n11296) );
  OAI222_X1 U13755 ( .A1(n11297), .A2(P3_U3151), .B1(n14787), .B2(n11296), 
        .C1(n11295), .C2(n12784), .ZN(P3_U3270) );
  INV_X1 U13756 ( .A(n13541), .ZN(n11330) );
  OAI222_X1 U13757 ( .A1(P1_U3086), .A2(n11298), .B1(n11699), .B2(n11330), 
        .C1(n13542), .C2(n14571), .ZN(P1_U3335) );
  OR2_X1 U13758 ( .A1(n13374), .A2(n11300), .ZN(n11301) );
  XNOR2_X1 U13759 ( .A(n11498), .B(n11307), .ZN(n11302) );
  AOI22_X1 U13760 ( .A1(n12979), .A2(n12963), .B1(n13095), .B2(n12981), .ZN(
        n11322) );
  OAI21_X1 U13761 ( .B1(n11302), .B2(n13247), .A(n11322), .ZN(n11442) );
  INV_X1 U13762 ( .A(n11442), .ZN(n11314) );
  AND2_X1 U13763 ( .A1(n13374), .A2(n12981), .ZN(n11303) );
  OR2_X1 U13764 ( .A1(n13374), .A2(n12981), .ZN(n11305) );
  NAND2_X1 U13765 ( .A1(n11307), .A2(n11306), .ZN(n11308) );
  AND2_X1 U13766 ( .A1(n11507), .A2(n11308), .ZN(n11444) );
  OAI211_X1 U13767 ( .C1(n7536), .C2(n11309), .A(n13294), .B(n11502), .ZN(
        n11441) );
  AOI22_X1 U13768 ( .A1(n13282), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11324), 
        .B2(n13273), .ZN(n11311) );
  NAND2_X1 U13769 ( .A1(n11505), .A2(n13240), .ZN(n11310) );
  OAI211_X1 U13770 ( .C1(n11441), .C2(n13206), .A(n11311), .B(n11310), .ZN(
        n11312) );
  AOI21_X1 U13771 ( .B1(n13280), .B2(n11444), .A(n11312), .ZN(n11313) );
  OAI21_X1 U13772 ( .B1(n11314), .B2(n13282), .A(n11313), .ZN(P2_U3251) );
  XNOR2_X1 U13773 ( .A(n11505), .B(n11315), .ZN(n11545) );
  NAND2_X1 U13774 ( .A1(n12980), .A2(n12824), .ZN(n11546) );
  XNOR2_X1 U13775 ( .A(n11545), .B(n11546), .ZN(n11320) );
  NAND3_X1 U13776 ( .A1(n11320), .A2(n11316), .A3(n11319), .ZN(n11549) );
  NAND3_X1 U13777 ( .A1(n11317), .A2(n12940), .A3(n12981), .ZN(n11318) );
  OAI21_X1 U13778 ( .B1(n11319), .B2(n12968), .A(n11318), .ZN(n11328) );
  INV_X1 U13779 ( .A(n11320), .ZN(n11327) );
  OAI22_X1 U13780 ( .A1(n12967), .A2(n11322), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11321), .ZN(n11323) );
  AOI21_X1 U13781 ( .B1(n12965), .B2(n11324), .A(n11323), .ZN(n11325) );
  OAI21_X1 U13782 ( .B1(n7536), .B2(n12957), .A(n11325), .ZN(n11326) );
  AOI21_X1 U13783 ( .B1(n11328), .B2(n11327), .A(n11326), .ZN(n11329) );
  OAI21_X1 U13784 ( .B1(n11549), .B2(n12968), .A(n11329), .ZN(P2_U3187) );
  OAI222_X1 U13785 ( .A1(n13417), .A2(n11331), .B1(P2_U3088), .B2(n7288), .C1(
        n13399), .C2(n11330), .ZN(P2_U3307) );
  NAND2_X1 U13786 ( .A1(n15304), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11335) );
  INV_X1 U13787 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11333) );
  INV_X1 U13788 ( .A(n11335), .ZN(n11332) );
  AOI21_X1 U13789 ( .B1(n11333), .B2(n11342), .A(n11332), .ZN(n15308) );
  OAI21_X1 U13790 ( .B1(n11341), .B2(n11586), .A(n11334), .ZN(n15309) );
  NAND2_X1 U13791 ( .A1(n15308), .A2(n15309), .ZN(n15307) );
  NAND2_X1 U13792 ( .A1(n11335), .A2(n15307), .ZN(n13009) );
  XNOR2_X1 U13793 ( .A(n13014), .B(n13009), .ZN(n11336) );
  NOR2_X1 U13794 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11336), .ZN(n13011) );
  AOI21_X1 U13795 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n11336), .A(n13011), 
        .ZN(n11349) );
  INV_X1 U13796 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n11338) );
  NAND2_X1 U13797 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n11337)
         );
  OAI21_X1 U13798 ( .B1(n15260), .B2(n11338), .A(n11337), .ZN(n11347) );
  XNOR2_X1 U13799 ( .A(n11342), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15302) );
  INV_X1 U13800 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11340) );
  OAI21_X1 U13801 ( .B1(n11341), .B2(n11340), .A(n11339), .ZN(n15303) );
  NAND2_X1 U13802 ( .A1(n15302), .A2(n15303), .ZN(n15301) );
  OAI21_X1 U13803 ( .B1(n11343), .B2(n11342), .A(n15301), .ZN(n13013) );
  XOR2_X1 U13804 ( .A(n13014), .B(n13013), .Z(n11344) );
  NAND2_X1 U13805 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11344), .ZN(n13016) );
  OAI21_X1 U13806 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n11344), .A(n13016), 
        .ZN(n11345) );
  NOR2_X1 U13807 ( .A1(n11345), .A2(n15265), .ZN(n11346) );
  AOI211_X1 U13808 ( .C1(n15305), .C2(n13014), .A(n11347), .B(n11346), .ZN(
        n11348) );
  OAI21_X1 U13809 ( .B1(n11349), .B2(n15270), .A(n11348), .ZN(P2_U3232) );
  XNOR2_X1 U13810 ( .A(n11350), .B(n11352), .ZN(n11356) );
  INV_X1 U13811 ( .A(n11352), .ZN(n11975) );
  XNOR2_X1 U13812 ( .A(n11351), .B(n11975), .ZN(n11354) );
  OAI22_X1 U13813 ( .A1(n11836), .A2(n12589), .B1(n11564), .B2(n12587), .ZN(
        n11353) );
  AOI21_X1 U13814 ( .B1(n11354), .B2(n12636), .A(n11353), .ZN(n11355) );
  OAI21_X1 U13815 ( .B1(n12433), .B2(n11356), .A(n11355), .ZN(n15589) );
  INV_X1 U13816 ( .A(n15589), .ZN(n11362) );
  INV_X1 U13817 ( .A(n11356), .ZN(n15592) );
  INV_X1 U13818 ( .A(n11357), .ZN(n12438) );
  INV_X1 U13819 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11359) );
  NOR2_X1 U13820 ( .A1(n11979), .A2(n12621), .ZN(n15590) );
  AOI22_X1 U13821 ( .A1(n11415), .A2(n15590), .B1(n12624), .B2(n11566), .ZN(
        n11358) );
  OAI21_X1 U13822 ( .B1(n11359), .B2(n14895), .A(n11358), .ZN(n11360) );
  AOI21_X1 U13823 ( .B1(n15592), .B2(n12438), .A(n11360), .ZN(n11361) );
  OAI21_X1 U13824 ( .B1(n11362), .B2(n12648), .A(n11361), .ZN(P3_U3224) );
  NAND2_X1 U13825 ( .A1(n11364), .A2(n11363), .ZN(n11365) );
  XOR2_X1 U13826 ( .A(n11969), .B(n11365), .Z(n11372) );
  OR2_X1 U13827 ( .A1(n11366), .A2(n11969), .ZN(n11367) );
  NAND2_X1 U13828 ( .A1(n11368), .A2(n11367), .ZN(n15587) );
  OAI22_X1 U13829 ( .A1(n11394), .A2(n12587), .B1(n11609), .B2(n12589), .ZN(
        n11369) );
  AOI21_X1 U13830 ( .B1(n15587), .B2(n11370), .A(n11369), .ZN(n11371) );
  OAI21_X1 U13831 ( .B1(n11372), .B2(n12584), .A(n11371), .ZN(n15585) );
  INV_X1 U13832 ( .A(n15585), .ZN(n11377) );
  INV_X1 U13833 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11374) );
  NOR2_X1 U13834 ( .A1(n11971), .A2(n12621), .ZN(n15586) );
  AOI22_X1 U13835 ( .A1(n11415), .A2(n15586), .B1(n12624), .B2(n11390), .ZN(
        n11373) );
  OAI21_X1 U13836 ( .B1(n11374), .B2(n14895), .A(n11373), .ZN(n11375) );
  AOI21_X1 U13837 ( .B1(n15587), .B2(n12438), .A(n11375), .ZN(n11376) );
  OAI21_X1 U13838 ( .B1(n11377), .B2(n12648), .A(n11376), .ZN(P3_U3225) );
  AOI21_X1 U13839 ( .B1(n15595), .B2(n11379), .A(n11378), .ZN(n11386) );
  INV_X1 U13840 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11380) );
  OAI22_X1 U13841 ( .A1(n11965), .A2(n12770), .B1(n15599), .B2(n11380), .ZN(
        n11381) );
  INV_X1 U13842 ( .A(n11381), .ZN(n11382) );
  OAI21_X1 U13843 ( .B1(n11386), .B2(n15601), .A(n11382), .ZN(P3_U3411) );
  INV_X1 U13844 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11383) );
  OAI22_X1 U13845 ( .A1(n12715), .A2(n11965), .B1(n15611), .B2(n11383), .ZN(
        n11384) );
  INV_X1 U13846 ( .A(n11384), .ZN(n11385) );
  OAI21_X1 U13847 ( .B1(n11386), .B2(n15608), .A(n11385), .ZN(P3_U3466) );
  INV_X1 U13848 ( .A(n13450), .ZN(n11389) );
  OAI222_X1 U13849 ( .A1(n13417), .A2(n11388), .B1(n13399), .B2(n11389), .C1(
        n11387), .C2(P2_U3088), .ZN(P2_U3306) );
  INV_X1 U13850 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n13451) );
  OAI222_X1 U13851 ( .A1(n13862), .A2(P1_U3086), .B1(n11699), .B2(n11389), 
        .C1(n13451), .C2(n14571), .ZN(P1_U3334) );
  INV_X1 U13852 ( .A(n11390), .ZN(n11398) );
  OAI211_X1 U13853 ( .C1(n11393), .C2(n11392), .A(n11391), .B(n11863), .ZN(
        n11397) );
  AND2_X1 U13854 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n12403) );
  OAI22_X1 U13855 ( .A1(n11394), .A2(n11848), .B1(n11875), .B2(n11971), .ZN(
        n11395) );
  AOI211_X1 U13856 ( .C1(n11845), .C2(n12100), .A(n12403), .B(n11395), .ZN(
        n11396) );
  OAI211_X1 U13857 ( .C1(n11398), .C2(n11613), .A(n11397), .B(n11396), .ZN(
        P3_U3161) );
  INV_X1 U13858 ( .A(n11399), .ZN(n11400) );
  OAI222_X1 U13859 ( .A1(P3_U3151), .A2(n11402), .B1(n12784), .B2(n11401), 
        .C1(n14787), .C2(n11400), .ZN(P3_U3269) );
  AOI222_X1 U13860 ( .A1(n11404), .A2(n13404), .B1(P1_DATAO_REG_22__SCAN_IN), 
        .B2(n13397), .C1(n11403), .C2(P2_STATE_REG_SCAN_IN), .ZN(n11405) );
  INV_X1 U13861 ( .A(n11405), .ZN(P2_U3305) );
  INV_X1 U13862 ( .A(n11917), .ZN(n11988) );
  XNOR2_X1 U13863 ( .A(n11406), .B(n11988), .ZN(n11408) );
  OAI22_X1 U13864 ( .A1(n11836), .A2(n12587), .B1(n11820), .B2(n12589), .ZN(
        n11407) );
  AOI21_X1 U13865 ( .B1(n11408), .B2(n12636), .A(n11407), .ZN(n14916) );
  NAND2_X1 U13866 ( .A1(n11409), .A2(n11410), .ZN(n11411) );
  NAND2_X1 U13867 ( .A1(n11411), .A2(n11917), .ZN(n11413) );
  NAND2_X1 U13868 ( .A1(n11413), .A2(n11412), .ZN(n14914) );
  INV_X1 U13869 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11417) );
  AND2_X1 U13870 ( .A1(n11414), .A2(n14898), .ZN(n14913) );
  AOI22_X1 U13871 ( .A1(n11415), .A2(n14913), .B1(n12624), .B2(n11838), .ZN(
        n11416) );
  OAI21_X1 U13872 ( .B1(n11417), .B2(n14895), .A(n11416), .ZN(n11418) );
  AOI21_X1 U13873 ( .B1(n14914), .B2(n12627), .A(n11418), .ZN(n11419) );
  OAI21_X1 U13874 ( .B1(n14916), .B2(n12648), .A(n11419), .ZN(P3_U3222) );
  NAND2_X1 U13875 ( .A1(n14797), .A2(n13929), .ZN(n11421) );
  NAND2_X1 U13876 ( .A1(n11422), .A2(n11615), .ZN(n11425) );
  AOI22_X1 U13877 ( .A1(n13524), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n13523), 
        .B2(n11423), .ZN(n11424) );
  XNOR2_X1 U13878 ( .A(n13934), .B(n14057), .ZN(n13821) );
  XNOR2_X1 U13879 ( .A(n11521), .B(n11520), .ZN(n14948) );
  INV_X1 U13880 ( .A(n14948), .ZN(n11440) );
  AOI211_X1 U13881 ( .C1(n11520), .C2(n6744), .A(n15178), .B(n11513), .ZN(
        n14946) );
  NAND2_X1 U13882 ( .A1(n13832), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11430) );
  OR2_X1 U13883 ( .A1(n13842), .A2(n11525), .ZN(n11429) );
  OR2_X1 U13884 ( .A1(n10037), .A2(n14942), .ZN(n11428) );
  INV_X1 U13885 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11528) );
  XNOR2_X1 U13886 ( .A(n11530), .B(n11528), .ZN(n13653) );
  OR2_X1 U13887 ( .A1(n13692), .A2(n13653), .ZN(n11427) );
  OR2_X1 U13888 ( .A1(n13485), .A2(n14156), .ZN(n11432) );
  OR2_X1 U13889 ( .A1(n13929), .A2(n14432), .ZN(n11431) );
  AND2_X1 U13890 ( .A1(n11432), .A2(n11431), .ZN(n14943) );
  INV_X1 U13891 ( .A(n14943), .ZN(n11433) );
  OAI21_X1 U13892 ( .B1(n14946), .B2(n11433), .A(n14379), .ZN(n11439) );
  OAI22_X1 U13893 ( .A1(n14379), .A2(n10058), .B1(n11689), .B2(n15080), .ZN(
        n11437) );
  INV_X1 U13894 ( .A(n13934), .ZN(n14945) );
  INV_X1 U13895 ( .A(n11434), .ZN(n11435) );
  OAI211_X1 U13896 ( .C1(n14945), .C2(n11435), .A(n15076), .B(n11518), .ZN(
        n14944) );
  NOR2_X1 U13897 ( .A1(n14944), .A2(n15087), .ZN(n11436) );
  AOI211_X1 U13898 ( .C1(n15085), .C2(n13934), .A(n11437), .B(n11436), .ZN(
        n11438) );
  OAI211_X1 U13899 ( .C1(n11440), .C2(n14418), .A(n11439), .B(n11438), .ZN(
        P1_U3280) );
  OAI21_X1 U13900 ( .B1(n7536), .B2(n15376), .A(n11441), .ZN(n11443) );
  AOI211_X1 U13901 ( .C1(n11444), .C2(n15373), .A(n11443), .B(n11442), .ZN(
        n11447) );
  NAND2_X1 U13902 ( .A1(n15381), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n11445) );
  OAI21_X1 U13903 ( .B1(n11447), .B2(n15381), .A(n11445), .ZN(P2_U3472) );
  NAND2_X1 U13904 ( .A1(n15390), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11446) );
  OAI21_X1 U13905 ( .B1(n11447), .B2(n15390), .A(n11446), .ZN(P2_U3513) );
  NAND2_X1 U13906 ( .A1(n11449), .A2(n11448), .ZN(n11450) );
  NAND2_X1 U13907 ( .A1(n11451), .A2(n11450), .ZN(n11458) );
  NOR2_X1 U13908 ( .A1(n13680), .A2(n11452), .ZN(n11453) );
  AOI21_X1 U13909 ( .B1(n13917), .B2(n13607), .A(n11453), .ZN(n11457) );
  NAND2_X1 U13910 ( .A1(n11458), .A2(n11457), .ZN(n11483) );
  NAND2_X1 U13911 ( .A1(n13917), .A2(n13627), .ZN(n11455) );
  NAND2_X1 U13912 ( .A1(n13607), .A2(n15050), .ZN(n11454) );
  NAND2_X1 U13913 ( .A1(n11455), .A2(n11454), .ZN(n11456) );
  XNOR2_X1 U13914 ( .A(n11456), .B(n13682), .ZN(n11481) );
  NAND2_X1 U13915 ( .A1(n15201), .A2(n13627), .ZN(n11460) );
  NAND2_X1 U13916 ( .A1(n13607), .A2(n14059), .ZN(n11459) );
  NAND2_X1 U13917 ( .A1(n11460), .A2(n11459), .ZN(n11461) );
  XNOR2_X1 U13918 ( .A(n11461), .B(n13517), .ZN(n11647) );
  NOR2_X1 U13919 ( .A1(n13680), .A2(n11654), .ZN(n11462) );
  AOI21_X1 U13920 ( .B1(n15201), .B2(n13607), .A(n11462), .ZN(n11644) );
  INV_X1 U13921 ( .A(n11644), .ZN(n11648) );
  XNOR2_X1 U13922 ( .A(n11647), .B(n11648), .ZN(n11463) );
  XNOR2_X1 U13923 ( .A(n11646), .B(n11463), .ZN(n11469) );
  AOI21_X1 U13924 ( .B1(n13777), .B2(n15050), .A(n11464), .ZN(n11466) );
  NAND2_X1 U13925 ( .A1(n13776), .A2(n15060), .ZN(n11465) );
  OAI211_X1 U13926 ( .C1(n13780), .C2(n15068), .A(n11466), .B(n11465), .ZN(
        n11467) );
  AOI21_X1 U13927 ( .B1(n13782), .B2(n15201), .A(n11467), .ZN(n11468) );
  OAI21_X1 U13928 ( .B1(n11469), .B2(n13784), .A(n11468), .ZN(P1_U3217) );
  XOR2_X1 U13929 ( .A(n11470), .B(n11980), .Z(n11471) );
  AOI222_X1 U13930 ( .A1(n12636), .A2(n11471), .B1(n12632), .B2(n12633), .C1(
        n12100), .C2(n12631), .ZN(n15598) );
  NAND2_X1 U13931 ( .A1(n11472), .A2(n14898), .ZN(n15597) );
  INV_X1 U13932 ( .A(n11473), .ZN(n11614) );
  OAI22_X1 U13933 ( .A1(n12641), .A2(n15597), .B1(n11614), .B2(n12639), .ZN(
        n11474) );
  AOI21_X1 U13934 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n12648), .A(n11474), 
        .ZN(n11477) );
  NAND2_X1 U13935 ( .A1(n11475), .A2(n11980), .ZN(n15594) );
  NAND3_X1 U13936 ( .A1(n11409), .A2(n12627), .A3(n15594), .ZN(n11476) );
  OAI211_X1 U13937 ( .C1(n15598), .C2(n12648), .A(n11477), .B(n11476), .ZN(
        P3_U3223) );
  INV_X1 U13938 ( .A(n11646), .ZN(n11484) );
  INV_X1 U13939 ( .A(n11478), .ZN(n11480) );
  NAND2_X1 U13940 ( .A1(n11480), .A2(n11479), .ZN(n11482) );
  AOI22_X1 U13941 ( .A1(n11484), .A2(n11483), .B1(n11482), .B2(n11481), .ZN(
        n11490) );
  AND2_X1 U13942 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n14116) );
  AOI21_X1 U13943 ( .B1(n13777), .B2(n14060), .A(n14116), .ZN(n11486) );
  NAND2_X1 U13944 ( .A1(n13776), .A2(n14059), .ZN(n11485) );
  OAI211_X1 U13945 ( .C1(n13780), .C2(n11487), .A(n11486), .B(n11485), .ZN(
        n11488) );
  AOI21_X1 U13946 ( .B1(n13782), .B2(n13917), .A(n11488), .ZN(n11489) );
  OAI21_X1 U13947 ( .B1(n11490), .B2(n13784), .A(n11489), .ZN(P1_U3231) );
  INV_X1 U13948 ( .A(n13564), .ZN(n11493) );
  AOI21_X1 U13949 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n13397), .A(n11491), 
        .ZN(n11492) );
  OAI21_X1 U13950 ( .B1(n11493), .B2(n13399), .A(n11492), .ZN(P2_U3304) );
  INV_X1 U13951 ( .A(n11494), .ZN(n11496) );
  OAI222_X1 U13952 ( .A1(P3_U3151), .A2(n14633), .B1(n14787), .B2(n11496), 
        .C1(n11495), .C2(n12784), .ZN(P3_U3268) );
  NOR2_X1 U13953 ( .A1(n11505), .A2(n11499), .ZN(n11497) );
  XNOR2_X1 U13954 ( .A(n11576), .B(n11575), .ZN(n11500) );
  OAI22_X1 U13955 ( .A1(n12908), .A2(n13031), .B1(n11499), .B2(n12916), .ZN(
        n11552) );
  AOI21_X1 U13956 ( .B1(n11500), .B2(n13264), .A(n11552), .ZN(n13370) );
  INV_X1 U13957 ( .A(n11585), .ZN(n11501) );
  AOI211_X1 U13958 ( .C1(n13369), .C2(n11502), .A(n13270), .B(n11501), .ZN(
        n13368) );
  INV_X1 U13959 ( .A(n11554), .ZN(n11503) );
  AOI22_X1 U13960 ( .A1(n13282), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11503), 
        .B2(n13273), .ZN(n11504) );
  OAI21_X1 U13961 ( .B1(n7539), .B2(n13277), .A(n11504), .ZN(n11511) );
  NAND2_X1 U13962 ( .A1(n11505), .A2(n12980), .ZN(n11506) );
  INV_X1 U13963 ( .A(n11571), .ZN(n11508) );
  AOI21_X1 U13964 ( .B1(n11575), .B2(n11509), .A(n11508), .ZN(n13372) );
  NOR2_X1 U13965 ( .A1(n13372), .A2(n13256), .ZN(n11510) );
  AOI211_X1 U13966 ( .C1(n13368), .C2(n13272), .A(n11511), .B(n11510), .ZN(
        n11512) );
  OAI21_X1 U13967 ( .B1(n13282), .B2(n13370), .A(n11512), .ZN(P2_U3250) );
  NAND2_X1 U13968 ( .A1(n11514), .A2(n11615), .ZN(n11517) );
  AOI22_X1 U13969 ( .A1(n13523), .A2(n11515), .B1(n13524), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11516) );
  XNOR2_X1 U13970 ( .A(n13648), .B(n14056), .ZN(n13951) );
  XNOR2_X1 U13971 ( .A(n11624), .B(n13951), .ZN(n14941) );
  AOI21_X1 U13972 ( .B1(n13648), .B2(n11518), .A(n15147), .ZN(n11519) );
  NAND2_X1 U13973 ( .A1(n11519), .A2(n11634), .ZN(n14936) );
  INV_X1 U13974 ( .A(n11524), .ZN(n11523) );
  NAND2_X1 U13975 ( .A1(n11524), .A2(n13951), .ZN(n14933) );
  NAND3_X1 U13976 ( .A1(n14934), .A2(n14933), .A3(n15065), .ZN(n11541) );
  NOR2_X1 U13977 ( .A1(n14379), .A2(n11525), .ZN(n11539) );
  NAND2_X1 U13978 ( .A1(n13832), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11535) );
  INV_X1 U13979 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11526) );
  OR2_X1 U13980 ( .A1(n13842), .A2(n11526), .ZN(n11534) );
  INV_X1 U13981 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11527) );
  OR2_X1 U13982 ( .A1(n10037), .A2(n11527), .ZN(n11533) );
  OAI21_X1 U13983 ( .B1(n11530), .B2(n11528), .A(n13793), .ZN(n11531) );
  NAND2_X1 U13984 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n11529) );
  NAND2_X1 U13985 ( .A1(n11531), .A2(n11625), .ZN(n11635) );
  OR2_X1 U13986 ( .A1(n13692), .A2(n11635), .ZN(n11532) );
  OR2_X1 U13987 ( .A1(n13726), .A2(n14156), .ZN(n11537) );
  NAND2_X1 U13988 ( .A1(n14057), .A2(n15049), .ZN(n11536) );
  NAND2_X1 U13989 ( .A1(n11537), .A2(n11536), .ZN(n13649) );
  INV_X1 U13990 ( .A(n13649), .ZN(n14938) );
  OAI22_X1 U13991 ( .A1(n15105), .A2(n14938), .B1(n13653), .B2(n15080), .ZN(
        n11538) );
  AOI211_X1 U13992 ( .C1(n13648), .C2(n15085), .A(n11539), .B(n11538), .ZN(
        n11540) );
  OAI211_X1 U13993 ( .C1(n14936), .C2(n15087), .A(n11541), .B(n11540), .ZN(
        n11542) );
  AOI21_X1 U13994 ( .B1(n14941), .B2(n15064), .A(n11542), .ZN(n11543) );
  INV_X1 U13995 ( .A(n11543), .ZN(P1_U3279) );
  INV_X1 U13996 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13565) );
  NAND2_X1 U13997 ( .A1(n13564), .A2(n14559), .ZN(n11544) );
  OAI211_X1 U13998 ( .C1(n13565), .C2(n14571), .A(n11544), .B(n14055), .ZN(
        P1_U3332) );
  INV_X1 U13999 ( .A(n11545), .ZN(n11547) );
  NAND2_X1 U14000 ( .A1(n11547), .A2(n11546), .ZN(n11548) );
  XNOR2_X1 U14001 ( .A(n13369), .B(n12869), .ZN(n12786) );
  AOI22_X1 U14002 ( .A1(n11551), .A2(n12961), .B1(n12940), .B2(n12979), .ZN(
        n11558) );
  AND2_X1 U14003 ( .A1(n12979), .A2(n12824), .ZN(n11550) );
  INV_X1 U14004 ( .A(n12789), .ZN(n11557) );
  AOI22_X1 U14005 ( .A1(n12925), .A2(n11552), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11553) );
  OAI21_X1 U14006 ( .B1(n12928), .B2(n11554), .A(n11553), .ZN(n11555) );
  AOI21_X1 U14007 ( .B1(n13369), .B2(n12972), .A(n11555), .ZN(n11556) );
  OAI21_X1 U14008 ( .B1(n11558), .B2(n11557), .A(n11556), .ZN(P2_U3213) );
  INV_X1 U14009 ( .A(n11559), .ZN(n11560) );
  AOI21_X1 U14010 ( .B1(n11562), .B2(n11561), .A(n11560), .ZN(n11569) );
  NOR2_X1 U14011 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11563), .ZN(n15470) );
  OAI22_X1 U14012 ( .A1(n11564), .A2(n11848), .B1(n11875), .B2(n11979), .ZN(
        n11565) );
  AOI211_X1 U14013 ( .C1(n11845), .C2(n12099), .A(n15470), .B(n11565), .ZN(
        n11568) );
  NAND2_X1 U14014 ( .A1(n11872), .A2(n11566), .ZN(n11567) );
  OAI211_X1 U14015 ( .C1(n11569), .C2(n11852), .A(n11568), .B(n11567), .ZN(
        P3_U3171) );
  OR2_X1 U14016 ( .A1(n13369), .A2(n12979), .ZN(n11570) );
  INV_X1 U14017 ( .A(n11572), .ZN(n11580) );
  AND2_X1 U14018 ( .A1(n11573), .A2(n11580), .ZN(n11574) );
  NAND2_X1 U14019 ( .A1(n11576), .A2(n11575), .ZN(n11579) );
  INV_X1 U14020 ( .A(n12979), .ZN(n11577) );
  NAND2_X1 U14021 ( .A1(n13369), .A2(n11577), .ZN(n11578) );
  XNOR2_X1 U14022 ( .A(n11591), .B(n11580), .ZN(n11583) );
  NAND2_X1 U14023 ( .A1(n13065), .A2(n12963), .ZN(n11582) );
  NAND2_X1 U14024 ( .A1(n12979), .A2(n13095), .ZN(n11581) );
  NAND2_X1 U14025 ( .A1(n11582), .A2(n11581), .ZN(n12895) );
  AOI21_X1 U14026 ( .B1(n11583), .B2(n13264), .A(n12895), .ZN(n13365) );
  OAI21_X1 U14027 ( .B1(n12898), .B2(n13236), .A(n13365), .ZN(n11584) );
  NAND2_X1 U14028 ( .A1(n11584), .A2(n13252), .ZN(n11589) );
  AOI211_X1 U14029 ( .C1(n13364), .C2(n11585), .A(n13270), .B(n11597), .ZN(
        n13363) );
  OAI22_X1 U14030 ( .A1(n7738), .A2(n13277), .B1(n11586), .B2(n13252), .ZN(
        n11587) );
  AOI21_X1 U14031 ( .B1(n13363), .B2(n13272), .A(n11587), .ZN(n11588) );
  OAI211_X1 U14032 ( .C1(n13367), .C2(n13256), .A(n11589), .B(n11588), .ZN(
        P2_U3249) );
  AND2_X1 U14033 ( .A1(n13364), .A2(n12908), .ZN(n11590) );
  XNOR2_X1 U14034 ( .A(n13067), .B(n11595), .ZN(n11593) );
  AND2_X1 U14035 ( .A1(n12978), .A2(n13095), .ZN(n11592) );
  AOI21_X1 U14036 ( .B1(n13042), .B2(n12963), .A(n11592), .ZN(n12903) );
  OAI21_X1 U14037 ( .B1(n11593), .B2(n13247), .A(n12903), .ZN(n13360) );
  INV_X1 U14038 ( .A(n13360), .ZN(n11603) );
  AOI21_X1 U14039 ( .B1(n11596), .B2(n11595), .A(n6631), .ZN(n13361) );
  INV_X1 U14040 ( .A(n13069), .ZN(n13358) );
  NAND2_X1 U14041 ( .A1(n11597), .A2(n13358), .ZN(n13271) );
  OAI211_X1 U14042 ( .C1(n11597), .C2(n13358), .A(n13294), .B(n13271), .ZN(
        n13357) );
  INV_X1 U14043 ( .A(n12906), .ZN(n11598) );
  OAI22_X1 U14044 ( .A1(n13252), .A2(n11333), .B1(n11598), .B2(n13236), .ZN(
        n11599) );
  AOI21_X1 U14045 ( .B1(n13069), .B2(n13240), .A(n11599), .ZN(n11600) );
  OAI21_X1 U14046 ( .B1(n13357), .B2(n13206), .A(n11600), .ZN(n11601) );
  AOI21_X1 U14047 ( .B1(n13361), .B2(n13280), .A(n11601), .ZN(n11602) );
  OAI21_X1 U14048 ( .B1(n13282), .B2(n11603), .A(n11602), .ZN(P2_U3248) );
  AOI21_X1 U14049 ( .B1(n11605), .B2(n11604), .A(n11852), .ZN(n11607) );
  NAND2_X1 U14050 ( .A1(n11607), .A2(n11606), .ZN(n11612) );
  AND2_X1 U14051 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n15483) );
  OAI22_X1 U14052 ( .A1(n11609), .A2(n11848), .B1(n11875), .B2(n11608), .ZN(
        n11610) );
  AOI211_X1 U14053 ( .C1(n11845), .C2(n12632), .A(n15483), .B(n11610), .ZN(
        n11611) );
  OAI211_X1 U14054 ( .C1(n11614), .C2(n11613), .A(n11612), .B(n11611), .ZN(
        P3_U3157) );
  NAND2_X1 U14055 ( .A1(n11616), .A2(n11615), .ZN(n11619) );
  AOI22_X1 U14056 ( .A1(n13524), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n13523), 
        .B2(n11617), .ZN(n11618) );
  NAND2_X1 U14057 ( .A1(n14534), .A2(n13726), .ZN(n13944) );
  NAND2_X1 U14058 ( .A1(n14166), .A2(n13944), .ZN(n13823) );
  NAND2_X1 U14059 ( .A1(n13648), .A2(n14056), .ZN(n11620) );
  INV_X1 U14060 ( .A(n14184), .ZN(n11621) );
  AOI21_X1 U14061 ( .B1(n14168), .B2(n11622), .A(n11621), .ZN(n14536) );
  OR2_X1 U14062 ( .A1(n13648), .A2(n13485), .ZN(n13933) );
  NAND2_X1 U14063 ( .A1(n13648), .A2(n13485), .ZN(n13942) );
  INV_X1 U14064 ( .A(n13942), .ZN(n11623) );
  XNOR2_X1 U14065 ( .A(n14169), .B(n14168), .ZN(n11633) );
  OR2_X1 U14066 ( .A1(n13485), .A2(n14432), .ZN(n11632) );
  AND2_X1 U14067 ( .A1(n11625), .A2(n12184), .ZN(n11626) );
  NOR2_X1 U14068 ( .A1(n13511), .A2(n11626), .ZN(n14410) );
  NAND2_X1 U14069 ( .A1(n14410), .A2(n13553), .ZN(n11630) );
  OR2_X1 U14070 ( .A1(n13842), .A2(n11170), .ZN(n11629) );
  NAND2_X1 U14071 ( .A1(n13688), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11628) );
  NAND2_X1 U14072 ( .A1(n13832), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11627) );
  NAND4_X1 U14073 ( .A1(n11630), .A2(n11629), .A3(n11628), .A4(n11627), .ZN(
        n14389) );
  NAND2_X1 U14074 ( .A1(n14389), .A2(n15059), .ZN(n11631) );
  AND2_X1 U14075 ( .A1(n11632), .A2(n11631), .ZN(n13794) );
  OAI21_X1 U14076 ( .B1(n11633), .B2(n15178), .A(n13794), .ZN(n14532) );
  NAND2_X1 U14077 ( .A1(n14532), .A2(n14379), .ZN(n11639) );
  AOI211_X1 U14078 ( .C1(n14534), .C2(n11634), .A(n15147), .B(n7597), .ZN(
        n14533) );
  INV_X1 U14079 ( .A(n14534), .ZN(n13802) );
  INV_X1 U14080 ( .A(n11635), .ZN(n13797) );
  AOI22_X1 U14081 ( .A1(n15093), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13797), 
        .B2(n15091), .ZN(n11636) );
  OAI21_X1 U14082 ( .B1(n13802), .B2(n15096), .A(n11636), .ZN(n11637) );
  AOI21_X1 U14083 ( .B1(n14533), .B2(n15063), .A(n11637), .ZN(n11638) );
  OAI211_X1 U14084 ( .C1(n14536), .C2(n14418), .A(n11639), .B(n11638), .ZN(
        P1_U3278) );
  NAND2_X1 U14085 ( .A1(n13924), .A2(n13627), .ZN(n11641) );
  NAND2_X1 U14086 ( .A1(n13607), .A2(n15060), .ZN(n11640) );
  NAND2_X1 U14087 ( .A1(n11641), .A2(n11640), .ZN(n11642) );
  XNOR2_X1 U14088 ( .A(n11642), .B(n13517), .ZN(n11663) );
  NOR2_X1 U14089 ( .A1(n13680), .A2(n13925), .ZN(n11643) );
  AOI21_X1 U14090 ( .B1(n13924), .B2(n13607), .A(n11643), .ZN(n11662) );
  XNOR2_X1 U14091 ( .A(n11663), .B(n11662), .ZN(n11653) );
  NAND2_X1 U14092 ( .A1(n11647), .A2(n11644), .ZN(n11645) );
  INV_X1 U14093 ( .A(n11647), .ZN(n11649) );
  NAND2_X1 U14094 ( .A1(n11649), .A2(n11648), .ZN(n11650) );
  INV_X1 U14095 ( .A(n11669), .ZN(n11651) );
  AOI21_X1 U14096 ( .B1(n11653), .B2(n11652), .A(n11651), .ZN(n11661) );
  INV_X1 U14097 ( .A(n13777), .ZN(n13735) );
  NOR2_X1 U14098 ( .A1(n13735), .A2(n11654), .ZN(n11655) );
  AOI211_X1 U14099 ( .C1(n13776), .C2(n14058), .A(n11656), .B(n11655), .ZN(
        n11657) );
  OAI21_X1 U14100 ( .B1(n13780), .B2(n11658), .A(n11657), .ZN(n11659) );
  AOI21_X1 U14101 ( .B1(n13782), .B2(n13924), .A(n11659), .ZN(n11660) );
  OAI21_X1 U14102 ( .B1(n11661), .B2(n13784), .A(n11660), .ZN(P1_U3236) );
  NAND2_X1 U14103 ( .A1(n11663), .A2(n11662), .ZN(n11667) );
  AND2_X1 U14104 ( .A1(n11669), .A2(n11667), .ZN(n11671) );
  OAI22_X1 U14105 ( .A1(n14797), .A2(n10072), .B1(n13929), .B2(n13681), .ZN(
        n11664) );
  XNOR2_X1 U14106 ( .A(n11664), .B(n13517), .ZN(n11678) );
  OR2_X1 U14107 ( .A1(n14797), .A2(n13681), .ZN(n11666) );
  NAND2_X1 U14108 ( .A1(n13626), .A2(n14058), .ZN(n11665) );
  NAND2_X1 U14109 ( .A1(n11666), .A2(n11665), .ZN(n11679) );
  XNOR2_X1 U14110 ( .A(n11678), .B(n11679), .ZN(n11670) );
  AND2_X1 U14111 ( .A1(n11670), .A2(n11667), .ZN(n11668) );
  NAND2_X1 U14112 ( .A1(n11669), .A2(n11668), .ZN(n11682) );
  OAI211_X1 U14113 ( .C1(n11671), .C2(n11670), .A(n13790), .B(n11682), .ZN(
        n11677) );
  NAND2_X1 U14114 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n15015)
         );
  INV_X1 U14115 ( .A(n15015), .ZN(n11674) );
  NOR2_X1 U14116 ( .A1(n13780), .A2(n11672), .ZN(n11673) );
  AOI211_X1 U14117 ( .C1(n13650), .C2(n11675), .A(n11674), .B(n11673), .ZN(
        n11676) );
  OAI211_X1 U14118 ( .C1(n14797), .C2(n13801), .A(n11677), .B(n11676), .ZN(
        P1_U3224) );
  INV_X1 U14119 ( .A(n11678), .ZN(n11680) );
  NAND2_X1 U14120 ( .A1(n11680), .A2(n11679), .ZN(n11681) );
  NAND2_X1 U14121 ( .A1(n13934), .A2(n13627), .ZN(n11684) );
  NAND2_X1 U14122 ( .A1(n13607), .A2(n14057), .ZN(n11683) );
  NAND2_X1 U14123 ( .A1(n11684), .A2(n11683), .ZN(n11685) );
  XNOR2_X1 U14124 ( .A(n11685), .B(n13682), .ZN(n13476) );
  INV_X1 U14125 ( .A(n14057), .ZN(n13935) );
  NOR2_X1 U14126 ( .A1(n13680), .A2(n13935), .ZN(n11686) );
  AOI21_X1 U14127 ( .B1(n13934), .B2(n13607), .A(n11686), .ZN(n13477) );
  XNOR2_X1 U14128 ( .A(n13476), .B(n13477), .ZN(n13480) );
  XNOR2_X1 U14129 ( .A(n13481), .B(n13480), .ZN(n11692) );
  NAND2_X1 U14130 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n15020)
         );
  OAI21_X1 U14131 ( .B1(n13735), .B2(n13929), .A(n15020), .ZN(n11687) );
  AOI21_X1 U14132 ( .B1(n13776), .B2(n14056), .A(n11687), .ZN(n11688) );
  OAI21_X1 U14133 ( .B1(n13780), .B2(n11689), .A(n11688), .ZN(n11690) );
  AOI21_X1 U14134 ( .B1(n13934), .B2(n13782), .A(n11690), .ZN(n11691) );
  OAI21_X1 U14135 ( .B1(n11692), .B2(n13784), .A(n11691), .ZN(P1_U3234) );
  INV_X1 U14136 ( .A(n13676), .ZN(n11693) );
  OAI222_X1 U14137 ( .A1(n11694), .A2(P1_U3086), .B1(n11699), .B2(n11693), 
        .C1(n13677), .C2(n14571), .ZN(P1_U3327) );
  INV_X1 U14138 ( .A(n11695), .ZN(n11696) );
  OAI222_X1 U14139 ( .A1(n12784), .A2(n11697), .B1(P3_U3151), .B2(n9254), .C1(
        n14787), .C2(n11696), .ZN(P3_U3267) );
  INV_X1 U14140 ( .A(n13848), .ZN(n13403) );
  OAI222_X1 U14141 ( .A1(P1_U3086), .A2(n11698), .B1(n11699), .B2(n13403), 
        .C1(n13849), .C2(n14571), .ZN(P1_U3326) );
  INV_X1 U14142 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13838) );
  OAI222_X1 U14143 ( .A1(P1_U3086), .A2(n9990), .B1(n11699), .B2(n13837), .C1(
        n13838), .C2(n14571), .ZN(P1_U3325) );
  INV_X1 U14144 ( .A(n11700), .ZN(n11701) );
  OAI222_X1 U14145 ( .A1(n8726), .A2(P3_U3151), .B1(n14787), .B2(n11701), .C1(
        n7624), .C2(n12784), .ZN(P3_U3271) );
  XNOR2_X1 U14146 ( .A(n12417), .B(n8803), .ZN(n11708) );
  INV_X1 U14147 ( .A(n11708), .ZN(n11702) );
  NAND2_X1 U14148 ( .A1(n11702), .A2(n11863), .ZN(n11714) );
  INV_X1 U14149 ( .A(n11703), .ZN(n11704) );
  NAND4_X1 U14150 ( .A1(n11713), .A2(n11863), .A3(n11704), .A4(n11708), .ZN(
        n11712) );
  AOI22_X1 U14151 ( .A1(n12094), .A2(n11868), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11706) );
  NAND2_X1 U14152 ( .A1(n12419), .A2(n11872), .ZN(n11705) );
  OAI211_X1 U14153 ( .C1(n12413), .C2(n11870), .A(n11706), .B(n11705), .ZN(
        n11710) );
  NOR4_X1 U14154 ( .A1(n11708), .A2(n11707), .A3(n11852), .A4(n12094), .ZN(
        n11709) );
  AOI211_X1 U14155 ( .C1(n12652), .C2(n11850), .A(n11710), .B(n11709), .ZN(
        n11711) );
  OAI211_X1 U14156 ( .C1(n11714), .C2(n11713), .A(n11712), .B(n11711), .ZN(
        P3_U3160) );
  INV_X1 U14157 ( .A(n11716), .ZN(n11720) );
  AOI22_X1 U14158 ( .A1(n12408), .A2(n12624), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n12648), .ZN(n11717) );
  OAI21_X1 U14159 ( .B1(n11718), .B2(n12595), .A(n11717), .ZN(n11719) );
  AOI21_X1 U14160 ( .B1(n11720), .B2(n12627), .A(n11719), .ZN(n11721) );
  OAI21_X1 U14161 ( .B1(n11715), .B2(n12648), .A(n11721), .ZN(P3_U3204) );
  NAND2_X1 U14162 ( .A1(n13849), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11724) );
  NAND2_X1 U14163 ( .A1(n11725), .A2(n11724), .ZN(n11884) );
  NAND2_X1 U14164 ( .A1(n11726), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11882) );
  NAND2_X1 U14165 ( .A1(n13838), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11727) );
  NAND2_X1 U14166 ( .A1(n11882), .A2(n11727), .ZN(n11883) );
  XNOR2_X1 U14167 ( .A(n11884), .B(n11883), .ZN(n11878) );
  INV_X1 U14168 ( .A(n11878), .ZN(n11728) );
  INV_X1 U14169 ( .A(SI_30_), .ZN(n11879) );
  OAI222_X1 U14170 ( .A1(P3_U3151), .A2(n8766), .B1(n14787), .B2(n11728), .C1(
        n11879), .C2(n12784), .ZN(P3_U3265) );
  XNOR2_X1 U14171 ( .A(n11729), .B(n12617), .ZN(n11730) );
  XNOR2_X1 U14172 ( .A(n11731), .B(n11730), .ZN(n11737) );
  NOR2_X1 U14173 ( .A1(n12769), .A2(n11875), .ZN(n11735) );
  INV_X1 U14174 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12358) );
  NOR2_X1 U14175 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12358), .ZN(n15556) );
  AOI21_X1 U14176 ( .B1(n11868), .B2(n12634), .A(n15556), .ZN(n11732) );
  OAI21_X1 U14177 ( .B1(n11733), .B2(n11870), .A(n11732), .ZN(n11734) );
  AOI211_X1 U14178 ( .C1(n12606), .C2(n11872), .A(n11735), .B(n11734), .ZN(
        n11736) );
  OAI21_X1 U14179 ( .B1(n11737), .B2(n11852), .A(n11736), .ZN(P3_U3155) );
  AOI21_X1 U14180 ( .B1(n9346), .B2(n11738), .A(n6641), .ZN(n11744) );
  AOI22_X1 U14181 ( .A1(n11868), .A2(n12507), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11740) );
  NAND2_X1 U14182 ( .A1(n11872), .A2(n12488), .ZN(n11739) );
  OAI211_X1 U14183 ( .C1(n12487), .C2(n11870), .A(n11740), .B(n11739), .ZN(
        n11741) );
  AOI21_X1 U14184 ( .B1(n11742), .B2(n11850), .A(n11741), .ZN(n11743) );
  OAI21_X1 U14185 ( .B1(n11744), .B2(n11852), .A(n11743), .ZN(P3_U3156) );
  XOR2_X1 U14186 ( .A(n11746), .B(n11745), .Z(n11747) );
  NAND2_X1 U14187 ( .A1(n11747), .A2(n11863), .ZN(n11751) );
  NAND2_X1 U14188 ( .A1(n11868), .A2(n12558), .ZN(n11748) );
  NAND2_X1 U14189 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n14598)
         );
  OAI211_X1 U14190 ( .C1(n11870), .C2(n12509), .A(n11748), .B(n14598), .ZN(
        n11749) );
  AOI21_X1 U14191 ( .B1(n12537), .B2(n11872), .A(n11749), .ZN(n11750) );
  OAI211_X1 U14192 ( .C1(n11875), .C2(n12755), .A(n11751), .B(n11750), .ZN(
        P3_U3159) );
  XNOR2_X1 U14193 ( .A(n11753), .B(n11752), .ZN(n11759) );
  NAND2_X1 U14194 ( .A1(n11872), .A2(n12512), .ZN(n11755) );
  AOI22_X1 U14195 ( .A1(n11868), .A2(n12534), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11754) );
  OAI211_X1 U14196 ( .C1(n11756), .C2(n11870), .A(n11755), .B(n11754), .ZN(
        n11757) );
  AOI21_X1 U14197 ( .B1(n12516), .B2(n11850), .A(n11757), .ZN(n11758) );
  OAI21_X1 U14198 ( .B1(n11759), .B2(n11852), .A(n11758), .ZN(P3_U3163) );
  XNOR2_X1 U14199 ( .A(n11760), .B(n11761), .ZN(n11833) );
  OAI22_X1 U14200 ( .A1(n11833), .A2(n12632), .B1(n11760), .B2(n11761), .ZN(
        n11764) );
  XNOR2_X1 U14201 ( .A(n11762), .B(n12616), .ZN(n11763) );
  XNOR2_X1 U14202 ( .A(n11764), .B(n11763), .ZN(n11769) );
  AND2_X1 U14203 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n15517) );
  OAI22_X1 U14204 ( .A1(n11832), .A2(n11848), .B1(n11875), .B2(n11765), .ZN(
        n11766) );
  AOI211_X1 U14205 ( .C1(n11845), .C2(n12634), .A(n15517), .B(n11766), .ZN(
        n11768) );
  NAND2_X1 U14206 ( .A1(n11872), .A2(n12638), .ZN(n11767) );
  OAI211_X1 U14207 ( .C1(n11769), .C2(n11852), .A(n11768), .B(n11767), .ZN(
        P3_U3164) );
  INV_X1 U14208 ( .A(n11770), .ZN(n11801) );
  INV_X1 U14209 ( .A(n11771), .ZN(n11773) );
  NOR3_X1 U14210 ( .A1(n11801), .A2(n11773), .A3(n11772), .ZN(n11776) );
  INV_X1 U14211 ( .A(n11774), .ZN(n11775) );
  NOR2_X1 U14212 ( .A1(n12487), .A2(n11848), .ZN(n11779) );
  OAI22_X1 U14213 ( .A1(n12456), .A2(n11870), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11777), .ZN(n11778) );
  AOI211_X1 U14214 ( .C1(n12461), .C2(n11872), .A(n11779), .B(n11778), .ZN(
        n11780) );
  OAI211_X1 U14215 ( .C1(n12731), .C2(n11875), .A(n11781), .B(n11780), .ZN(
        P3_U3165) );
  XNOR2_X1 U14216 ( .A(n11782), .B(n12588), .ZN(n11783) );
  XNOR2_X1 U14217 ( .A(n11784), .B(n11783), .ZN(n11789) );
  NAND2_X1 U14218 ( .A1(n11872), .A2(n12577), .ZN(n11786) );
  NOR2_X1 U14219 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9033), .ZN(n14843) );
  AOI21_X1 U14220 ( .B1(n11868), .B2(n12603), .A(n14843), .ZN(n11785) );
  OAI211_X1 U14221 ( .C1(n12548), .C2(n11870), .A(n11786), .B(n11785), .ZN(
        n11787) );
  AOI21_X1 U14222 ( .B1(n12701), .B2(n11850), .A(n11787), .ZN(n11788) );
  OAI21_X1 U14223 ( .B1(n11789), .B2(n11852), .A(n11788), .ZN(P3_U3166) );
  XNOR2_X1 U14224 ( .A(n11790), .B(n12570), .ZN(n11791) );
  XNOR2_X1 U14225 ( .A(n11792), .B(n11791), .ZN(n11797) );
  NAND2_X1 U14226 ( .A1(n11872), .A2(n12563), .ZN(n11794) );
  NOR2_X1 U14227 ( .A1(n12256), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14872) );
  AOI21_X1 U14228 ( .B1(n11845), .B2(n12558), .A(n14872), .ZN(n11793) );
  OAI211_X1 U14229 ( .C1(n12588), .C2(n11848), .A(n11794), .B(n11793), .ZN(
        n11795) );
  AOI21_X1 U14230 ( .B1(n12697), .B2(n11850), .A(n11795), .ZN(n11796) );
  OAI21_X1 U14231 ( .B1(n11797), .B2(n11852), .A(n11796), .ZN(P3_U3168) );
  INV_X1 U14232 ( .A(n11798), .ZN(n11800) );
  NOR3_X1 U14233 ( .A1(n6641), .A2(n11800), .A3(n11799), .ZN(n11802) );
  OAI21_X1 U14234 ( .B1(n11802), .B2(n11801), .A(n11863), .ZN(n11806) );
  AOI22_X1 U14235 ( .A1(n12096), .A2(n11845), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11803) );
  OAI21_X1 U14236 ( .B1(n12495), .B2(n11848), .A(n11803), .ZN(n11804) );
  AOI21_X1 U14237 ( .B1(n12474), .B2(n11872), .A(n11804), .ZN(n11805) );
  OAI211_X1 U14238 ( .C1(n12735), .C2(n11875), .A(n11806), .B(n11805), .ZN(
        P3_U3169) );
  XNOR2_X1 U14239 ( .A(n11808), .B(n11807), .ZN(n11814) );
  OAI22_X1 U14240 ( .A1(n11870), .A2(n12522), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11809), .ZN(n11811) );
  NOR2_X1 U14241 ( .A1(n11848), .A2(n12549), .ZN(n11810) );
  AOI211_X1 U14242 ( .C1(n12525), .C2(n11872), .A(n11811), .B(n11810), .ZN(
        n11813) );
  NAND2_X1 U14243 ( .A1(n12524), .A2(n11850), .ZN(n11812) );
  OAI211_X1 U14244 ( .C1(n11814), .C2(n11852), .A(n11813), .B(n11812), .ZN(
        P3_U3173) );
  XNOR2_X1 U14245 ( .A(n11815), .B(n12634), .ZN(n11816) );
  XNOR2_X1 U14246 ( .A(n11817), .B(n11816), .ZN(n11824) );
  NOR2_X1 U14247 ( .A1(n11875), .A2(n12622), .ZN(n11822) );
  NOR2_X1 U14248 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11818), .ZN(n15534) );
  AOI21_X1 U14249 ( .B1(n11845), .B2(n12617), .A(n15534), .ZN(n11819) );
  OAI21_X1 U14250 ( .B1(n11820), .B2(n11848), .A(n11819), .ZN(n11821) );
  AOI211_X1 U14251 ( .C1(n12623), .C2(n11872), .A(n11822), .B(n11821), .ZN(
        n11823) );
  OAI21_X1 U14252 ( .B1(n11824), .B2(n11852), .A(n11823), .ZN(P3_U3174) );
  AOI21_X1 U14253 ( .B1(n12507), .B2(n11825), .A(n6737), .ZN(n11831) );
  NAND2_X1 U14254 ( .A1(n11872), .A2(n12498), .ZN(n11827) );
  INV_X1 U14255 ( .A(n12522), .ZN(n12097) );
  AOI22_X1 U14256 ( .A1(n12097), .A2(n11868), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11826) );
  OAI211_X1 U14257 ( .C1(n12495), .C2(n11870), .A(n11827), .B(n11826), .ZN(
        n11828) );
  AOI21_X1 U14258 ( .B1(n11829), .B2(n11850), .A(n11828), .ZN(n11830) );
  OAI21_X1 U14259 ( .B1(n11831), .B2(n11852), .A(n11830), .ZN(P3_U3175) );
  XNOR2_X1 U14260 ( .A(n11833), .B(n11832), .ZN(n11841) );
  INV_X1 U14261 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11834) );
  NOR2_X1 U14262 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11834), .ZN(n15499) );
  OAI22_X1 U14263 ( .A1(n11836), .A2(n11848), .B1(n11875), .B2(n11835), .ZN(
        n11837) );
  AOI211_X1 U14264 ( .C1(n11845), .C2(n12616), .A(n15499), .B(n11837), .ZN(
        n11840) );
  NAND2_X1 U14265 ( .A1(n11872), .A2(n11838), .ZN(n11839) );
  OAI211_X1 U14266 ( .C1(n11841), .C2(n11852), .A(n11840), .B(n11839), .ZN(
        P3_U3176) );
  XNOR2_X1 U14267 ( .A(n11842), .B(n12558), .ZN(n11843) );
  XNOR2_X1 U14268 ( .A(n11844), .B(n11843), .ZN(n11853) );
  NAND2_X1 U14269 ( .A1(n11872), .A2(n12551), .ZN(n11847) );
  AND2_X1 U14270 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14879) );
  AOI21_X1 U14271 ( .B1(n11845), .B2(n12098), .A(n14879), .ZN(n11846) );
  OAI211_X1 U14272 ( .C1(n12548), .C2(n11848), .A(n11847), .B(n11846), .ZN(
        n11849) );
  AOI21_X1 U14273 ( .B1(n12550), .B2(n11850), .A(n11849), .ZN(n11851) );
  OAI21_X1 U14274 ( .B1(n11853), .B2(n11852), .A(n11851), .ZN(P3_U3178) );
  OAI21_X1 U14275 ( .B1(n11856), .B2(n11855), .A(n11854), .ZN(n11857) );
  AOI22_X1 U14276 ( .A1(n12096), .A2(n11868), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11859) );
  OAI21_X1 U14277 ( .B1(n12443), .B2(n11870), .A(n11859), .ZN(n11860) );
  AOI21_X1 U14278 ( .B1(n12446), .B2(n11872), .A(n11860), .ZN(n11861) );
  INV_X1 U14279 ( .A(n11862), .ZN(n12765) );
  OAI211_X1 U14280 ( .C1(n11866), .C2(n11865), .A(n11864), .B(n11863), .ZN(
        n11874) );
  INV_X1 U14281 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n11867) );
  NOR2_X1 U14282 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11867), .ZN(n14825) );
  AOI21_X1 U14283 ( .B1(n11868), .B2(n12617), .A(n14825), .ZN(n11869) );
  OAI21_X1 U14284 ( .B1(n12588), .B2(n11870), .A(n11869), .ZN(n11871) );
  AOI21_X1 U14285 ( .B1(n12593), .B2(n11872), .A(n11871), .ZN(n11873) );
  OAI211_X1 U14286 ( .C1(n12765), .C2(n11875), .A(n11874), .B(n11873), .ZN(
        P3_U3181) );
  INV_X1 U14287 ( .A(n11876), .ZN(n12067) );
  NAND2_X1 U14288 ( .A1(n11877), .A2(n12067), .ZN(n11897) );
  NAND2_X1 U14289 ( .A1(n11878), .A2(n11887), .ZN(n11881) );
  OR2_X1 U14290 ( .A1(n6570), .A2(n11879), .ZN(n11880) );
  NAND2_X1 U14291 ( .A1(n11881), .A2(n11880), .ZN(n14899) );
  XNOR2_X1 U14292 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n11885) );
  XNOR2_X1 U14293 ( .A(n11886), .B(n11885), .ZN(n12778) );
  NAND2_X1 U14294 ( .A1(n12778), .A2(n11887), .ZN(n11889) );
  INV_X1 U14295 ( .A(SI_31_), .ZN(n12775) );
  OR2_X1 U14296 ( .A1(n6569), .A2(n12775), .ZN(n11888) );
  NAND2_X1 U14297 ( .A1(n11889), .A2(n11888), .ZN(n11902) );
  NAND2_X1 U14298 ( .A1(n8790), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11892) );
  NAND2_X1 U14299 ( .A1(n9354), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11891) );
  NAND2_X1 U14300 ( .A1(n8788), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11890) );
  AND3_X1 U14301 ( .A1(n11892), .A2(n11891), .A3(n11890), .ZN(n11893) );
  INV_X1 U14302 ( .A(n14899), .ZN(n11899) );
  INV_X1 U14303 ( .A(n12407), .ZN(n12090) );
  NAND2_X1 U14304 ( .A1(n14899), .A2(n12407), .ZN(n11896) );
  NAND3_X1 U14305 ( .A1(n11897), .A2(n12072), .A3(n11896), .ZN(n11903) );
  NAND2_X1 U14306 ( .A1(n11902), .A2(n12407), .ZN(n11901) );
  INV_X1 U14307 ( .A(n11898), .ZN(n12091) );
  NAND2_X1 U14308 ( .A1(n11899), .A2(n12091), .ZN(n11900) );
  INV_X1 U14309 ( .A(n11902), .ZN(n12719) );
  NAND2_X1 U14310 ( .A1(n11903), .A2(n7885), .ZN(n11904) );
  XNOR2_X1 U14311 ( .A(n11904), .B(n11927), .ZN(n12082) );
  INV_X1 U14312 ( .A(n11905), .ZN(n12081) );
  INV_X1 U14313 ( .A(n11906), .ZN(n12071) );
  INV_X1 U14314 ( .A(n12058), .ZN(n12066) );
  INV_X1 U14315 ( .A(n11908), .ZN(n12038) );
  AND4_X1 U14316 ( .A1(n11910), .A2(n9309), .A3(n7430), .A4(n11909), .ZN(
        n11915) );
  NOR2_X1 U14317 ( .A1(n9305), .A2(n11911), .ZN(n11914) );
  NOR2_X1 U14318 ( .A1(n11980), .A2(n11912), .ZN(n11913) );
  NAND4_X1 U14319 ( .A1(n11915), .A2(n11930), .A3(n11914), .A4(n11913), .ZN(
        n11919) );
  NAND3_X1 U14320 ( .A1(n12630), .A2(n11975), .A3(n11969), .ZN(n11918) );
  OR2_X1 U14321 ( .A1(n7440), .A2(n11998), .ZN(n11997) );
  NOR4_X1 U14322 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11997), .ZN(
        n11920) );
  NAND4_X1 U14323 ( .A1(n12573), .A2(n11920), .A3(n12600), .A4(n12591), .ZN(
        n11921) );
  NOR3_X1 U14324 ( .A1(n9340), .A2(n12013), .A3(n11921), .ZN(n11922) );
  NAND4_X1 U14325 ( .A1(n9344), .A2(n7860), .A3(n12531), .A4(n11922), .ZN(
        n11923) );
  NOR4_X1 U14326 ( .A1(n12469), .A2(n12483), .A3(n12496), .A4(n11923), .ZN(
        n11925) );
  XNOR2_X1 U14327 ( .A(n12727), .B(n12095), .ZN(n12444) );
  INV_X1 U14328 ( .A(n12444), .ZN(n11924) );
  NAND4_X1 U14329 ( .A1(n12067), .A2(n7080), .A3(n11925), .A4(n11924), .ZN(
        n11926) );
  XNOR2_X1 U14330 ( .A(n11928), .B(n11927), .ZN(n12078) );
  NAND3_X1 U14331 ( .A1(n11930), .A2(n12086), .A3(n11929), .ZN(n11934) );
  OAI211_X1 U14332 ( .C1(n11931), .C2(n11932), .A(n12044), .B(n11936), .ZN(
        n11933) );
  AOI22_X1 U14333 ( .A1(n11934), .A2(n11933), .B1(n10315), .B2(n11932), .ZN(
        n11940) );
  INV_X1 U14334 ( .A(n11935), .ZN(n11938) );
  INV_X1 U14335 ( .A(n11936), .ZN(n11937) );
  MUX2_X1 U14336 ( .A(n11938), .B(n11937), .S(n12070), .Z(n11939) );
  NOR3_X1 U14337 ( .A1(n11940), .A2(n11939), .A3(n9305), .ZN(n11950) );
  NAND2_X1 U14338 ( .A1(n11946), .A2(n11941), .ZN(n11944) );
  NAND2_X1 U14339 ( .A1(n11945), .A2(n11942), .ZN(n11943) );
  MUX2_X1 U14340 ( .A(n11944), .B(n11943), .S(n12044), .Z(n11949) );
  MUX2_X1 U14341 ( .A(n11946), .B(n11945), .S(n12070), .Z(n11947) );
  OAI211_X1 U14342 ( .C1(n11950), .C2(n11949), .A(n11948), .B(n11947), .ZN(
        n11954) );
  MUX2_X1 U14343 ( .A(n11952), .B(n11951), .S(n12044), .Z(n11953) );
  AND3_X1 U14344 ( .A1(n11954), .A2(n7430), .A3(n11953), .ZN(n11964) );
  NAND2_X1 U14345 ( .A1(n11960), .A2(n11955), .ZN(n11958) );
  NAND2_X1 U14346 ( .A1(n11959), .A2(n11956), .ZN(n11957) );
  MUX2_X1 U14347 ( .A(n11958), .B(n11957), .S(n12070), .Z(n11963) );
  MUX2_X1 U14348 ( .A(n11960), .B(n11959), .S(n12044), .Z(n11961) );
  OAI211_X1 U14349 ( .C1(n11964), .C2(n11963), .A(n11962), .B(n11961), .ZN(
        n11970) );
  NAND2_X1 U14350 ( .A1(n12102), .A2(n11965), .ZN(n11967) );
  MUX2_X1 U14351 ( .A(n11967), .B(n11966), .S(n12070), .Z(n11968) );
  NAND3_X1 U14352 ( .A1(n11970), .A2(n11969), .A3(n11968), .ZN(n11976) );
  NAND2_X1 U14353 ( .A1(n12101), .A2(n11971), .ZN(n11972) );
  MUX2_X1 U14354 ( .A(n11973), .B(n11972), .S(n12070), .Z(n11974) );
  NAND3_X1 U14355 ( .A1(n11976), .A2(n11975), .A3(n11974), .ZN(n11982) );
  MUX2_X1 U14356 ( .A(n11977), .B(n12044), .S(n12100), .Z(n11978) );
  OAI21_X1 U14357 ( .B1(n12070), .B2(n11979), .A(n11978), .ZN(n11981) );
  AOI21_X1 U14358 ( .B1(n11982), .B2(n11981), .A(n11980), .ZN(n11992) );
  INV_X1 U14359 ( .A(n11983), .ZN(n11985) );
  OAI211_X1 U14360 ( .C1(n11992), .C2(n11985), .A(n11993), .B(n11984), .ZN(
        n11986) );
  NAND2_X1 U14361 ( .A1(n11986), .A2(n11989), .ZN(n11996) );
  NAND2_X1 U14362 ( .A1(n11988), .A2(n11987), .ZN(n11991) );
  OAI211_X1 U14363 ( .C1(n11992), .C2(n11991), .A(n11990), .B(n11989), .ZN(
        n11994) );
  NAND2_X1 U14364 ( .A1(n11994), .A2(n11993), .ZN(n11995) );
  MUX2_X1 U14365 ( .A(n11996), .B(n11995), .S(n12070), .Z(n12000) );
  INV_X1 U14366 ( .A(n11997), .ZN(n12620) );
  MUX2_X1 U14367 ( .A(n7440), .B(n11998), .S(n12070), .Z(n11999) );
  AOI211_X1 U14368 ( .C1(n12000), .C2(n12620), .A(n11999), .B(n12611), .ZN(
        n12010) );
  MUX2_X1 U14369 ( .A(n12002), .B(n12001), .S(n12044), .Z(n12003) );
  NAND2_X1 U14370 ( .A1(n12591), .A2(n12003), .ZN(n12009) );
  AND2_X1 U14371 ( .A1(n12012), .A2(n12004), .ZN(n12007) );
  AND2_X1 U14372 ( .A1(n12011), .A2(n12005), .ZN(n12006) );
  MUX2_X1 U14373 ( .A(n12007), .B(n12006), .S(n12044), .Z(n12008) );
  OAI21_X1 U14374 ( .B1(n12010), .B2(n12009), .A(n12008), .ZN(n12015) );
  MUX2_X1 U14375 ( .A(n12012), .B(n12011), .S(n12070), .Z(n12014) );
  AOI211_X1 U14376 ( .C1(n12015), .C2(n12014), .A(n12013), .B(n9340), .ZN(
        n12028) );
  INV_X1 U14377 ( .A(n12019), .ZN(n12017) );
  OAI211_X1 U14378 ( .C1(n12017), .C2(n12016), .A(n12025), .B(n12018), .ZN(
        n12023) );
  INV_X1 U14379 ( .A(n12018), .ZN(n12021) );
  OAI211_X1 U14380 ( .C1(n12021), .C2(n12020), .A(n12024), .B(n12019), .ZN(
        n12022) );
  MUX2_X1 U14381 ( .A(n12023), .B(n12022), .S(n12044), .Z(n12027) );
  MUX2_X1 U14382 ( .A(n12025), .B(n12024), .S(n12070), .Z(n12026) );
  OAI21_X1 U14383 ( .B1(n12028), .B2(n12027), .A(n12026), .ZN(n12032) );
  MUX2_X1 U14384 ( .A(n12030), .B(n12029), .S(n12070), .Z(n12031) );
  OAI211_X1 U14385 ( .C1(n12032), .C2(n12519), .A(n9344), .B(n12031), .ZN(
        n12037) );
  INV_X1 U14386 ( .A(n12496), .ZN(n12036) );
  MUX2_X1 U14387 ( .A(n12034), .B(n12033), .S(n12044), .Z(n12035) );
  AND3_X1 U14388 ( .A1(n12037), .A2(n12036), .A3(n12035), .ZN(n12041) );
  MUX2_X1 U14389 ( .A(n12039), .B(n12038), .S(n12044), .Z(n12040) );
  OAI33_X1 U14390 ( .A1(n12044), .A2(n12739), .A3(n9346), .B1(n12483), .B2(
        n12041), .B3(n12040), .ZN(n12049) );
  INV_X1 U14391 ( .A(n12469), .ZN(n12048) );
  AOI21_X1 U14392 ( .B1(n12043), .B2(n12042), .A(n12046), .ZN(n12045) );
  MUX2_X1 U14393 ( .A(n12046), .B(n12045), .S(n12044), .Z(n12047) );
  AOI211_X1 U14394 ( .C1(n12049), .C2(n12048), .A(n12047), .B(n12458), .ZN(
        n12054) );
  INV_X1 U14395 ( .A(n12050), .ZN(n12051) );
  MUX2_X1 U14396 ( .A(n12052), .B(n12051), .S(n12070), .Z(n12053) );
  NOR3_X1 U14397 ( .A1(n12054), .A2(n12444), .A3(n12053), .ZN(n12060) );
  INV_X1 U14398 ( .A(n12055), .ZN(n12056) );
  MUX2_X1 U14399 ( .A(n12057), .B(n12056), .S(n12070), .Z(n12059) );
  OAI21_X1 U14400 ( .B1(n12060), .B2(n12059), .A(n12058), .ZN(n12069) );
  INV_X1 U14401 ( .A(n12061), .ZN(n12062) );
  AOI21_X1 U14402 ( .B1(n12064), .B2(n12063), .A(n12062), .ZN(n12065) );
  OAI211_X1 U14403 ( .C1(n12070), .C2(n12066), .A(n12069), .B(n12065), .ZN(
        n12068) );
  OAI211_X1 U14404 ( .C1(n12070), .C2(n12069), .A(n12068), .B(n12067), .ZN(
        n12073) );
  AOI22_X1 U14405 ( .A1(n12073), .A2(n12072), .B1(n7409), .B2(n12071), .ZN(
        n12074) );
  MUX2_X1 U14406 ( .A(n12076), .B(n12075), .S(n12074), .Z(n12077) );
  OAI21_X1 U14407 ( .B1(n12079), .B2(n12078), .A(n12077), .ZN(n12080) );
  AOI21_X1 U14408 ( .B1(n12082), .B2(n12081), .A(n12080), .ZN(n12089) );
  NAND3_X1 U14409 ( .A1(n12631), .A2(n12084), .A3(n12083), .ZN(n12085) );
  OAI211_X1 U14410 ( .C1(n12086), .C2(n12088), .A(n12085), .B(P3_B_REG_SCAN_IN), .ZN(n12087) );
  OAI21_X1 U14411 ( .B1(n12089), .B2(n12088), .A(n12087), .ZN(P3_U3296) );
  MUX2_X1 U14412 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12090), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14413 ( .A(n12091), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12107), .Z(
        P3_U3521) );
  MUX2_X1 U14414 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12092), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14415 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12093), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14416 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12094), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14417 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12095), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14418 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12096), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14419 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12453), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14420 ( .A(n9346), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12107), .Z(
        P3_U3514) );
  MUX2_X1 U14421 ( .A(n12507), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12107), .Z(
        P3_U3513) );
  MUX2_X1 U14422 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12097), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14423 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12534), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14424 ( .A(n12098), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12107), .Z(
        P3_U3510) );
  MUX2_X1 U14425 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12558), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14426 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12570), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14427 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12557), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14428 ( .A(n12603), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12107), .Z(
        P3_U3506) );
  MUX2_X1 U14429 ( .A(n12617), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12107), .Z(
        P3_U3505) );
  MUX2_X1 U14430 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12634), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14431 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12616), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14432 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12632), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14433 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12099), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14434 ( .A(n12100), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12107), .Z(
        P3_U3500) );
  MUX2_X1 U14435 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12101), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14436 ( .A(n12102), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12107), .Z(
        P3_U3498) );
  MUX2_X1 U14437 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12103), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14438 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12104), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14439 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12105), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14440 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n9268), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14441 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12106), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14442 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n8806), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14443 ( .A(n12108), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12107), .Z(
        P3_U3491) );
  NAND2_X1 U14444 ( .A1(keyinput35), .A2(keyinput84), .ZN(n12109) );
  NOR3_X1 U14445 ( .A1(keyinput68), .A2(keyinput89), .A3(n12109), .ZN(n12169)
         );
  NAND2_X1 U14446 ( .A1(keyinput8), .A2(keyinput112), .ZN(n12110) );
  NOR3_X1 U14447 ( .A1(keyinput73), .A2(keyinput104), .A3(n12110), .ZN(n12168)
         );
  NAND2_X1 U14448 ( .A1(keyinput72), .A2(keyinput29), .ZN(n12111) );
  NOR3_X1 U14449 ( .A1(keyinput70), .A2(keyinput10), .A3(n12111), .ZN(n12112)
         );
  NAND3_X1 U14450 ( .A1(keyinput65), .A2(keyinput63), .A3(n12112), .ZN(n12119)
         );
  OR4_X1 U14451 ( .A1(keyinput38), .A2(keyinput88), .A3(keyinput76), .A4(
        keyinput33), .ZN(n12113) );
  NOR4_X1 U14452 ( .A1(keyinput75), .A2(keyinput83), .A3(keyinput121), .A4(
        n12113), .ZN(n12117) );
  NOR2_X1 U14453 ( .A1(keyinput69), .A2(keyinput91), .ZN(n12114) );
  NAND3_X1 U14454 ( .A1(keyinput25), .A2(keyinput56), .A3(n12114), .ZN(n12115)
         );
  NOR3_X1 U14455 ( .A1(keyinput66), .A2(keyinput113), .A3(n12115), .ZN(n12116)
         );
  NAND4_X1 U14456 ( .A1(n12117), .A2(keyinput126), .A3(keyinput47), .A4(n12116), .ZN(n12118) );
  NOR4_X1 U14457 ( .A1(keyinput32), .A2(keyinput97), .A3(n12119), .A4(n12118), 
        .ZN(n12167) );
  INV_X1 U14458 ( .A(keyinput93), .ZN(n12122) );
  NOR2_X1 U14459 ( .A1(keyinput31), .A2(keyinput107), .ZN(n12120) );
  NAND3_X1 U14460 ( .A1(keyinput59), .A2(keyinput36), .A3(n12120), .ZN(n12121)
         );
  NOR3_X1 U14461 ( .A1(keyinput20), .A2(n12122), .A3(n12121), .ZN(n12133) );
  NOR4_X1 U14462 ( .A1(keyinput78), .A2(keyinput39), .A3(keyinput30), .A4(
        keyinput24), .ZN(n12123) );
  NAND3_X1 U14463 ( .A1(keyinput41), .A2(keyinput111), .A3(n12123), .ZN(n12131) );
  NAND3_X1 U14464 ( .A1(keyinput7), .A2(keyinput11), .A3(keyinput3), .ZN(
        n12124) );
  NOR2_X1 U14465 ( .A1(keyinput98), .A2(n12124), .ZN(n12129) );
  NOR4_X1 U14466 ( .A1(keyinput81), .A2(keyinput12), .A3(keyinput120), .A4(
        keyinput1), .ZN(n12128) );
  NOR4_X1 U14467 ( .A1(keyinput50), .A2(keyinput119), .A3(keyinput18), .A4(
        keyinput17), .ZN(n12127) );
  NAND2_X1 U14468 ( .A1(keyinput53), .A2(keyinput43), .ZN(n12125) );
  NOR3_X1 U14469 ( .A1(keyinput116), .A2(keyinput99), .A3(n12125), .ZN(n12126)
         );
  NAND4_X1 U14470 ( .A1(n12129), .A2(n12128), .A3(n12127), .A4(n12126), .ZN(
        n12130) );
  NOR4_X1 U14471 ( .A1(keyinput100), .A2(keyinput28), .A3(n12131), .A4(n12130), 
        .ZN(n12132) );
  NAND4_X1 U14472 ( .A1(keyinput21), .A2(keyinput127), .A3(n12133), .A4(n12132), .ZN(n12165) );
  NOR2_X1 U14473 ( .A1(keyinput74), .A2(keyinput115), .ZN(n12134) );
  NAND3_X1 U14474 ( .A1(keyinput49), .A2(keyinput110), .A3(n12134), .ZN(n12140) );
  INV_X1 U14475 ( .A(keyinput51), .ZN(n12135) );
  NAND4_X1 U14476 ( .A1(keyinput45), .A2(keyinput9), .A3(keyinput103), .A4(
        n12135), .ZN(n12139) );
  NOR2_X1 U14477 ( .A1(keyinput86), .A2(keyinput87), .ZN(n12136) );
  NAND3_X1 U14478 ( .A1(keyinput61), .A2(keyinput34), .A3(n12136), .ZN(n12138)
         );
  NAND4_X1 U14479 ( .A1(keyinput85), .A2(keyinput105), .A3(keyinput58), .A4(
        keyinput118), .ZN(n12137) );
  OR4_X1 U14480 ( .A1(n12140), .A2(n12139), .A3(n12138), .A4(n12137), .ZN(
        n12164) );
  NOR4_X1 U14481 ( .A1(keyinput46), .A2(keyinput37), .A3(keyinput54), .A4(
        keyinput92), .ZN(n12147) );
  NAND2_X1 U14482 ( .A1(keyinput96), .A2(keyinput44), .ZN(n12141) );
  NOR3_X1 U14483 ( .A1(keyinput80), .A2(keyinput124), .A3(n12141), .ZN(n12146)
         );
  INV_X1 U14484 ( .A(keyinput42), .ZN(n12142) );
  NOR4_X1 U14485 ( .A1(keyinput0), .A2(keyinput4), .A3(keyinput108), .A4(
        n12142), .ZN(n12145) );
  NAND2_X1 U14486 ( .A1(keyinput52), .A2(keyinput14), .ZN(n12143) );
  NOR3_X1 U14487 ( .A1(keyinput114), .A2(keyinput67), .A3(n12143), .ZN(n12144)
         );
  NAND4_X1 U14488 ( .A1(n12147), .A2(n12146), .A3(n12145), .A4(n12144), .ZN(
        n12163) );
  INV_X1 U14489 ( .A(keyinput19), .ZN(n12148) );
  NAND4_X1 U14490 ( .A1(keyinput77), .A2(keyinput79), .A3(keyinput94), .A4(
        n12148), .ZN(n12149) );
  NOR3_X1 U14491 ( .A1(keyinput117), .A2(keyinput109), .A3(n12149), .ZN(n12161) );
  NAND2_X1 U14492 ( .A1(keyinput15), .A2(keyinput55), .ZN(n12150) );
  NOR3_X1 U14493 ( .A1(keyinput40), .A2(keyinput5), .A3(n12150), .ZN(n12151)
         );
  NAND3_X1 U14494 ( .A1(keyinput82), .A2(keyinput60), .A3(n12151), .ZN(n12158)
         );
  NOR4_X1 U14495 ( .A1(keyinput101), .A2(keyinput57), .A3(keyinput123), .A4(
        keyinput2), .ZN(n12156) );
  NAND2_X1 U14496 ( .A1(keyinput62), .A2(keyinput23), .ZN(n12152) );
  NOR3_X1 U14497 ( .A1(keyinput6), .A2(keyinput90), .A3(n12152), .ZN(n12155)
         );
  AND4_X1 U14498 ( .A1(keyinput64), .A2(keyinput26), .A3(keyinput13), .A4(
        keyinput27), .ZN(n12154) );
  NOR4_X1 U14499 ( .A1(keyinput95), .A2(keyinput125), .A3(keyinput16), .A4(
        keyinput122), .ZN(n12153) );
  NAND4_X1 U14500 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n12157) );
  NOR4_X1 U14501 ( .A1(keyinput106), .A2(keyinput102), .A3(n12158), .A4(n12157), .ZN(n12160) );
  INV_X1 U14502 ( .A(keyinput22), .ZN(n12159) );
  NAND4_X1 U14503 ( .A1(keyinput71), .A2(n12161), .A3(n12160), .A4(n12159), 
        .ZN(n12162) );
  NOR4_X1 U14504 ( .A1(n12165), .A2(n12164), .A3(n12163), .A4(n12162), .ZN(
        n12166) );
  NAND4_X1 U14505 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n12170) );
  AND2_X1 U14506 ( .A1(n12170), .A2(keyinput48), .ZN(n12379) );
  INV_X1 U14507 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15121) );
  AOI22_X1 U14508 ( .A1(n13545), .A2(keyinput37), .B1(n15121), .B2(keyinput54), 
        .ZN(n12171) );
  OAI221_X1 U14509 ( .B1(n13545), .B2(keyinput37), .C1(n15121), .C2(keyinput54), .A(n12171), .ZN(n12182) );
  AOI22_X1 U14510 ( .A1(n12174), .A2(keyinput124), .B1(n12173), .B2(keyinput45), .ZN(n12172) );
  OAI221_X1 U14511 ( .B1(n12174), .B2(keyinput124), .C1(n12173), .C2(
        keyinput45), .A(n12172), .ZN(n12181) );
  INV_X1 U14512 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n13551) );
  AOI22_X1 U14513 ( .A1(n12176), .A2(keyinput44), .B1(n13551), .B2(keyinput46), 
        .ZN(n12175) );
  OAI221_X1 U14514 ( .B1(n12176), .B2(keyinput44), .C1(n13551), .C2(keyinput46), .A(n12175), .ZN(n12180) );
  XNOR2_X1 U14515 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput92), .ZN(n12178) );
  XNOR2_X1 U14516 ( .A(P3_REG3_REG_9__SCAN_IN), .B(keyinput96), .ZN(n12177) );
  NAND2_X1 U14517 ( .A1(n12178), .A2(n12177), .ZN(n12179) );
  NOR4_X1 U14518 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(
        n12218) );
  AOI22_X1 U14519 ( .A1(n11374), .A2(keyinput51), .B1(keyinput9), .B2(n12184), 
        .ZN(n12183) );
  OAI221_X1 U14520 ( .B1(n11374), .B2(keyinput51), .C1(n12184), .C2(keyinput9), 
        .A(n12183), .ZN(n12194) );
  INV_X1 U14521 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U14522 ( .A1(n7910), .A2(keyinput49), .B1(keyinput115), .B2(n12186), 
        .ZN(n12185) );
  OAI221_X1 U14523 ( .B1(n7910), .B2(keyinput49), .C1(n12186), .C2(keyinput115), .A(n12185), .ZN(n12193) );
  XNOR2_X1 U14524 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput85), .ZN(n12189) );
  XNOR2_X1 U14525 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput74), .ZN(n12188) );
  XNOR2_X1 U14526 ( .A(P3_IR_REG_16__SCAN_IN), .B(keyinput103), .ZN(n12187) );
  NAND3_X1 U14527 ( .A1(n12189), .A2(n12188), .A3(n12187), .ZN(n12192) );
  XNOR2_X1 U14528 ( .A(n12190), .B(keyinput110), .ZN(n12191) );
  NOR4_X1 U14529 ( .A1(n12194), .A2(n12193), .A3(n12192), .A4(n12191), .ZN(
        n12217) );
  INV_X1 U14530 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15130) );
  INV_X1 U14531 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14802) );
  AOI22_X1 U14532 ( .A1(n15130), .A2(keyinput105), .B1(keyinput86), .B2(n14802), .ZN(n12195) );
  OAI221_X1 U14533 ( .B1(n15130), .B2(keyinput105), .C1(n14802), .C2(
        keyinput86), .A(n12195), .ZN(n12203) );
  INV_X1 U14534 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12708) );
  INV_X1 U14535 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n13689) );
  AOI22_X1 U14536 ( .A1(n12708), .A2(keyinput61), .B1(keyinput34), .B2(n13689), 
        .ZN(n12196) );
  OAI221_X1 U14537 ( .B1(n12708), .B2(keyinput61), .C1(n13689), .C2(keyinput34), .A(n12196), .ZN(n12202) );
  INV_X1 U14538 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15116) );
  INV_X1 U14539 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15316) );
  AOI22_X1 U14540 ( .A1(n15116), .A2(keyinput87), .B1(keyinput58), .B2(n15316), 
        .ZN(n12197) );
  OAI221_X1 U14541 ( .B1(n15116), .B2(keyinput87), .C1(n15316), .C2(keyinput58), .A(n12197), .ZN(n12201) );
  AOI22_X1 U14542 ( .A1(n12199), .A2(keyinput118), .B1(keyinput14), .B2(n14691), .ZN(n12198) );
  OAI221_X1 U14543 ( .B1(n12199), .B2(keyinput118), .C1(n14691), .C2(
        keyinput14), .A(n12198), .ZN(n12200) );
  NOR4_X1 U14544 ( .A1(n12203), .A2(n12202), .A3(n12201), .A4(n12200), .ZN(
        n12216) );
  INV_X1 U14545 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n13585) );
  AOI22_X1 U14546 ( .A1(n9962), .A2(keyinput108), .B1(keyinput22), .B2(n13585), 
        .ZN(n12204) );
  OAI221_X1 U14547 ( .B1(n9962), .B2(keyinput108), .C1(n13585), .C2(keyinput22), .A(n12204), .ZN(n12214) );
  INV_X1 U14548 ( .A(keyinput4), .ZN(n12205) );
  XOR2_X1 U14549 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12205), .Z(n12210) );
  XOR2_X1 U14550 ( .A(n12206), .B(keyinput67), .Z(n12209) );
  XNOR2_X1 U14551 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput114), .ZN(n12208) );
  XNOR2_X1 U14552 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput42), .ZN(n12207) );
  NAND4_X1 U14553 ( .A1(n12210), .A2(n12209), .A3(n12208), .A4(n12207), .ZN(
        n12213) );
  INV_X1 U14554 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13468) );
  AOI22_X1 U14555 ( .A1(n12476), .A2(keyinput52), .B1(keyinput0), .B2(n13468), 
        .ZN(n12211) );
  OAI221_X1 U14556 ( .B1(n12476), .B2(keyinput52), .C1(n13468), .C2(keyinput0), 
        .A(n12211), .ZN(n12212) );
  NOR3_X1 U14557 ( .A1(n12214), .A2(n12213), .A3(n12212), .ZN(n12215) );
  NAND4_X1 U14558 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12376) );
  INV_X1 U14559 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15125) );
  INV_X1 U14560 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14698) );
  AOI22_X1 U14561 ( .A1(n15125), .A2(keyinput71), .B1(keyinput19), .B2(n14698), 
        .ZN(n12219) );
  OAI221_X1 U14562 ( .B1(n15125), .B2(keyinput71), .C1(n14698), .C2(keyinput19), .A(n12219), .ZN(n12229) );
  INV_X1 U14563 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U14564 ( .A1(n7468), .A2(keyinput94), .B1(n12221), .B2(keyinput117), 
        .ZN(n12220) );
  OAI221_X1 U14565 ( .B1(n7468), .B2(keyinput94), .C1(n12221), .C2(keyinput117), .A(n12220), .ZN(n12228) );
  AOI22_X1 U14566 ( .A1(n13410), .A2(keyinput109), .B1(keyinput6), .B2(n12223), 
        .ZN(n12222) );
  OAI221_X1 U14567 ( .B1(n13410), .B2(keyinput109), .C1(n12223), .C2(keyinput6), .A(n12222), .ZN(n12227) );
  XNOR2_X1 U14568 ( .A(P3_REG2_REG_2__SCAN_IN), .B(keyinput79), .ZN(n12225) );
  XNOR2_X1 U14569 ( .A(P3_IR_REG_3__SCAN_IN), .B(keyinput77), .ZN(n12224) );
  NAND2_X1 U14570 ( .A1(n12225), .A2(n12224), .ZN(n12226) );
  NOR4_X1 U14571 ( .A1(n12229), .A2(n12228), .A3(n12227), .A4(n12226), .ZN(
        n12267) );
  INV_X1 U14572 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14809) );
  AOI22_X1 U14573 ( .A1(n14809), .A2(keyinput23), .B1(n10861), .B2(keyinput101), .ZN(n12230) );
  OAI221_X1 U14574 ( .B1(n14809), .B2(keyinput23), .C1(n10861), .C2(
        keyinput101), .A(n12230), .ZN(n12239) );
  INV_X1 U14575 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15318) );
  INV_X1 U14576 ( .A(keyinput62), .ZN(n12232) );
  AOI22_X1 U14577 ( .A1(n15318), .A2(keyinput57), .B1(P3_DATAO_REG_30__SCAN_IN), .B2(n12232), .ZN(n12231) );
  OAI221_X1 U14578 ( .B1(n15318), .B2(keyinput57), .C1(n12232), .C2(
        P3_DATAO_REG_30__SCAN_IN), .A(n12231), .ZN(n12238) );
  INV_X1 U14579 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15315) );
  AOI22_X1 U14580 ( .A1(n15315), .A2(keyinput90), .B1(keyinput123), .B2(n12234), .ZN(n12233) );
  OAI221_X1 U14581 ( .B1(n15315), .B2(keyinput90), .C1(n12234), .C2(
        keyinput123), .A(n12233), .ZN(n12237) );
  INV_X1 U14582 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15144) );
  AOI22_X1 U14583 ( .A1(n15144), .A2(keyinput2), .B1(keyinput95), .B2(n9507), 
        .ZN(n12235) );
  OAI221_X1 U14584 ( .B1(n15144), .B2(keyinput2), .C1(n9507), .C2(keyinput95), 
        .A(n12235), .ZN(n12236) );
  NOR4_X1 U14585 ( .A1(n12239), .A2(n12238), .A3(n12237), .A4(n12236), .ZN(
        n12266) );
  INV_X1 U14586 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U14587 ( .A1(n12241), .A2(keyinput27), .B1(n15219), .B2(keyinput16), 
        .ZN(n12240) );
  OAI221_X1 U14588 ( .B1(n12241), .B2(keyinput27), .C1(n15219), .C2(keyinput16), .A(n12240), .ZN(n12251) );
  AOI22_X1 U14589 ( .A1(n14725), .A2(keyinput125), .B1(n12243), .B2(keyinput64), .ZN(n12242) );
  OAI221_X1 U14590 ( .B1(n14725), .B2(keyinput125), .C1(n12243), .C2(
        keyinput64), .A(n12242), .ZN(n12250) );
  INV_X1 U14591 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12245) );
  INV_X1 U14592 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n13835) );
  AOI22_X1 U14593 ( .A1(n12245), .A2(keyinput122), .B1(keyinput40), .B2(n13835), .ZN(n12244) );
  OAI221_X1 U14594 ( .B1(n12245), .B2(keyinput122), .C1(n13835), .C2(
        keyinput40), .A(n12244), .ZN(n12249) );
  INV_X1 U14595 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14734) );
  XOR2_X1 U14596 ( .A(n14734), .B(keyinput13), .Z(n12247) );
  XNOR2_X1 U14597 ( .A(P3_IR_REG_20__SCAN_IN), .B(keyinput26), .ZN(n12246) );
  NAND2_X1 U14598 ( .A1(n12247), .A2(n12246), .ZN(n12248) );
  NOR4_X1 U14599 ( .A1(n12251), .A2(n12250), .A3(n12249), .A4(n12248), .ZN(
        n12265) );
  INV_X1 U14600 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14777) );
  AOI22_X1 U14601 ( .A1(n13413), .A2(keyinput55), .B1(keyinput82), .B2(n14777), 
        .ZN(n12252) );
  OAI221_X1 U14602 ( .B1(n13413), .B2(keyinput55), .C1(n14777), .C2(keyinput82), .A(n12252), .ZN(n12263) );
  AOI22_X1 U14603 ( .A1(n12254), .A2(keyinput60), .B1(keyinput5), .B2(n13849), 
        .ZN(n12253) );
  OAI221_X1 U14604 ( .B1(n12254), .B2(keyinput60), .C1(n13849), .C2(keyinput5), 
        .A(n12253), .ZN(n12262) );
  AOI22_X1 U14605 ( .A1(n12257), .A2(keyinput15), .B1(n12256), .B2(keyinput106), .ZN(n12255) );
  OAI221_X1 U14606 ( .B1(n12257), .B2(keyinput15), .C1(n12256), .C2(
        keyinput106), .A(n12255), .ZN(n12261) );
  XNOR2_X1 U14607 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput102), .ZN(n12259) );
  XNOR2_X1 U14608 ( .A(keyinput75), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U14609 ( .A1(n12259), .A2(n12258), .ZN(n12260) );
  NOR4_X1 U14610 ( .A1(n12263), .A2(n12262), .A3(n12261), .A4(n12260), .ZN(
        n12264) );
  NAND4_X1 U14611 ( .A1(n12267), .A2(n12266), .A3(n12265), .A4(n12264), .ZN(
        n12375) );
  AOI22_X1 U14612 ( .A1(n12269), .A2(keyinput17), .B1(keyinput100), .B2(n10438), .ZN(n12268) );
  OAI221_X1 U14613 ( .B1(n12269), .B2(keyinput17), .C1(n10438), .C2(
        keyinput100), .A(n12268), .ZN(n12277) );
  INV_X1 U14614 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15109) );
  INV_X1 U14615 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15319) );
  AOI22_X1 U14616 ( .A1(n15109), .A2(keyinput99), .B1(keyinput50), .B2(n15319), 
        .ZN(n12270) );
  OAI221_X1 U14617 ( .B1(n15109), .B2(keyinput99), .C1(n15319), .C2(keyinput50), .A(n12270), .ZN(n12276) );
  INV_X1 U14618 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14694) );
  INV_X1 U14619 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n13636) );
  AOI22_X1 U14620 ( .A1(n14694), .A2(keyinput119), .B1(n13636), .B2(keyinput18), .ZN(n12271) );
  OAI221_X1 U14621 ( .B1(n14694), .B2(keyinput119), .C1(n13636), .C2(
        keyinput18), .A(n12271), .ZN(n12275) );
  XNOR2_X1 U14622 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput116), .ZN(n12273) );
  XNOR2_X1 U14623 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput53), .ZN(n12272)
         );
  NAND2_X1 U14624 ( .A1(n12273), .A2(n12272), .ZN(n12274) );
  NOR4_X1 U14625 ( .A1(n12277), .A2(n12276), .A3(n12275), .A4(n12274), .ZN(
        n12316) );
  INV_X1 U14626 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15113) );
  AOI22_X1 U14627 ( .A1(n15113), .A2(keyinput12), .B1(n12279), .B2(keyinput98), 
        .ZN(n12278) );
  OAI221_X1 U14628 ( .B1(n15113), .B2(keyinput12), .C1(n12279), .C2(keyinput98), .A(n12278), .ZN(n12287) );
  AOI22_X1 U14629 ( .A1(n14949), .A2(keyinput3), .B1(n9033), .B2(keyinput120), 
        .ZN(n12280) );
  OAI221_X1 U14630 ( .B1(n14949), .B2(keyinput3), .C1(n9033), .C2(keyinput120), 
        .A(n12280), .ZN(n12286) );
  XNOR2_X1 U14631 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput43), .ZN(n12284) );
  XNOR2_X1 U14632 ( .A(P3_REG2_REG_30__SCAN_IN), .B(keyinput7), .ZN(n12283) );
  XNOR2_X1 U14633 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput11), .ZN(n12282)
         );
  XNOR2_X1 U14634 ( .A(keyinput1), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n12281) );
  NAND4_X1 U14635 ( .A1(n12284), .A2(n12283), .A3(n12282), .A4(n12281), .ZN(
        n12285) );
  NOR3_X1 U14636 ( .A1(n12287), .A2(n12286), .A3(n12285), .ZN(n12315) );
  INV_X1 U14637 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n13428) );
  AOI22_X1 U14638 ( .A1(n13428), .A2(keyinput93), .B1(n13408), .B2(keyinput59), 
        .ZN(n12288) );
  OAI221_X1 U14639 ( .B1(n13428), .B2(keyinput93), .C1(n13408), .C2(keyinput59), .A(n12288), .ZN(n12299) );
  INV_X1 U14640 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U14641 ( .A1(n12290), .A2(keyinput127), .B1(n15082), .B2(keyinput20), .ZN(n12289) );
  OAI221_X1 U14642 ( .B1(n12290), .B2(keyinput127), .C1(n15082), .C2(
        keyinput20), .A(n12289), .ZN(n12298) );
  INV_X1 U14643 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U14644 ( .A1(n12293), .A2(keyinput36), .B1(n12292), .B2(keyinput80), 
        .ZN(n12291) );
  OAI221_X1 U14645 ( .B1(n12293), .B2(keyinput36), .C1(n12292), .C2(keyinput80), .A(n12291), .ZN(n12297) );
  INV_X1 U14646 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U14647 ( .A1(n12295), .A2(keyinput107), .B1(n10367), .B2(keyinput31), .ZN(n12294) );
  OAI221_X1 U14648 ( .B1(n12295), .B2(keyinput107), .C1(n10367), .C2(
        keyinput31), .A(n12294), .ZN(n12296) );
  NOR4_X1 U14649 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12314) );
  INV_X1 U14650 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U14651 ( .A1(n14435), .A2(keyinput111), .B1(keyinput21), .B2(n12301), .ZN(n12300) );
  OAI221_X1 U14652 ( .B1(n14435), .B2(keyinput111), .C1(n12301), .C2(
        keyinput21), .A(n12300), .ZN(n12305) );
  XOR2_X1 U14653 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput28), .Z(n12304) );
  XOR2_X1 U14654 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput30), .Z(n12303) );
  XNOR2_X1 U14655 ( .A(keyinput39), .B(n10080), .ZN(n12302) );
  OR4_X1 U14656 ( .A1(n12305), .A2(n12304), .A3(n12303), .A4(n12302), .ZN(
        n12312) );
  XNOR2_X1 U14657 ( .A(n12306), .B(keyinput41), .ZN(n12311) );
  XNOR2_X1 U14658 ( .A(n12307), .B(keyinput24), .ZN(n12310) );
  INV_X1 U14659 ( .A(keyinput78), .ZN(n12308) );
  XNOR2_X1 U14660 ( .A(n12308), .B(P3_DATAO_REG_8__SCAN_IN), .ZN(n12309) );
  NOR4_X1 U14661 ( .A1(n12312), .A2(n12311), .A3(n12310), .A4(n12309), .ZN(
        n12313) );
  NAND4_X1 U14662 ( .A1(n12316), .A2(n12315), .A3(n12314), .A4(n12313), .ZN(
        n12374) );
  INV_X1 U14663 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15117) );
  AOI22_X1 U14664 ( .A1(n15117), .A2(keyinput63), .B1(keyinput32), .B2(n8567), 
        .ZN(n12317) );
  OAI221_X1 U14665 ( .B1(n15117), .B2(keyinput63), .C1(n8567), .C2(keyinput32), 
        .A(n12317), .ZN(n12328) );
  INV_X1 U14666 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12680) );
  INV_X1 U14667 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U14668 ( .A1(n12680), .A2(keyinput72), .B1(keyinput65), .B2(n12319), 
        .ZN(n12318) );
  OAI221_X1 U14669 ( .B1(n12680), .B2(keyinput72), .C1(n12319), .C2(keyinput65), .A(n12318), .ZN(n12327) );
  INV_X1 U14670 ( .A(keyinput70), .ZN(n12321) );
  AOI22_X1 U14671 ( .A1(n12322), .A2(keyinput10), .B1(P3_DATAO_REG_25__SCAN_IN), .B2(n12321), .ZN(n12320) );
  OAI221_X1 U14672 ( .B1(n12322), .B2(keyinput10), .C1(n12321), .C2(
        P3_DATAO_REG_25__SCAN_IN), .A(n12320), .ZN(n12326) );
  XOR2_X1 U14673 ( .A(n7911), .B(keyinput97), .Z(n12324) );
  XNOR2_X1 U14674 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput112), .ZN(n12323) );
  NAND2_X1 U14675 ( .A1(n12324), .A2(n12323), .ZN(n12325) );
  NOR4_X1 U14676 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n12325), .ZN(
        n12372) );
  XNOR2_X1 U14677 ( .A(n12329), .B(keyinput121), .ZN(n12330) );
  AOI21_X1 U14678 ( .B1(keyinput48), .B2(n12378), .A(n12330), .ZN(n12334) );
  INV_X1 U14679 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12331) );
  XOR2_X1 U14680 ( .A(n12331), .B(keyinput38), .Z(n12333) );
  INV_X1 U14681 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15609) );
  XOR2_X1 U14682 ( .A(n15609), .B(keyinput83), .Z(n12332) );
  NAND3_X1 U14683 ( .A1(n12334), .A2(n12333), .A3(n12332), .ZN(n12343) );
  INV_X1 U14684 ( .A(keyinput88), .ZN(n12337) );
  INV_X1 U14685 ( .A(keyinput76), .ZN(n12336) );
  AOI22_X1 U14686 ( .A1(n12337), .A2(P3_DATAO_REG_29__SCAN_IN), .B1(
        P3_RD_REG_SCAN_IN), .B2(n12336), .ZN(n12335) );
  OAI221_X1 U14687 ( .B1(n12337), .B2(P3_DATAO_REG_29__SCAN_IN), .C1(n12336), 
        .C2(P3_RD_REG_SCAN_IN), .A(n12335), .ZN(n12342) );
  AOI22_X1 U14688 ( .A1(n12340), .A2(keyinput33), .B1(n12339), .B2(keyinput29), 
        .ZN(n12338) );
  OAI221_X1 U14689 ( .B1(n12340), .B2(keyinput33), .C1(n12339), .C2(keyinput29), .A(n12338), .ZN(n12341) );
  NOR3_X1 U14690 ( .A1(n12343), .A2(n12342), .A3(n12341), .ZN(n12371) );
  INV_X1 U14691 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12676) );
  AOI22_X1 U14692 ( .A1(n12345), .A2(keyinput47), .B1(n12676), .B2(keyinput56), 
        .ZN(n12344) );
  OAI221_X1 U14693 ( .B1(n12345), .B2(keyinput47), .C1(n12676), .C2(keyinput56), .A(n12344), .ZN(n12355) );
  AOI22_X1 U14694 ( .A1(n14668), .A2(keyinput25), .B1(n12347), .B2(keyinput126), .ZN(n12346) );
  OAI221_X1 U14695 ( .B1(n14668), .B2(keyinput25), .C1(n12347), .C2(
        keyinput126), .A(n12346), .ZN(n12354) );
  INV_X1 U14696 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U14697 ( .A1(n13416), .A2(keyinput113), .B1(keyinput81), .B2(n12349), .ZN(n12348) );
  OAI221_X1 U14698 ( .B1(n13416), .B2(keyinput113), .C1(n12349), .C2(
        keyinput81), .A(n12348), .ZN(n12353) );
  INV_X1 U14699 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U14700 ( .A1(n12351), .A2(keyinput91), .B1(n12775), .B2(keyinput66), 
        .ZN(n12350) );
  OAI221_X1 U14701 ( .B1(n12351), .B2(keyinput91), .C1(n12775), .C2(keyinput66), .A(n12350), .ZN(n12352) );
  NOR4_X1 U14702 ( .A1(n12355), .A2(n12354), .A3(n12353), .A4(n12352), .ZN(
        n12370) );
  INV_X1 U14703 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U14704 ( .A1(n12358), .A2(keyinput104), .B1(keyinput68), .B2(n12357), .ZN(n12356) );
  OAI221_X1 U14705 ( .B1(n12358), .B2(keyinput104), .C1(n12357), .C2(
        keyinput68), .A(n12356), .ZN(n12368) );
  INV_X1 U14706 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15317) );
  AOI22_X1 U14707 ( .A1(n12360), .A2(keyinput73), .B1(keyinput8), .B2(n15317), 
        .ZN(n12359) );
  OAI221_X1 U14708 ( .B1(n12360), .B2(keyinput73), .C1(n15317), .C2(keyinput8), 
        .A(n12359), .ZN(n12367) );
  AOI22_X1 U14709 ( .A1(n12362), .A2(keyinput35), .B1(n13451), .B2(keyinput69), 
        .ZN(n12361) );
  OAI221_X1 U14710 ( .B1(n12362), .B2(keyinput35), .C1(n13451), .C2(keyinput69), .A(n12361), .ZN(n12366) );
  INV_X1 U14711 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15579) );
  INV_X1 U14712 ( .A(keyinput84), .ZN(n12364) );
  AOI22_X1 U14713 ( .A1(n15579), .A2(keyinput89), .B1(P3_DATAO_REG_7__SCAN_IN), 
        .B2(n12364), .ZN(n12363) );
  OAI221_X1 U14714 ( .B1(n15579), .B2(keyinput89), .C1(n12364), .C2(
        P3_DATAO_REG_7__SCAN_IN), .A(n12363), .ZN(n12365) );
  NOR4_X1 U14715 ( .A1(n12368), .A2(n12367), .A3(n12366), .A4(n12365), .ZN(
        n12369) );
  NAND4_X1 U14716 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12373) );
  NOR4_X1 U14717 ( .A1(n12376), .A2(n12375), .A3(n12374), .A4(n12373), .ZN(
        n12377) );
  OAI21_X1 U14718 ( .B1(n12379), .B2(n12378), .A(n12377), .ZN(n12405) );
  NOR2_X1 U14719 ( .A1(n12381), .A2(n12380), .ZN(n12383) );
  AOI22_X1 U14720 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n14640), .B1(n14601), 
        .B2(n11374), .ZN(n12384) );
  AOI21_X1 U14721 ( .B1(n12385), .B2(n12384), .A(n14578), .ZN(n12401) );
  INV_X1 U14722 ( .A(n15555), .ZN(n15419) );
  MUX2_X1 U14723 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n14633), .Z(n14602) );
  XNOR2_X1 U14724 ( .A(n14602), .B(n14640), .ZN(n12390) );
  OR2_X1 U14725 ( .A1(n12386), .A2(n12393), .ZN(n12388) );
  NAND2_X1 U14726 ( .A1(n12388), .A2(n12387), .ZN(n12389) );
  NAND2_X1 U14727 ( .A1(n12390), .A2(n12389), .ZN(n14603) );
  OAI21_X1 U14728 ( .B1(n12390), .B2(n12389), .A(n14603), .ZN(n12391) );
  AOI22_X1 U14729 ( .A1(n15419), .A2(n14640), .B1(n15543), .B2(n12391), .ZN(
        n12400) );
  NAND2_X1 U14730 ( .A1(n12393), .A2(n12392), .ZN(n12395) );
  INV_X1 U14731 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15604) );
  AOI22_X1 U14732 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n14601), .B1(n14640), 
        .B2(n15604), .ZN(n12396) );
  NAND2_X1 U14733 ( .A1(n12396), .A2(n12397), .ZN(n14639) );
  OAI21_X1 U14734 ( .B1(n12397), .B2(n12396), .A(n14639), .ZN(n12398) );
  NAND2_X1 U14735 ( .A1(n12398), .A2(n15562), .ZN(n12399) );
  OAI211_X1 U14736 ( .C1(n12401), .C2(n15571), .A(n12400), .B(n12399), .ZN(
        n12402) );
  AOI211_X1 U14737 ( .C1(n15535), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n12403), .B(
        n12402), .ZN(n12404) );
  XOR2_X1 U14738 ( .A(n12405), .B(n12404), .Z(P3_U3190) );
  NOR2_X1 U14739 ( .A1(n12407), .A2(n12406), .ZN(n14897) );
  AND2_X1 U14740 ( .A1(n12624), .A2(n12408), .ZN(n12409) );
  OR2_X1 U14741 ( .A1(n14897), .A2(n12409), .ZN(n12410) );
  NAND2_X1 U14742 ( .A1(n12410), .A2(n14895), .ZN(n14891) );
  NAND2_X1 U14743 ( .A1(n12648), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12411) );
  OAI211_X1 U14744 ( .C1(n12719), .C2(n12595), .A(n14891), .B(n12411), .ZN(
        P3_U3202) );
  AOI21_X1 U14745 ( .B1(n12412), .B2(n12417), .A(n12584), .ZN(n12416) );
  OAI22_X1 U14746 ( .A1(n12413), .A2(n12589), .B1(n12443), .B2(n12587), .ZN(
        n12414) );
  AOI21_X1 U14747 ( .B1(n12416), .B2(n12415), .A(n12414), .ZN(n12654) );
  XNOR2_X1 U14748 ( .A(n12418), .B(n12417), .ZN(n12655) );
  INV_X1 U14749 ( .A(n12655), .ZN(n12423) );
  INV_X1 U14750 ( .A(n12652), .ZN(n12421) );
  AOI22_X1 U14751 ( .A1(n12419), .A2(n12624), .B1(n12648), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12420) );
  OAI21_X1 U14752 ( .B1(n12421), .B2(n12595), .A(n12420), .ZN(n12422) );
  AOI21_X1 U14753 ( .B1(n12423), .B2(n12627), .A(n12422), .ZN(n12424) );
  OAI21_X1 U14754 ( .B1(n12654), .B2(n12648), .A(n12424), .ZN(P3_U3205) );
  XNOR2_X1 U14755 ( .A(n12425), .B(n12428), .ZN(n12434) );
  OAI22_X1 U14756 ( .A1(n6575), .A2(n12589), .B1(n12456), .B2(n12587), .ZN(
        n12430) );
  INV_X1 U14757 ( .A(n12657), .ZN(n12440) );
  INV_X1 U14758 ( .A(n12434), .ZN(n12658) );
  AOI22_X1 U14759 ( .A1(n12435), .A2(n12624), .B1(n12648), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12436) );
  OAI21_X1 U14760 ( .B1(n12723), .B2(n12595), .A(n12436), .ZN(n12437) );
  AOI21_X1 U14761 ( .B1(n12658), .B2(n12438), .A(n12437), .ZN(n12439) );
  OAI21_X1 U14762 ( .B1(n12440), .B2(n12648), .A(n12439), .ZN(P3_U3206) );
  XNOR2_X1 U14763 ( .A(n12441), .B(n12444), .ZN(n12442) );
  OAI222_X1 U14764 ( .A1(n12587), .A2(n12473), .B1(n12589), .B2(n12443), .C1(
        n12584), .C2(n12442), .ZN(n12661) );
  INV_X1 U14765 ( .A(n12661), .ZN(n12450) );
  XNOR2_X1 U14766 ( .A(n12445), .B(n12444), .ZN(n12662) );
  AOI22_X1 U14767 ( .A1(n12648), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n12446), 
        .B2(n12624), .ZN(n12447) );
  OAI21_X1 U14768 ( .B1(n12727), .B2(n12595), .A(n12447), .ZN(n12448) );
  AOI21_X1 U14769 ( .B1(n12662), .B2(n12627), .A(n12448), .ZN(n12449) );
  OAI21_X1 U14770 ( .B1(n12450), .B2(n12648), .A(n12449), .ZN(P3_U3207) );
  OAI211_X1 U14771 ( .C1(n12452), .C2(n12458), .A(n12451), .B(n12636), .ZN(
        n12455) );
  NAND2_X1 U14772 ( .A1(n12453), .A2(n12631), .ZN(n12454) );
  OAI211_X1 U14773 ( .C1(n12456), .C2(n12589), .A(n12455), .B(n12454), .ZN(
        n12665) );
  INV_X1 U14774 ( .A(n12665), .ZN(n12465) );
  AOI21_X1 U14775 ( .B1(n12459), .B2(n12458), .A(n12457), .ZN(n12460) );
  INV_X1 U14776 ( .A(n12460), .ZN(n12666) );
  AOI22_X1 U14777 ( .A1(n12648), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n12624), 
        .B2(n12461), .ZN(n12462) );
  OAI21_X1 U14778 ( .B1(n12731), .B2(n12595), .A(n12462), .ZN(n12463) );
  AOI21_X1 U14779 ( .B1(n12666), .B2(n12627), .A(n12463), .ZN(n12464) );
  OAI21_X1 U14780 ( .B1(n12465), .B2(n12648), .A(n12464), .ZN(P3_U3208) );
  AOI21_X1 U14781 ( .B1(n12469), .B2(n12467), .A(n12466), .ZN(n12669) );
  OAI211_X1 U14782 ( .C1(n12470), .C2(n12469), .A(n12468), .B(n12636), .ZN(
        n12472) );
  NAND2_X1 U14783 ( .A1(n9346), .A2(n12631), .ZN(n12471) );
  OAI211_X1 U14784 ( .C1(n12473), .C2(n12589), .A(n12472), .B(n12471), .ZN(
        n12670) );
  NAND2_X1 U14785 ( .A1(n12670), .A2(n14895), .ZN(n12480) );
  INV_X1 U14786 ( .A(n12474), .ZN(n12475) );
  OAI22_X1 U14787 ( .A1(n14895), .A2(n12476), .B1(n12475), .B2(n12639), .ZN(
        n12477) );
  AOI21_X1 U14788 ( .B1(n12478), .B2(n14893), .A(n12477), .ZN(n12479) );
  OAI211_X1 U14789 ( .C1(n12644), .C2(n12669), .A(n12480), .B(n12479), .ZN(
        P3_U3209) );
  XOR2_X1 U14790 ( .A(n12483), .B(n12481), .Z(n12675) );
  INV_X1 U14791 ( .A(n12675), .ZN(n12492) );
  OAI211_X1 U14792 ( .C1(n12484), .C2(n12483), .A(n12482), .B(n12636), .ZN(
        n12486) );
  NAND2_X1 U14793 ( .A1(n12507), .A2(n12631), .ZN(n12485) );
  OAI211_X1 U14794 ( .C1(n12487), .C2(n12589), .A(n12486), .B(n12485), .ZN(
        n12674) );
  AOI22_X1 U14795 ( .A1(n12648), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12624), 
        .B2(n12488), .ZN(n12489) );
  OAI21_X1 U14796 ( .B1(n12739), .B2(n12595), .A(n12489), .ZN(n12490) );
  AOI21_X1 U14797 ( .B1(n12674), .B2(n14895), .A(n12490), .ZN(n12491) );
  OAI21_X1 U14798 ( .B1(n12644), .B2(n12492), .A(n12491), .ZN(P3_U3210) );
  XNOR2_X1 U14799 ( .A(n12493), .B(n12496), .ZN(n12494) );
  OAI222_X1 U14800 ( .A1(n12589), .A2(n12495), .B1(n12587), .B2(n12522), .C1(
        n12584), .C2(n12494), .ZN(n12678) );
  INV_X1 U14801 ( .A(n12678), .ZN(n12502) );
  XNOR2_X1 U14802 ( .A(n12497), .B(n12496), .ZN(n12679) );
  AOI22_X1 U14803 ( .A1(n12648), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12624), 
        .B2(n12498), .ZN(n12499) );
  OAI21_X1 U14804 ( .B1(n12743), .B2(n12595), .A(n12499), .ZN(n12500) );
  AOI21_X1 U14805 ( .B1(n12679), .B2(n12627), .A(n12500), .ZN(n12501) );
  OAI21_X1 U14806 ( .B1(n12502), .B2(n12648), .A(n12501), .ZN(P3_U3211) );
  NOR2_X1 U14807 ( .A1(n12504), .A2(n12503), .ZN(n12505) );
  OR2_X1 U14808 ( .A1(n12506), .A2(n12505), .ZN(n12511) );
  NAND2_X1 U14809 ( .A1(n12507), .A2(n12633), .ZN(n12508) );
  OAI21_X1 U14810 ( .B1(n12509), .B2(n12587), .A(n12508), .ZN(n12510) );
  AOI21_X1 U14811 ( .B1(n12511), .B2(n12636), .A(n12510), .ZN(n12684) );
  INV_X1 U14812 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12514) );
  INV_X1 U14813 ( .A(n12512), .ZN(n12513) );
  OAI22_X1 U14814 ( .A1(n14895), .A2(n12514), .B1(n12513), .B2(n12639), .ZN(
        n12515) );
  AOI21_X1 U14815 ( .B1(n12516), .B2(n14893), .A(n12515), .ZN(n12518) );
  XNOR2_X1 U14816 ( .A(n6635), .B(n9344), .ZN(n12682) );
  NAND2_X1 U14817 ( .A1(n12682), .A2(n12627), .ZN(n12517) );
  OAI211_X1 U14818 ( .C1(n12684), .C2(n12648), .A(n12518), .B(n12517), .ZN(
        P3_U3212) );
  XNOR2_X1 U14819 ( .A(n12520), .B(n12519), .ZN(n12521) );
  OAI222_X1 U14820 ( .A1(n12589), .A2(n12522), .B1(n12587), .B2(n12549), .C1(
        n12521), .C2(n12584), .ZN(n12687) );
  INV_X1 U14821 ( .A(n12687), .ZN(n12529) );
  XNOR2_X1 U14822 ( .A(n12523), .B(n7860), .ZN(n12688) );
  INV_X1 U14823 ( .A(n12524), .ZN(n12751) );
  AOI22_X1 U14824 ( .A1(n12648), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n12624), 
        .B2(n12525), .ZN(n12526) );
  OAI21_X1 U14825 ( .B1(n12751), .B2(n12595), .A(n12526), .ZN(n12527) );
  AOI21_X1 U14826 ( .B1(n12688), .B2(n12627), .A(n12527), .ZN(n12528) );
  OAI21_X1 U14827 ( .B1(n12529), .B2(n12648), .A(n12528), .ZN(P3_U3213) );
  XOR2_X1 U14828 ( .A(n12530), .B(n12531), .Z(n12692) );
  INV_X1 U14829 ( .A(n12692), .ZN(n12541) );
  OAI211_X1 U14830 ( .C1(n12533), .C2(n9342), .A(n12636), .B(n12532), .ZN(
        n12536) );
  AOI22_X1 U14831 ( .A1(n12631), .A2(n12558), .B1(n12534), .B2(n12633), .ZN(
        n12535) );
  NAND2_X1 U14832 ( .A1(n12536), .A2(n12535), .ZN(n12691) );
  AOI22_X1 U14833 ( .A1(n12648), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n12624), 
        .B2(n12537), .ZN(n12538) );
  OAI21_X1 U14834 ( .B1(n12755), .B2(n12595), .A(n12538), .ZN(n12539) );
  AOI21_X1 U14835 ( .B1(n12691), .B2(n14895), .A(n12539), .ZN(n12540) );
  OAI21_X1 U14836 ( .B1(n12541), .B2(n12644), .A(n12540), .ZN(P3_U3214) );
  XNOR2_X1 U14837 ( .A(n12542), .B(n12546), .ZN(n12695) );
  INV_X1 U14838 ( .A(n12695), .ZN(n12555) );
  INV_X1 U14839 ( .A(n12543), .ZN(n12544) );
  AOI21_X1 U14840 ( .B1(n12546), .B2(n12545), .A(n12544), .ZN(n12547) );
  OAI222_X1 U14841 ( .A1(n12589), .A2(n12549), .B1(n12587), .B2(n12548), .C1(
        n12584), .C2(n12547), .ZN(n12694) );
  INV_X1 U14842 ( .A(n12550), .ZN(n12759) );
  AOI22_X1 U14843 ( .A1(n12648), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n12624), 
        .B2(n12551), .ZN(n12552) );
  OAI21_X1 U14844 ( .B1(n12759), .B2(n12595), .A(n12552), .ZN(n12553) );
  AOI21_X1 U14845 ( .B1(n12694), .B2(n14895), .A(n12553), .ZN(n12554) );
  OAI21_X1 U14846 ( .B1(n12644), .B2(n12555), .A(n12554), .ZN(P3_U3215) );
  XNOR2_X1 U14847 ( .A(n12556), .B(n12561), .ZN(n12559) );
  AOI222_X1 U14848 ( .A1(n12636), .A2(n12559), .B1(n12558), .B2(n12633), .C1(
        n12557), .C2(n12631), .ZN(n12700) );
  OAI21_X1 U14849 ( .B1(n12562), .B2(n12561), .A(n12560), .ZN(n12698) );
  INV_X1 U14850 ( .A(n12697), .ZN(n12565) );
  AOI22_X1 U14851 ( .A1(n12648), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n12624), 
        .B2(n12563), .ZN(n12564) );
  OAI21_X1 U14852 ( .B1(n12565), .B2(n12595), .A(n12564), .ZN(n12566) );
  AOI21_X1 U14853 ( .B1(n12698), .B2(n12627), .A(n12566), .ZN(n12567) );
  OAI21_X1 U14854 ( .B1(n12700), .B2(n12648), .A(n12567), .ZN(P3_U3216) );
  XNOR2_X1 U14855 ( .A(n12568), .B(n12573), .ZN(n12569) );
  NAND2_X1 U14856 ( .A1(n12569), .A2(n12636), .ZN(n12572) );
  AOI22_X1 U14857 ( .A1(n12570), .A2(n12633), .B1(n12631), .B2(n12603), .ZN(
        n12571) );
  NAND2_X1 U14858 ( .A1(n12572), .A2(n12571), .ZN(n12705) );
  INV_X1 U14859 ( .A(n12705), .ZN(n12582) );
  OR2_X1 U14860 ( .A1(n12574), .A2(n12573), .ZN(n12575) );
  NAND2_X1 U14861 ( .A1(n12576), .A2(n12575), .ZN(n12702) );
  INV_X1 U14862 ( .A(n12701), .ZN(n12579) );
  AOI22_X1 U14863 ( .A1(n12648), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12624), 
        .B2(n12577), .ZN(n12578) );
  OAI21_X1 U14864 ( .B1(n12579), .B2(n12595), .A(n12578), .ZN(n12580) );
  AOI21_X1 U14865 ( .B1(n12702), .B2(n12627), .A(n12580), .ZN(n12581) );
  OAI21_X1 U14866 ( .B1(n12582), .B2(n12648), .A(n12581), .ZN(P3_U3217) );
  XOR2_X1 U14867 ( .A(n12583), .B(n12591), .Z(n12585) );
  OAI222_X1 U14868 ( .A1(n12589), .A2(n12588), .B1(n12587), .B2(n12586), .C1(
        n12585), .C2(n12584), .ZN(n12706) );
  INV_X1 U14869 ( .A(n12706), .ZN(n12598) );
  OAI21_X1 U14870 ( .B1(n12592), .B2(n12591), .A(n12590), .ZN(n12707) );
  AOI22_X1 U14871 ( .A1(n12648), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12624), 
        .B2(n12593), .ZN(n12594) );
  OAI21_X1 U14872 ( .B1(n12595), .B2(n12765), .A(n12594), .ZN(n12596) );
  AOI21_X1 U14873 ( .B1(n12707), .B2(n12627), .A(n12596), .ZN(n12597) );
  OAI21_X1 U14874 ( .B1(n12598), .B2(n12648), .A(n12597), .ZN(P3_U3218) );
  NAND2_X1 U14875 ( .A1(n12599), .A2(n12600), .ZN(n12601) );
  NAND3_X1 U14876 ( .A1(n12602), .A2(n12636), .A3(n12601), .ZN(n12605) );
  AOI22_X1 U14877 ( .A1(n12634), .A2(n12631), .B1(n12633), .B2(n12603), .ZN(
        n12604) );
  INV_X1 U14878 ( .A(n12769), .ZN(n12610) );
  INV_X1 U14879 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12608) );
  INV_X1 U14880 ( .A(n12606), .ZN(n12607) );
  OAI22_X1 U14881 ( .A1(n14895), .A2(n12608), .B1(n12607), .B2(n12639), .ZN(
        n12609) );
  AOI21_X1 U14882 ( .B1(n14893), .B2(n12610), .A(n12609), .ZN(n12614) );
  XNOR2_X1 U14883 ( .A(n12612), .B(n12611), .ZN(n12710) );
  NAND2_X1 U14884 ( .A1(n12710), .A2(n12627), .ZN(n12613) );
  OAI211_X1 U14885 ( .C1(n12712), .C2(n12648), .A(n12614), .B(n12613), .ZN(
        P3_U3219) );
  XNOR2_X1 U14886 ( .A(n12615), .B(n12620), .ZN(n12618) );
  AOI222_X1 U14887 ( .A1(n12636), .A2(n12618), .B1(n12617), .B2(n12633), .C1(
        n12616), .C2(n12631), .ZN(n14902) );
  XNOR2_X1 U14888 ( .A(n12619), .B(n12620), .ZN(n14905) );
  OR2_X1 U14889 ( .A1(n12622), .A2(n12621), .ZN(n14901) );
  AOI22_X1 U14890 ( .A1(n12648), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n12624), 
        .B2(n12623), .ZN(n12625) );
  OAI21_X1 U14891 ( .B1(n12641), .B2(n14901), .A(n12625), .ZN(n12626) );
  AOI21_X1 U14892 ( .B1(n14905), .B2(n12627), .A(n12626), .ZN(n12628) );
  OAI21_X1 U14893 ( .B1(n14902), .B2(n12648), .A(n12628), .ZN(P3_U3220) );
  XNOR2_X1 U14894 ( .A(n12629), .B(n12630), .ZN(n12635) );
  AOI222_X1 U14895 ( .A1(n12636), .A2(n12635), .B1(n12634), .B2(n12633), .C1(
        n12632), .C2(n12631), .ZN(n14908) );
  NAND2_X1 U14896 ( .A1(n12637), .A2(n14898), .ZN(n14907) );
  INV_X1 U14897 ( .A(n12638), .ZN(n12640) );
  OAI22_X1 U14898 ( .A1(n12641), .A2(n14907), .B1(n12640), .B2(n12639), .ZN(
        n12646) );
  XNOR2_X1 U14899 ( .A(n12643), .B(n12642), .ZN(n14909) );
  NOR2_X1 U14900 ( .A1(n14909), .A2(n12644), .ZN(n12645) );
  AOI211_X1 U14901 ( .C1(n12648), .C2(P3_REG2_REG_12__SCAN_IN), .A(n12646), 
        .B(n12645), .ZN(n12647) );
  OAI21_X1 U14902 ( .B1(n12648), .B2(n14908), .A(n12647), .ZN(P3_U3221) );
  INV_X1 U14903 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12649) );
  NOR2_X1 U14904 ( .A1(n15611), .A2(n12649), .ZN(n12650) );
  AOI21_X1 U14905 ( .B1(n14897), .B2(n15611), .A(n12650), .ZN(n12651) );
  OAI21_X1 U14906 ( .B1(n12719), .B2(n12715), .A(n12651), .ZN(P3_U3490) );
  NAND2_X1 U14907 ( .A1(n12652), .A2(n14898), .ZN(n12653) );
  OAI211_X1 U14908 ( .C1(n14910), .C2(n12655), .A(n12654), .B(n12653), .ZN(
        n12720) );
  MUX2_X1 U14909 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n12720), .S(n15611), .Z(
        P3_U3487) );
  INV_X1 U14910 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12659) );
  INV_X1 U14911 ( .A(n12656), .ZN(n15591) );
  AOI21_X1 U14912 ( .B1(n15591), .B2(n12658), .A(n12657), .ZN(n12721) );
  MUX2_X1 U14913 ( .A(n12659), .B(n12721), .S(n15611), .Z(n12660) );
  INV_X1 U14914 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12663) );
  AOI21_X1 U14915 ( .B1(n15595), .B2(n12662), .A(n12661), .ZN(n12724) );
  MUX2_X1 U14916 ( .A(n12663), .B(n12724), .S(n15611), .Z(n12664) );
  OAI21_X1 U14917 ( .B1(n12727), .B2(n12715), .A(n12664), .ZN(P3_U3485) );
  INV_X1 U14918 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12667) );
  AOI21_X1 U14919 ( .B1(n15595), .B2(n12666), .A(n12665), .ZN(n12728) );
  MUX2_X1 U14920 ( .A(n12667), .B(n12728), .S(n15611), .Z(n12668) );
  OAI21_X1 U14921 ( .B1(n12731), .B2(n12715), .A(n12668), .ZN(P3_U3484) );
  INV_X1 U14922 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12672) );
  INV_X1 U14923 ( .A(n12669), .ZN(n12671) );
  AOI21_X1 U14924 ( .B1(n15595), .B2(n12671), .A(n12670), .ZN(n12732) );
  MUX2_X1 U14925 ( .A(n12672), .B(n12732), .S(n15611), .Z(n12673) );
  OAI21_X1 U14926 ( .B1(n12735), .B2(n12715), .A(n12673), .ZN(P3_U3483) );
  AOI21_X1 U14927 ( .B1(n15595), .B2(n12675), .A(n12674), .ZN(n12736) );
  MUX2_X1 U14928 ( .A(n12676), .B(n12736), .S(n15611), .Z(n12677) );
  OAI21_X1 U14929 ( .B1(n12739), .B2(n12715), .A(n12677), .ZN(P3_U3482) );
  AOI21_X1 U14930 ( .B1(n15595), .B2(n12679), .A(n12678), .ZN(n12740) );
  MUX2_X1 U14931 ( .A(n12680), .B(n12740), .S(n15611), .Z(n12681) );
  OAI21_X1 U14932 ( .B1(n12743), .B2(n12715), .A(n12681), .ZN(P3_U3481) );
  INV_X1 U14933 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12685) );
  NAND2_X1 U14934 ( .A1(n12682), .A2(n15595), .ZN(n12683) );
  AND2_X1 U14935 ( .A1(n12684), .A2(n12683), .ZN(n12744) );
  MUX2_X1 U14936 ( .A(n12685), .B(n12744), .S(n15611), .Z(n12686) );
  OAI21_X1 U14937 ( .B1(n12747), .B2(n12715), .A(n12686), .ZN(P3_U3480) );
  INV_X1 U14938 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12689) );
  AOI21_X1 U14939 ( .B1(n12688), .B2(n15595), .A(n12687), .ZN(n12748) );
  MUX2_X1 U14940 ( .A(n12689), .B(n12748), .S(n15611), .Z(n12690) );
  OAI21_X1 U14941 ( .B1(n12751), .B2(n12715), .A(n12690), .ZN(P3_U3479) );
  INV_X1 U14942 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n14632) );
  AOI21_X1 U14943 ( .B1(n12692), .B2(n15595), .A(n12691), .ZN(n12752) );
  MUX2_X1 U14944 ( .A(n14632), .B(n12752), .S(n15611), .Z(n12693) );
  OAI21_X1 U14945 ( .B1(n12715), .B2(n12755), .A(n12693), .ZN(P3_U3478) );
  INV_X1 U14946 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n14659) );
  AOI21_X1 U14947 ( .B1(n12695), .B2(n15595), .A(n12694), .ZN(n12756) );
  MUX2_X1 U14948 ( .A(n14659), .B(n12756), .S(n15611), .Z(n12696) );
  OAI21_X1 U14949 ( .B1(n12759), .B2(n12715), .A(n12696), .ZN(P3_U3477) );
  AOI22_X1 U14950 ( .A1(n12698), .A2(n15595), .B1(n14898), .B2(n12697), .ZN(
        n12699) );
  NAND2_X1 U14951 ( .A1(n12700), .A2(n12699), .ZN(n12760) );
  MUX2_X1 U14952 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12760), .S(n15611), .Z(
        P3_U3476) );
  AND2_X1 U14953 ( .A1(n12701), .A2(n14898), .ZN(n12704) );
  AND2_X1 U14954 ( .A1(n12702), .A2(n15595), .ZN(n12703) );
  MUX2_X1 U14955 ( .A(n12761), .B(P3_REG1_REG_16__SCAN_IN), .S(n15608), .Z(
        P3_U3475) );
  AOI21_X1 U14956 ( .B1(n15595), .B2(n12707), .A(n12706), .ZN(n12762) );
  MUX2_X1 U14957 ( .A(n12708), .B(n12762), .S(n15611), .Z(n12709) );
  OAI21_X1 U14958 ( .B1(n12765), .B2(n12715), .A(n12709), .ZN(P3_U3474) );
  NAND2_X1 U14959 ( .A1(n12710), .A2(n15595), .ZN(n12711) );
  NAND2_X1 U14960 ( .A1(n12712), .A2(n12711), .ZN(n12766) );
  MUX2_X1 U14961 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n12766), .S(n15611), .Z(
        n12713) );
  INV_X1 U14962 ( .A(n12713), .ZN(n12714) );
  OAI21_X1 U14963 ( .B1(n12715), .B2(n12769), .A(n12714), .ZN(P3_U3473) );
  INV_X1 U14964 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12716) );
  NOR2_X1 U14965 ( .A1(n15599), .A2(n12716), .ZN(n12717) );
  AOI21_X1 U14966 ( .B1(n14897), .B2(n15599), .A(n12717), .ZN(n12718) );
  OAI21_X1 U14967 ( .B1(n12719), .B2(n12770), .A(n12718), .ZN(P3_U3458) );
  MUX2_X1 U14968 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n12720), .S(n15599), .Z(
        P3_U3455) );
  MUX2_X1 U14969 ( .A(n12725), .B(n12724), .S(n15599), .Z(n12726) );
  OAI21_X1 U14970 ( .B1(n12727), .B2(n12770), .A(n12726), .ZN(P3_U3453) );
  MUX2_X1 U14971 ( .A(n12729), .B(n12728), .S(n15599), .Z(n12730) );
  OAI21_X1 U14972 ( .B1(n12731), .B2(n12770), .A(n12730), .ZN(P3_U3452) );
  INV_X1 U14973 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12733) );
  MUX2_X1 U14974 ( .A(n12733), .B(n12732), .S(n15599), .Z(n12734) );
  OAI21_X1 U14975 ( .B1(n12735), .B2(n12770), .A(n12734), .ZN(P3_U3451) );
  INV_X1 U14976 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12737) );
  MUX2_X1 U14977 ( .A(n12737), .B(n12736), .S(n15599), .Z(n12738) );
  OAI21_X1 U14978 ( .B1(n12739), .B2(n12770), .A(n12738), .ZN(P3_U3450) );
  INV_X1 U14979 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12741) );
  MUX2_X1 U14980 ( .A(n12741), .B(n12740), .S(n15599), .Z(n12742) );
  OAI21_X1 U14981 ( .B1(n12743), .B2(n12770), .A(n12742), .ZN(P3_U3449) );
  INV_X1 U14982 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12745) );
  MUX2_X1 U14983 ( .A(n12745), .B(n12744), .S(n15599), .Z(n12746) );
  OAI21_X1 U14984 ( .B1(n12747), .B2(n12770), .A(n12746), .ZN(P3_U3448) );
  INV_X1 U14985 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12749) );
  MUX2_X1 U14986 ( .A(n12749), .B(n12748), .S(n15599), .Z(n12750) );
  OAI21_X1 U14987 ( .B1(n12751), .B2(n12770), .A(n12750), .ZN(P3_U3447) );
  INV_X1 U14988 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12753) );
  MUX2_X1 U14989 ( .A(n12753), .B(n12752), .S(n15599), .Z(n12754) );
  OAI21_X1 U14990 ( .B1(n12770), .B2(n12755), .A(n12754), .ZN(P3_U3446) );
  INV_X1 U14991 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12757) );
  MUX2_X1 U14992 ( .A(n12757), .B(n12756), .S(n15599), .Z(n12758) );
  OAI21_X1 U14993 ( .B1(n12759), .B2(n12770), .A(n12758), .ZN(P3_U3444) );
  MUX2_X1 U14994 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12760), .S(n15599), .Z(
        P3_U3441) );
  MUX2_X1 U14995 ( .A(n12761), .B(P3_REG0_REG_16__SCAN_IN), .S(n15601), .Z(
        P3_U3438) );
  INV_X1 U14996 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12763) );
  MUX2_X1 U14997 ( .A(n12763), .B(n12762), .S(n15599), .Z(n12764) );
  OAI21_X1 U14998 ( .B1(n12765), .B2(n12770), .A(n12764), .ZN(P3_U3435) );
  MUX2_X1 U14999 ( .A(n12766), .B(P3_REG0_REG_14__SCAN_IN), .S(n15601), .Z(
        n12767) );
  INV_X1 U15000 ( .A(n12767), .ZN(n12768) );
  OAI21_X1 U15001 ( .B1(n12770), .B2(n12769), .A(n12768), .ZN(P3_U3432) );
  MUX2_X1 U15002 ( .A(P3_D_REG_1__SCAN_IN), .B(n12771), .S(n12772), .Z(
        P3_U3377) );
  MUX2_X1 U15003 ( .A(P3_D_REG_0__SCAN_IN), .B(n12773), .S(n12772), .Z(
        P3_U3376) );
  NAND3_X1 U15004 ( .A1(n12774), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n12776) );
  OAI22_X1 U15005 ( .A1(n8762), .A2(n12776), .B1(n12775), .B2(n12784), .ZN(
        n12777) );
  AOI21_X1 U15006 ( .B1(n12778), .B2(n14780), .A(n12777), .ZN(n12779) );
  INV_X1 U15007 ( .A(n12779), .ZN(P3_U3264) );
  INV_X1 U15008 ( .A(n12780), .ZN(n12782) );
  OAI222_X1 U15009 ( .A1(n12784), .A2(n12783), .B1(n14787), .B2(n12782), .C1(
        n12781), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U15010 ( .A(n13301), .ZN(n13090) );
  INV_X1 U15011 ( .A(n12785), .ZN(n12787) );
  NAND2_X1 U15012 ( .A1(n12787), .A2(n12786), .ZN(n12788) );
  XNOR2_X1 U15013 ( .A(n13364), .B(n12806), .ZN(n12909) );
  NAND2_X1 U15014 ( .A1(n12978), .A2(n12824), .ZN(n12790) );
  XNOR2_X1 U15015 ( .A(n12909), .B(n12790), .ZN(n12894) );
  NAND2_X1 U15016 ( .A1(n12909), .A2(n12790), .ZN(n12791) );
  XNOR2_X1 U15017 ( .A(n13069), .B(n12869), .ZN(n12792) );
  NAND2_X1 U15018 ( .A1(n13065), .A2(n12824), .ZN(n12793) );
  XNOR2_X1 U15019 ( .A(n12792), .B(n12793), .ZN(n12907) );
  INV_X1 U15020 ( .A(n12792), .ZN(n12794) );
  XNOR2_X1 U15021 ( .A(n13353), .B(n12869), .ZN(n12795) );
  AND2_X1 U15022 ( .A1(n13042), .A2(n12824), .ZN(n12796) );
  NAND2_X1 U15023 ( .A1(n12795), .A2(n12796), .ZN(n12799) );
  INV_X1 U15024 ( .A(n12795), .ZN(n12858) );
  INV_X1 U15025 ( .A(n12796), .ZN(n12797) );
  NAND2_X1 U15026 ( .A1(n12858), .A2(n12797), .ZN(n12798) );
  AND2_X1 U15027 ( .A1(n12799), .A2(n12798), .ZN(n12950) );
  XNOR2_X1 U15028 ( .A(n13348), .B(n12869), .ZN(n12929) );
  NAND2_X1 U15029 ( .A1(n13043), .A2(n12824), .ZN(n12801) );
  XNOR2_X1 U15030 ( .A(n12929), .B(n12801), .ZN(n12865) );
  AND2_X1 U15031 ( .A1(n12865), .A2(n12799), .ZN(n12800) );
  INV_X1 U15032 ( .A(n12929), .ZN(n12802) );
  XNOR2_X1 U15033 ( .A(n13343), .B(n12869), .ZN(n12803) );
  NAND2_X1 U15034 ( .A1(n13047), .A2(n12824), .ZN(n12804) );
  XNOR2_X1 U15035 ( .A(n12803), .B(n12804), .ZN(n12930) );
  INV_X1 U15036 ( .A(n12803), .ZN(n12805) );
  XNOR2_X1 U15037 ( .A(n13337), .B(n12806), .ZN(n12807) );
  NAND2_X1 U15038 ( .A1(n13048), .A2(n12824), .ZN(n12808) );
  XNOR2_X1 U15039 ( .A(n12807), .B(n12808), .ZN(n12876) );
  INV_X1 U15040 ( .A(n12807), .ZN(n12810) );
  INV_X1 U15041 ( .A(n12808), .ZN(n12809) );
  NAND2_X1 U15042 ( .A1(n12810), .A2(n12809), .ZN(n12936) );
  XNOR2_X1 U15043 ( .A(n13330), .B(n12806), .ZN(n12938) );
  NAND2_X1 U15044 ( .A1(n12977), .A2(n12824), .ZN(n12941) );
  NAND2_X1 U15045 ( .A1(n12938), .A2(n12941), .ZN(n12812) );
  NAND2_X1 U15046 ( .A1(n12813), .A2(n12812), .ZN(n12816) );
  XNOR2_X1 U15047 ( .A(n13325), .B(n12869), .ZN(n12814) );
  XNOR2_X1 U15048 ( .A(n12816), .B(n12814), .ZN(n12849) );
  NAND2_X1 U15049 ( .A1(n13051), .A2(n12824), .ZN(n12848) );
  NAND2_X1 U15050 ( .A1(n12849), .A2(n12848), .ZN(n12818) );
  INV_X1 U15051 ( .A(n12814), .ZN(n12815) );
  NAND2_X1 U15052 ( .A1(n12816), .A2(n12815), .ZN(n12817) );
  XNOR2_X1 U15053 ( .A(n13318), .B(n12869), .ZN(n12819) );
  AND2_X1 U15054 ( .A1(n13052), .A2(n12824), .ZN(n12820) );
  NAND2_X1 U15055 ( .A1(n12819), .A2(n12820), .ZN(n12823) );
  INV_X1 U15056 ( .A(n12819), .ZN(n12882) );
  INV_X1 U15057 ( .A(n12820), .ZN(n12821) );
  NAND2_X1 U15058 ( .A1(n12882), .A2(n12821), .ZN(n12822) );
  NAND2_X1 U15059 ( .A1(n12823), .A2(n12822), .ZN(n12921) );
  XNOR2_X1 U15060 ( .A(n13313), .B(n12869), .ZN(n12825) );
  AND2_X1 U15061 ( .A1(n13053), .A2(n12824), .ZN(n12826) );
  NAND2_X1 U15062 ( .A1(n12825), .A2(n12826), .ZN(n12829) );
  INV_X1 U15063 ( .A(n12825), .ZN(n12959) );
  INV_X1 U15064 ( .A(n12826), .ZN(n12827) );
  NAND2_X1 U15065 ( .A1(n12959), .A2(n12827), .ZN(n12828) );
  AND2_X1 U15066 ( .A1(n12829), .A2(n12828), .ZN(n12880) );
  XNOR2_X1 U15067 ( .A(n13307), .B(n12869), .ZN(n12831) );
  NAND2_X1 U15068 ( .A1(n13087), .A2(n12824), .ZN(n12832) );
  XNOR2_X1 U15069 ( .A(n12831), .B(n12832), .ZN(n12974) );
  AND2_X1 U15070 ( .A1(n12974), .A2(n12829), .ZN(n12830) );
  NAND2_X1 U15071 ( .A1(n12883), .A2(n12830), .ZN(n12969) );
  INV_X1 U15072 ( .A(n12831), .ZN(n12833) );
  NAND2_X1 U15073 ( .A1(n12833), .A2(n12832), .ZN(n12834) );
  XNOR2_X1 U15074 ( .A(n13301), .B(n12869), .ZN(n12835) );
  AND2_X1 U15075 ( .A1(n13089), .A2(n12824), .ZN(n12836) );
  NAND2_X1 U15076 ( .A1(n12835), .A2(n12836), .ZN(n12867) );
  INV_X1 U15077 ( .A(n12835), .ZN(n12838) );
  INV_X1 U15078 ( .A(n12836), .ZN(n12837) );
  NAND2_X1 U15079 ( .A1(n12838), .A2(n12837), .ZN(n12839) );
  NAND2_X1 U15080 ( .A1(n12867), .A2(n12839), .ZN(n12841) );
  AOI21_X1 U15081 ( .B1(n12840), .B2(n12841), .A(n12968), .ZN(n12842) );
  NAND2_X1 U15082 ( .A1(n12842), .A2(n12868), .ZN(n12847) );
  OAI22_X1 U15083 ( .A1(n13058), .A2(n13031), .B1(n13088), .B2(n12916), .ZN(
        n13123) );
  INV_X1 U15084 ( .A(n13129), .ZN(n12844) );
  OAI22_X1 U15085 ( .A1(n12844), .A2(n12928), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12843), .ZN(n12845) );
  AOI21_X1 U15086 ( .B1(n13123), .B2(n12925), .A(n12845), .ZN(n12846) );
  OAI211_X1 U15087 ( .C1(n13090), .C2(n12957), .A(n12847), .B(n12846), .ZN(
        P2_U3186) );
  INV_X1 U15088 ( .A(n13325), .ZN(n13190) );
  NAND2_X1 U15089 ( .A1(n13051), .A2(n12940), .ZN(n12851) );
  NAND2_X1 U15090 ( .A1(n12848), .A2(n12961), .ZN(n12850) );
  MUX2_X1 U15091 ( .A(n12851), .B(n12850), .S(n12849), .Z(n12857) );
  INV_X1 U15092 ( .A(n13188), .ZN(n12855) );
  AND2_X1 U15093 ( .A1(n12977), .A2(n13095), .ZN(n12852) );
  AOI21_X1 U15094 ( .B1(n13052), .B2(n12963), .A(n12852), .ZN(n13323) );
  OAI22_X1 U15095 ( .A1(n13323), .A2(n12967), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12853), .ZN(n12854) );
  AOI21_X1 U15096 ( .B1(n12855), .B2(n12965), .A(n12854), .ZN(n12856) );
  OAI211_X1 U15097 ( .C1(n13190), .C2(n12957), .A(n12857), .B(n12856), .ZN(
        P2_U3188) );
  INV_X1 U15098 ( .A(n12949), .ZN(n12860) );
  NOR3_X1 U15099 ( .A1(n12858), .A2(n13071), .A3(n12958), .ZN(n12859) );
  AOI21_X1 U15100 ( .B1(n12860), .B2(n12961), .A(n12859), .ZN(n12866) );
  AND2_X1 U15101 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13027) );
  AOI22_X1 U15102 ( .A1(n13047), .A2(n12963), .B1(n13095), .B2(n13042), .ZN(
        n13246) );
  NOR2_X1 U15103 ( .A1(n13246), .A2(n12967), .ZN(n12861) );
  AOI211_X1 U15104 ( .C1(n12965), .C2(n13249), .A(n13027), .B(n12861), .ZN(
        n12862) );
  OAI21_X1 U15105 ( .B1(n7533), .B2(n12957), .A(n12862), .ZN(n12863) );
  AOI21_X1 U15106 ( .B1(n6727), .B2(n12961), .A(n12863), .ZN(n12864) );
  OAI21_X1 U15107 ( .B1(n12866), .B2(n12865), .A(n12864), .ZN(P2_U3191) );
  AOI22_X1 U15108 ( .A1(n12976), .A2(n12963), .B1(n13095), .B2(n13089), .ZN(
        n13111) );
  INV_X1 U15109 ( .A(n12824), .ZN(n13117) );
  NOR2_X1 U15110 ( .A1(n13058), .A2(n13117), .ZN(n12870) );
  INV_X1 U15111 ( .A(n12871), .ZN(n13116) );
  AOI22_X1 U15112 ( .A1(n13116), .A2(n12965), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12872) );
  INV_X1 U15113 ( .A(n12977), .ZN(n13081) );
  OAI22_X1 U15114 ( .A1(n13081), .A2(n13031), .B1(n13044), .B2(n12916), .ZN(
        n13215) );
  AOI22_X1 U15115 ( .A1(n13215), .A2(n12925), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12873) );
  OAI21_X1 U15116 ( .B1(n13219), .B2(n12928), .A(n12873), .ZN(n12878) );
  INV_X1 U15117 ( .A(n12937), .ZN(n12874) );
  AOI211_X1 U15118 ( .C1(n12876), .C2(n12875), .A(n12968), .B(n12874), .ZN(
        n12877) );
  AOI211_X1 U15119 ( .C1(n13337), .C2(n12972), .A(n12878), .B(n12877), .ZN(
        n12879) );
  INV_X1 U15120 ( .A(n12879), .ZN(P2_U3195) );
  INV_X1 U15121 ( .A(n13313), .ZN(n13054) );
  INV_X1 U15122 ( .A(n12880), .ZN(n12881) );
  AOI21_X1 U15123 ( .B1(n12918), .B2(n12881), .A(n12968), .ZN(n12885) );
  NOR3_X1 U15124 ( .A1(n12882), .A2(n12886), .A3(n12958), .ZN(n12884) );
  OAI21_X1 U15125 ( .B1(n12885), .B2(n12884), .A(n12883), .ZN(n12891) );
  OAI22_X1 U15126 ( .A1(n13088), .A2(n13031), .B1(n12886), .B2(n12916), .ZN(
        n13156) );
  INV_X1 U15127 ( .A(n13162), .ZN(n12888) );
  OAI22_X1 U15128 ( .A1(n12888), .A2(n12928), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12887), .ZN(n12889) );
  AOI21_X1 U15129 ( .B1(n13156), .B2(n12925), .A(n12889), .ZN(n12890) );
  OAI211_X1 U15130 ( .C1(n13054), .C2(n12957), .A(n12891), .B(n12890), .ZN(
        P2_U3197) );
  INV_X1 U15131 ( .A(n12912), .ZN(n12892) );
  AOI21_X1 U15132 ( .B1(n12894), .B2(n12893), .A(n12892), .ZN(n12901) );
  NAND2_X1 U15133 ( .A1(n12925), .A2(n12895), .ZN(n12896) );
  OAI211_X1 U15134 ( .C1(n12928), .C2(n12898), .A(n12897), .B(n12896), .ZN(
        n12899) );
  AOI21_X1 U15135 ( .B1(n13364), .B2(n12972), .A(n12899), .ZN(n12900) );
  OAI21_X1 U15136 ( .B1(n12901), .B2(n12968), .A(n12900), .ZN(P2_U3198) );
  OAI22_X1 U15137 ( .A1(n12903), .A2(n12967), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12902), .ZN(n12905) );
  NOR2_X1 U15138 ( .A1(n13358), .A2(n12957), .ZN(n12904) );
  AOI211_X1 U15139 ( .C1(n12965), .C2(n12906), .A(n12905), .B(n12904), .ZN(
        n12914) );
  INV_X1 U15140 ( .A(n12907), .ZN(n12911) );
  OAI22_X1 U15141 ( .A1(n12909), .A2(n12968), .B1(n12908), .B2(n12958), .ZN(
        n12910) );
  NAND3_X1 U15142 ( .A1(n12912), .A2(n12911), .A3(n12910), .ZN(n12913) );
  OAI211_X1 U15143 ( .C1(n12915), .C2(n12968), .A(n12914), .B(n12913), .ZN(
        P2_U3200) );
  INV_X1 U15144 ( .A(n13051), .ZN(n13083) );
  OAI22_X1 U15145 ( .A1(n13086), .A2(n13031), .B1(n13083), .B2(n12916), .ZN(
        n13171) );
  AOI22_X1 U15146 ( .A1(n13171), .A2(n12925), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12917) );
  OAI21_X1 U15147 ( .B1(n13177), .B2(n12928), .A(n12917), .ZN(n12923) );
  INV_X1 U15148 ( .A(n12918), .ZN(n12919) );
  AOI211_X1 U15149 ( .C1(n12921), .C2(n12920), .A(n12968), .B(n12919), .ZN(
        n12922) );
  AOI211_X1 U15150 ( .C1(n13318), .C2(n12972), .A(n12923), .B(n12922), .ZN(
        n12924) );
  INV_X1 U15151 ( .A(n12924), .ZN(P2_U3201) );
  AOI22_X1 U15152 ( .A1(n13048), .A2(n12963), .B1(n13095), .B2(n13043), .ZN(
        n13232) );
  INV_X1 U15153 ( .A(n13232), .ZN(n12926) );
  AOI22_X1 U15154 ( .A1(n12926), .A2(n12925), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12927) );
  OAI21_X1 U15155 ( .B1(n13237), .B2(n12928), .A(n12927), .ZN(n12933) );
  AOI22_X1 U15156 ( .A1(n12929), .A2(n12961), .B1(n12940), .B2(n13043), .ZN(
        n12931) );
  NOR3_X1 U15157 ( .A1(n6727), .A2(n12931), .A3(n12930), .ZN(n12932) );
  AOI211_X1 U15158 ( .C1(n13343), .C2(n12972), .A(n12933), .B(n12932), .ZN(
        n12934) );
  OAI21_X1 U15159 ( .B1(n12935), .B2(n12968), .A(n12934), .ZN(P2_U3205) );
  NAND2_X1 U15160 ( .A1(n12937), .A2(n12936), .ZN(n12939) );
  XNOR2_X1 U15161 ( .A(n12939), .B(n12938), .ZN(n12948) );
  NAND2_X1 U15162 ( .A1(n12977), .A2(n12940), .ZN(n12947) );
  NAND3_X1 U15163 ( .A1(n12948), .A2(n12961), .A3(n12941), .ZN(n12946) );
  AOI22_X1 U15164 ( .A1(n13051), .A2(n12963), .B1(n13095), .B2(n13048), .ZN(
        n13198) );
  OAI22_X1 U15165 ( .A1(n13198), .A2(n12967), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12942), .ZN(n12944) );
  INV_X1 U15166 ( .A(n13330), .ZN(n13050) );
  NOR2_X1 U15167 ( .A1(n13050), .A2(n12957), .ZN(n12943) );
  AOI211_X1 U15168 ( .C1(n12965), .C2(n13203), .A(n12944), .B(n12943), .ZN(
        n12945) );
  OAI211_X1 U15169 ( .C1(n12948), .C2(n12947), .A(n12946), .B(n12945), .ZN(
        P2_U3207) );
  INV_X1 U15170 ( .A(n13353), .ZN(n13278) );
  OAI211_X1 U15171 ( .C1(n12951), .C2(n12950), .A(n12949), .B(n12961), .ZN(
        n12956) );
  INV_X1 U15172 ( .A(n12952), .ZN(n13274) );
  AOI22_X1 U15173 ( .A1(n13043), .A2(n12963), .B1(n13095), .B2(n13065), .ZN(
        n13262) );
  OAI22_X1 U15174 ( .A1(n13262), .A2(n12967), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12953), .ZN(n12954) );
  AOI21_X1 U15175 ( .B1(n13274), .B2(n12965), .A(n12954), .ZN(n12955) );
  OAI211_X1 U15176 ( .C1(n13278), .C2(n12957), .A(n12956), .B(n12955), .ZN(
        P2_U3210) );
  INV_X1 U15177 ( .A(n12883), .ZN(n12962) );
  NOR3_X1 U15178 ( .A1(n12959), .A2(n13086), .A3(n12958), .ZN(n12960) );
  AOI21_X1 U15179 ( .B1(n12962), .B2(n12961), .A(n12960), .ZN(n12975) );
  AOI22_X1 U15180 ( .A1(n13089), .A2(n12963), .B1(n13095), .B2(n13053), .ZN(
        n13138) );
  INV_X1 U15181 ( .A(n12964), .ZN(n13144) );
  AOI22_X1 U15182 ( .A1(n13144), .A2(n12965), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12966) );
  OAI21_X1 U15183 ( .B1(n13138), .B2(n12967), .A(n12966), .ZN(n12971) );
  NOR2_X1 U15184 ( .A1(n12969), .A2(n12968), .ZN(n12970) );
  AOI211_X1 U15185 ( .C1(n13307), .C2(n12972), .A(n12971), .B(n12970), .ZN(
        n12973) );
  OAI21_X1 U15186 ( .B1(n12975), .B2(n12974), .A(n12973), .ZN(P2_U3212) );
  MUX2_X1 U15187 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13033), .S(n12993), .Z(
        P2_U3562) );
  MUX2_X1 U15188 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13097), .S(n12993), .Z(
        P2_U3561) );
  MUX2_X1 U15189 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n12976), .S(n12993), .Z(
        P2_U3560) );
  MUX2_X1 U15190 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13096), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15191 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13089), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15192 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13087), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15193 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13053), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15194 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13052), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15195 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13051), .S(n12993), .Z(
        P2_U3554) );
  MUX2_X1 U15196 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n12977), .S(n12993), .Z(
        P2_U3553) );
  MUX2_X1 U15197 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13048), .S(n12993), .Z(
        P2_U3552) );
  MUX2_X1 U15198 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13047), .S(n12993), .Z(
        P2_U3551) );
  MUX2_X1 U15199 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13043), .S(n12993), .Z(
        P2_U3550) );
  MUX2_X1 U15200 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13042), .S(n12993), .Z(
        P2_U3549) );
  MUX2_X1 U15201 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13065), .S(n12993), .Z(
        P2_U3548) );
  MUX2_X1 U15202 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n12978), .S(n12993), .Z(
        P2_U3547) );
  MUX2_X1 U15203 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n12979), .S(n12993), .Z(
        P2_U3546) );
  MUX2_X1 U15204 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n12980), .S(n12993), .Z(
        P2_U3545) );
  MUX2_X1 U15205 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n12981), .S(n12993), .Z(
        P2_U3544) );
  MUX2_X1 U15206 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n12982), .S(n12993), .Z(
        P2_U3543) );
  MUX2_X1 U15207 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n12983), .S(n12993), .Z(
        P2_U3542) );
  MUX2_X1 U15208 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n12984), .S(n12993), .Z(
        P2_U3541) );
  MUX2_X1 U15209 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n12985), .S(n12993), .Z(
        P2_U3540) );
  MUX2_X1 U15210 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n12986), .S(n12993), .Z(
        P2_U3539) );
  MUX2_X1 U15211 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n12987), .S(n12993), .Z(
        P2_U3538) );
  MUX2_X1 U15212 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n12988), .S(n12993), .Z(
        P2_U3537) );
  MUX2_X1 U15213 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n12989), .S(n12993), .Z(
        P2_U3536) );
  MUX2_X1 U15214 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n12990), .S(n12993), .Z(
        P2_U3535) );
  MUX2_X1 U15215 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n12991), .S(n12993), .Z(
        P2_U3534) );
  MUX2_X1 U15216 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n12992), .S(n12993), .Z(
        P2_U3533) );
  MUX2_X1 U15217 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n12994), .S(n12993), .Z(
        P2_U3532) );
  NOR2_X1 U15218 ( .A1(n15262), .A2(n13001), .ZN(n12995) );
  AOI211_X1 U15219 ( .C1(n15299), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n12996), .B(
        n12995), .ZN(n13008) );
  MUX2_X1 U15220 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9630), .S(n13001), .Z(
        n12997) );
  NAND3_X1 U15221 ( .A1(n15233), .A2(n12998), .A3(n12997), .ZN(n12999) );
  NAND3_X1 U15222 ( .A1(n13000), .A2(n15300), .A3(n12999), .ZN(n13007) );
  MUX2_X1 U15223 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10484), .S(n13001), .Z(
        n13002) );
  NAND3_X1 U15224 ( .A1(n15236), .A2(n13003), .A3(n13002), .ZN(n13004) );
  NAND3_X1 U15225 ( .A1(n13005), .A2(n15306), .A3(n13004), .ZN(n13006) );
  NAND3_X1 U15226 ( .A1(n13008), .A2(n13007), .A3(n13006), .ZN(P2_U3222) );
  NOR2_X1 U15227 ( .A1(n13014), .A2(n13009), .ZN(n13010) );
  NOR2_X1 U15228 ( .A1(n13011), .A2(n13010), .ZN(n13012) );
  XOR2_X1 U15229 ( .A(n13012), .B(n13253), .Z(n13023) );
  NAND2_X1 U15230 ( .A1(n13014), .A2(n13013), .ZN(n13015) );
  NAND2_X1 U15231 ( .A1(n13016), .A2(n13015), .ZN(n13018) );
  XOR2_X1 U15232 ( .A(n13018), .B(n13017), .Z(n13020) );
  OAI22_X1 U15233 ( .A1(n13023), .A2(n15270), .B1(n13020), .B2(n15265), .ZN(
        n13019) );
  INV_X1 U15234 ( .A(n13019), .ZN(n13026) );
  NAND2_X1 U15235 ( .A1(n13020), .A2(n15300), .ZN(n13021) );
  NAND2_X1 U15236 ( .A1(n13021), .A2(n15262), .ZN(n13022) );
  AOI21_X1 U15237 ( .B1(n13023), .B2(n15306), .A(n13022), .ZN(n13025) );
  MUX2_X1 U15238 ( .A(n13026), .B(n13025), .S(n13024), .Z(n13029) );
  AOI21_X1 U15239 ( .B1(n15299), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n13027), 
        .ZN(n13028) );
  NAND2_X1 U15240 ( .A1(n13029), .A2(n13028), .ZN(P2_U3233) );
  NAND2_X1 U15241 ( .A1(n13200), .A2(n13190), .ZN(n13189) );
  NAND2_X1 U15242 ( .A1(n13059), .A2(n13287), .ZN(n13036) );
  XNOR2_X1 U15243 ( .A(n13036), .B(n13284), .ZN(n13030) );
  AOI21_X1 U15244 ( .B1(n13032), .B2(P2_B_REG_SCAN_IN), .A(n13031), .ZN(n13098) );
  NAND2_X1 U15245 ( .A1(n13098), .A2(n13033), .ZN(n13285) );
  NOR2_X1 U15246 ( .A1(n13282), .A2(n13285), .ZN(n13038) );
  NOR2_X1 U15247 ( .A1(n13284), .A2(n13277), .ZN(n13034) );
  AOI211_X1 U15248 ( .C1(n13282), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13038), 
        .B(n13034), .ZN(n13035) );
  OAI21_X1 U15249 ( .B1(n13283), .B2(n13206), .A(n13035), .ZN(P2_U3234) );
  OAI211_X1 U15250 ( .C1(n13059), .C2(n13287), .A(n13294), .B(n13036), .ZN(
        n13286) );
  NOR2_X1 U15251 ( .A1(n13252), .A2(n13037), .ZN(n13039) );
  AOI211_X1 U15252 ( .C1(n13040), .C2(n13240), .A(n13039), .B(n13038), .ZN(
        n13041) );
  OAI21_X1 U15253 ( .B1(n13286), .B2(n13206), .A(n13041), .ZN(P2_U3235) );
  INV_X1 U15254 ( .A(n13089), .ZN(n13056) );
  INV_X1 U15255 ( .A(n13343), .ZN(n13045) );
  OAI21_X1 U15256 ( .B1(n13047), .B2(n13343), .A(n13046), .ZN(n13223) );
  INV_X1 U15257 ( .A(n13222), .ZN(n13049) );
  INV_X1 U15258 ( .A(n13048), .ZN(n13078) );
  INV_X1 U15259 ( .A(n13196), .ZN(n13208) );
  INV_X1 U15260 ( .A(n13057), .ZN(n13110) );
  NAND2_X1 U15261 ( .A1(n13106), .A2(n13110), .ZN(n13105) );
  AOI211_X1 U15262 ( .C1(n13289), .C2(n13115), .A(n13270), .B(n13059), .ZN(
        n13288) );
  INV_X1 U15263 ( .A(n13060), .ZN(n13061) );
  AOI22_X1 U15264 ( .A1(n13061), .A2(n13273), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13282), .ZN(n13062) );
  OAI21_X1 U15265 ( .B1(n13063), .B2(n13277), .A(n13062), .ZN(n13064) );
  AOI21_X1 U15266 ( .B1(n13288), .B2(n13272), .A(n13064), .ZN(n13104) );
  INV_X1 U15267 ( .A(n13065), .ZN(n13068) );
  NOR2_X1 U15268 ( .A1(n13069), .A2(n13068), .ZN(n13066) );
  OR2_X1 U15269 ( .A1(n13353), .A2(n13071), .ZN(n13070) );
  NAND2_X1 U15270 ( .A1(n13261), .A2(n13070), .ZN(n13073) );
  NAND2_X1 U15271 ( .A1(n13353), .A2(n13071), .ZN(n13072) );
  AND2_X1 U15272 ( .A1(n13348), .A2(n13075), .ZN(n13074) );
  OR2_X1 U15273 ( .A1(n13348), .A2(n13075), .ZN(n13076) );
  OR2_X1 U15274 ( .A1(n13337), .A2(n13078), .ZN(n13079) );
  OR2_X1 U15275 ( .A1(n13330), .A2(n13081), .ZN(n13082) );
  NOR2_X1 U15276 ( .A1(n13109), .A2(n13110), .ZN(n13108) );
  NOR2_X1 U15277 ( .A1(n13108), .A2(n13091), .ZN(n13094) );
  NAND2_X1 U15278 ( .A1(n13096), .A2(n13095), .ZN(n13100) );
  INV_X1 U15279 ( .A(n13290), .ZN(n13102) );
  NAND2_X1 U15280 ( .A1(n13102), .A2(n13252), .ZN(n13103) );
  OAI211_X1 U15281 ( .C1(n13291), .C2(n13256), .A(n13104), .B(n13103), .ZN(
        P2_U3236) );
  OAI21_X1 U15282 ( .B1(n13106), .B2(n13110), .A(n13105), .ZN(n13298) );
  AOI22_X1 U15283 ( .A1(n13107), .A2(n13240), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n13282), .ZN(n13121) );
  AOI211_X1 U15284 ( .C1(n13110), .C2(n13109), .A(n13247), .B(n13108), .ZN(
        n13113) );
  INV_X1 U15285 ( .A(n13111), .ZN(n13112) );
  NOR2_X1 U15286 ( .A1(n13113), .A2(n13112), .ZN(n13297) );
  OR2_X1 U15287 ( .A1(n13292), .A2(n13126), .ZN(n13114) );
  AND2_X1 U15288 ( .A1(n13115), .A2(n13114), .ZN(n13295) );
  AOI22_X1 U15289 ( .A1(n13295), .A2(n13117), .B1(n13116), .B2(n13273), .ZN(
        n13118) );
  AOI21_X1 U15290 ( .B1(n13297), .B2(n13118), .A(n13282), .ZN(n13119) );
  INV_X1 U15291 ( .A(n13119), .ZN(n13120) );
  OAI211_X1 U15292 ( .C1(n13298), .C2(n13256), .A(n13121), .B(n13120), .ZN(
        P2_U3237) );
  XNOR2_X1 U15293 ( .A(n13122), .B(n13127), .ZN(n13124) );
  AOI21_X1 U15294 ( .B1(n13124), .B2(n13264), .A(n13123), .ZN(n13304) );
  AND2_X1 U15295 ( .A1(n13301), .A2(n13141), .ZN(n13125) );
  OR3_X1 U15296 ( .A1(n13126), .A2(n13125), .A3(n13270), .ZN(n13303) );
  OR2_X1 U15297 ( .A1(n13128), .A2(n13127), .ZN(n13300) );
  NAND3_X1 U15298 ( .A1(n13300), .A2(n13299), .A3(n13280), .ZN(n13134) );
  NAND2_X1 U15299 ( .A1(n13129), .A2(n13273), .ZN(n13130) );
  OAI21_X1 U15300 ( .B1(n13252), .B2(n13131), .A(n13130), .ZN(n13132) );
  AOI21_X1 U15301 ( .B1(n13301), .B2(n13240), .A(n13132), .ZN(n13133) );
  OAI211_X1 U15302 ( .C1(n13303), .C2(n13206), .A(n13134), .B(n13133), .ZN(
        n13135) );
  INV_X1 U15303 ( .A(n13135), .ZN(n13136) );
  OAI21_X1 U15304 ( .B1(n13282), .B2(n13304), .A(n13136), .ZN(P2_U3238) );
  XOR2_X1 U15305 ( .A(n13148), .B(n13137), .Z(n13140) );
  INV_X1 U15306 ( .A(n13138), .ZN(n13139) );
  AOI21_X1 U15307 ( .B1(n13140), .B2(n13264), .A(n13139), .ZN(n13309) );
  INV_X1 U15308 ( .A(n13161), .ZN(n13143) );
  INV_X1 U15309 ( .A(n13141), .ZN(n13142) );
  AOI211_X1 U15310 ( .C1(n13307), .C2(n13143), .A(n13270), .B(n13142), .ZN(
        n13306) );
  AOI22_X1 U15311 ( .A1(n13144), .A2(n13273), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13282), .ZN(n13145) );
  OAI21_X1 U15312 ( .B1(n13146), .B2(n13277), .A(n13145), .ZN(n13150) );
  XOR2_X1 U15313 ( .A(n13148), .B(n13147), .Z(n13310) );
  NOR2_X1 U15314 ( .A1(n13310), .A2(n13256), .ZN(n13149) );
  AOI211_X1 U15315 ( .C1(n13306), .C2(n13272), .A(n13150), .B(n13149), .ZN(
        n13151) );
  OAI21_X1 U15316 ( .B1(n13282), .B2(n13309), .A(n13151), .ZN(P2_U3239) );
  XOR2_X1 U15317 ( .A(n13154), .B(n13152), .Z(n13315) );
  AOI21_X1 U15318 ( .B1(n13155), .B2(n13154), .A(n13153), .ZN(n13158) );
  INV_X1 U15319 ( .A(n13156), .ZN(n13157) );
  OAI21_X1 U15320 ( .B1(n13158), .B2(n13247), .A(n13157), .ZN(n13311) );
  NAND2_X1 U15321 ( .A1(n13313), .A2(n6602), .ZN(n13159) );
  NAND2_X1 U15322 ( .A1(n13159), .A2(n13294), .ZN(n13160) );
  NOR2_X1 U15323 ( .A1(n13161), .A2(n13160), .ZN(n13312) );
  NAND2_X1 U15324 ( .A1(n13312), .A2(n13272), .ZN(n13167) );
  NAND2_X1 U15325 ( .A1(n13162), .A2(n13273), .ZN(n13163) );
  OAI21_X1 U15326 ( .B1(n13252), .B2(n13164), .A(n13163), .ZN(n13165) );
  AOI21_X1 U15327 ( .B1(n13313), .B2(n13240), .A(n13165), .ZN(n13166) );
  NAND2_X1 U15328 ( .A1(n13167), .A2(n13166), .ZN(n13168) );
  AOI21_X1 U15329 ( .B1(n13311), .B2(n13252), .A(n13168), .ZN(n13169) );
  OAI21_X1 U15330 ( .B1(n13315), .B2(n13256), .A(n13169), .ZN(P2_U3240) );
  OAI21_X1 U15331 ( .B1(n6658), .B2(n7346), .A(n13170), .ZN(n13172) );
  AOI21_X1 U15332 ( .B1(n13172), .B2(n13264), .A(n13171), .ZN(n13320) );
  AOI21_X1 U15333 ( .B1(n7346), .B2(n13174), .A(n13173), .ZN(n13316) );
  AOI21_X1 U15334 ( .B1(n13318), .B2(n13189), .A(n13270), .ZN(n13175) );
  AND2_X1 U15335 ( .A1(n13175), .A2(n6602), .ZN(n13317) );
  NAND2_X1 U15336 ( .A1(n13317), .A2(n13272), .ZN(n13180) );
  OAI22_X1 U15337 ( .A1(n13177), .A2(n13236), .B1(n13176), .B2(n13252), .ZN(
        n13178) );
  AOI21_X1 U15338 ( .B1(n13318), .B2(n13240), .A(n13178), .ZN(n13179) );
  NAND2_X1 U15339 ( .A1(n13180), .A2(n13179), .ZN(n13181) );
  AOI21_X1 U15340 ( .B1(n13316), .B2(n13280), .A(n13181), .ZN(n13182) );
  OAI21_X1 U15341 ( .B1(n13282), .B2(n13320), .A(n13182), .ZN(P2_U3241) );
  XNOR2_X1 U15342 ( .A(n13183), .B(n13184), .ZN(n13322) );
  INV_X1 U15343 ( .A(n13322), .ZN(n13195) );
  INV_X1 U15344 ( .A(n13184), .ZN(n13185) );
  XNOR2_X1 U15345 ( .A(n13186), .B(n13185), .ZN(n13187) );
  NAND2_X1 U15346 ( .A1(n13187), .A2(n13264), .ZN(n13327) );
  OAI211_X1 U15347 ( .C1(n13236), .C2(n13188), .A(n13327), .B(n13323), .ZN(
        n13193) );
  OAI211_X1 U15348 ( .C1(n13200), .C2(n13190), .A(n13294), .B(n13189), .ZN(
        n13326) );
  AOI22_X1 U15349 ( .A1(n13325), .A2(n13240), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n13282), .ZN(n13191) );
  OAI21_X1 U15350 ( .B1(n13326), .B2(n13206), .A(n13191), .ZN(n13192) );
  AOI21_X1 U15351 ( .B1(n13193), .B2(n13252), .A(n13192), .ZN(n13194) );
  OAI21_X1 U15352 ( .B1(n13195), .B2(n13256), .A(n13194), .ZN(P2_U3242) );
  XNOR2_X1 U15353 ( .A(n13197), .B(n13196), .ZN(n13199) );
  OAI21_X1 U15354 ( .B1(n13199), .B2(n13247), .A(n13198), .ZN(n13334) );
  INV_X1 U15355 ( .A(n13200), .ZN(n13202) );
  AOI21_X1 U15356 ( .B1(n13217), .B2(n13330), .A(n13270), .ZN(n13201) );
  NAND2_X1 U15357 ( .A1(n13202), .A2(n13201), .ZN(n13332) );
  AOI22_X1 U15358 ( .A1(n13282), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13203), 
        .B2(n13273), .ZN(n13205) );
  NAND2_X1 U15359 ( .A1(n13330), .A2(n13240), .ZN(n13204) );
  OAI211_X1 U15360 ( .C1(n13332), .C2(n13206), .A(n13205), .B(n13204), .ZN(
        n13211) );
  OAI21_X1 U15361 ( .B1(n13209), .B2(n13208), .A(n13207), .ZN(n13333) );
  NOR2_X1 U15362 ( .A1(n13333), .A2(n13256), .ZN(n13210) );
  AOI211_X1 U15363 ( .C1(n13252), .C2(n13334), .A(n13211), .B(n13210), .ZN(
        n13212) );
  INV_X1 U15364 ( .A(n13212), .ZN(P2_U3243) );
  OR2_X1 U15365 ( .A1(n13230), .A2(n13231), .ZN(n13228) );
  NAND2_X1 U15366 ( .A1(n13228), .A2(n13213), .ZN(n13214) );
  XNOR2_X1 U15367 ( .A(n13214), .B(n13222), .ZN(n13216) );
  AOI21_X1 U15368 ( .B1(n13216), .B2(n13264), .A(n13215), .ZN(n13339) );
  INV_X1 U15369 ( .A(n13217), .ZN(n13218) );
  AOI211_X1 U15370 ( .C1(n13337), .C2(n13234), .A(n13270), .B(n13218), .ZN(
        n13336) );
  INV_X1 U15371 ( .A(n13219), .ZN(n13220) );
  AOI22_X1 U15372 ( .A1(n13282), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13220), 
        .B2(n13273), .ZN(n13221) );
  OAI21_X1 U15373 ( .B1(n7531), .B2(n13277), .A(n13221), .ZN(n13225) );
  XNOR2_X1 U15374 ( .A(n13223), .B(n13222), .ZN(n13340) );
  NOR2_X1 U15375 ( .A1(n13340), .A2(n13256), .ZN(n13224) );
  AOI211_X1 U15376 ( .C1(n13336), .C2(n13272), .A(n13225), .B(n13224), .ZN(
        n13226) );
  OAI21_X1 U15377 ( .B1(n13282), .B2(n13339), .A(n13226), .ZN(P2_U3244) );
  XOR2_X1 U15378 ( .A(n13231), .B(n13227), .Z(n13345) );
  INV_X1 U15379 ( .A(n13228), .ZN(n13229) );
  AOI21_X1 U15380 ( .B1(n13231), .B2(n13230), .A(n13229), .ZN(n13233) );
  OAI21_X1 U15381 ( .B1(n13233), .B2(n13247), .A(n13232), .ZN(n13341) );
  AOI21_X1 U15382 ( .B1(n13343), .B2(n13250), .A(n13270), .ZN(n13235) );
  AND2_X1 U15383 ( .A1(n13235), .A2(n13234), .ZN(n13342) );
  NAND2_X1 U15384 ( .A1(n13342), .A2(n13272), .ZN(n13242) );
  OAI22_X1 U15385 ( .A1(n13252), .A2(n13238), .B1(n13237), .B2(n13236), .ZN(
        n13239) );
  AOI21_X1 U15386 ( .B1(n13343), .B2(n13240), .A(n13239), .ZN(n13241) );
  NAND2_X1 U15387 ( .A1(n13242), .A2(n13241), .ZN(n13243) );
  AOI21_X1 U15388 ( .B1(n13341), .B2(n13252), .A(n13243), .ZN(n13244) );
  OAI21_X1 U15389 ( .B1(n13345), .B2(n13256), .A(n13244), .ZN(P2_U3245) );
  XNOR2_X1 U15390 ( .A(n13245), .B(n13255), .ZN(n13248) );
  OAI21_X1 U15391 ( .B1(n13248), .B2(n13247), .A(n13246), .ZN(n13346) );
  AOI21_X1 U15392 ( .B1(n13249), .B2(n13273), .A(n13346), .ZN(n13260) );
  INV_X1 U15393 ( .A(n13250), .ZN(n13251) );
  AOI211_X1 U15394 ( .C1(n13348), .C2(n13269), .A(n13270), .B(n13251), .ZN(
        n13347) );
  OAI22_X1 U15395 ( .A1(n7533), .A2(n13277), .B1(n13253), .B2(n13252), .ZN(
        n13258) );
  XOR2_X1 U15396 ( .A(n13255), .B(n13254), .Z(n13350) );
  NOR2_X1 U15397 ( .A1(n13350), .A2(n13256), .ZN(n13257) );
  AOI211_X1 U15398 ( .C1(n13347), .C2(n13272), .A(n13258), .B(n13257), .ZN(
        n13259) );
  OAI21_X1 U15399 ( .B1(n13282), .B2(n13260), .A(n13259), .ZN(P2_U3246) );
  XOR2_X1 U15400 ( .A(n13261), .B(n13267), .Z(n13265) );
  INV_X1 U15401 ( .A(n13262), .ZN(n13263) );
  AOI21_X1 U15402 ( .B1(n13265), .B2(n13264), .A(n13263), .ZN(n13355) );
  OAI21_X1 U15403 ( .B1(n13268), .B2(n13267), .A(n13266), .ZN(n13351) );
  AOI211_X1 U15404 ( .C1(n13353), .C2(n13271), .A(n13270), .B(n7534), .ZN(
        n13352) );
  NAND2_X1 U15405 ( .A1(n13352), .A2(n13272), .ZN(n13276) );
  AOI22_X1 U15406 ( .A1(n13282), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13274), 
        .B2(n13273), .ZN(n13275) );
  OAI211_X1 U15407 ( .C1(n13278), .C2(n13277), .A(n13276), .B(n13275), .ZN(
        n13279) );
  AOI21_X1 U15408 ( .B1(n13351), .B2(n13280), .A(n13279), .ZN(n13281) );
  OAI21_X1 U15409 ( .B1(n13282), .B2(n13355), .A(n13281), .ZN(P2_U3247) );
  OAI211_X1 U15410 ( .C1(n13284), .C2(n15376), .A(n13283), .B(n13285), .ZN(
        n13378) );
  MUX2_X1 U15411 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13378), .S(n15392), .Z(
        P2_U3530) );
  OAI211_X1 U15412 ( .C1(n13287), .C2(n15376), .A(n13286), .B(n13285), .ZN(
        n13379) );
  MUX2_X1 U15413 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13379), .S(n15392), .Z(
        P2_U3529) );
  NOR2_X1 U15414 ( .A1(n13292), .A2(n15376), .ZN(n13293) );
  AOI21_X1 U15415 ( .B1(n13295), .B2(n13294), .A(n13293), .ZN(n13296) );
  OAI211_X1 U15416 ( .C1(n13298), .C2(n15352), .A(n13297), .B(n13296), .ZN(
        n13380) );
  MUX2_X1 U15417 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13380), .S(n15392), .Z(
        P2_U3527) );
  NAND3_X1 U15418 ( .A1(n13300), .A2(n13299), .A3(n15373), .ZN(n13305) );
  NAND2_X1 U15419 ( .A1(n13301), .A2(n15366), .ZN(n13302) );
  NAND4_X1 U15420 ( .A1(n13305), .A2(n13304), .A3(n13303), .A4(n13302), .ZN(
        n13381) );
  MUX2_X1 U15421 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13381), .S(n15392), .Z(
        P2_U3526) );
  AOI21_X1 U15422 ( .B1(n15366), .B2(n13307), .A(n13306), .ZN(n13308) );
  OAI211_X1 U15423 ( .C1(n13310), .C2(n15352), .A(n13309), .B(n13308), .ZN(
        n13382) );
  MUX2_X1 U15424 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13382), .S(n15392), .Z(
        P2_U3525) );
  AOI211_X1 U15425 ( .C1(n15366), .C2(n13313), .A(n13312), .B(n13311), .ZN(
        n13314) );
  OAI21_X1 U15426 ( .B1(n13315), .B2(n15352), .A(n13314), .ZN(n13383) );
  MUX2_X1 U15427 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13383), .S(n15392), .Z(
        P2_U3524) );
  INV_X1 U15428 ( .A(n13316), .ZN(n13321) );
  AOI21_X1 U15429 ( .B1(n15366), .B2(n13318), .A(n13317), .ZN(n13319) );
  OAI211_X1 U15430 ( .C1(n13321), .C2(n15352), .A(n13320), .B(n13319), .ZN(
        n13384) );
  MUX2_X1 U15431 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13384), .S(n15392), .Z(
        P2_U3523) );
  NAND2_X1 U15432 ( .A1(n13322), .A2(n15373), .ZN(n13329) );
  INV_X1 U15433 ( .A(n13323), .ZN(n13324) );
  AOI21_X1 U15434 ( .B1(n13325), .B2(n15366), .A(n13324), .ZN(n13328) );
  NAND4_X1 U15435 ( .A1(n13329), .A2(n13328), .A3(n13327), .A4(n13326), .ZN(
        n13385) );
  MUX2_X1 U15436 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13385), .S(n15392), .Z(
        P2_U3522) );
  NAND2_X1 U15437 ( .A1(n13330), .A2(n15366), .ZN(n13331) );
  OAI211_X1 U15438 ( .C1(n13333), .C2(n15352), .A(n13332), .B(n13331), .ZN(
        n13335) );
  MUX2_X1 U15439 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13386), .S(n15392), .Z(
        P2_U3521) );
  AOI21_X1 U15440 ( .B1(n15366), .B2(n13337), .A(n13336), .ZN(n13338) );
  OAI211_X1 U15441 ( .C1(n13340), .C2(n15352), .A(n13339), .B(n13338), .ZN(
        n13387) );
  MUX2_X1 U15442 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13387), .S(n15392), .Z(
        P2_U3520) );
  AOI211_X1 U15443 ( .C1(n15366), .C2(n13343), .A(n13342), .B(n13341), .ZN(
        n13344) );
  OAI21_X1 U15444 ( .B1(n13345), .B2(n15352), .A(n13344), .ZN(n13388) );
  MUX2_X1 U15445 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13388), .S(n15392), .Z(
        P2_U3519) );
  AOI211_X1 U15446 ( .C1(n15366), .C2(n13348), .A(n13347), .B(n13346), .ZN(
        n13349) );
  OAI21_X1 U15447 ( .B1(n13350), .B2(n15352), .A(n13349), .ZN(n13389) );
  MUX2_X1 U15448 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13389), .S(n15392), .Z(
        P2_U3518) );
  INV_X1 U15449 ( .A(n13351), .ZN(n13356) );
  AOI21_X1 U15450 ( .B1(n15366), .B2(n13353), .A(n13352), .ZN(n13354) );
  OAI211_X1 U15451 ( .C1(n13356), .C2(n15352), .A(n13355), .B(n13354), .ZN(
        n13390) );
  MUX2_X1 U15452 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13390), .S(n15392), .Z(
        P2_U3517) );
  OAI21_X1 U15453 ( .B1(n13358), .B2(n15376), .A(n13357), .ZN(n13359) );
  AOI211_X1 U15454 ( .C1(n13361), .C2(n15373), .A(n13360), .B(n13359), .ZN(
        n13362) );
  INV_X1 U15455 ( .A(n13362), .ZN(n13391) );
  MUX2_X1 U15456 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13391), .S(n15392), .Z(
        P2_U3516) );
  AOI21_X1 U15457 ( .B1(n15366), .B2(n13364), .A(n13363), .ZN(n13366) );
  OAI211_X1 U15458 ( .C1(n15352), .C2(n13367), .A(n13366), .B(n13365), .ZN(
        n13392) );
  MUX2_X1 U15459 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13392), .S(n15392), .Z(
        P2_U3515) );
  AOI21_X1 U15460 ( .B1(n15366), .B2(n13369), .A(n13368), .ZN(n13371) );
  OAI211_X1 U15461 ( .C1(n15352), .C2(n13372), .A(n13371), .B(n13370), .ZN(
        n13393) );
  MUX2_X1 U15462 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13393), .S(n15392), .Z(
        P2_U3514) );
  AOI21_X1 U15463 ( .B1(n15366), .B2(n13374), .A(n13373), .ZN(n13375) );
  OAI211_X1 U15464 ( .C1(n15352), .C2(n13377), .A(n13376), .B(n13375), .ZN(
        n13394) );
  MUX2_X1 U15465 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13394), .S(n15392), .Z(
        P2_U3512) );
  MUX2_X1 U15466 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13378), .S(n15383), .Z(
        P2_U3498) );
  MUX2_X1 U15467 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13379), .S(n15383), .Z(
        P2_U3497) );
  MUX2_X1 U15468 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13380), .S(n15383), .Z(
        P2_U3495) );
  MUX2_X1 U15469 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13381), .S(n15383), .Z(
        P2_U3494) );
  MUX2_X1 U15470 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13382), .S(n15383), .Z(
        P2_U3493) );
  MUX2_X1 U15471 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13383), .S(n15383), .Z(
        P2_U3492) );
  MUX2_X1 U15472 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13384), .S(n15383), .Z(
        P2_U3491) );
  MUX2_X1 U15473 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13385), .S(n15383), .Z(
        P2_U3490) );
  MUX2_X1 U15474 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13386), .S(n15383), .Z(
        P2_U3489) );
  MUX2_X1 U15475 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13387), .S(n15383), .Z(
        P2_U3488) );
  MUX2_X1 U15476 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13388), .S(n15383), .Z(
        P2_U3487) );
  MUX2_X1 U15477 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13389), .S(n15383), .Z(
        P2_U3486) );
  MUX2_X1 U15478 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13390), .S(n15383), .Z(
        P2_U3484) );
  MUX2_X1 U15479 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13391), .S(n15383), .Z(
        P2_U3481) );
  MUX2_X1 U15480 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13392), .S(n15383), .Z(
        P2_U3478) );
  MUX2_X1 U15481 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13393), .S(n15383), .Z(
        P2_U3475) );
  MUX2_X1 U15482 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13394), .S(n15383), .Z(
        P2_U3469) );
  INV_X1 U15483 ( .A(n14560), .ZN(n13400) );
  NOR4_X1 U15484 ( .A1(n13395), .A2(P2_IR_REG_30__SCAN_IN), .A3(n7991), .A4(
        P2_U3088), .ZN(n13396) );
  AOI21_X1 U15485 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13397), .A(n13396), 
        .ZN(n13398) );
  OAI21_X1 U15486 ( .B1(n13400), .B2(n13399), .A(n13398), .ZN(P2_U3296) );
  OAI222_X1 U15487 ( .A1(n13399), .A2(n13403), .B1(P2_U3088), .B2(n13402), 
        .C1(n13401), .C2(n13417), .ZN(P2_U3298) );
  NAND2_X1 U15488 ( .A1(n13676), .A2(n13404), .ZN(n13406) );
  OAI211_X1 U15489 ( .C1(n13417), .C2(n13407), .A(n13406), .B(n13405), .ZN(
        P2_U3299) );
  INV_X1 U15490 ( .A(n13420), .ZN(n14563) );
  OAI222_X1 U15491 ( .A1(n13409), .A2(P2_U3088), .B1(n13399), .B2(n14563), 
        .C1(n13408), .C2(n13417), .ZN(P2_U3300) );
  INV_X1 U15492 ( .A(n13614), .ZN(n14566) );
  OAI222_X1 U15493 ( .A1(n13411), .A2(P2_U3088), .B1(n13399), .B2(n14566), 
        .C1(n13410), .C2(n13417), .ZN(P2_U3301) );
  INV_X1 U15494 ( .A(n13598), .ZN(n14569) );
  OAI222_X1 U15495 ( .A1(n13417), .A2(n13413), .B1(n13399), .B2(n14569), .C1(
        n13412), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U15496 ( .A(n13582), .ZN(n14573) );
  INV_X1 U15497 ( .A(n13414), .ZN(n13415) );
  OAI222_X1 U15498 ( .A1(n13417), .A2(n13416), .B1(n13399), .B2(n14573), .C1(
        n13415), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U15499 ( .A(n13418), .ZN(n13419) );
  MUX2_X1 U15500 ( .A(n13419), .B(n15229), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  NAND2_X1 U15501 ( .A1(n13420), .A2(n11615), .ZN(n13422) );
  OR2_X1 U15502 ( .A1(n13850), .A2(n14562), .ZN(n13421) );
  NAND2_X1 U15503 ( .A1(n14460), .A2(n13627), .ZN(n13434) );
  NAND2_X1 U15504 ( .A1(n13831), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n13432) );
  INV_X1 U15505 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n13423) );
  OR2_X1 U15506 ( .A1(n10037), .A2(n13423), .ZN(n13431) );
  NAND2_X1 U15507 ( .A1(n13527), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13529) );
  NAND2_X1 U15508 ( .A1(n13455), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n13439) );
  INV_X1 U15509 ( .A(n13439), .ZN(n13570) );
  NAND2_X1 U15510 ( .A1(n13570), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n13569) );
  INV_X1 U15511 ( .A(n13569), .ZN(n13587) );
  NAND2_X1 U15512 ( .A1(n13587), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n13586) );
  INV_X1 U15513 ( .A(n13586), .ZN(n13602) );
  NAND2_X1 U15514 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n13602), .ZN(n13618) );
  INV_X1 U15515 ( .A(n13618), .ZN(n13424) );
  NAND2_X1 U15516 ( .A1(n13424), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n13620) );
  INV_X1 U15517 ( .A(n13620), .ZN(n13425) );
  NAND2_X1 U15518 ( .A1(n13425), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n13690) );
  INV_X1 U15519 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13426) );
  NAND2_X1 U15520 ( .A1(n13620), .A2(n13426), .ZN(n13427) );
  NAND2_X1 U15521 ( .A1(n13690), .A2(n13427), .ZN(n14237) );
  OR2_X1 U15522 ( .A1(n13692), .A2(n14237), .ZN(n13430) );
  OR2_X1 U15523 ( .A1(n13844), .A2(n13428), .ZN(n13429) );
  NAND4_X1 U15524 ( .A1(n13432), .A2(n13431), .A3(n13430), .A4(n13429), .ZN(
        n14246) );
  NAND2_X1 U15525 ( .A1(n13607), .A2(n14246), .ZN(n13433) );
  NAND2_X1 U15526 ( .A1(n13434), .A2(n13433), .ZN(n13435) );
  XNOR2_X1 U15527 ( .A(n13435), .B(n13682), .ZN(n13671) );
  AOI22_X1 U15528 ( .A1(n14460), .A2(n13607), .B1(n13626), .B2(n14246), .ZN(
        n13672) );
  XNOR2_X1 U15529 ( .A(n13671), .B(n13672), .ZN(n13674) );
  OR2_X1 U15530 ( .A1(n13437), .A2(n13436), .ZN(n13438) );
  XNOR2_X1 U15531 ( .A(n13438), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14575) );
  OR2_X1 U15532 ( .A1(n13455), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n13440) );
  AND2_X1 U15533 ( .A1(n13440), .A2(n13439), .ZN(n14313) );
  NAND2_X1 U15534 ( .A1(n14313), .A2(n13553), .ZN(n13446) );
  INV_X1 U15535 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n13443) );
  NAND2_X1 U15536 ( .A1(n13831), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n13442) );
  NAND2_X1 U15537 ( .A1(n13832), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n13441) );
  OAI211_X1 U15538 ( .C1(n10037), .C2(n13443), .A(n13442), .B(n13441), .ZN(
        n13444) );
  INV_X1 U15539 ( .A(n13444), .ZN(n13445) );
  AOI22_X1 U15540 ( .A1(n14314), .A2(n13607), .B1(n13626), .B2(n14326), .ZN(
        n13561) );
  INV_X1 U15541 ( .A(n13561), .ZN(n13563) );
  NAND2_X1 U15542 ( .A1(n14314), .A2(n13627), .ZN(n13448) );
  NAND2_X1 U15543 ( .A1(n14326), .A2(n13607), .ZN(n13447) );
  NAND2_X1 U15544 ( .A1(n13448), .A2(n13447), .ZN(n13449) );
  XNOR2_X1 U15545 ( .A(n13449), .B(n13682), .ZN(n13562) );
  NAND2_X1 U15546 ( .A1(n13450), .A2(n11615), .ZN(n13453) );
  OR2_X1 U15547 ( .A1(n13850), .A2(n13451), .ZN(n13452) );
  NOR2_X1 U15548 ( .A1(n13547), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n13454) );
  OR2_X1 U15549 ( .A1(n13455), .A2(n13454), .ZN(n13707) );
  NAND2_X1 U15550 ( .A1(n13688), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n13457) );
  NAND2_X1 U15551 ( .A1(n13832), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n13456) );
  OAI211_X1 U15552 ( .C1(n13842), .C2(n12293), .A(n13457), .B(n13456), .ZN(
        n13458) );
  INV_X1 U15553 ( .A(n13458), .ZN(n13459) );
  AOI22_X1 U15554 ( .A1(n14496), .A2(n13607), .B1(n13626), .B2(n14347), .ZN(
        n13558) );
  INV_X1 U15555 ( .A(n13558), .ZN(n13560) );
  AOI22_X1 U15556 ( .A1(n14496), .A2(n13627), .B1(n13607), .B2(n14347), .ZN(
        n13460) );
  XNOR2_X1 U15557 ( .A(n13460), .B(n13682), .ZN(n13557) );
  INV_X1 U15558 ( .A(n13557), .ZN(n13559) );
  NAND2_X1 U15559 ( .A1(n13461), .A2(n11615), .ZN(n13464) );
  AOI22_X1 U15560 ( .A1(n13524), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13462), 
        .B2(n13523), .ZN(n13463) );
  NAND2_X1 U15561 ( .A1(n13529), .A2(n13667), .ZN(n13465) );
  AND2_X1 U15562 ( .A1(n13546), .A2(n13465), .ZN(n14359) );
  NAND2_X1 U15563 ( .A1(n14359), .A2(n13553), .ZN(n13471) );
  NAND2_X1 U15564 ( .A1(n13831), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n13467) );
  NAND2_X1 U15565 ( .A1(n13832), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n13466) );
  OAI211_X1 U15566 ( .C1(n10037), .C2(n13468), .A(n13467), .B(n13466), .ZN(
        n13469) );
  INV_X1 U15567 ( .A(n13469), .ZN(n13470) );
  NAND2_X1 U15568 ( .A1(n13471), .A2(n13470), .ZN(n14345) );
  INV_X1 U15569 ( .A(n14345), .ZN(n14172) );
  NOR2_X1 U15570 ( .A1(n14172), .A2(n13680), .ZN(n13472) );
  AOI21_X1 U15571 ( .B1(n14358), .B2(n13607), .A(n13472), .ZN(n13538) );
  INV_X1 U15572 ( .A(n13538), .ZN(n13540) );
  NAND2_X1 U15573 ( .A1(n14358), .A2(n13627), .ZN(n13474) );
  NAND2_X1 U15574 ( .A1(n14345), .A2(n13607), .ZN(n13473) );
  NAND2_X1 U15575 ( .A1(n13474), .A2(n13473), .ZN(n13475) );
  XNOR2_X1 U15576 ( .A(n13475), .B(n13682), .ZN(n13539) );
  INV_X1 U15577 ( .A(n13476), .ZN(n13478) );
  NOR2_X1 U15578 ( .A1(n13478), .A2(n13477), .ZN(n13479) );
  NAND2_X1 U15579 ( .A1(n13648), .A2(n13627), .ZN(n13483) );
  NAND2_X1 U15580 ( .A1(n13607), .A2(n14056), .ZN(n13482) );
  NAND2_X1 U15581 ( .A1(n13483), .A2(n13482), .ZN(n13484) );
  XNOR2_X1 U15582 ( .A(n13484), .B(n13682), .ZN(n13487) );
  NOR2_X1 U15583 ( .A1(n13680), .A2(n13485), .ZN(n13486) );
  AOI21_X1 U15584 ( .B1(n13648), .B2(n13607), .A(n13486), .ZN(n13488) );
  XNOR2_X1 U15585 ( .A(n13487), .B(n13488), .ZN(n13647) );
  INV_X1 U15586 ( .A(n13487), .ZN(n13489) );
  NAND2_X1 U15587 ( .A1(n14534), .A2(n13627), .ZN(n13491) );
  INV_X1 U15588 ( .A(n13726), .ZN(n14409) );
  NAND2_X1 U15589 ( .A1(n13607), .A2(n14409), .ZN(n13490) );
  NAND2_X1 U15590 ( .A1(n13491), .A2(n13490), .ZN(n13492) );
  XNOR2_X1 U15591 ( .A(n13492), .B(n13682), .ZN(n13494) );
  NOR2_X1 U15592 ( .A1(n13680), .A2(n13726), .ZN(n13493) );
  AOI21_X1 U15593 ( .B1(n14534), .B2(n13607), .A(n13493), .ZN(n13787) );
  NAND2_X1 U15594 ( .A1(n13495), .A2(n11615), .ZN(n13498) );
  AOI22_X1 U15595 ( .A1(n13524), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n13523), 
        .B2(n13496), .ZN(n13497) );
  NAND2_X1 U15596 ( .A1(n14414), .A2(n13627), .ZN(n13500) );
  NAND2_X1 U15597 ( .A1(n13607), .A2(n14389), .ZN(n13499) );
  NAND2_X1 U15598 ( .A1(n13500), .A2(n13499), .ZN(n13501) );
  XNOR2_X1 U15599 ( .A(n13501), .B(n13682), .ZN(n13505) );
  INV_X1 U15600 ( .A(n14389), .ZN(n14170) );
  NOR2_X1 U15601 ( .A1(n13680), .A2(n14170), .ZN(n13502) );
  AOI21_X1 U15602 ( .B1(n14414), .B2(n13607), .A(n13502), .ZN(n13503) );
  XNOR2_X1 U15603 ( .A(n13505), .B(n13503), .ZN(n13721) );
  INV_X1 U15604 ( .A(n13503), .ZN(n13504) );
  NAND2_X1 U15605 ( .A1(n13507), .A2(n11615), .ZN(n13510) );
  AOI22_X1 U15606 ( .A1(n13524), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n13523), 
        .B2(n13508), .ZN(n13509) );
  NAND2_X1 U15607 ( .A1(n14522), .A2(n13627), .ZN(n13516) );
  NOR2_X1 U15608 ( .A1(n13511), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13512) );
  OR2_X1 U15609 ( .A1(n13527), .A2(n13512), .ZN(n14398) );
  AOI22_X1 U15610 ( .A1(n13688), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n13832), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n13514) );
  OR2_X1 U15611 ( .A1(n13842), .A2(n12245), .ZN(n13513) );
  OAI211_X1 U15612 ( .C1(n14398), .C2(n13692), .A(n13514), .B(n13513), .ZN(
        n14408) );
  NAND2_X1 U15613 ( .A1(n13607), .A2(n14408), .ZN(n13515) );
  NAND2_X1 U15614 ( .A1(n13516), .A2(n13515), .ZN(n13518) );
  XNOR2_X1 U15615 ( .A(n13518), .B(n13517), .ZN(n13521) );
  INV_X1 U15616 ( .A(n14408), .ZN(n14171) );
  NOR2_X1 U15617 ( .A1(n13680), .A2(n14171), .ZN(n13519) );
  AOI21_X1 U15618 ( .B1(n14522), .B2(n13607), .A(n13519), .ZN(n13520) );
  OR2_X1 U15619 ( .A1(n13521), .A2(n13520), .ZN(n13731) );
  AND2_X1 U15620 ( .A1(n13521), .A2(n13520), .ZN(n13730) );
  NAND2_X1 U15621 ( .A1(n13522), .A2(n11615), .ZN(n13526) );
  AOI22_X1 U15622 ( .A1(n13524), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n13523), 
        .B2(n14139), .ZN(n13525) );
  OR2_X1 U15623 ( .A1(n13527), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13528) );
  NAND2_X1 U15624 ( .A1(n13529), .A2(n13528), .ZN(n14377) );
  AOI22_X1 U15625 ( .A1(n13688), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n13831), 
        .B2(P1_REG2_REG_18__SCAN_IN), .ZN(n13531) );
  NAND2_X1 U15626 ( .A1(n13832), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n13530) );
  OAI211_X1 U15627 ( .C1(n14377), .C2(n13692), .A(n13531), .B(n13530), .ZN(
        n14390) );
  AOI22_X1 U15628 ( .A1(n14375), .A2(n13607), .B1(n13626), .B2(n14390), .ZN(
        n13535) );
  NAND2_X1 U15629 ( .A1(n14375), .A2(n13627), .ZN(n13533) );
  NAND2_X1 U15630 ( .A1(n13607), .A2(n14390), .ZN(n13532) );
  NAND2_X1 U15631 ( .A1(n13533), .A2(n13532), .ZN(n13534) );
  XNOR2_X1 U15632 ( .A(n13534), .B(n13682), .ZN(n13537) );
  XOR2_X1 U15633 ( .A(n13535), .B(n13537), .Z(n13768) );
  INV_X1 U15634 ( .A(n13535), .ZN(n13536) );
  XOR2_X1 U15635 ( .A(n13538), .B(n13539), .Z(n13665) );
  NAND2_X1 U15636 ( .A1(n13541), .A2(n11615), .ZN(n13544) );
  OR2_X1 U15637 ( .A1(n13850), .A2(n13542), .ZN(n13543) );
  AND2_X1 U15638 ( .A1(n13546), .A2(n13545), .ZN(n13548) );
  OR2_X1 U15639 ( .A1(n13548), .A2(n13547), .ZN(n13750) );
  INV_X1 U15640 ( .A(n13750), .ZN(n14348) );
  NAND2_X1 U15641 ( .A1(n13831), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n13550) );
  NAND2_X1 U15642 ( .A1(n13688), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n13549) );
  OAI211_X1 U15643 ( .C1(n13551), .C2(n13844), .A(n13550), .B(n13549), .ZN(
        n13552) );
  AOI21_X1 U15644 ( .B1(n14348), .B2(n13553), .A(n13552), .ZN(n14195) );
  OAI22_X1 U15645 ( .A1(n14502), .A2(n10072), .B1(n14195), .B2(n13681), .ZN(
        n13554) );
  XNOR2_X1 U15646 ( .A(n13554), .B(n13682), .ZN(n13556) );
  OAI22_X1 U15647 ( .A1(n14502), .A2(n13681), .B1(n14195), .B2(n13680), .ZN(
        n13555) );
  XNOR2_X1 U15648 ( .A(n13556), .B(n13555), .ZN(n13752) );
  XOR2_X1 U15649 ( .A(n13558), .B(n13557), .Z(n13705) );
  OAI21_X1 U15650 ( .B1(n13560), .B2(n13559), .A(n13703), .ZN(n13758) );
  XNOR2_X1 U15651 ( .A(n13562), .B(n13561), .ZN(n13759) );
  NAND2_X1 U15652 ( .A1(n13758), .A2(n13759), .ZN(n13757) );
  OAI21_X1 U15653 ( .B1(n13563), .B2(n13562), .A(n13757), .ZN(n13657) );
  NAND2_X1 U15654 ( .A1(n13564), .A2(n11615), .ZN(n13567) );
  OR2_X1 U15655 ( .A1(n13850), .A2(n13565), .ZN(n13566) );
  NAND2_X1 U15656 ( .A1(n14304), .A2(n13627), .ZN(n13577) );
  NAND2_X1 U15657 ( .A1(n13688), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n13575) );
  INV_X1 U15658 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n13568) );
  OR2_X1 U15659 ( .A1(n13844), .A2(n13568), .ZN(n13574) );
  OAI21_X1 U15660 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n13570), .A(n13569), 
        .ZN(n14302) );
  OR2_X1 U15661 ( .A1(n13692), .A2(n14302), .ZN(n13573) );
  INV_X1 U15662 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n13571) );
  OR2_X1 U15663 ( .A1(n13842), .A2(n13571), .ZN(n13572) );
  NAND4_X1 U15664 ( .A1(n13575), .A2(n13574), .A3(n13573), .A4(n13572), .ZN(
        n14318) );
  NAND2_X1 U15665 ( .A1(n13607), .A2(n14318), .ZN(n13576) );
  NAND2_X1 U15666 ( .A1(n13577), .A2(n13576), .ZN(n13578) );
  XNOR2_X1 U15667 ( .A(n13578), .B(n13682), .ZN(n13579) );
  AOI22_X1 U15668 ( .A1(n14304), .A2(n13607), .B1(n13626), .B2(n14318), .ZN(
        n13580) );
  XNOR2_X1 U15669 ( .A(n13579), .B(n13580), .ZN(n13658) );
  INV_X1 U15670 ( .A(n13579), .ZN(n13581) );
  NAND2_X1 U15671 ( .A1(n13582), .A2(n11615), .ZN(n13584) );
  OR2_X1 U15672 ( .A1(n13850), .A2(n14572), .ZN(n13583) );
  NAND2_X1 U15673 ( .A1(n13688), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n13591) );
  OR2_X1 U15674 ( .A1(n13844), .A2(n13585), .ZN(n13590) );
  OAI21_X1 U15675 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n13587), .A(n13586), 
        .ZN(n14285) );
  OR2_X1 U15676 ( .A1(n13692), .A2(n14285), .ZN(n13589) );
  INV_X1 U15677 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14286) );
  OR2_X1 U15678 ( .A1(n13842), .A2(n14286), .ZN(n13588) );
  NAND4_X1 U15679 ( .A1(n13591), .A2(n13590), .A3(n13589), .A4(n13588), .ZN(
        n14295) );
  AOI22_X1 U15680 ( .A1(n14284), .A2(n13607), .B1(n13626), .B2(n14295), .ZN(
        n13595) );
  NAND2_X1 U15681 ( .A1(n14284), .A2(n13627), .ZN(n13593) );
  NAND2_X1 U15682 ( .A1(n13607), .A2(n14295), .ZN(n13592) );
  NAND2_X1 U15683 ( .A1(n13593), .A2(n13592), .ZN(n13594) );
  XNOR2_X1 U15684 ( .A(n13594), .B(n13682), .ZN(n13597) );
  XOR2_X1 U15685 ( .A(n13595), .B(n13597), .Z(n13742) );
  INV_X1 U15686 ( .A(n13595), .ZN(n13596) );
  NAND2_X1 U15687 ( .A1(n13598), .A2(n11615), .ZN(n13600) );
  OR2_X1 U15688 ( .A1(n13850), .A2(n14568), .ZN(n13599) );
  NAND2_X1 U15689 ( .A1(n14472), .A2(n13627), .ZN(n13609) );
  NAND2_X1 U15690 ( .A1(n13688), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n13606) );
  INV_X1 U15691 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n13601) );
  OR2_X1 U15692 ( .A1(n13844), .A2(n13601), .ZN(n13605) );
  OAI21_X1 U15693 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n13602), .A(n13618), 
        .ZN(n14266) );
  OR2_X1 U15694 ( .A1(n13692), .A2(n14266), .ZN(n13604) );
  INV_X1 U15695 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14267) );
  OR2_X1 U15696 ( .A1(n13842), .A2(n14267), .ZN(n13603) );
  NAND4_X1 U15697 ( .A1(n13606), .A2(n13605), .A3(n13604), .A4(n13603), .ZN(
        n14278) );
  NAND2_X1 U15698 ( .A1(n13607), .A2(n14278), .ZN(n13608) );
  NAND2_X1 U15699 ( .A1(n13609), .A2(n13608), .ZN(n13610) );
  XNOR2_X1 U15700 ( .A(n13610), .B(n13682), .ZN(n13611) );
  AOI22_X1 U15701 ( .A1(n14472), .A2(n13607), .B1(n13626), .B2(n14278), .ZN(
        n13612) );
  XNOR2_X1 U15702 ( .A(n13611), .B(n13612), .ZN(n13714) );
  INV_X1 U15703 ( .A(n13611), .ZN(n13613) );
  NAND2_X1 U15704 ( .A1(n13614), .A2(n11615), .ZN(n13616) );
  OR2_X1 U15705 ( .A1(n13850), .A2(n14565), .ZN(n13615) );
  NAND2_X1 U15706 ( .A1(n13688), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n13625) );
  OR2_X1 U15707 ( .A1(n13842), .A2(n12319), .ZN(n13624) );
  INV_X1 U15708 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13617) );
  NAND2_X1 U15709 ( .A1(n13618), .A2(n13617), .ZN(n13619) );
  NAND2_X1 U15710 ( .A1(n13620), .A2(n13619), .ZN(n14252) );
  OR2_X1 U15711 ( .A1(n13692), .A2(n14252), .ZN(n13623) );
  INV_X1 U15712 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n13621) );
  OR2_X1 U15713 ( .A1(n13844), .A2(n13621), .ZN(n13622) );
  NAND4_X1 U15714 ( .A1(n13625), .A2(n13624), .A3(n13623), .A4(n13622), .ZN(
        n14262) );
  AOI22_X1 U15715 ( .A1(n14254), .A2(n13607), .B1(n13626), .B2(n14262), .ZN(
        n13631) );
  NAND2_X1 U15716 ( .A1(n14254), .A2(n13627), .ZN(n13629) );
  NAND2_X1 U15717 ( .A1(n13607), .A2(n14262), .ZN(n13628) );
  NAND2_X1 U15718 ( .A1(n13629), .A2(n13628), .ZN(n13630) );
  XNOR2_X1 U15719 ( .A(n13630), .B(n13682), .ZN(n13633) );
  XOR2_X1 U15720 ( .A(n13631), .B(n13633), .Z(n13775) );
  INV_X1 U15721 ( .A(n13631), .ZN(n13632) );
  XOR2_X1 U15722 ( .A(n13674), .B(n13675), .Z(n13645) );
  NAND2_X1 U15723 ( .A1(n13831), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n13640) );
  INV_X1 U15724 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n13634) );
  OR2_X1 U15725 ( .A1(n10037), .A2(n13634), .ZN(n13639) );
  INV_X1 U15726 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13635) );
  XNOR2_X1 U15727 ( .A(n13690), .B(n13635), .ZN(n14222) );
  OR2_X1 U15728 ( .A1(n13692), .A2(n14222), .ZN(n13638) );
  OR2_X1 U15729 ( .A1(n13844), .A2(n13636), .ZN(n13637) );
  NAND4_X1 U15730 ( .A1(n13640), .A2(n13639), .A3(n13638), .A4(n13637), .ZN(
        n14233) );
  AOI22_X1 U15731 ( .A1(n13776), .A2(n14233), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13642) );
  NAND2_X1 U15732 ( .A1(n13777), .A2(n14262), .ZN(n13641) );
  OAI211_X1 U15733 ( .C1(n13780), .C2(n14237), .A(n13642), .B(n13641), .ZN(
        n13643) );
  AOI21_X1 U15734 ( .B1(n14460), .B2(n13782), .A(n13643), .ZN(n13644) );
  OAI21_X1 U15735 ( .B1(n13645), .B2(n13784), .A(n13644), .ZN(P1_U3214) );
  XOR2_X1 U15736 ( .A(n13647), .B(n13646), .Z(n13656) );
  NOR2_X1 U15737 ( .A1(n7598), .A2(n15191), .ZN(n14935) );
  NAND2_X1 U15738 ( .A1(n13650), .A2(n13649), .ZN(n13651) );
  OAI211_X1 U15739 ( .C1(n13780), .C2(n13653), .A(n13652), .B(n13651), .ZN(
        n13654) );
  AOI21_X1 U15740 ( .B1(n14935), .B2(n13772), .A(n13654), .ZN(n13655) );
  OAI21_X1 U15741 ( .B1(n13656), .B2(n13784), .A(n13655), .ZN(P1_U3215) );
  XOR2_X1 U15742 ( .A(n13658), .B(n13657), .Z(n13663) );
  AND2_X1 U15743 ( .A1(n14304), .A2(n15200), .ZN(n14483) );
  AOI22_X1 U15744 ( .A1(n13776), .A2(n14295), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13660) );
  NAND2_X1 U15745 ( .A1(n13777), .A2(n14326), .ZN(n13659) );
  OAI211_X1 U15746 ( .C1(n13780), .C2(n14302), .A(n13660), .B(n13659), .ZN(
        n13661) );
  AOI21_X1 U15747 ( .B1(n14483), .B2(n13772), .A(n13661), .ZN(n13662) );
  OAI21_X1 U15748 ( .B1(n13663), .B2(n13784), .A(n13662), .ZN(P1_U3216) );
  INV_X1 U15749 ( .A(n14358), .ZN(n14508) );
  AOI211_X1 U15750 ( .C1(n13665), .C2(n13664), .A(n13784), .B(n6661), .ZN(
        n13666) );
  INV_X1 U15751 ( .A(n13666), .ZN(n13670) );
  AOI22_X1 U15752 ( .A1(n14173), .A2(n15059), .B1(n15049), .B2(n14390), .ZN(
        n14507) );
  OAI22_X1 U15753 ( .A1(n13795), .A2(n14507), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13667), .ZN(n13668) );
  AOI21_X1 U15754 ( .B1(n13798), .B2(n14359), .A(n13668), .ZN(n13669) );
  OAI211_X1 U15755 ( .C1(n14508), .C2(n13801), .A(n13670), .B(n13669), .ZN(
        P1_U3219) );
  INV_X1 U15756 ( .A(n13671), .ZN(n13673) );
  AOI22_X1 U15757 ( .A1(n13675), .A2(n13674), .B1(n13673), .B2(n13672), .ZN(
        n13687) );
  NAND2_X1 U15758 ( .A1(n13676), .A2(n11615), .ZN(n13679) );
  OR2_X1 U15759 ( .A1(n13850), .A2(n13677), .ZN(n13678) );
  OAI22_X1 U15760 ( .A1(n14182), .A2(n13681), .B1(n14181), .B2(n13680), .ZN(
        n13685) );
  OAI22_X1 U15761 ( .A1(n14182), .A2(n10072), .B1(n14181), .B2(n13681), .ZN(
        n13683) );
  XNOR2_X1 U15762 ( .A(n13683), .B(n13682), .ZN(n13684) );
  XOR2_X1 U15763 ( .A(n13685), .B(n13684), .Z(n13686) );
  XNOR2_X1 U15764 ( .A(n13687), .B(n13686), .ZN(n13702) );
  NAND2_X1 U15765 ( .A1(n13688), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n13697) );
  OR2_X1 U15766 ( .A1(n13842), .A2(n13689), .ZN(n13696) );
  INV_X1 U15767 ( .A(n13690), .ZN(n13691) );
  NAND2_X1 U15768 ( .A1(n13691), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14205) );
  OR2_X1 U15769 ( .A1(n13692), .A2(n14205), .ZN(n13695) );
  INV_X1 U15770 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n13693) );
  OR2_X1 U15771 ( .A1(n13844), .A2(n13693), .ZN(n13694) );
  NAND4_X1 U15772 ( .A1(n13697), .A2(n13696), .A3(n13695), .A4(n13694), .ZN(
        n14215) );
  AOI22_X1 U15773 ( .A1(n13776), .A2(n14215), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13699) );
  NAND2_X1 U15774 ( .A1(n13777), .A2(n14246), .ZN(n13698) );
  OAI211_X1 U15775 ( .C1(n13780), .C2(n14222), .A(n13699), .B(n13698), .ZN(
        n13700) );
  AOI21_X1 U15776 ( .B1(n14452), .B2(n13782), .A(n13700), .ZN(n13701) );
  OAI21_X1 U15777 ( .B1(n13702), .B2(n13784), .A(n13701), .ZN(P1_U3220) );
  INV_X1 U15778 ( .A(n14496), .ZN(n14330) );
  OAI21_X1 U15779 ( .B1(n13705), .B2(n13704), .A(n13703), .ZN(n13706) );
  NAND2_X1 U15780 ( .A1(n13706), .A2(n13790), .ZN(n13712) );
  INV_X1 U15781 ( .A(n13707), .ZN(n14328) );
  INV_X1 U15782 ( .A(n14326), .ZN(n13709) );
  AOI22_X1 U15783 ( .A1(n13777), .A2(n14173), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13708) );
  OAI21_X1 U15784 ( .B1(n13709), .B2(n13762), .A(n13708), .ZN(n13710) );
  AOI21_X1 U15785 ( .B1(n14328), .B2(n13798), .A(n13710), .ZN(n13711) );
  OAI211_X1 U15786 ( .C1(n14330), .C2(n13801), .A(n13712), .B(n13711), .ZN(
        P1_U3223) );
  XOR2_X1 U15787 ( .A(n13714), .B(n13713), .Z(n13719) );
  AOI22_X1 U15788 ( .A1(n13776), .A2(n14262), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13716) );
  NAND2_X1 U15789 ( .A1(n13777), .A2(n14295), .ZN(n13715) );
  OAI211_X1 U15790 ( .C1(n13780), .C2(n14266), .A(n13716), .B(n13715), .ZN(
        n13717) );
  AOI21_X1 U15791 ( .B1(n14472), .B2(n13782), .A(n13717), .ZN(n13718) );
  OAI21_X1 U15792 ( .B1(n13719), .B2(n13784), .A(n13718), .ZN(P1_U3225) );
  INV_X1 U15793 ( .A(n14414), .ZN(n14527) );
  INV_X1 U15794 ( .A(n13720), .ZN(n13723) );
  AOI21_X1 U15795 ( .B1(n13792), .B2(n13786), .A(n13721), .ZN(n13722) );
  OAI21_X1 U15796 ( .B1(n13723), .B2(n13722), .A(n13790), .ZN(n13729) );
  NAND2_X1 U15797 ( .A1(n13776), .A2(n14408), .ZN(n13724) );
  OAI211_X1 U15798 ( .C1(n13735), .C2(n13726), .A(n13725), .B(n13724), .ZN(
        n13727) );
  AOI21_X1 U15799 ( .B1(n14410), .B2(n13798), .A(n13727), .ZN(n13728) );
  OAI211_X1 U15800 ( .C1(n14527), .C2(n13801), .A(n13729), .B(n13728), .ZN(
        P1_U3226) );
  NAND2_X1 U15801 ( .A1(n7506), .A2(n13731), .ZN(n13732) );
  XNOR2_X1 U15802 ( .A(n13733), .B(n13732), .ZN(n13740) );
  OAI21_X1 U15803 ( .B1(n13735), .B2(n14170), .A(n13734), .ZN(n13736) );
  AOI21_X1 U15804 ( .B1(n13776), .B2(n14390), .A(n13736), .ZN(n13737) );
  OAI21_X1 U15805 ( .B1(n13780), .B2(n14398), .A(n13737), .ZN(n13738) );
  AOI21_X1 U15806 ( .B1(n14522), .B2(n13782), .A(n13738), .ZN(n13739) );
  OAI21_X1 U15807 ( .B1(n13740), .B2(n13784), .A(n13739), .ZN(P1_U3228) );
  XOR2_X1 U15808 ( .A(n13742), .B(n13741), .Z(n13747) );
  AND2_X1 U15809 ( .A1(n14284), .A2(n15200), .ZN(n14478) );
  AOI22_X1 U15810 ( .A1(n13776), .A2(n14278), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13744) );
  NAND2_X1 U15811 ( .A1(n13777), .A2(n14318), .ZN(n13743) );
  OAI211_X1 U15812 ( .C1(n13780), .C2(n14285), .A(n13744), .B(n13743), .ZN(
        n13745) );
  AOI21_X1 U15813 ( .B1(n14478), .B2(n13772), .A(n13745), .ZN(n13746) );
  OAI21_X1 U15814 ( .B1(n13747), .B2(n13784), .A(n13746), .ZN(P1_U3229) );
  AOI22_X1 U15815 ( .A1(n13777), .A2(n14345), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13749) );
  NAND2_X1 U15816 ( .A1(n13776), .A2(n14347), .ZN(n13748) );
  OAI211_X1 U15817 ( .C1(n13780), .C2(n13750), .A(n13749), .B(n13748), .ZN(
        n13755) );
  AOI211_X1 U15818 ( .C1(n13753), .C2(n13752), .A(n13784), .B(n13751), .ZN(
        n13754) );
  AOI211_X1 U15819 ( .C1(n13782), .C2(n7272), .A(n13755), .B(n13754), .ZN(
        n13756) );
  INV_X1 U15820 ( .A(n13756), .ZN(P1_U3233) );
  NAND2_X1 U15821 ( .A1(n14314), .A2(n15200), .ZN(n14492) );
  OAI21_X1 U15822 ( .B1(n13759), .B2(n13758), .A(n13757), .ZN(n13760) );
  NAND2_X1 U15823 ( .A1(n13760), .A2(n13790), .ZN(n13765) );
  INV_X1 U15824 ( .A(n14318), .ZN(n14176) );
  AOI22_X1 U15825 ( .A1(n13777), .A2(n14347), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13761) );
  OAI21_X1 U15826 ( .B1(n14176), .B2(n13762), .A(n13761), .ZN(n13763) );
  AOI21_X1 U15827 ( .B1(n14313), .B2(n13798), .A(n13763), .ZN(n13764) );
  OAI211_X1 U15828 ( .C1(n14492), .C2(n13766), .A(n13765), .B(n13764), .ZN(
        P1_U3235) );
  XOR2_X1 U15829 ( .A(n13768), .B(n13767), .Z(n13774) );
  INV_X1 U15830 ( .A(n14375), .ZN(n14376) );
  NOR2_X1 U15831 ( .A1(n14376), .A2(n15191), .ZN(n14515) );
  NAND2_X1 U15832 ( .A1(n14345), .A2(n15059), .ZN(n14371) );
  NAND2_X1 U15833 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15045)
         );
  OAI21_X1 U15834 ( .B1(n13795), .B2(n14371), .A(n15045), .ZN(n13769) );
  AOI21_X1 U15835 ( .B1(n13777), .B2(n14408), .A(n13769), .ZN(n13770) );
  OAI21_X1 U15836 ( .B1(n13780), .B2(n14377), .A(n13770), .ZN(n13771) );
  AOI21_X1 U15837 ( .B1(n14515), .B2(n13772), .A(n13771), .ZN(n13773) );
  OAI21_X1 U15838 ( .B1(n13774), .B2(n13784), .A(n13773), .ZN(P1_U3238) );
  AOI22_X1 U15839 ( .A1(n13776), .A2(n14246), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13779) );
  NAND2_X1 U15840 ( .A1(n13777), .A2(n14278), .ZN(n13778) );
  OAI211_X1 U15841 ( .C1(n13780), .C2(n14252), .A(n13779), .B(n13778), .ZN(
        n13781) );
  AOI21_X1 U15842 ( .B1(n14254), .B2(n13782), .A(n13781), .ZN(n13783) );
  OAI21_X1 U15843 ( .B1(n13785), .B2(n13784), .A(n13783), .ZN(P1_U3240) );
  INV_X1 U15844 ( .A(n13786), .ZN(n13791) );
  OAI21_X1 U15845 ( .B1(n13788), .B2(n13791), .A(n13787), .ZN(n13789) );
  OAI211_X1 U15846 ( .C1(n13792), .C2(n13791), .A(n13790), .B(n13789), .ZN(
        n13800) );
  OAI22_X1 U15847 ( .A1(n13795), .A2(n13794), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13793), .ZN(n13796) );
  AOI21_X1 U15848 ( .B1(n13798), .B2(n13797), .A(n13796), .ZN(n13799) );
  OAI211_X1 U15849 ( .C1(n13802), .C2(n13801), .A(n13800), .B(n13799), .ZN(
        P1_U3241) );
  INV_X1 U15850 ( .A(n14032), .ZN(n14049) );
  NOR2_X1 U15851 ( .A1(n14182), .A2(n14181), .ZN(n14200) );
  AOI21_X1 U15852 ( .B1(n14181), .B2(n14182), .A(n14200), .ZN(n14213) );
  INV_X1 U15853 ( .A(n14246), .ZN(n14180) );
  XNOR2_X1 U15854 ( .A(n14460), .B(n14180), .ZN(n14231) );
  INV_X1 U15855 ( .A(n14278), .ZN(n13803) );
  XNOR2_X1 U15856 ( .A(n14472), .B(n13803), .ZN(n14199) );
  INV_X1 U15857 ( .A(n14262), .ZN(n13804) );
  NAND2_X1 U15858 ( .A1(n14254), .A2(n13804), .ZN(n14179) );
  OR2_X1 U15859 ( .A1(n14254), .A2(n13804), .ZN(n13805) );
  INV_X1 U15860 ( .A(n14314), .ZN(n13806) );
  NAND2_X1 U15861 ( .A1(n13806), .A2(n14326), .ZN(n13807) );
  NAND2_X1 U15862 ( .A1(n14292), .A2(n13807), .ZN(n14309) );
  XNOR2_X1 U15863 ( .A(n14496), .B(n14175), .ZN(n14323) );
  XNOR2_X1 U15864 ( .A(n7272), .B(n14195), .ZN(n14339) );
  NOR2_X1 U15865 ( .A1(n14522), .A2(n14408), .ZN(n14188) );
  INV_X1 U15866 ( .A(n14188), .ZN(n13808) );
  NAND2_X1 U15867 ( .A1(n14522), .A2(n14408), .ZN(n14189) );
  NAND2_X1 U15868 ( .A1(n13808), .A2(n14189), .ZN(n14387) );
  NAND4_X1 U15869 ( .A1(n13810), .A2(n15137), .A3(n13885), .A4(n13809), .ZN(
        n13811) );
  NOR4_X1 U15870 ( .A1(n13813), .A2(n13812), .A3(n7821), .A4(n13811), .ZN(
        n13816) );
  NAND4_X1 U15871 ( .A1(n13817), .A2(n13816), .A3(n13815), .A4(n13814), .ZN(
        n13818) );
  NOR4_X1 U15872 ( .A1(n13820), .A2(n13819), .A3(n15054), .A4(n13818), .ZN(
        n13822) );
  XNOR2_X1 U15873 ( .A(n14414), .B(n14389), .ZN(n14404) );
  NAND4_X1 U15874 ( .A1(n14387), .A2(n13822), .A3(n14404), .A4(n13821), .ZN(
        n13824) );
  NOR2_X1 U15875 ( .A1(n13824), .A2(n13823), .ZN(n13825) );
  XNOR2_X1 U15876 ( .A(n14375), .B(n14390), .ZN(n14368) );
  NAND4_X1 U15877 ( .A1(n14356), .A2(n13825), .A3(n14368), .A4(n13951), .ZN(
        n13826) );
  NOR4_X1 U15878 ( .A1(n14309), .A2(n14323), .A3(n14339), .A4(n13826), .ZN(
        n13827) );
  XNOR2_X1 U15879 ( .A(n14304), .B(n14318), .ZN(n14299) );
  XNOR2_X1 U15880 ( .A(n14284), .B(n14295), .ZN(n14276) );
  NAND4_X1 U15881 ( .A1(n14248), .A2(n13827), .A3(n14299), .A4(n14276), .ZN(
        n13828) );
  NOR4_X1 U15882 ( .A1(n14213), .A2(n14231), .A3(n14199), .A4(n13828), .ZN(
        n13854) );
  NAND2_X1 U15883 ( .A1(n14560), .A2(n11615), .ZN(n13830) );
  INV_X1 U15884 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14555) );
  OR2_X1 U15885 ( .A1(n13850), .A2(n14555), .ZN(n13829) );
  NAND2_X1 U15886 ( .A1(n13830), .A2(n13829), .ZN(n14158) );
  NAND2_X1 U15887 ( .A1(n13831), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n13834) );
  NAND2_X1 U15888 ( .A1(n13832), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n13833) );
  OAI211_X1 U15889 ( .C1(n10037), .C2(n13835), .A(n13834), .B(n13833), .ZN(
        n14157) );
  XNOR2_X1 U15890 ( .A(n14158), .B(n14157), .ZN(n14037) );
  OR2_X1 U15891 ( .A1(n13850), .A2(n13838), .ZN(n13839) );
  INV_X1 U15892 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n13841) );
  OR2_X1 U15893 ( .A1(n10037), .A2(n13841), .ZN(n13847) );
  OR2_X1 U15894 ( .A1(n13842), .A2(n12290), .ZN(n13846) );
  INV_X1 U15895 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n13843) );
  OR2_X1 U15896 ( .A1(n13844), .A2(n13843), .ZN(n13845) );
  AND3_X1 U15897 ( .A1(n13847), .A2(n13846), .A3(n13845), .ZN(n14018) );
  INV_X1 U15898 ( .A(n14018), .ZN(n14204) );
  XNOR2_X1 U15899 ( .A(n14162), .B(n14204), .ZN(n13853) );
  NAND2_X1 U15900 ( .A1(n13848), .A2(n11615), .ZN(n13852) );
  OR2_X1 U15901 ( .A1(n13850), .A2(n13849), .ZN(n13851) );
  NAND2_X1 U15902 ( .A1(n13852), .A2(n13851), .ZN(n14151) );
  XNOR2_X1 U15903 ( .A(n14151), .B(n14215), .ZN(n14201) );
  NAND4_X1 U15904 ( .A1(n13854), .A2(n14037), .A3(n13853), .A4(n14201), .ZN(
        n13855) );
  XOR2_X1 U15905 ( .A(n14265), .B(n13855), .Z(n14048) );
  NAND2_X1 U15906 ( .A1(n13857), .A2(n13856), .ZN(n13860) );
  NAND2_X1 U15907 ( .A1(n10212), .A2(n15140), .ZN(n13858) );
  NAND2_X1 U15908 ( .A1(n13860), .A2(n13859), .ZN(n13867) );
  NAND2_X1 U15909 ( .A1(n13865), .A2(n13862), .ZN(n14019) );
  NAND2_X1 U15910 ( .A1(n13865), .A2(n13864), .ZN(n13866) );
  NAND2_X1 U15911 ( .A1(n13867), .A2(n14021), .ZN(n13870) );
  NAND2_X1 U15912 ( .A1(n13868), .A2(n14029), .ZN(n13869) );
  NAND2_X1 U15913 ( .A1(n13870), .A2(n13869), .ZN(n13874) );
  MUX2_X1 U15914 ( .A(n13872), .B(n13871), .S(n14029), .Z(n13873) );
  NAND2_X1 U15915 ( .A1(n13874), .A2(n13873), .ZN(n13881) );
  NAND2_X1 U15916 ( .A1(n13881), .A2(n13879), .ZN(n13878) );
  MUX2_X1 U15917 ( .A(n13876), .B(n15156), .S(n14021), .Z(n13877) );
  NAND2_X1 U15918 ( .A1(n13878), .A2(n13877), .ZN(n13886) );
  INV_X1 U15919 ( .A(n13879), .ZN(n13883) );
  NOR2_X1 U15920 ( .A1(n13881), .A2(n15156), .ZN(n13882) );
  NAND2_X1 U15921 ( .A1(n13883), .A2(n13882), .ZN(n13884) );
  NAND3_X1 U15922 ( .A1(n13886), .A2(n13885), .A3(n13884), .ZN(n13890) );
  NAND2_X1 U15923 ( .A1(n15163), .A2(n14065), .ZN(n13887) );
  MUX2_X1 U15924 ( .A(n13888), .B(n13887), .S(n14029), .Z(n13889) );
  MUX2_X1 U15925 ( .A(n13892), .B(n13891), .S(n14021), .Z(n13894) );
  MUX2_X1 U15926 ( .A(n14064), .B(n7261), .S(n14021), .Z(n13893) );
  NAND3_X1 U15927 ( .A1(n13897), .A2(n13896), .A3(n13895), .ZN(n13902) );
  AND2_X1 U15928 ( .A1(n14021), .A2(n14063), .ZN(n13900) );
  OAI21_X1 U15929 ( .B1(n14063), .B2(n14021), .A(n13899), .ZN(n13898) );
  OAI21_X1 U15930 ( .B1(n13900), .B2(n13899), .A(n13898), .ZN(n13901) );
  MUX2_X1 U15931 ( .A(n14062), .B(n15084), .S(n14029), .Z(n13904) );
  MUX2_X1 U15932 ( .A(n14062), .B(n15084), .S(n14021), .Z(n13903) );
  MUX2_X1 U15933 ( .A(n14061), .B(n13906), .S(n14021), .Z(n13909) );
  MUX2_X1 U15934 ( .A(n13906), .B(n14061), .S(n14021), .Z(n13907) );
  NAND2_X1 U15935 ( .A1(n13908), .A2(n13907), .ZN(n13912) );
  INV_X1 U15936 ( .A(n13909), .ZN(n13910) );
  MUX2_X1 U15937 ( .A(n14060), .B(n13913), .S(n14029), .Z(n13915) );
  MUX2_X1 U15938 ( .A(n14060), .B(n13913), .S(n14021), .Z(n13914) );
  MUX2_X1 U15939 ( .A(n15050), .B(n13917), .S(n14021), .Z(n13919) );
  MUX2_X1 U15940 ( .A(n15050), .B(n13917), .S(n14029), .Z(n13918) );
  INV_X1 U15941 ( .A(n13919), .ZN(n13920) );
  MUX2_X1 U15942 ( .A(n14059), .B(n15201), .S(n14029), .Z(n13923) );
  MUX2_X1 U15943 ( .A(n14059), .B(n15201), .S(n14021), .Z(n13921) );
  MUX2_X1 U15944 ( .A(n15060), .B(n13924), .S(n14021), .Z(n13927) );
  MUX2_X1 U15945 ( .A(n13925), .B(n14952), .S(n14029), .Z(n13926) );
  MUX2_X1 U15946 ( .A(n13929), .B(n14797), .S(n14021), .Z(n13937) );
  MUX2_X1 U15947 ( .A(n14058), .B(n13930), .S(n14029), .Z(n13936) );
  AND2_X1 U15948 ( .A1(n14166), .A2(n13933), .ZN(n13953) );
  MUX2_X1 U15949 ( .A(n14057), .B(n13934), .S(n14021), .Z(n13945) );
  OR2_X1 U15950 ( .A1(n13934), .A2(n14021), .ZN(n13946) );
  NAND2_X1 U15951 ( .A1(n14021), .A2(n13935), .ZN(n13949) );
  NAND2_X1 U15952 ( .A1(n13946), .A2(n13949), .ZN(n13940) );
  INV_X1 U15953 ( .A(n13936), .ZN(n13939) );
  INV_X1 U15954 ( .A(n13937), .ZN(n13938) );
  OAI22_X1 U15955 ( .A1(n13945), .A2(n13940), .B1(n13939), .B2(n13938), .ZN(
        n13941) );
  INV_X1 U15956 ( .A(n13941), .ZN(n13943) );
  AND2_X1 U15957 ( .A1(n13944), .A2(n13942), .ZN(n13947) );
  MUX2_X1 U15958 ( .A(n13944), .B(n14166), .S(n14029), .Z(n13956) );
  INV_X1 U15959 ( .A(n13945), .ZN(n13950) );
  OAI22_X1 U15960 ( .A1(n13951), .A2(n14021), .B1(n13950), .B2(n13946), .ZN(
        n13948) );
  NAND2_X1 U15961 ( .A1(n13948), .A2(n13947), .ZN(n13955) );
  OAI22_X1 U15962 ( .A1(n13951), .A2(n14029), .B1(n13950), .B2(n13949), .ZN(
        n13952) );
  NAND2_X1 U15963 ( .A1(n13953), .A2(n13952), .ZN(n13954) );
  MUX2_X1 U15964 ( .A(n14389), .B(n14414), .S(n14021), .Z(n13960) );
  MUX2_X1 U15965 ( .A(n14389), .B(n14414), .S(n14029), .Z(n13957) );
  NAND2_X1 U15966 ( .A1(n13958), .A2(n13957), .ZN(n13964) );
  INV_X1 U15967 ( .A(n13960), .ZN(n13961) );
  INV_X1 U15968 ( .A(n14522), .ZN(n14397) );
  MUX2_X1 U15969 ( .A(n14171), .B(n14397), .S(n14029), .Z(n13965) );
  XNOR2_X1 U15970 ( .A(n14390), .B(n14029), .ZN(n13967) );
  XNOR2_X1 U15971 ( .A(n14375), .B(n14021), .ZN(n13966) );
  OAI21_X1 U15972 ( .B1(n13968), .B2(n13967), .A(n13966), .ZN(n13970) );
  NAND2_X1 U15973 ( .A1(n13968), .A2(n13967), .ZN(n13969) );
  OR2_X1 U15974 ( .A1(n14358), .A2(n14029), .ZN(n13972) );
  NAND2_X1 U15975 ( .A1(n14358), .A2(n14029), .ZN(n13971) );
  MUX2_X1 U15976 ( .A(n13972), .B(n13971), .S(n14172), .Z(n13973) );
  MUX2_X1 U15977 ( .A(n14195), .B(n14502), .S(n14021), .Z(n13975) );
  MUX2_X1 U15978 ( .A(n7272), .B(n14173), .S(n14021), .Z(n13974) );
  MUX2_X1 U15979 ( .A(n14347), .B(n14496), .S(n14029), .Z(n13977) );
  MUX2_X1 U15980 ( .A(n14347), .B(n14496), .S(n14021), .Z(n13976) );
  MUX2_X1 U15981 ( .A(n14326), .B(n14314), .S(n14021), .Z(n13979) );
  MUX2_X1 U15982 ( .A(n14326), .B(n14314), .S(n14029), .Z(n13978) );
  MUX2_X1 U15983 ( .A(n14318), .B(n14304), .S(n14029), .Z(n13981) );
  MUX2_X1 U15984 ( .A(n14318), .B(n14304), .S(n14021), .Z(n13980) );
  MUX2_X1 U15985 ( .A(n14295), .B(n14284), .S(n14021), .Z(n13986) );
  MUX2_X1 U15986 ( .A(n14295), .B(n14284), .S(n14029), .Z(n13983) );
  NAND2_X1 U15987 ( .A1(n13984), .A2(n13983), .ZN(n13990) );
  INV_X1 U15988 ( .A(n13985), .ZN(n13988) );
  INV_X1 U15989 ( .A(n13986), .ZN(n13987) );
  MUX2_X1 U15990 ( .A(n14278), .B(n14472), .S(n14029), .Z(n13992) );
  MUX2_X1 U15991 ( .A(n14278), .B(n14472), .S(n14021), .Z(n13991) );
  MUX2_X1 U15992 ( .A(n14262), .B(n14254), .S(n14021), .Z(n13994) );
  MUX2_X1 U15993 ( .A(n14262), .B(n14254), .S(n14029), .Z(n13993) );
  INV_X1 U15994 ( .A(n13994), .ZN(n13995) );
  MUX2_X1 U15995 ( .A(n14246), .B(n14460), .S(n14029), .Z(n13999) );
  NAND2_X1 U15996 ( .A1(n13998), .A2(n13999), .ZN(n13997) );
  MUX2_X1 U15997 ( .A(n14246), .B(n14460), .S(n14021), .Z(n13996) );
  NAND2_X1 U15998 ( .A1(n13997), .A2(n13996), .ZN(n14003) );
  INV_X1 U15999 ( .A(n13999), .ZN(n14000) );
  NAND2_X1 U16000 ( .A1(n14001), .A2(n14000), .ZN(n14002) );
  MUX2_X1 U16001 ( .A(n14233), .B(n14452), .S(n14021), .Z(n14005) );
  MUX2_X1 U16002 ( .A(n14233), .B(n14452), .S(n14029), .Z(n14004) );
  INV_X1 U16003 ( .A(n14005), .ZN(n14006) );
  MUX2_X1 U16004 ( .A(n14215), .B(n14151), .S(n14029), .Z(n14010) );
  NAND2_X1 U16005 ( .A1(n14009), .A2(n14010), .ZN(n14008) );
  MUX2_X1 U16006 ( .A(n14215), .B(n14151), .S(n14021), .Z(n14007) );
  INV_X1 U16007 ( .A(n14009), .ZN(n14012) );
  INV_X1 U16008 ( .A(n14010), .ZN(n14011) );
  INV_X1 U16009 ( .A(n14157), .ZN(n14017) );
  AOI21_X1 U16010 ( .B1(n14017), .B2(n14015), .A(n14018), .ZN(n14016) );
  MUX2_X1 U16011 ( .A(n14016), .B(n14162), .S(n14029), .Z(n14028) );
  OR2_X1 U16012 ( .A1(n14021), .A2(n14017), .ZN(n14031) );
  AOI21_X1 U16013 ( .B1(n14031), .B2(n14019), .A(n14018), .ZN(n14020) );
  AOI21_X1 U16014 ( .B1(n14162), .B2(n14021), .A(n14020), .ZN(n14027) );
  NAND2_X1 U16015 ( .A1(n14023), .A2(n14022), .ZN(n14025) );
  AND2_X1 U16016 ( .A1(n14025), .A2(n14024), .ZN(n14040) );
  NAND2_X1 U16017 ( .A1(n14037), .A2(n14040), .ZN(n14043) );
  INV_X1 U16018 ( .A(n14043), .ZN(n14026) );
  OR2_X1 U16019 ( .A1(n14028), .A2(n14027), .ZN(n14042) );
  INV_X1 U16020 ( .A(n14042), .ZN(n14034) );
  INV_X1 U16021 ( .A(n14040), .ZN(n14033) );
  AND2_X1 U16022 ( .A1(n14033), .A2(n14032), .ZN(n14035) );
  NAND2_X1 U16023 ( .A1(n14038), .A2(n14035), .ZN(n14044) );
  INV_X1 U16024 ( .A(n14035), .ZN(n14036) );
  NOR2_X1 U16025 ( .A1(n14037), .A2(n14036), .ZN(n14039) );
  MUX2_X1 U16026 ( .A(n14040), .B(n14039), .S(n14038), .Z(n14041) );
  INV_X1 U16027 ( .A(n14041), .ZN(n14047) );
  OAI22_X1 U16028 ( .A1(n14044), .A2(n6623), .B1(n14043), .B2(n14042), .ZN(
        n14045) );
  INV_X1 U16029 ( .A(n14045), .ZN(n14046) );
  NAND4_X1 U16030 ( .A1(n14052), .A2(n14051), .A3(n15049), .A4(n14050), .ZN(
        n14053) );
  OAI211_X1 U16031 ( .C1(n13861), .C2(n14055), .A(n14053), .B(P1_B_REG_SCAN_IN), .ZN(n14054) );
  OAI21_X1 U16032 ( .B1(n6706), .B2(n14055), .A(n14054), .ZN(P1_U3242) );
  MUX2_X1 U16033 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14157), .S(n14081), .Z(
        P1_U3591) );
  MUX2_X1 U16034 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14204), .S(n14081), .Z(
        P1_U3590) );
  MUX2_X1 U16035 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14215), .S(n14081), .Z(
        P1_U3589) );
  MUX2_X1 U16036 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14233), .S(n14081), .Z(
        P1_U3588) );
  MUX2_X1 U16037 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14246), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16038 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14262), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16039 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14278), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16040 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14295), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16041 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14318), .S(n14081), .Z(
        P1_U3583) );
  MUX2_X1 U16042 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14326), .S(n14081), .Z(
        P1_U3582) );
  MUX2_X1 U16043 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14347), .S(n14081), .Z(
        P1_U3581) );
  MUX2_X1 U16044 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14173), .S(n14081), .Z(
        P1_U3580) );
  MUX2_X1 U16045 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14345), .S(n14081), .Z(
        P1_U3579) );
  MUX2_X1 U16046 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14390), .S(n14081), .Z(
        P1_U3578) );
  MUX2_X1 U16047 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14408), .S(n14081), .Z(
        P1_U3577) );
  MUX2_X1 U16048 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14389), .S(n14081), .Z(
        P1_U3576) );
  MUX2_X1 U16049 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14409), .S(n14081), .Z(
        P1_U3575) );
  MUX2_X1 U16050 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14056), .S(n14081), .Z(
        P1_U3574) );
  MUX2_X1 U16051 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14057), .S(n14081), .Z(
        P1_U3573) );
  MUX2_X1 U16052 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14058), .S(n14081), .Z(
        P1_U3572) );
  MUX2_X1 U16053 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15060), .S(n14081), .Z(
        P1_U3571) );
  MUX2_X1 U16054 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14059), .S(n14081), .Z(
        P1_U3570) );
  MUX2_X1 U16055 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n15050), .S(n14081), .Z(
        P1_U3569) );
  MUX2_X1 U16056 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14060), .S(n14081), .Z(
        P1_U3568) );
  MUX2_X1 U16057 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14061), .S(n14081), .Z(
        P1_U3567) );
  MUX2_X1 U16058 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14062), .S(n14081), .Z(
        P1_U3566) );
  MUX2_X1 U16059 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14063), .S(n14081), .Z(
        P1_U3565) );
  MUX2_X1 U16060 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14064), .S(n14081), .Z(
        P1_U3564) );
  MUX2_X1 U16061 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14065), .S(n14081), .Z(
        P1_U3563) );
  MUX2_X1 U16062 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14434), .S(n14081), .Z(
        P1_U3562) );
  MUX2_X1 U16063 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14066), .S(n14081), .Z(
        P1_U3561) );
  MUX2_X1 U16064 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n10212), .S(n14081), .Z(
        P1_U3560) );
  INV_X1 U16065 ( .A(n14069), .ZN(n14068) );
  OAI22_X1 U16066 ( .A1(n15047), .A2(n14668), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7471), .ZN(n14067) );
  AOI21_X1 U16067 ( .B1(n14068), .B2(n15012), .A(n14067), .ZN(n14076) );
  MUX2_X1 U16068 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10015), .S(n14069), .Z(
        n14070) );
  OAI21_X1 U16069 ( .B1(n9992), .B2(n14071), .A(n14070), .ZN(n14072) );
  NAND3_X1 U16070 ( .A1(n15028), .A2(n14090), .A3(n14072), .ZN(n14075) );
  OAI211_X1 U16071 ( .C1(n14078), .C2(n14073), .A(n15024), .B(n14084), .ZN(
        n14074) );
  NAND3_X1 U16072 ( .A1(n14076), .A2(n14075), .A3(n14074), .ZN(P1_U3244) );
  MUX2_X1 U16073 ( .A(n14078), .B(n14077), .S(n6573), .Z(n14080) );
  NAND2_X1 U16074 ( .A1(n14080), .A2(n14079), .ZN(n14082) );
  OAI211_X1 U16075 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n6761), .A(n14082), .B(
        n14081), .ZN(n15000) );
  AOI22_X1 U16076 ( .A1(n15018), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14095) );
  MUX2_X1 U16077 ( .A(n10039), .B(P1_REG2_REG_2__SCAN_IN), .S(n14088), .Z(
        n14085) );
  NAND3_X1 U16078 ( .A1(n14085), .A2(n14084), .A3(n14083), .ZN(n14086) );
  AND3_X1 U16079 ( .A1(n15024), .A2(n14104), .A3(n14086), .ZN(n14087) );
  AOI21_X1 U16080 ( .B1(n15012), .B2(n14088), .A(n14087), .ZN(n14094) );
  MUX2_X1 U16081 ( .A(n9754), .B(P1_REG1_REG_2__SCAN_IN), .S(n14088), .Z(
        n14091) );
  NAND3_X1 U16082 ( .A1(n14091), .A2(n14090), .A3(n14089), .ZN(n14092) );
  NAND3_X1 U16083 ( .A1(n15028), .A2(n14099), .A3(n14092), .ZN(n14093) );
  NAND4_X1 U16084 ( .A1(n15000), .A2(n14095), .A3(n14094), .A4(n14093), .ZN(
        P1_U3245) );
  OAI22_X1 U16085 ( .A1(n15047), .A2(n14712), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14096), .ZN(n14097) );
  AOI21_X1 U16086 ( .B1(n14102), .B2(n15012), .A(n14097), .ZN(n14109) );
  MUX2_X1 U16087 ( .A(n10079), .B(P1_REG1_REG_3__SCAN_IN), .S(n14102), .Z(
        n14100) );
  NAND3_X1 U16088 ( .A1(n14100), .A2(n14099), .A3(n14098), .ZN(n14101) );
  NAND3_X1 U16089 ( .A1(n15028), .A2(n14991), .A3(n14101), .ZN(n14108) );
  MUX2_X1 U16090 ( .A(n10080), .B(P1_REG2_REG_3__SCAN_IN), .S(n14102), .Z(
        n14105) );
  NAND3_X1 U16091 ( .A1(n14105), .A2(n14104), .A3(n14103), .ZN(n14106) );
  NAND3_X1 U16092 ( .A1(n15024), .A2(n14985), .A3(n14106), .ZN(n14107) );
  NAND3_X1 U16093 ( .A1(n14109), .A2(n14108), .A3(n14107), .ZN(P1_U3246) );
  INV_X1 U16094 ( .A(n14110), .ZN(n14115) );
  NOR3_X1 U16095 ( .A1(n14113), .A2(n14112), .A3(n14111), .ZN(n14114) );
  OAI21_X1 U16096 ( .B1(n14115), .B2(n14114), .A(n15028), .ZN(n14126) );
  AOI21_X1 U16097 ( .B1(n15018), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n14116), .ZN(
        n14125) );
  MUX2_X1 U16098 ( .A(n11051), .B(P1_REG2_REG_9__SCAN_IN), .S(n14122), .Z(
        n14117) );
  NAND3_X1 U16099 ( .A1(n14119), .A2(n14118), .A3(n14117), .ZN(n14120) );
  NAND3_X1 U16100 ( .A1(n15024), .A2(n14121), .A3(n14120), .ZN(n14124) );
  NAND2_X1 U16101 ( .A1(n15012), .A2(n14122), .ZN(n14123) );
  NAND4_X1 U16102 ( .A1(n14126), .A2(n14125), .A3(n14124), .A4(n14123), .ZN(
        P1_U3252) );
  INV_X1 U16103 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14129) );
  OAI21_X1 U16104 ( .B1(n14129), .B2(n14128), .A(n14127), .ZN(n14130) );
  XOR2_X1 U16105 ( .A(n14139), .B(n14130), .Z(n15035) );
  NAND2_X1 U16106 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n15035), .ZN(n15034) );
  NAND2_X1 U16107 ( .A1(n14139), .A2(n14130), .ZN(n14131) );
  NAND2_X1 U16108 ( .A1(n15034), .A2(n14131), .ZN(n14132) );
  XOR2_X1 U16109 ( .A(n14132), .B(P1_REG1_REG_19__SCAN_IN), .Z(n14146) );
  INV_X1 U16110 ( .A(n14133), .ZN(n14134) );
  NAND2_X1 U16111 ( .A1(n14135), .A2(n14134), .ZN(n14136) );
  NAND2_X1 U16112 ( .A1(n14137), .A2(n14136), .ZN(n14138) );
  NAND2_X1 U16113 ( .A1(n14139), .A2(n14138), .ZN(n14140) );
  XOR2_X1 U16114 ( .A(n14139), .B(n14138), .Z(n15037) );
  NAND2_X1 U16115 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n15037), .ZN(n15036) );
  NAND2_X1 U16116 ( .A1(n14140), .A2(n15036), .ZN(n14141) );
  XOR2_X1 U16117 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14141), .Z(n14145) );
  INV_X1 U16118 ( .A(n14145), .ZN(n14142) );
  NAND2_X1 U16119 ( .A1(n14142), .A2(n15024), .ZN(n14143) );
  OAI211_X1 U16120 ( .C1(n14146), .C2(n15041), .A(n14143), .B(n15043), .ZN(
        n14144) );
  INV_X1 U16121 ( .A(n14144), .ZN(n14148) );
  AOI22_X1 U16122 ( .A1(n14146), .A2(n15028), .B1(n15024), .B2(n14145), .ZN(
        n14147) );
  MUX2_X1 U16123 ( .A(n14148), .B(n14147), .S(n14265), .Z(n14150) );
  NAND2_X1 U16124 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n14149)
         );
  OAI211_X1 U16125 ( .C1(n7911), .C2(n15047), .A(n14150), .B(n14149), .ZN(
        P1_U3262) );
  INV_X1 U16126 ( .A(n14254), .ZN(n14465) );
  NAND2_X1 U16127 ( .A1(n14447), .A2(n14218), .ZN(n14202) );
  NOR2_X1 U16128 ( .A1(n14202), .A2(n14162), .ZN(n14152) );
  XNOR2_X1 U16129 ( .A(n14152), .B(n14158), .ZN(n14153) );
  NAND2_X1 U16130 ( .A1(n14153), .A2(n15076), .ZN(n14439) );
  INV_X1 U16131 ( .A(P1_B_REG_SCAN_IN), .ZN(n14154) );
  NOR2_X1 U16132 ( .A1(n6573), .A2(n14154), .ZN(n14155) );
  NOR2_X1 U16133 ( .A1(n14156), .A2(n14155), .ZN(n14203) );
  NAND2_X1 U16134 ( .A1(n14203), .A2(n14157), .ZN(n14441) );
  NOR2_X1 U16135 ( .A1(n15093), .A2(n14441), .ZN(n14164) );
  INV_X1 U16136 ( .A(n14158), .ZN(n14440) );
  NOR2_X1 U16137 ( .A1(n14440), .A2(n15096), .ZN(n14159) );
  AOI211_X1 U16138 ( .C1(n15105), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14164), 
        .B(n14159), .ZN(n14160) );
  OAI21_X1 U16139 ( .B1(n14439), .B2(n15087), .A(n14160), .ZN(P1_U3263) );
  XOR2_X1 U16140 ( .A(n14162), .B(n14202), .Z(n14161) );
  NAND2_X1 U16141 ( .A1(n14161), .A2(n15076), .ZN(n14442) );
  INV_X1 U16142 ( .A(n14162), .ZN(n14443) );
  NOR2_X1 U16143 ( .A1(n14443), .A2(n15096), .ZN(n14163) );
  AOI211_X1 U16144 ( .C1(n15105), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14164), 
        .B(n14163), .ZN(n14165) );
  OAI21_X1 U16145 ( .B1(n15087), .B2(n14442), .A(n14165), .ZN(P1_U3264) );
  INV_X1 U16146 ( .A(n14295), .ZN(n14177) );
  INV_X1 U16147 ( .A(n14166), .ZN(n14167) );
  INV_X1 U16148 ( .A(n14339), .ZN(n14341) );
  NAND2_X1 U16149 ( .A1(n14502), .A2(n14173), .ZN(n14174) );
  INV_X1 U16150 ( .A(n14323), .ZN(n14334) );
  INV_X1 U16151 ( .A(n14299), .ZN(n14293) );
  INV_X1 U16152 ( .A(n14472), .ZN(n14178) );
  OR2_X1 U16153 ( .A1(n14534), .A2(n14409), .ZN(n14183) );
  INV_X1 U16154 ( .A(n14404), .ZN(n14185) );
  OR2_X1 U16155 ( .A1(n14414), .A2(n14389), .ZN(n14186) );
  AND2_X1 U16156 ( .A1(n14375), .A2(n14390), .ZN(n14191) );
  OR2_X1 U16157 ( .A1(n14375), .A2(n14390), .ZN(n14190) );
  INV_X1 U16158 ( .A(n14356), .ZN(n14192) );
  NAND2_X1 U16159 ( .A1(n14355), .A2(n14192), .ZN(n14194) );
  OR2_X1 U16160 ( .A1(n14358), .A2(n14345), .ZN(n14193) );
  OR2_X1 U16161 ( .A1(n14502), .A2(n14195), .ZN(n14196) );
  OR2_X1 U16162 ( .A1(n14496), .A2(n14347), .ZN(n14197) );
  NAND2_X1 U16163 ( .A1(n14304), .A2(n14318), .ZN(n14198) );
  INV_X1 U16164 ( .A(n14213), .ZN(n14219) );
  OAI21_X1 U16165 ( .B1(n14447), .B2(n14218), .A(n14202), .ZN(n14444) );
  NOR2_X1 U16166 ( .A1(n14444), .A2(n14422), .ZN(n14211) );
  NAND2_X1 U16167 ( .A1(n14204), .A2(n14203), .ZN(n14446) );
  OAI22_X1 U16168 ( .A1(n14206), .A2(n14446), .B1(n14205), .B2(n15080), .ZN(
        n14208) );
  NAND2_X1 U16169 ( .A1(n14233), .A2(n15049), .ZN(n14445) );
  NOR2_X1 U16170 ( .A1(n15093), .A2(n14445), .ZN(n14207) );
  AOI211_X1 U16171 ( .C1(n15105), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14208), 
        .B(n14207), .ZN(n14209) );
  OAI21_X1 U16172 ( .B1(n14447), .B2(n15096), .A(n14209), .ZN(n14210) );
  OAI21_X1 U16173 ( .B1(n14449), .B2(n14273), .A(n14212), .ZN(P1_U3356) );
  XNOR2_X1 U16174 ( .A(n14214), .B(n14213), .ZN(n14216) );
  AND2_X1 U16175 ( .A1(n14452), .A2(n14236), .ZN(n14217) );
  OR3_X1 U16176 ( .A1(n14218), .A2(n14217), .A3(n15147), .ZN(n14454) );
  NAND2_X1 U16177 ( .A1(n14220), .A2(n14219), .ZN(n14453) );
  NAND3_X1 U16178 ( .A1(n6612), .A2(n15065), .A3(n14453), .ZN(n14225) );
  NAND2_X1 U16179 ( .A1(n15093), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14221) );
  OAI21_X1 U16180 ( .B1(n15080), .B2(n14222), .A(n14221), .ZN(n14223) );
  AOI21_X1 U16181 ( .B1(n14452), .B2(n15085), .A(n14223), .ZN(n14224) );
  OAI211_X1 U16182 ( .C1(n15087), .C2(n14454), .A(n14225), .B(n14224), .ZN(
        n14226) );
  INV_X1 U16183 ( .A(n14226), .ZN(n14227) );
  OAI21_X1 U16184 ( .B1(n14457), .B2(n15093), .A(n14227), .ZN(P1_U3265) );
  OAI21_X1 U16185 ( .B1(n14229), .B2(n14231), .A(n14228), .ZN(n14458) );
  AOI21_X1 U16186 ( .B1(n14232), .B2(n14231), .A(n14230), .ZN(n14235) );
  AOI22_X1 U16187 ( .A1(n15049), .A2(n14262), .B1(n14233), .B2(n15059), .ZN(
        n14234) );
  INV_X1 U16188 ( .A(n14460), .ZN(n14241) );
  AOI211_X1 U16189 ( .C1(n14460), .C2(n14250), .A(n15147), .B(n7258), .ZN(
        n14459) );
  NAND2_X1 U16190 ( .A1(n14459), .A2(n15063), .ZN(n14240) );
  INV_X1 U16191 ( .A(n14237), .ZN(n14238) );
  AOI22_X1 U16192 ( .A1(n15093), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14238), 
        .B2(n15091), .ZN(n14239) );
  OAI211_X1 U16193 ( .C1(n14241), .C2(n15096), .A(n14240), .B(n14239), .ZN(
        n14242) );
  AOI21_X1 U16194 ( .B1(n14458), .B2(n15100), .A(n14242), .ZN(n14243) );
  OAI21_X1 U16195 ( .B1(n14462), .B2(n15093), .A(n14243), .ZN(P1_U3266) );
  OAI21_X1 U16196 ( .B1(n14248), .B2(n14245), .A(n14244), .ZN(n14247) );
  AOI222_X1 U16197 ( .A1(n14247), .A2(n15196), .B1(n14246), .B2(n15059), .C1(
        n14278), .C2(n15049), .ZN(n14469) );
  AOI21_X1 U16198 ( .B1(n14249), .B2(n14248), .A(n6670), .ZN(n14467) );
  OAI211_X1 U16199 ( .C1(n14465), .C2(n14261), .A(n15076), .B(n14250), .ZN(
        n14464) );
  NAND2_X1 U16200 ( .A1(n15105), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n14251) );
  OAI21_X1 U16201 ( .B1(n15080), .B2(n14252), .A(n14251), .ZN(n14253) );
  AOI21_X1 U16202 ( .B1(n14254), .B2(n15085), .A(n14253), .ZN(n14255) );
  OAI21_X1 U16203 ( .B1(n14464), .B2(n15087), .A(n14255), .ZN(n14256) );
  AOI21_X1 U16204 ( .B1(n14467), .B2(n15065), .A(n14256), .ZN(n14257) );
  OAI21_X1 U16205 ( .B1(n14469), .B2(n15093), .A(n14257), .ZN(P1_U3267) );
  XNOR2_X1 U16206 ( .A(n14258), .B(n14260), .ZN(n14476) );
  AOI21_X1 U16207 ( .B1(n14260), .B2(n14259), .A(n6669), .ZN(n14473) );
  AOI211_X1 U16208 ( .C1(n14472), .C2(n14282), .A(n15147), .B(n14261), .ZN(
        n14470) );
  NAND2_X1 U16209 ( .A1(n14295), .A2(n15049), .ZN(n14264) );
  NAND2_X1 U16210 ( .A1(n14262), .A2(n15059), .ZN(n14263) );
  NAND2_X1 U16211 ( .A1(n14264), .A2(n14263), .ZN(n14471) );
  AOI21_X1 U16212 ( .B1(n14470), .B2(n14265), .A(n14471), .ZN(n14270) );
  OAI22_X1 U16213 ( .A1(n14379), .A2(n14267), .B1(n14266), .B2(n15080), .ZN(
        n14268) );
  AOI21_X1 U16214 ( .B1(n14472), .B2(n15085), .A(n14268), .ZN(n14269) );
  OAI21_X1 U16215 ( .B1(n14270), .B2(n15093), .A(n14269), .ZN(n14271) );
  AOI21_X1 U16216 ( .B1(n14473), .B2(n15065), .A(n14271), .ZN(n14272) );
  OAI21_X1 U16217 ( .B1(n14476), .B2(n14273), .A(n14272), .ZN(P1_U3268) );
  XNOR2_X1 U16218 ( .A(n14274), .B(n14276), .ZN(n14477) );
  OAI211_X1 U16219 ( .C1(n14277), .C2(n14276), .A(n14275), .B(n15196), .ZN(
        n14280) );
  AOI22_X1 U16220 ( .A1(n15049), .A2(n14318), .B1(n14278), .B2(n15059), .ZN(
        n14279) );
  NAND2_X1 U16221 ( .A1(n14280), .A2(n14279), .ZN(n14281) );
  AOI21_X1 U16222 ( .B1(n15074), .B2(n14477), .A(n14281), .ZN(n14481) );
  INV_X1 U16223 ( .A(n14282), .ZN(n14283) );
  AOI211_X1 U16224 ( .C1(n14284), .C2(n14297), .A(n15147), .B(n14283), .ZN(
        n14479) );
  NOR2_X1 U16225 ( .A1(n7600), .A2(n15096), .ZN(n14288) );
  OAI22_X1 U16226 ( .A1(n14379), .A2(n14286), .B1(n14285), .B2(n15080), .ZN(
        n14287) );
  AOI211_X1 U16227 ( .C1(n14479), .C2(n15063), .A(n14288), .B(n14287), .ZN(
        n14290) );
  NAND2_X1 U16228 ( .A1(n14477), .A2(n15100), .ZN(n14289) );
  OAI211_X1 U16229 ( .C1(n14481), .C2(n15093), .A(n14290), .B(n14289), .ZN(
        P1_U3269) );
  NAND3_X1 U16230 ( .A1(n14291), .A2(n14293), .A3(n14292), .ZN(n14294) );
  NAND2_X1 U16231 ( .A1(n6676), .A2(n14294), .ZN(n14296) );
  AOI222_X1 U16232 ( .A1(n14296), .A2(n15196), .B1(n14295), .B2(n15059), .C1(
        n14326), .C2(n15049), .ZN(n14489) );
  AOI21_X1 U16233 ( .B1(n14311), .B2(n14304), .A(n15147), .ZN(n14298) );
  NAND2_X1 U16234 ( .A1(n14298), .A2(n14297), .ZN(n14486) );
  NAND2_X1 U16235 ( .A1(n14300), .A2(n14299), .ZN(n14484) );
  NAND3_X1 U16236 ( .A1(n14485), .A2(n14484), .A3(n15065), .ZN(n14306) );
  NAND2_X1 U16237 ( .A1(n15105), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n14301) );
  OAI21_X1 U16238 ( .B1(n15080), .B2(n14302), .A(n14301), .ZN(n14303) );
  AOI21_X1 U16239 ( .B1(n14304), .B2(n15085), .A(n14303), .ZN(n14305) );
  OAI211_X1 U16240 ( .C1(n14486), .C2(n15087), .A(n14306), .B(n14305), .ZN(
        n14307) );
  INV_X1 U16241 ( .A(n14307), .ZN(n14308) );
  OAI21_X1 U16242 ( .B1(n14489), .B2(n15093), .A(n14308), .ZN(P1_U3270) );
  XNOR2_X1 U16243 ( .A(n14310), .B(n14309), .ZN(n14490) );
  AOI21_X1 U16244 ( .B1(n14327), .B2(n14314), .A(n15147), .ZN(n14312) );
  NAND2_X1 U16245 ( .A1(n14312), .A2(n14311), .ZN(n14491) );
  AOI22_X1 U16246 ( .A1(n15093), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14313), 
        .B2(n15091), .ZN(n14316) );
  NAND2_X1 U16247 ( .A1(n14314), .A2(n15085), .ZN(n14315) );
  OAI211_X1 U16248 ( .C1(n14491), .C2(n15087), .A(n14316), .B(n14315), .ZN(
        n14321) );
  OAI21_X1 U16249 ( .B1(n6947), .B2(n14317), .A(n14291), .ZN(n14319) );
  AOI222_X1 U16250 ( .A1(n14319), .A2(n15196), .B1(n14318), .B2(n15059), .C1(
        n14347), .C2(n15049), .ZN(n14494) );
  NOR2_X1 U16251 ( .A1(n14494), .A2(n15093), .ZN(n14320) );
  AOI211_X1 U16252 ( .C1(n15065), .C2(n14490), .A(n14321), .B(n14320), .ZN(
        n14322) );
  INV_X1 U16253 ( .A(n14322), .ZN(P1_U3271) );
  XNOR2_X1 U16254 ( .A(n14324), .B(n14323), .ZN(n14325) );
  AOI222_X1 U16255 ( .A1(n14326), .A2(n15059), .B1(n14173), .B2(n15049), .C1(
        n15196), .C2(n14325), .ZN(n14498) );
  AOI211_X1 U16256 ( .C1(n14496), .C2(n14344), .A(n15147), .B(n7602), .ZN(
        n14495) );
  AOI22_X1 U16257 ( .A1(n15105), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14328), 
        .B2(n15091), .ZN(n14329) );
  OAI21_X1 U16258 ( .B1(n14330), .B2(n15096), .A(n14329), .ZN(n14336) );
  INV_X1 U16259 ( .A(n14331), .ZN(n14332) );
  AOI21_X1 U16260 ( .B1(n14334), .B2(n14333), .A(n14332), .ZN(n14499) );
  NOR2_X1 U16261 ( .A1(n14499), .A2(n14418), .ZN(n14335) );
  AOI211_X1 U16262 ( .C1(n14495), .C2(n15063), .A(n14336), .B(n14335), .ZN(
        n14337) );
  OAI21_X1 U16263 ( .B1(n14498), .B2(n15093), .A(n14337), .ZN(P1_U3272) );
  OAI21_X1 U16264 ( .B1(n6735), .B2(n14339), .A(n14338), .ZN(n14506) );
  OAI21_X1 U16265 ( .B1(n14342), .B2(n14341), .A(n14340), .ZN(n14343) );
  INV_X1 U16266 ( .A(n14343), .ZN(n14504) );
  OAI211_X1 U16267 ( .C1(n14502), .C2(n6728), .A(n15076), .B(n14344), .ZN(
        n14501) );
  AND2_X1 U16268 ( .A1(n14345), .A2(n15049), .ZN(n14346) );
  AOI21_X1 U16269 ( .B1(n14347), .B2(n15059), .A(n14346), .ZN(n14500) );
  NAND2_X1 U16270 ( .A1(n15105), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n14350) );
  NAND2_X1 U16271 ( .A1(n15091), .A2(n14348), .ZN(n14349) );
  OAI211_X1 U16272 ( .C1(n15105), .C2(n14500), .A(n14350), .B(n14349), .ZN(
        n14351) );
  AOI21_X1 U16273 ( .B1(n7272), .B2(n15085), .A(n14351), .ZN(n14352) );
  OAI21_X1 U16274 ( .B1(n14501), .B2(n15087), .A(n14352), .ZN(n14353) );
  AOI21_X1 U16275 ( .B1(n14504), .B2(n15064), .A(n14353), .ZN(n14354) );
  OAI21_X1 U16276 ( .B1(n14418), .B2(n14506), .A(n14354), .ZN(P1_U3273) );
  XNOR2_X1 U16277 ( .A(n14355), .B(n14356), .ZN(n14513) );
  XNOR2_X1 U16278 ( .A(n14357), .B(n14356), .ZN(n14511) );
  AOI211_X1 U16279 ( .C1(n14358), .C2(n14373), .A(n15147), .B(n6728), .ZN(
        n14510) );
  NAND2_X1 U16280 ( .A1(n14510), .A2(n15063), .ZN(n14363) );
  NAND2_X1 U16281 ( .A1(n15091), .A2(n14359), .ZN(n14360) );
  AOI21_X1 U16282 ( .B1(n14507), .B2(n14360), .A(n15093), .ZN(n14361) );
  AOI21_X1 U16283 ( .B1(n15105), .B2(P1_REG2_REG_19__SCAN_IN), .A(n14361), 
        .ZN(n14362) );
  OAI211_X1 U16284 ( .C1(n14508), .C2(n15096), .A(n14363), .B(n14362), .ZN(
        n14364) );
  AOI21_X1 U16285 ( .B1(n14511), .B2(n15064), .A(n14364), .ZN(n14365) );
  OAI21_X1 U16286 ( .B1(n14418), .B2(n14513), .A(n14365), .ZN(P1_U3274) );
  XNOR2_X1 U16287 ( .A(n14366), .B(n14368), .ZN(n14370) );
  INV_X1 U16288 ( .A(n14370), .ZN(n14519) );
  XOR2_X1 U16289 ( .A(n14368), .B(n14367), .Z(n14369) );
  AOI222_X1 U16290 ( .A1(n14370), .A2(n15074), .B1(n14408), .B2(n15049), .C1(
        n15196), .C2(n14369), .ZN(n14518) );
  INV_X1 U16291 ( .A(n14518), .ZN(n14372) );
  INV_X1 U16292 ( .A(n14371), .ZN(n14514) );
  OAI21_X1 U16293 ( .B1(n14372), .B2(n14514), .A(n14379), .ZN(n14383) );
  INV_X1 U16294 ( .A(n14373), .ZN(n14374) );
  AOI211_X1 U16295 ( .C1(n14375), .C2(n14394), .A(n15147), .B(n14374), .ZN(
        n14516) );
  NOR2_X1 U16296 ( .A1(n14376), .A2(n15096), .ZN(n14381) );
  INV_X1 U16297 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14378) );
  OAI22_X1 U16298 ( .A1(n14379), .A2(n14378), .B1(n14377), .B2(n15080), .ZN(
        n14380) );
  AOI211_X1 U16299 ( .C1(n14516), .C2(n15063), .A(n14381), .B(n14380), .ZN(
        n14382) );
  OAI211_X1 U16300 ( .C1(n14519), .C2(n14384), .A(n14383), .B(n14382), .ZN(
        P1_U3275) );
  XNOR2_X1 U16301 ( .A(n14385), .B(n14387), .ZN(n14524) );
  OAI211_X1 U16302 ( .C1(n14388), .C2(n14387), .A(n14386), .B(n15196), .ZN(
        n14392) );
  AOI22_X1 U16303 ( .A1(n14390), .A2(n15059), .B1(n15049), .B2(n14389), .ZN(
        n14391) );
  NAND2_X1 U16304 ( .A1(n14392), .A2(n14391), .ZN(n14520) );
  NAND2_X1 U16305 ( .A1(n14520), .A2(n14379), .ZN(n14402) );
  INV_X1 U16306 ( .A(n14393), .ZN(n14396) );
  INV_X1 U16307 ( .A(n14394), .ZN(n14395) );
  AOI211_X1 U16308 ( .C1(n14522), .C2(n14396), .A(n15147), .B(n14395), .ZN(
        n14521) );
  NOR2_X1 U16309 ( .A1(n14397), .A2(n15096), .ZN(n14400) );
  OAI22_X1 U16310 ( .A1(n14379), .A2(n12245), .B1(n14398), .B2(n15080), .ZN(
        n14399) );
  AOI211_X1 U16311 ( .C1(n14521), .C2(n15063), .A(n14400), .B(n14399), .ZN(
        n14401) );
  OAI211_X1 U16312 ( .C1(n14524), .C2(n14418), .A(n14402), .B(n14401), .ZN(
        P1_U3276) );
  XNOR2_X1 U16313 ( .A(n14403), .B(n14404), .ZN(n14531) );
  XNOR2_X1 U16314 ( .A(n14405), .B(n14404), .ZN(n14529) );
  XNOR2_X1 U16315 ( .A(n14406), .B(n14527), .ZN(n14407) );
  NAND2_X1 U16316 ( .A1(n14407), .A2(n15076), .ZN(n14526) );
  NOR2_X1 U16317 ( .A1(n14379), .A2(n11170), .ZN(n14413) );
  AOI22_X1 U16318 ( .A1(n14409), .A2(n15049), .B1(n14408), .B2(n15059), .ZN(
        n14525) );
  NAND2_X1 U16319 ( .A1(n15091), .A2(n14410), .ZN(n14411) );
  AOI21_X1 U16320 ( .B1(n14525), .B2(n14411), .A(n15093), .ZN(n14412) );
  AOI211_X1 U16321 ( .C1(n14414), .C2(n15085), .A(n14413), .B(n14412), .ZN(
        n14415) );
  OAI21_X1 U16322 ( .B1(n14526), .B2(n15087), .A(n14415), .ZN(n14416) );
  AOI21_X1 U16323 ( .B1(n14529), .B2(n15064), .A(n14416), .ZN(n14417) );
  OAI21_X1 U16324 ( .B1(n14418), .B2(n14531), .A(n14417), .ZN(P1_U3277) );
  OAI21_X1 U16325 ( .B1(n14427), .B2(n14420), .A(n14419), .ZN(n15152) );
  AOI22_X1 U16326 ( .A1(n15065), .A2(n15152), .B1(n15085), .B2(n14421), .ZN(
        n14438) );
  INV_X1 U16327 ( .A(n14422), .ZN(n15099) );
  NOR2_X1 U16328 ( .A1(n14423), .A2(n15140), .ZN(n14424) );
  NOR2_X1 U16329 ( .A1(n14425), .A2(n14424), .ZN(n15145) );
  AOI22_X1 U16330 ( .A1(n15099), .A2(n15145), .B1(n15091), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n14437) );
  OAI21_X1 U16331 ( .B1(n14427), .B2(n14426), .A(n15196), .ZN(n14431) );
  XNOR2_X1 U16332 ( .A(n15145), .B(n14428), .ZN(n14429) );
  AOI21_X1 U16333 ( .B1(n14429), .B2(n15196), .A(n10212), .ZN(n14430) );
  AOI21_X1 U16334 ( .B1(n14432), .B2(n14431), .A(n14430), .ZN(n14433) );
  AOI21_X1 U16335 ( .B1(n15059), .B2(n14434), .A(n14433), .ZN(n15149) );
  MUX2_X1 U16336 ( .A(n15149), .B(n14435), .S(n15105), .Z(n14436) );
  NAND3_X1 U16337 ( .A1(n14438), .A2(n14437), .A3(n14436), .ZN(P1_U3292) );
  OAI211_X1 U16338 ( .C1(n14440), .C2(n15191), .A(n14439), .B(n14441), .ZN(
        n14537) );
  MUX2_X1 U16339 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14537), .S(n15224), .Z(
        P1_U3559) );
  OAI211_X1 U16340 ( .C1(n14443), .C2(n15191), .A(n14442), .B(n14441), .ZN(
        n14538) );
  MUX2_X1 U16341 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14538), .S(n15224), .Z(
        P1_U3558) );
  OAI211_X1 U16342 ( .C1(n14447), .C2(n15191), .A(n14446), .B(n14445), .ZN(
        n14448) );
  NAND2_X1 U16343 ( .A1(n14452), .A2(n15200), .ZN(n14456) );
  NAND3_X1 U16344 ( .A1(n6612), .A2(n15207), .A3(n14453), .ZN(n14455) );
  MUX2_X1 U16345 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14540), .S(n15224), .Z(
        P1_U3556) );
  INV_X1 U16346 ( .A(n14458), .ZN(n14463) );
  AOI21_X1 U16347 ( .B1(n14460), .B2(n15200), .A(n14459), .ZN(n14461) );
  MUX2_X1 U16348 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14541), .S(n15224), .Z(
        P1_U3555) );
  OAI21_X1 U16349 ( .B1(n14465), .B2(n15191), .A(n14464), .ZN(n14466) );
  AOI21_X1 U16350 ( .B1(n14467), .B2(n15207), .A(n14466), .ZN(n14468) );
  NAND2_X1 U16351 ( .A1(n14469), .A2(n14468), .ZN(n14542) );
  MUX2_X1 U16352 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14542), .S(n15224), .Z(
        P1_U3554) );
  AOI211_X1 U16353 ( .C1(n14472), .C2(n15200), .A(n14471), .B(n14470), .ZN(
        n14475) );
  NAND2_X1 U16354 ( .A1(n14473), .A2(n15207), .ZN(n14474) );
  OAI211_X1 U16355 ( .C1(n14476), .C2(n15178), .A(n14475), .B(n14474), .ZN(
        n14543) );
  MUX2_X1 U16356 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14543), .S(n15224), .Z(
        P1_U3553) );
  INV_X1 U16357 ( .A(n14477), .ZN(n14482) );
  NOR2_X1 U16358 ( .A1(n14479), .A2(n14478), .ZN(n14480) );
  OAI211_X1 U16359 ( .C1(n14482), .C2(n14795), .A(n14481), .B(n14480), .ZN(
        n14544) );
  MUX2_X1 U16360 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14544), .S(n15224), .Z(
        P1_U3552) );
  INV_X1 U16361 ( .A(n14483), .ZN(n14488) );
  NAND3_X1 U16362 ( .A1(n14485), .A2(n14484), .A3(n15207), .ZN(n14487) );
  NAND4_X1 U16363 ( .A1(n14489), .A2(n14488), .A3(n14487), .A4(n14486), .ZN(
        n14545) );
  MUX2_X1 U16364 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14545), .S(n15224), .Z(
        P1_U3551) );
  NAND2_X1 U16365 ( .A1(n14490), .A2(n15207), .ZN(n14493) );
  NAND4_X1 U16366 ( .A1(n14494), .A2(n14493), .A3(n14492), .A4(n14491), .ZN(
        n14546) );
  MUX2_X1 U16367 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14546), .S(n15224), .Z(
        P1_U3550) );
  AOI21_X1 U16368 ( .B1(n14496), .B2(n15200), .A(n14495), .ZN(n14497) );
  OAI211_X1 U16369 ( .C1(n14450), .C2(n14499), .A(n14498), .B(n14497), .ZN(
        n14547) );
  MUX2_X1 U16370 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14547), .S(n15224), .Z(
        P1_U3549) );
  OAI211_X1 U16371 ( .C1(n14502), .C2(n15191), .A(n14501), .B(n14500), .ZN(
        n14503) );
  AOI21_X1 U16372 ( .B1(n14504), .B2(n15196), .A(n14503), .ZN(n14505) );
  OAI21_X1 U16373 ( .B1(n14450), .B2(n14506), .A(n14505), .ZN(n14548) );
  MUX2_X1 U16374 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14548), .S(n15224), .Z(
        P1_U3548) );
  OAI21_X1 U16375 ( .B1(n14508), .B2(n15191), .A(n14507), .ZN(n14509) );
  AOI211_X1 U16376 ( .C1(n14511), .C2(n15196), .A(n14510), .B(n14509), .ZN(
        n14512) );
  OAI21_X1 U16377 ( .B1(n14450), .B2(n14513), .A(n14512), .ZN(n14549) );
  MUX2_X1 U16378 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14549), .S(n15224), .Z(
        P1_U3547) );
  NOR3_X1 U16379 ( .A1(n14516), .A2(n14515), .A3(n14514), .ZN(n14517) );
  OAI211_X1 U16380 ( .C1(n14519), .C2(n14795), .A(n14518), .B(n14517), .ZN(
        n14550) );
  MUX2_X1 U16381 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14550), .S(n15224), .Z(
        P1_U3546) );
  AOI211_X1 U16382 ( .C1(n14522), .C2(n15200), .A(n14521), .B(n14520), .ZN(
        n14523) );
  OAI21_X1 U16383 ( .B1(n14450), .B2(n14524), .A(n14523), .ZN(n14551) );
  MUX2_X1 U16384 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14551), .S(n15224), .Z(
        P1_U3545) );
  OAI211_X1 U16385 ( .C1(n14527), .C2(n15191), .A(n14526), .B(n14525), .ZN(
        n14528) );
  AOI21_X1 U16386 ( .B1(n14529), .B2(n15196), .A(n14528), .ZN(n14530) );
  OAI21_X1 U16387 ( .B1(n14450), .B2(n14531), .A(n14530), .ZN(n14552) );
  MUX2_X1 U16388 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14552), .S(n15224), .Z(
        P1_U3544) );
  AOI211_X1 U16389 ( .C1(n14534), .C2(n15200), .A(n14533), .B(n14532), .ZN(
        n14535) );
  OAI21_X1 U16390 ( .B1(n14450), .B2(n14536), .A(n14535), .ZN(n14553) );
  MUX2_X1 U16391 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14553), .S(n15224), .Z(
        P1_U3543) );
  MUX2_X1 U16392 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14537), .S(n15209), .Z(
        P1_U3527) );
  MUX2_X1 U16393 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14538), .S(n15209), .Z(
        P1_U3526) );
  MUX2_X1 U16394 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14540), .S(n15209), .Z(
        P1_U3524) );
  MUX2_X1 U16395 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14542), .S(n15209), .Z(
        P1_U3522) );
  MUX2_X1 U16396 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14543), .S(n15209), .Z(
        P1_U3521) );
  MUX2_X1 U16397 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14544), .S(n15209), .Z(
        P1_U3520) );
  MUX2_X1 U16398 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14545), .S(n15209), .Z(
        P1_U3519) );
  MUX2_X1 U16399 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14546), .S(n15209), .Z(
        P1_U3518) );
  MUX2_X1 U16400 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14547), .S(n15209), .Z(
        P1_U3517) );
  MUX2_X1 U16401 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14548), .S(n15209), .Z(
        P1_U3516) );
  MUX2_X1 U16402 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14549), .S(n15209), .Z(
        P1_U3515) );
  MUX2_X1 U16403 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14550), .S(n15209), .Z(
        P1_U3513) );
  MUX2_X1 U16404 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14551), .S(n15209), .Z(
        P1_U3510) );
  MUX2_X1 U16405 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14552), .S(n15209), .Z(
        P1_U3507) );
  MUX2_X1 U16406 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14553), .S(n15209), .Z(
        P1_U3504) );
  NAND3_X1 U16407 ( .A1(n14554), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n14556) );
  OAI22_X1 U16408 ( .A1(n14557), .A2(n14556), .B1(n14555), .B2(n14571), .ZN(
        n14558) );
  AOI21_X1 U16409 ( .B1(n14560), .B2(n14559), .A(n14558), .ZN(n14561) );
  INV_X1 U16410 ( .A(n14561), .ZN(P1_U3324) );
  OAI222_X1 U16411 ( .A1(P1_U3086), .A2(n6573), .B1(n11699), .B2(n14563), .C1(
        n14562), .C2(n14571), .ZN(P1_U3328) );
  OAI222_X1 U16412 ( .A1(n14567), .A2(P1_U3086), .B1(n11699), .B2(n14566), 
        .C1(n14565), .C2(n14571), .ZN(P1_U3329) );
  OAI222_X1 U16413 ( .A1(P1_U3086), .A2(n14570), .B1(n11699), .B2(n14569), 
        .C1(n14568), .C2(n14571), .ZN(P1_U3330) );
  OAI222_X1 U16414 ( .A1(P1_U3086), .A2(n14574), .B1(n11699), .B2(n14573), 
        .C1(n14572), .C2(n14571), .ZN(P1_U3331) );
  MUX2_X1 U16415 ( .A(n14575), .B(n13861), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16416 ( .A(n14576), .ZN(n14577) );
  MUX2_X1 U16417 ( .A(n14577), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16418 ( .A(n14660), .ZN(n14877) );
  NAND2_X1 U16419 ( .A1(n15554), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n14620) );
  INV_X1 U16420 ( .A(n15537), .ZN(n14650) );
  NOR2_X1 U16421 ( .A1(n14642), .A2(n6715), .ZN(n14579) );
  INV_X1 U16422 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n14580) );
  AOI22_X1 U16423 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n14644), .B1(n15485), 
        .B2(n14580), .ZN(n15478) );
  NOR2_X1 U16424 ( .A1(n14646), .A2(n14581), .ZN(n14582) );
  INV_X1 U16425 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n14583) );
  AOI22_X1 U16426 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n14648), .B1(n15519), 
        .B2(n14583), .ZN(n15512) );
  NOR2_X1 U16427 ( .A1(n14650), .A2(n14584), .ZN(n14585) );
  INV_X1 U16428 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15531) );
  OR2_X1 U16429 ( .A1(n15554), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n14586) );
  NAND2_X1 U16430 ( .A1(n14620), .A2(n14586), .ZN(n15549) );
  AND2_X1 U16431 ( .A1(n14827), .A2(n14587), .ZN(n14588) );
  INV_X1 U16432 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14822) );
  INV_X1 U16433 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n14589) );
  NAND2_X1 U16434 ( .A1(n14845), .A2(n14589), .ZN(n14591) );
  NAND2_X1 U16435 ( .A1(n14655), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n14590) );
  AND2_X1 U16436 ( .A1(n14591), .A2(n14590), .ZN(n14839) );
  NAND2_X1 U16437 ( .A1(n14845), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n14592) );
  INV_X1 U16438 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14859) );
  INV_X1 U16439 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n14595) );
  AOI22_X1 U16440 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14660), .B1(n14877), 
        .B2(n14595), .ZN(n14876) );
  INV_X1 U16441 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n14596) );
  MUX2_X1 U16442 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n14596), .S(n14638), .Z(
        n14634) );
  XNOR2_X1 U16443 ( .A(n14597), .B(n14634), .ZN(n14666) );
  INV_X1 U16444 ( .A(n14598), .ZN(n14599) );
  AOI21_X1 U16445 ( .B1(n15535), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n14599), 
        .ZN(n14637) );
  MUX2_X1 U16446 ( .A(n14595), .B(n14659), .S(n14633), .Z(n14884) );
  INV_X1 U16447 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n14600) );
  MUX2_X1 U16448 ( .A(n14859), .B(n14600), .S(n14633), .Z(n14627) );
  NOR2_X1 U16449 ( .A1(n14627), .A2(n14628), .ZN(n14629) );
  INV_X1 U16450 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15606) );
  MUX2_X1 U16451 ( .A(n11359), .B(n15606), .S(n14633), .Z(n14605) );
  OR2_X1 U16452 ( .A1(n14605), .A2(n14642), .ZN(n15463) );
  OR2_X1 U16453 ( .A1(n14602), .A2(n14601), .ZN(n14604) );
  NAND2_X1 U16454 ( .A1(n14604), .A2(n14603), .ZN(n15466) );
  NAND2_X1 U16455 ( .A1(n15463), .A2(n15466), .ZN(n14606) );
  NAND2_X1 U16456 ( .A1(n14605), .A2(n14642), .ZN(n15464) );
  NAND2_X1 U16457 ( .A1(n14606), .A2(n15464), .ZN(n15490) );
  MUX2_X1 U16458 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n14633), .Z(n14607) );
  XNOR2_X1 U16459 ( .A(n14607), .B(n14644), .ZN(n15489) );
  NAND2_X1 U16460 ( .A1(n15490), .A2(n15489), .ZN(n15488) );
  INV_X1 U16461 ( .A(n14607), .ZN(n14608) );
  NAND2_X1 U16462 ( .A1(n14608), .A2(n14644), .ZN(n14609) );
  NAND2_X1 U16463 ( .A1(n15488), .A2(n14609), .ZN(n15506) );
  MUX2_X1 U16464 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n14633), .Z(n14610) );
  XNOR2_X1 U16465 ( .A(n14610), .B(n14646), .ZN(n15505) );
  NAND2_X1 U16466 ( .A1(n15506), .A2(n15505), .ZN(n15504) );
  INV_X1 U16467 ( .A(n14610), .ZN(n14611) );
  NAND2_X1 U16468 ( .A1(n14611), .A2(n14646), .ZN(n14612) );
  MUX2_X1 U16469 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n14633), .Z(n14613) );
  XNOR2_X1 U16470 ( .A(n14613), .B(n15519), .ZN(n15522) );
  NAND2_X1 U16471 ( .A1(n14613), .A2(n15519), .ZN(n14614) );
  MUX2_X1 U16472 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n14633), .Z(n14615) );
  XNOR2_X1 U16473 ( .A(n14615), .B(n14650), .ZN(n15541) );
  INV_X1 U16474 ( .A(n14615), .ZN(n14616) );
  NAND2_X1 U16475 ( .A1(n14616), .A2(n14650), .ZN(n14617) );
  NAND2_X1 U16476 ( .A1(n15540), .A2(n14617), .ZN(n15566) );
  OR2_X1 U16477 ( .A1(n15554), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n14618) );
  NAND2_X1 U16478 ( .A1(n15554), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n14652) );
  AND2_X1 U16479 ( .A1(n14618), .A2(n14652), .ZN(n15553) );
  INV_X1 U16480 ( .A(n15553), .ZN(n14619) );
  MUX2_X1 U16481 ( .A(n15549), .B(n14619), .S(n14633), .Z(n15565) );
  MUX2_X1 U16482 ( .A(n14620), .B(n14652), .S(n14633), .Z(n14621) );
  NAND2_X1 U16483 ( .A1(n15567), .A2(n14621), .ZN(n14622) );
  INV_X1 U16484 ( .A(n14622), .ZN(n14624) );
  MUX2_X1 U16485 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n14633), .Z(n14832) );
  MUX2_X1 U16486 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n14633), .Z(n14625) );
  NAND2_X1 U16487 ( .A1(n14625), .A2(n14845), .ZN(n14848) );
  NOR2_X1 U16488 ( .A1(n14625), .A2(n14845), .ZN(n14850) );
  AOI21_X1 U16489 ( .B1(n14626), .B2(n14848), .A(n14850), .ZN(n14864) );
  AOI21_X1 U16490 ( .B1(n14628), .B2(n14627), .A(n14629), .ZN(n14863) );
  NAND2_X1 U16491 ( .A1(n14884), .A2(n14885), .ZN(n14883) );
  NAND2_X1 U16492 ( .A1(n14660), .A2(n14630), .ZN(n14631) );
  NAND2_X1 U16493 ( .A1(n14883), .A2(n14631), .ZN(n14636) );
  XNOR2_X1 U16494 ( .A(n14638), .B(n14632), .ZN(n14661) );
  MUX2_X1 U16495 ( .A(n14634), .B(n14661), .S(n14633), .Z(n14635) );
  AOI22_X1 U16496 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n14877), .B1(n14660), 
        .B2(n14659), .ZN(n14882) );
  INV_X1 U16497 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14912) );
  AOI22_X1 U16498 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n15519), .B1(n14648), 
        .B2(n14912), .ZN(n15516) );
  AOI22_X1 U16499 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n15485), .B1(n14644), 
        .B2(n15609), .ZN(n15482) );
  OAI21_X1 U16500 ( .B1(n14640), .B2(n15604), .A(n14639), .ZN(n14641) );
  NAND2_X1 U16501 ( .A1(n15467), .A2(n14641), .ZN(n14643) );
  XNOR2_X1 U16502 ( .A(n14642), .B(n14641), .ZN(n15472) );
  NAND2_X1 U16503 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15472), .ZN(n15471) );
  NAND2_X1 U16504 ( .A1(n15501), .A2(n14645), .ZN(n14647) );
  NAND2_X1 U16505 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n15498), .ZN(n15497) );
  NAND2_X1 U16506 ( .A1(n14647), .A2(n15497), .ZN(n15515) );
  NAND2_X1 U16507 ( .A1(n15537), .A2(n14649), .ZN(n14651) );
  NAND2_X1 U16508 ( .A1(n14651), .A2(n15532), .ZN(n15552) );
  NAND2_X1 U16509 ( .A1(n15553), .A2(n15552), .ZN(n15551) );
  NAND2_X1 U16510 ( .A1(n14827), .A2(n14653), .ZN(n14654) );
  XNOR2_X1 U16511 ( .A(n14655), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n14841) );
  AOI22_X1 U16512 ( .A1(n14842), .A2(n14841), .B1(P3_REG1_REG_16__SCAN_IN), 
        .B2(n14845), .ZN(n14657) );
  INV_X1 U16513 ( .A(n14657), .ZN(n14656) );
  NAND2_X1 U16514 ( .A1(n14868), .A2(n14656), .ZN(n14658) );
  XNOR2_X1 U16515 ( .A(n14657), .B(n14868), .ZN(n14861) );
  NAND2_X1 U16516 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14861), .ZN(n14860) );
  NAND2_X1 U16517 ( .A1(n14658), .A2(n14860), .ZN(n14881) );
  NAND2_X1 U16518 ( .A1(n14882), .A2(n14881), .ZN(n14880) );
  OAI21_X1 U16519 ( .B1(n14660), .B2(n14659), .A(n14880), .ZN(n14662) );
  XNOR2_X1 U16520 ( .A(n14662), .B(n14661), .ZN(n14663) );
  NAND2_X1 U16521 ( .A1(n14663), .A2(n15562), .ZN(n14664) );
  OAI211_X1 U16522 ( .C1(n14666), .C2(n15571), .A(n14665), .B(n14664), .ZN(
        P3_U3201) );
  INV_X1 U16523 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14699) );
  INV_X1 U16524 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14667) );
  XNOR2_X1 U16525 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(n14667), .ZN(n14701) );
  INV_X1 U16526 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14696) );
  INV_X1 U16527 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n15017) );
  XNOR2_X1 U16528 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n15017), .ZN(n14705) );
  INV_X1 U16529 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14687) );
  XOR2_X1 U16530 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Z(
        n14709) );
  XOR2_X1 U16531 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n14685), .Z(n14739) );
  XOR2_X1 U16532 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n14670), .Z(n14714) );
  NAND2_X1 U16533 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14671), .ZN(n14673) );
  NAND2_X1 U16534 ( .A1(n14713), .A2(n14712), .ZN(n14672) );
  NAND2_X1 U16535 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14674), .ZN(n14675) );
  NAND2_X1 U16536 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14676), .ZN(n14678) );
  NAND2_X1 U16537 ( .A1(n14726), .A2(n14725), .ZN(n14677) );
  NAND2_X1 U16538 ( .A1(n14678), .A2(n14677), .ZN(n14733) );
  INV_X1 U16539 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14680) );
  NAND2_X1 U16540 ( .A1(n14681), .A2(n14680), .ZN(n14683) );
  XOR2_X1 U16541 ( .A(n14681), .B(n14680), .Z(n14735) );
  NAND2_X1 U16542 ( .A1(n14735), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14682) );
  NAND2_X1 U16543 ( .A1(n14683), .A2(n14682), .ZN(n14738) );
  NAND2_X1 U16544 ( .A1(n14739), .A2(n14738), .ZN(n14684) );
  NOR2_X1 U16545 ( .A1(n14709), .A2(n14708), .ZN(n14686) );
  NAND2_X1 U16546 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14706), .ZN(n14689) );
  NOR2_X1 U16547 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14706), .ZN(n14688) );
  XOR2_X1 U16548 ( .A(n14691), .B(P3_ADDR_REG_11__SCAN_IN), .Z(n14745) );
  NAND2_X1 U16549 ( .A1(n14746), .A2(n14745), .ZN(n14690) );
  NOR2_X1 U16550 ( .A1(n14705), .A2(n14704), .ZN(n14692) );
  XNOR2_X1 U16551 ( .A(n14694), .B(P3_ADDR_REG_13__SCAN_IN), .ZN(n14748) );
  NOR2_X1 U16552 ( .A1(n14749), .A2(n14748), .ZN(n14693) );
  AOI21_X1 U16553 ( .B1(P3_ADDR_REG_13__SCAN_IN), .B2(n14694), .A(n14693), 
        .ZN(n14703) );
  XOR2_X1 U16554 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n14696), .Z(n14702) );
  NAND2_X1 U16555 ( .A1(n14703), .A2(n14702), .ZN(n14695) );
  NOR2_X1 U16556 ( .A1(n14701), .A2(n14700), .ZN(n14697) );
  AOI21_X1 U16557 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n14698), .A(n14697), 
        .ZN(n14754) );
  XNOR2_X1 U16558 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n14754), .ZN(n14755) );
  XOR2_X1 U16559 ( .A(n14699), .B(n14755), .Z(n14981) );
  XOR2_X1 U16560 ( .A(n14701), .B(n14700), .Z(n14977) );
  XNOR2_X1 U16561 ( .A(n14703), .B(n14702), .ZN(n14974) );
  XOR2_X1 U16562 ( .A(n14705), .B(n14704), .Z(n14967) );
  XNOR2_X1 U16563 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n14706), .ZN(n14707) );
  XNOR2_X1 U16564 ( .A(n14707), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n14792) );
  XOR2_X1 U16565 ( .A(n14709), .B(n14708), .Z(n14785) );
  XNOR2_X1 U16566 ( .A(n14711), .B(n14710), .ZN(n14723) );
  AND2_X1 U16567 ( .A1(n14723), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n14724) );
  XOR2_X1 U16568 ( .A(n14713), .B(n14712), .Z(n15624) );
  XOR2_X1 U16569 ( .A(n14715), .B(n14714), .Z(n14771) );
  NOR2_X1 U16570 ( .A1(n14720), .A2(n6908), .ZN(n14721) );
  AOI21_X1 U16571 ( .B1(n14718), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n14717), .ZN(
        n14719) );
  INV_X1 U16572 ( .A(n14719), .ZN(n15618) );
  NAND2_X1 U16573 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15618), .ZN(n15628) );
  NOR2_X1 U16574 ( .A1(n15628), .A2(n15627), .ZN(n15626) );
  NAND2_X1 U16575 ( .A1(n14771), .A2(n14770), .ZN(n14769) );
  NAND2_X1 U16576 ( .A1(n15624), .A2(n15623), .ZN(n14722) );
  XNOR2_X1 U16577 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n14723), .ZN(n15613) );
  NAND2_X1 U16578 ( .A1(n14728), .A2(n14727), .ZN(n14729) );
  NAND2_X1 U16579 ( .A1(n14729), .A2(n15615), .ZN(n14730) );
  XNOR2_X1 U16580 ( .A(n14731), .B(P3_ADDR_REG_6__SCAN_IN), .ZN(n14732) );
  XNOR2_X1 U16581 ( .A(n14733), .B(n14732), .ZN(n14774) );
  NOR2_X1 U16582 ( .A1(n14736), .A2(n14734), .ZN(n14737) );
  XNOR2_X1 U16583 ( .A(n14735), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15621) );
  XNOR2_X1 U16584 ( .A(n14739), .B(n14738), .ZN(n14741) );
  NAND2_X1 U16585 ( .A1(n14740), .A2(n14741), .ZN(n14742) );
  NAND2_X1 U16586 ( .A1(n14785), .A2(n14784), .ZN(n14743) );
  NAND2_X1 U16587 ( .A1(n14792), .A2(n14793), .ZN(n14744) );
  NOR2_X1 U16588 ( .A1(n14792), .A2(n14793), .ZN(n14791) );
  XNOR2_X1 U16589 ( .A(n14746), .B(n14745), .ZN(n14962) );
  NAND2_X1 U16590 ( .A1(n14963), .A2(n14962), .ZN(n14747) );
  NOR2_X1 U16591 ( .A1(n14963), .A2(n14962), .ZN(n14961) );
  XOR2_X1 U16592 ( .A(n14749), .B(n14748), .Z(n14750) );
  INV_X1 U16593 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14970) );
  NAND2_X1 U16594 ( .A1(n14751), .A2(n14750), .ZN(n14752) );
  NOR2_X1 U16595 ( .A1(n14977), .A2(n14978), .ZN(n14753) );
  NAND2_X1 U16596 ( .A1(n14977), .A2(n14978), .ZN(n14976) );
  NAND2_X1 U16597 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14754), .ZN(n14757) );
  OR2_X1 U16598 ( .A1(n14755), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n14756) );
  NAND2_X1 U16599 ( .A1(n14757), .A2(n14756), .ZN(n14760) );
  XNOR2_X1 U16600 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14760), .ZN(n14761) );
  XOR2_X1 U16601 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14761), .Z(n14758) );
  INV_X1 U16602 ( .A(n14806), .ZN(n14807) );
  NAND2_X1 U16603 ( .A1(n14809), .A2(n14808), .ZN(n14805) );
  INV_X1 U16604 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14815) );
  XOR2_X1 U16605 ( .A(n14815), .B(P1_ADDR_REG_18__SCAN_IN), .Z(n14764) );
  NOR2_X1 U16606 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14760), .ZN(n14763) );
  INV_X1 U16607 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14867) );
  NOR2_X1 U16608 ( .A1(n14867), .A2(n14761), .ZN(n14762) );
  NOR2_X1 U16609 ( .A1(n14763), .A2(n14762), .ZN(n14814) );
  XNOR2_X1 U16610 ( .A(n14764), .B(n14814), .ZN(n14810) );
  NAND2_X1 U16611 ( .A1(n14811), .A2(n14810), .ZN(n14812) );
  OAI21_X1 U16612 ( .B1(n14811), .B2(n14810), .A(n14812), .ZN(n14765) );
  XNOR2_X1 U16613 ( .A(n14765), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16614 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14766) );
  OAI21_X1 U16615 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14766), 
        .ZN(U28) );
  AOI221_X1 U16616 ( .B1(n14767), .B2(n7910), .C1(P2_RD_REG_SCAN_IN), .C2(
        P1_RD_REG_SCAN_IN), .A(P3_RD_REG_SCAN_IN), .ZN(n14768) );
  INV_X1 U16617 ( .A(n14768), .ZN(U29) );
  OAI21_X1 U16618 ( .B1(n14771), .B2(n14770), .A(n14769), .ZN(n14772) );
  XNOR2_X1 U16619 ( .A(n14772), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16620 ( .B1(n14775), .B2(n14774), .A(n14773), .ZN(SUB_1596_U57) );
  OAI21_X1 U16621 ( .B1(n14778), .B2(n14777), .A(n14776), .ZN(SUB_1596_U55) );
  AOI22_X1 U16622 ( .A1(n14781), .A2(n14780), .B1(SI_18_), .B2(n14779), .ZN(
        n14782) );
  OAI21_X1 U16623 ( .B1(P3_U3151), .B2(n14877), .A(n14782), .ZN(P3_U3277) );
  AOI21_X1 U16624 ( .B1(n14785), .B2(n14784), .A(n14783), .ZN(n14786) );
  XOR2_X1 U16625 ( .A(n14786), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  OAI22_X1 U16626 ( .A1(n14788), .A2(n14787), .B1(SI_22_), .B2(n12784), .ZN(
        n14789) );
  AOI21_X1 U16627 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n14790), .A(n14789), .ZN(
        P3_U3273) );
  AOI21_X1 U16628 ( .B1(n14793), .B2(n14792), .A(n14791), .ZN(n14794) );
  XOR2_X1 U16629 ( .A(n14794), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  INV_X1 U16630 ( .A(n14795), .ZN(n15195) );
  OAI21_X1 U16631 ( .B1(n14797), .B2(n15191), .A(n14796), .ZN(n14798) );
  AOI21_X1 U16632 ( .B1(n14799), .B2(n15195), .A(n14798), .ZN(n14800) );
  AND2_X1 U16633 ( .A1(n14801), .A2(n14800), .ZN(n14804) );
  AOI22_X1 U16634 ( .A1(n15209), .A2(n14804), .B1(n14802), .B2(n15208), .ZN(
        P1_U3495) );
  AOI22_X1 U16635 ( .A1(n15224), .A2(n14804), .B1(n14803), .B2(n15221), .ZN(
        P1_U3540) );
  OAI222_X1 U16636 ( .A1(n14809), .A2(n14808), .B1(n14809), .B2(n14807), .C1(
        n14806), .C2(n14805), .ZN(SUB_1596_U63) );
  INV_X1 U16637 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15048) );
  NOR2_X1 U16638 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n15048), .ZN(n14813) );
  OAI22_X1 U16639 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14815), .B1(n14814), 
        .B2(n14813), .ZN(n14816) );
  INV_X1 U16640 ( .A(n14816), .ZN(n14818) );
  XNOR2_X1 U16641 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14817) );
  AOI21_X1 U16642 ( .B1(n14822), .B2(n14821), .A(n14820), .ZN(n14836) );
  OAI21_X1 U16643 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14824), .A(n14823), 
        .ZN(n14829) );
  AOI21_X1 U16644 ( .B1(n15535), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n14825), 
        .ZN(n14826) );
  OAI21_X1 U16645 ( .B1(n15555), .B2(n14827), .A(n14826), .ZN(n14828) );
  AOI21_X1 U16646 ( .B1(n14829), .B2(n15562), .A(n14828), .ZN(n14835) );
  AOI21_X1 U16647 ( .B1(n14832), .B2(n14831), .A(n14830), .ZN(n14833) );
  OR2_X1 U16648 ( .A1(n14833), .A2(n15564), .ZN(n14834) );
  OAI211_X1 U16649 ( .C1(n14836), .C2(n15571), .A(n14835), .B(n14834), .ZN(
        P3_U3197) );
  INV_X1 U16650 ( .A(n14837), .ZN(n14838) );
  AOI21_X1 U16651 ( .B1(n14840), .B2(n14839), .A(n14838), .ZN(n14856) );
  XNOR2_X1 U16652 ( .A(n14842), .B(n14841), .ZN(n14847) );
  AOI21_X1 U16653 ( .B1(n15535), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n14843), 
        .ZN(n14844) );
  OAI21_X1 U16654 ( .B1(n15555), .B2(n14845), .A(n14844), .ZN(n14846) );
  AOI21_X1 U16655 ( .B1(n14847), .B2(n15562), .A(n14846), .ZN(n14855) );
  INV_X1 U16656 ( .A(n14848), .ZN(n14849) );
  NOR2_X1 U16657 ( .A1(n14850), .A2(n14849), .ZN(n14852) );
  AOI21_X1 U16658 ( .B1(n14853), .B2(n14852), .A(n15564), .ZN(n14851) );
  OAI21_X1 U16659 ( .B1(n14853), .B2(n14852), .A(n14851), .ZN(n14854) );
  OAI211_X1 U16660 ( .C1(n14856), .C2(n15571), .A(n14855), .B(n14854), .ZN(
        P3_U3198) );
  AOI21_X1 U16661 ( .B1(n14859), .B2(n14858), .A(n14857), .ZN(n14874) );
  OAI21_X1 U16662 ( .B1(n14861), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14860), 
        .ZN(n14862) );
  AND2_X1 U16663 ( .A1(n14862), .A2(n15562), .ZN(n14871) );
  OAI21_X1 U16664 ( .B1(n14864), .B2(n14863), .A(n15543), .ZN(n14866) );
  NOR2_X1 U16665 ( .A1(n14866), .A2(n14865), .ZN(n14870) );
  INV_X1 U16666 ( .A(n15535), .ZN(n15559) );
  OAI22_X1 U16667 ( .A1(n15555), .A2(n14868), .B1(n15559), .B2(n14867), .ZN(
        n14869) );
  NOR4_X1 U16668 ( .A1(n14872), .A2(n14871), .A3(n14870), .A4(n14869), .ZN(
        n14873) );
  OAI21_X1 U16669 ( .B1(n14874), .B2(n15571), .A(n14873), .ZN(P3_U3199) );
  AOI21_X1 U16670 ( .B1(n6718), .B2(n14876), .A(n14875), .ZN(n14890) );
  NOR2_X1 U16671 ( .A1(n15555), .A2(n14877), .ZN(n14878) );
  AOI211_X1 U16672 ( .C1(n15535), .C2(P3_ADDR_REG_18__SCAN_IN), .A(n14879), 
        .B(n14878), .ZN(n14889) );
  OAI21_X1 U16673 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n14887) );
  OAI21_X1 U16674 ( .B1(n14885), .B2(n14884), .A(n14883), .ZN(n14886) );
  AOI22_X1 U16675 ( .A1(n14887), .A2(n15562), .B1(n15543), .B2(n14886), .ZN(
        n14888) );
  OAI211_X1 U16676 ( .C1(n14890), .C2(n15571), .A(n14889), .B(n14888), .ZN(
        P3_U3200) );
  INV_X1 U16677 ( .A(n14891), .ZN(n14892) );
  AOI21_X1 U16678 ( .B1(n14899), .B2(n14893), .A(n14892), .ZN(n14894) );
  OAI21_X1 U16679 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(P3_U3203) );
  AOI21_X1 U16680 ( .B1(n14899), .B2(n14898), .A(n14897), .ZN(n14918) );
  INV_X1 U16681 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14900) );
  AOI22_X1 U16682 ( .A1(n15611), .A2(n14918), .B1(n14900), .B2(n15608), .ZN(
        P3_U3489) );
  INV_X1 U16683 ( .A(n14901), .ZN(n14904) );
  INV_X1 U16684 ( .A(n14902), .ZN(n14903) );
  AOI211_X1 U16685 ( .C1(n14905), .C2(n15595), .A(n14904), .B(n14903), .ZN(
        n14920) );
  INV_X1 U16686 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14906) );
  AOI22_X1 U16687 ( .A1(n15611), .A2(n14920), .B1(n14906), .B2(n15608), .ZN(
        P3_U3472) );
  OAI211_X1 U16688 ( .C1(n14910), .C2(n14909), .A(n14908), .B(n14907), .ZN(
        n14911) );
  INV_X1 U16689 ( .A(n14911), .ZN(n14922) );
  AOI22_X1 U16690 ( .A1(n15611), .A2(n14922), .B1(n14912), .B2(n15608), .ZN(
        P3_U3471) );
  AOI21_X1 U16691 ( .B1(n14914), .B2(n15595), .A(n14913), .ZN(n14915) );
  AND2_X1 U16692 ( .A1(n14916), .A2(n14915), .ZN(n14924) );
  INV_X1 U16693 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14917) );
  AOI22_X1 U16694 ( .A1(n15611), .A2(n14924), .B1(n14917), .B2(n15608), .ZN(
        P3_U3470) );
  INV_X1 U16695 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14919) );
  AOI22_X1 U16696 ( .A1(n15601), .A2(n14919), .B1(n14918), .B2(n15599), .ZN(
        P3_U3457) );
  INV_X1 U16697 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14921) );
  AOI22_X1 U16698 ( .A1(n15601), .A2(n14921), .B1(n14920), .B2(n15599), .ZN(
        P3_U3429) );
  INV_X1 U16699 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14923) );
  AOI22_X1 U16700 ( .A1(n15601), .A2(n14923), .B1(n14922), .B2(n15599), .ZN(
        P3_U3426) );
  INV_X1 U16701 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14925) );
  AOI22_X1 U16702 ( .A1(n15601), .A2(n14925), .B1(n14924), .B2(n15599), .ZN(
        P3_U3423) );
  OAI21_X1 U16703 ( .B1(n14927), .B2(n15376), .A(n14926), .ZN(n14929) );
  AOI211_X1 U16704 ( .C1(n14930), .C2(n15373), .A(n14929), .B(n14928), .ZN(
        n14932) );
  AOI22_X1 U16705 ( .A1(n15392), .A2(n14932), .B1(n10809), .B2(n15390), .ZN(
        P2_U3511) );
  INV_X1 U16706 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14931) );
  AOI22_X1 U16707 ( .A1(n15383), .A2(n14932), .B1(n14931), .B2(n15381), .ZN(
        P2_U3466) );
  NAND3_X1 U16708 ( .A1(n14934), .A2(n14933), .A3(n15207), .ZN(n14939) );
  INV_X1 U16709 ( .A(n14935), .ZN(n14937) );
  NAND4_X1 U16710 ( .A1(n14939), .A2(n14938), .A3(n14937), .A4(n14936), .ZN(
        n14940) );
  AOI21_X1 U16711 ( .B1(n14941), .B2(n15196), .A(n14940), .ZN(n14957) );
  AOI22_X1 U16712 ( .A1(n15224), .A2(n14957), .B1(n14942), .B2(n15221), .ZN(
        P1_U3542) );
  OAI211_X1 U16713 ( .C1(n14945), .C2(n15191), .A(n14944), .B(n14943), .ZN(
        n14947) );
  AOI211_X1 U16714 ( .C1(n14948), .C2(n15207), .A(n14947), .B(n14946), .ZN(
        n14959) );
  AOI22_X1 U16715 ( .A1(n15224), .A2(n14959), .B1(n14949), .B2(n15221), .ZN(
        P1_U3541) );
  OAI211_X1 U16716 ( .C1(n14952), .C2(n15191), .A(n14951), .B(n14950), .ZN(
        n14953) );
  AOI21_X1 U16717 ( .B1(n14954), .B2(n15207), .A(n14953), .ZN(n14960) );
  AOI22_X1 U16718 ( .A1(n15224), .A2(n14960), .B1(n14955), .B2(n15221), .ZN(
        P1_U3539) );
  INV_X1 U16719 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14956) );
  AOI22_X1 U16720 ( .A1(n15209), .A2(n14957), .B1(n14956), .B2(n15208), .ZN(
        P1_U3501) );
  INV_X1 U16721 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14958) );
  AOI22_X1 U16722 ( .A1(n15209), .A2(n14959), .B1(n14958), .B2(n15208), .ZN(
        P1_U3498) );
  AOI22_X1 U16723 ( .A1(n15209), .A2(n14960), .B1(n11154), .B2(n15208), .ZN(
        P1_U3492) );
  AOI21_X1 U16724 ( .B1(n14963), .B2(n14962), .A(n14961), .ZN(n14964) );
  XOR2_X1 U16725 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14964), .Z(SUB_1596_U69)
         );
  AOI21_X1 U16726 ( .B1(n14967), .B2(n14966), .A(n14965), .ZN(n14968) );
  XNOR2_X1 U16727 ( .A(n7455), .B(n14968), .ZN(SUB_1596_U68) );
  OAI21_X1 U16728 ( .B1(n14971), .B2(n14970), .A(n14969), .ZN(SUB_1596_U67) );
  OAI21_X1 U16729 ( .B1(n14974), .B2(n14973), .A(n14972), .ZN(n14975) );
  XNOR2_X1 U16730 ( .A(n14975), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI21_X1 U16731 ( .B1(n14978), .B2(n14977), .A(n14976), .ZN(n14979) );
  XNOR2_X1 U16732 ( .A(n14979), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  AOI21_X1 U16733 ( .B1(n14981), .B2(n14980), .A(n6708), .ZN(n14982) );
  XOR2_X1 U16734 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14982), .Z(SUB_1596_U64)
         );
  MUX2_X1 U16735 ( .A(n10219), .B(P1_REG2_REG_4__SCAN_IN), .S(n14994), .Z(
        n14983) );
  NAND3_X1 U16736 ( .A1(n14985), .A2(n14984), .A3(n14983), .ZN(n14986) );
  NAND3_X1 U16737 ( .A1(n15024), .A2(n14987), .A3(n14986), .ZN(n14999) );
  INV_X1 U16738 ( .A(n14988), .ZN(n14993) );
  NAND3_X1 U16739 ( .A1(n14991), .A2(n14990), .A3(n14989), .ZN(n14992) );
  NAND3_X1 U16740 ( .A1(n15028), .A2(n14993), .A3(n14992), .ZN(n14998) );
  NAND2_X1 U16741 ( .A1(n15012), .A2(n14994), .ZN(n14997) );
  AOI21_X1 U16742 ( .B1(n15018), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14995), .ZN(
        n14996) );
  AND4_X1 U16743 ( .A1(n14999), .A2(n14998), .A3(n14997), .A4(n14996), .ZN(
        n15001) );
  NAND2_X1 U16744 ( .A1(n15001), .A2(n15000), .ZN(P1_U3247) );
  OAI21_X1 U16745 ( .B1(n15004), .B2(n15003), .A(n15002), .ZN(n15014) );
  INV_X1 U16746 ( .A(n15005), .ZN(n15010) );
  NAND3_X1 U16747 ( .A1(n15008), .A2(n15007), .A3(n15006), .ZN(n15009) );
  NAND2_X1 U16748 ( .A1(n15010), .A2(n15009), .ZN(n15011) );
  AOI222_X1 U16749 ( .A1(n15014), .A2(n15024), .B1(n15013), .B2(n15012), .C1(
        n15011), .C2(n15028), .ZN(n15016) );
  OAI211_X1 U16750 ( .C1(n15017), .C2(n15047), .A(n15016), .B(n15015), .ZN(
        P1_U3255) );
  NAND2_X1 U16751 ( .A1(n15018), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n15019) );
  OAI211_X1 U16752 ( .C1(n15043), .C2(n15021), .A(n15020), .B(n15019), .ZN(
        n15022) );
  INV_X1 U16753 ( .A(n15022), .ZN(n15033) );
  OAI211_X1 U16754 ( .C1(n15026), .C2(n15025), .A(n15024), .B(n15023), .ZN(
        n15032) );
  OAI211_X1 U16755 ( .C1(n15030), .C2(n15029), .A(n15028), .B(n15027), .ZN(
        n15031) );
  NAND3_X1 U16756 ( .A1(n15033), .A2(n15032), .A3(n15031), .ZN(P1_U3256) );
  OAI21_X1 U16757 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n15035), .A(n15034), 
        .ZN(n15040) );
  OAI21_X1 U16758 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n15037), .A(n15036), 
        .ZN(n15038) );
  OAI222_X1 U16759 ( .A1(n15043), .A2(n15042), .B1(n15041), .B2(n15040), .C1(
        n15039), .C2(n15038), .ZN(n15044) );
  INV_X1 U16760 ( .A(n15044), .ZN(n15046) );
  OAI211_X1 U16761 ( .C1(n15048), .C2(n15047), .A(n15046), .B(n15045), .ZN(
        P1_U3261) );
  AND2_X1 U16762 ( .A1(n15050), .A2(n15049), .ZN(n15199) );
  MUX2_X1 U16763 ( .A(n15199), .B(P1_REG2_REG_10__SCAN_IN), .S(n15105), .Z(
        n15051) );
  AOI21_X1 U16764 ( .B1(n15085), .B2(n15201), .A(n15051), .ZN(n15067) );
  OAI21_X1 U16765 ( .B1(n15053), .B2(n15054), .A(n15052), .ZN(n15206) );
  NAND2_X1 U16766 ( .A1(n15055), .A2(n15054), .ZN(n15056) );
  AND2_X1 U16767 ( .A1(n15057), .A2(n15056), .ZN(n15197) );
  XNOR2_X1 U16768 ( .A(n7264), .B(n15201), .ZN(n15058) );
  NAND2_X1 U16769 ( .A1(n15058), .A2(n15076), .ZN(n15062) );
  NAND2_X1 U16770 ( .A1(n15060), .A2(n15059), .ZN(n15061) );
  NAND2_X1 U16771 ( .A1(n15062), .A2(n15061), .ZN(n15198) );
  AOI222_X1 U16772 ( .A1(n15206), .A2(n15065), .B1(n15064), .B2(n15197), .C1(
        n15198), .C2(n15063), .ZN(n15066) );
  OAI211_X1 U16773 ( .C1(n15068), .C2(n15080), .A(n15067), .B(n15066), .ZN(
        P1_U3283) );
  OAI21_X1 U16774 ( .B1(n15070), .B2(n6864), .A(n15069), .ZN(n15174) );
  INV_X1 U16775 ( .A(n15170), .ZN(n15073) );
  XNOR2_X1 U16776 ( .A(n15071), .B(n6864), .ZN(n15072) );
  NOR2_X1 U16777 ( .A1(n15072), .A2(n15178), .ZN(n15172) );
  AOI211_X1 U16778 ( .C1(n15074), .C2(n15174), .A(n15073), .B(n15172), .ZN(
        n15090) );
  NAND2_X1 U16779 ( .A1(n15075), .A2(n15084), .ZN(n15077) );
  NAND2_X1 U16780 ( .A1(n15077), .A2(n15076), .ZN(n15078) );
  OR2_X1 U16781 ( .A1(n15079), .A2(n15078), .ZN(n15169) );
  OAI22_X1 U16782 ( .A1(n14379), .A2(n15082), .B1(n15081), .B2(n15080), .ZN(
        n15083) );
  AOI21_X1 U16783 ( .B1(n15085), .B2(n15084), .A(n15083), .ZN(n15086) );
  OAI21_X1 U16784 ( .B1(n15087), .B2(n15169), .A(n15086), .ZN(n15088) );
  AOI21_X1 U16785 ( .B1(n15100), .B2(n15174), .A(n15088), .ZN(n15089) );
  OAI21_X1 U16786 ( .B1(n15105), .B2(n15090), .A(n15089), .ZN(P1_U3287) );
  AOI22_X1 U16787 ( .A1(n15093), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n15092), 
        .B2(n15091), .ZN(n15094) );
  OAI21_X1 U16788 ( .B1(n15096), .B2(n15095), .A(n15094), .ZN(n15097) );
  INV_X1 U16789 ( .A(n15097), .ZN(n15103) );
  AOI22_X1 U16790 ( .A1(n15101), .A2(n15100), .B1(n15099), .B2(n15098), .ZN(
        n15102) );
  OAI211_X1 U16791 ( .C1(n15105), .C2(n15104), .A(n15103), .B(n15102), .ZN(
        P1_U3288) );
  INV_X1 U16792 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15106) );
  NOR2_X1 U16793 ( .A1(n15136), .A2(n15106), .ZN(P1_U3294) );
  INV_X1 U16794 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15107) );
  NOR2_X1 U16795 ( .A1(n15136), .A2(n15107), .ZN(P1_U3295) );
  INV_X1 U16796 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15108) );
  NOR2_X1 U16797 ( .A1(n15136), .A2(n15108), .ZN(P1_U3296) );
  NOR2_X1 U16798 ( .A1(n15136), .A2(n15109), .ZN(P1_U3297) );
  INV_X1 U16799 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15110) );
  NOR2_X1 U16800 ( .A1(n15136), .A2(n15110), .ZN(P1_U3298) );
  INV_X1 U16801 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15111) );
  NOR2_X1 U16802 ( .A1(n15136), .A2(n15111), .ZN(P1_U3299) );
  INV_X1 U16803 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15112) );
  NOR2_X1 U16804 ( .A1(n15136), .A2(n15112), .ZN(P1_U3300) );
  NOR2_X1 U16805 ( .A1(n15136), .A2(n15113), .ZN(P1_U3301) );
  INV_X1 U16806 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15114) );
  NOR2_X1 U16807 ( .A1(n15136), .A2(n15114), .ZN(P1_U3302) );
  INV_X1 U16808 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15115) );
  NOR2_X1 U16809 ( .A1(n15136), .A2(n15115), .ZN(P1_U3303) );
  NOR2_X1 U16810 ( .A1(n15136), .A2(n15116), .ZN(P1_U3304) );
  NOR2_X1 U16811 ( .A1(n15136), .A2(n15117), .ZN(P1_U3305) );
  INV_X1 U16812 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15118) );
  NOR2_X1 U16813 ( .A1(n15136), .A2(n15118), .ZN(P1_U3306) );
  INV_X1 U16814 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15119) );
  NOR2_X1 U16815 ( .A1(n15136), .A2(n15119), .ZN(P1_U3307) );
  INV_X1 U16816 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15120) );
  NOR2_X1 U16817 ( .A1(n15136), .A2(n15120), .ZN(P1_U3308) );
  NOR2_X1 U16818 ( .A1(n15136), .A2(n15121), .ZN(P1_U3309) );
  INV_X1 U16819 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15122) );
  NOR2_X1 U16820 ( .A1(n15136), .A2(n15122), .ZN(P1_U3310) );
  INV_X1 U16821 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15123) );
  NOR2_X1 U16822 ( .A1(n15136), .A2(n15123), .ZN(P1_U3311) );
  INV_X1 U16823 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15124) );
  NOR2_X1 U16824 ( .A1(n15136), .A2(n15124), .ZN(P1_U3312) );
  NOR2_X1 U16825 ( .A1(n15136), .A2(n15125), .ZN(P1_U3313) );
  INV_X1 U16826 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15126) );
  NOR2_X1 U16827 ( .A1(n15136), .A2(n15126), .ZN(P1_U3314) );
  INV_X1 U16828 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15127) );
  NOR2_X1 U16829 ( .A1(n15136), .A2(n15127), .ZN(P1_U3315) );
  INV_X1 U16830 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15128) );
  NOR2_X1 U16831 ( .A1(n15136), .A2(n15128), .ZN(P1_U3316) );
  INV_X1 U16832 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15129) );
  NOR2_X1 U16833 ( .A1(n15136), .A2(n15129), .ZN(P1_U3317) );
  NOR2_X1 U16834 ( .A1(n15136), .A2(n15130), .ZN(P1_U3318) );
  INV_X1 U16835 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15131) );
  NOR2_X1 U16836 ( .A1(n15136), .A2(n15131), .ZN(P1_U3319) );
  INV_X1 U16837 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15132) );
  NOR2_X1 U16838 ( .A1(n15136), .A2(n15132), .ZN(P1_U3320) );
  INV_X1 U16839 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15133) );
  NOR2_X1 U16840 ( .A1(n15136), .A2(n15133), .ZN(P1_U3321) );
  INV_X1 U16841 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15134) );
  NOR2_X1 U16842 ( .A1(n15136), .A2(n15134), .ZN(P1_U3322) );
  INV_X1 U16843 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15135) );
  NOR2_X1 U16844 ( .A1(n15136), .A2(n15135), .ZN(P1_U3323) );
  AOI21_X1 U16845 ( .B1(n15178), .B2(n14450), .A(n15137), .ZN(n15143) );
  INV_X1 U16846 ( .A(n15138), .ZN(n15142) );
  NOR3_X1 U16847 ( .A1(n15140), .A2(n15139), .A3(n13861), .ZN(n15141) );
  NOR3_X1 U16848 ( .A1(n15143), .A2(n15142), .A3(n15141), .ZN(n15210) );
  AOI22_X1 U16849 ( .A1(n15209), .A2(n15210), .B1(n15144), .B2(n15208), .ZN(
        P1_U3459) );
  INV_X1 U16850 ( .A(n15145), .ZN(n15148) );
  OAI21_X1 U16851 ( .B1(n15148), .B2(n15147), .A(n15146), .ZN(n15151) );
  INV_X1 U16852 ( .A(n15149), .ZN(n15150) );
  AOI211_X1 U16853 ( .C1(n15207), .C2(n15152), .A(n15151), .B(n15150), .ZN(
        n15211) );
  AOI22_X1 U16854 ( .A1(n15209), .A2(n15211), .B1(n10014), .B2(n15208), .ZN(
        P1_U3462) );
  INV_X1 U16855 ( .A(n15153), .ZN(n15155) );
  OAI211_X1 U16856 ( .C1(n15156), .C2(n15191), .A(n15155), .B(n15154), .ZN(
        n15159) );
  NOR2_X1 U16857 ( .A1(n15157), .A2(n15178), .ZN(n15158) );
  AOI211_X1 U16858 ( .C1(n15160), .C2(n15207), .A(n15159), .B(n15158), .ZN(
        n15212) );
  AOI22_X1 U16859 ( .A1(n15209), .A2(n15212), .B1(n10038), .B2(n15208), .ZN(
        P1_U3465) );
  INV_X1 U16860 ( .A(n15161), .ZN(n15162) );
  OAI21_X1 U16861 ( .B1(n15163), .B2(n15191), .A(n15162), .ZN(n15165) );
  AOI211_X1 U16862 ( .C1(n15195), .C2(n15166), .A(n15165), .B(n15164), .ZN(
        n15213) );
  INV_X1 U16863 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15167) );
  AOI22_X1 U16864 ( .A1(n15209), .A2(n15213), .B1(n15167), .B2(n15208), .ZN(
        P1_U3468) );
  INV_X1 U16865 ( .A(n15168), .ZN(n15171) );
  NAND3_X1 U16866 ( .A1(n15171), .A2(n15170), .A3(n15169), .ZN(n15173) );
  AOI211_X1 U16867 ( .C1(n15207), .C2(n15174), .A(n15173), .B(n15172), .ZN(
        n15215) );
  AOI22_X1 U16868 ( .A1(n15209), .A2(n15215), .B1(n10416), .B2(n15208), .ZN(
        P1_U3477) );
  OAI211_X1 U16869 ( .C1(n15177), .C2(n15191), .A(n15176), .B(n15175), .ZN(
        n15181) );
  NOR2_X1 U16870 ( .A1(n15179), .A2(n15178), .ZN(n15180) );
  AOI211_X1 U16871 ( .C1(n15207), .C2(n15182), .A(n15181), .B(n15180), .ZN(
        n15217) );
  AOI22_X1 U16872 ( .A1(n15209), .A2(n15217), .B1(n10864), .B2(n15208), .ZN(
        P1_U3480) );
  OR3_X1 U16873 ( .A1(n15185), .A2(n15184), .A3(n15183), .ZN(n15187) );
  AOI211_X1 U16874 ( .C1(n15207), .C2(n15188), .A(n15187), .B(n15186), .ZN(
        n15218) );
  INV_X1 U16875 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15189) );
  AOI22_X1 U16876 ( .A1(n15209), .A2(n15218), .B1(n15189), .B2(n15208), .ZN(
        P1_U3483) );
  OAI21_X1 U16877 ( .B1(n7265), .B2(n15191), .A(n15190), .ZN(n15193) );
  AOI211_X1 U16878 ( .C1(n15195), .C2(n15194), .A(n15193), .B(n15192), .ZN(
        n15220) );
  AOI22_X1 U16879 ( .A1(n15209), .A2(n15220), .B1(n10899), .B2(n15208), .ZN(
        P1_U3486) );
  NAND2_X1 U16880 ( .A1(n15197), .A2(n15196), .ZN(n15204) );
  INV_X1 U16881 ( .A(n15198), .ZN(n15203) );
  AOI21_X1 U16882 ( .B1(n15201), .B2(n15200), .A(n15199), .ZN(n15202) );
  NAND3_X1 U16883 ( .A1(n15204), .A2(n15203), .A3(n15202), .ZN(n15205) );
  AOI21_X1 U16884 ( .B1(n15207), .B2(n15206), .A(n15205), .ZN(n15223) );
  AOI22_X1 U16885 ( .A1(n15209), .A2(n15223), .B1(n11042), .B2(n15208), .ZN(
        P1_U3489) );
  AOI22_X1 U16886 ( .A1(n15224), .A2(n15210), .B1(n9992), .B2(n15221), .ZN(
        P1_U3528) );
  AOI22_X1 U16887 ( .A1(n15224), .A2(n15211), .B1(n10015), .B2(n15221), .ZN(
        P1_U3529) );
  AOI22_X1 U16888 ( .A1(n15224), .A2(n15212), .B1(n9754), .B2(n15221), .ZN(
        P1_U3530) );
  AOI22_X1 U16889 ( .A1(n15224), .A2(n15213), .B1(n10079), .B2(n15221), .ZN(
        P1_U3531) );
  AOI22_X1 U16890 ( .A1(n15224), .A2(n15215), .B1(n15214), .B2(n15221), .ZN(
        P1_U3534) );
  AOI22_X1 U16891 ( .A1(n15224), .A2(n15217), .B1(n15216), .B2(n15221), .ZN(
        P1_U3535) );
  AOI22_X1 U16892 ( .A1(n15224), .A2(n15218), .B1(n10874), .B2(n15221), .ZN(
        P1_U3536) );
  AOI22_X1 U16893 ( .A1(n15224), .A2(n15220), .B1(n15219), .B2(n15221), .ZN(
        P1_U3537) );
  AOI22_X1 U16894 ( .A1(n15224), .A2(n15223), .B1(n15222), .B2(n15221), .ZN(
        P1_U3538) );
  NOR2_X1 U16895 ( .A1(n15299), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16896 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15306), .B1(n15300), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n15228) );
  AOI22_X1 U16897 ( .A1(n15299), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15227) );
  OAI22_X1 U16898 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15265), .B1(n15270), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n15225) );
  OAI21_X1 U16899 ( .B1(n15305), .B2(n15225), .A(n15229), .ZN(n15226) );
  OAI211_X1 U16900 ( .C1(n15229), .C2(n15228), .A(n15227), .B(n15226), .ZN(
        P2_U3214) );
  OAI21_X1 U16901 ( .B1(n15260), .B2(n14734), .A(n15230), .ZN(n15231) );
  AOI21_X1 U16902 ( .B1(n15232), .B2(n15305), .A(n15231), .ZN(n15241) );
  OAI211_X1 U16903 ( .C1(n15235), .C2(n15234), .A(n15233), .B(n15300), .ZN(
        n15240) );
  OAI211_X1 U16904 ( .C1(n15238), .C2(n15237), .A(n15236), .B(n15306), .ZN(
        n15239) );
  NAND3_X1 U16905 ( .A1(n15241), .A2(n15240), .A3(n15239), .ZN(P2_U3221) );
  INV_X1 U16906 ( .A(n15242), .ZN(n15244) );
  NAND3_X1 U16907 ( .A1(n15245), .A2(n15244), .A3(n15243), .ZN(n15246) );
  NAND2_X1 U16908 ( .A1(n15247), .A2(n15246), .ZN(n15248) );
  NAND2_X1 U16909 ( .A1(n15248), .A2(n15306), .ZN(n15255) );
  NAND2_X1 U16910 ( .A1(n15250), .A2(n15249), .ZN(n15251) );
  NAND2_X1 U16911 ( .A1(n15252), .A2(n15251), .ZN(n15253) );
  NAND2_X1 U16912 ( .A1(n15253), .A2(n15300), .ZN(n15254) );
  OAI211_X1 U16913 ( .C1(n15262), .C2(n15256), .A(n15255), .B(n15254), .ZN(
        n15257) );
  INV_X1 U16914 ( .A(n15257), .ZN(n15259) );
  OAI211_X1 U16915 ( .C1(n7455), .C2(n15260), .A(n15259), .B(n15258), .ZN(
        P2_U3226) );
  OAI22_X1 U16916 ( .A1(n15262), .A2(n15261), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11225), .ZN(n15263) );
  AOI21_X1 U16917 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(n15299), .A(n15263), 
        .ZN(n15276) );
  AOI211_X1 U16918 ( .C1(n15267), .C2(n15266), .A(n15265), .B(n15264), .ZN(
        n15268) );
  INV_X1 U16919 ( .A(n15268), .ZN(n15275) );
  AOI211_X1 U16920 ( .C1(n15272), .C2(n15271), .A(n15270), .B(n15269), .ZN(
        n15273) );
  INV_X1 U16921 ( .A(n15273), .ZN(n15274) );
  NAND3_X1 U16922 ( .A1(n15276), .A2(n15275), .A3(n15274), .ZN(P2_U3227) );
  INV_X1 U16923 ( .A(n15277), .ZN(n15279) );
  OAI21_X1 U16924 ( .B1(n15279), .B2(n15278), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15280) );
  OAI21_X1 U16925 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15280), .ZN(n15289) );
  OAI211_X1 U16926 ( .C1(n15282), .C2(P2_REG2_REG_14__SCAN_IN), .A(n15281), 
        .B(n15306), .ZN(n15288) );
  XOR2_X1 U16927 ( .A(n15284), .B(n15283), .Z(n15285) );
  NAND2_X1 U16928 ( .A1(n15285), .A2(n15300), .ZN(n15287) );
  NAND2_X1 U16929 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n15299), .ZN(n15286) );
  NAND4_X1 U16930 ( .A1(n15289), .A2(n15288), .A3(n15287), .A4(n15286), .ZN(
        P2_U3228) );
  AOI22_X1 U16931 ( .A1(n15299), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n15298) );
  NAND2_X1 U16932 ( .A1(n15305), .A2(n15290), .ZN(n15297) );
  OAI211_X1 U16933 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15292), .A(n15306), 
        .B(n15291), .ZN(n15296) );
  OAI211_X1 U16934 ( .C1(n15294), .C2(P2_REG1_REG_15__SCAN_IN), .A(n15300), 
        .B(n15293), .ZN(n15295) );
  NAND4_X1 U16935 ( .A1(n15298), .A2(n15297), .A3(n15296), .A4(n15295), .ZN(
        P2_U3229) );
  AOI22_X1 U16936 ( .A1(n15299), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n15313) );
  OAI211_X1 U16937 ( .C1(n15303), .C2(n15302), .A(n15301), .B(n15300), .ZN(
        n15312) );
  NAND2_X1 U16938 ( .A1(n15305), .A2(n15304), .ZN(n15311) );
  OAI211_X1 U16939 ( .C1(n15309), .C2(n15308), .A(n15307), .B(n15306), .ZN(
        n15310) );
  NAND4_X1 U16940 ( .A1(n15313), .A2(n15312), .A3(n15311), .A4(n15310), .ZN(
        P2_U3231) );
  INV_X1 U16941 ( .A(n15320), .ZN(n15321) );
  AND2_X1 U16942 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15321), .ZN(P2_U3266) );
  AND2_X1 U16943 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15321), .ZN(P2_U3267) );
  AND2_X1 U16944 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15321), .ZN(P2_U3268) );
  NOR2_X1 U16945 ( .A1(n15320), .A2(n15315), .ZN(P2_U3269) );
  AND2_X1 U16946 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15321), .ZN(P2_U3270) );
  AND2_X1 U16947 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15321), .ZN(P2_U3271) );
  AND2_X1 U16948 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15321), .ZN(P2_U3272) );
  AND2_X1 U16949 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15321), .ZN(P2_U3273) );
  AND2_X1 U16950 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15321), .ZN(P2_U3274) );
  AND2_X1 U16951 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15321), .ZN(P2_U3275) );
  AND2_X1 U16952 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15321), .ZN(P2_U3276) );
  AND2_X1 U16953 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15321), .ZN(P2_U3277) );
  AND2_X1 U16954 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15321), .ZN(P2_U3278) );
  AND2_X1 U16955 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15321), .ZN(P2_U3279) );
  AND2_X1 U16956 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15321), .ZN(P2_U3280) );
  AND2_X1 U16957 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15321), .ZN(P2_U3281) );
  AND2_X1 U16958 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15321), .ZN(P2_U3282) );
  AND2_X1 U16959 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15321), .ZN(P2_U3283) );
  AND2_X1 U16960 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15321), .ZN(P2_U3284) );
  AND2_X1 U16961 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15321), .ZN(P2_U3285) );
  AND2_X1 U16962 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15321), .ZN(P2_U3286) );
  NOR2_X1 U16963 ( .A1(n15320), .A2(n15316), .ZN(P2_U3287) );
  AND2_X1 U16964 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15321), .ZN(P2_U3288) );
  AND2_X1 U16965 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15321), .ZN(P2_U3289) );
  AND2_X1 U16966 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15321), .ZN(P2_U3290) );
  NOR2_X1 U16967 ( .A1(n15320), .A2(n15317), .ZN(P2_U3291) );
  NOR2_X1 U16968 ( .A1(n15320), .A2(n15318), .ZN(P2_U3292) );
  NOR2_X1 U16969 ( .A1(n15320), .A2(n15319), .ZN(P2_U3293) );
  AND2_X1 U16970 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15321), .ZN(P2_U3294) );
  AND2_X1 U16971 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15321), .ZN(P2_U3295) );
  OAI21_X1 U16972 ( .B1(n15323), .B2(n15327), .A(n15322), .ZN(P2_U3416) );
  AOI22_X1 U16973 ( .A1(n15327), .A2(n15326), .B1(n15325), .B2(n15324), .ZN(
        P2_U3417) );
  INV_X1 U16974 ( .A(n15328), .ZN(n15330) );
  AOI211_X1 U16975 ( .C1(n7308), .C2(n15331), .A(n15330), .B(n15329), .ZN(
        n15384) );
  INV_X1 U16976 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15332) );
  AOI22_X1 U16977 ( .A1(n15383), .A2(n15384), .B1(n15332), .B2(n15381), .ZN(
        P2_U3430) );
  AOI21_X1 U16978 ( .B1(n15366), .B2(n6574), .A(n15333), .ZN(n15335) );
  OAI211_X1 U16979 ( .C1(n15352), .C2(n15336), .A(n15335), .B(n15334), .ZN(
        n15337) );
  INV_X1 U16980 ( .A(n15337), .ZN(n15385) );
  INV_X1 U16981 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15338) );
  AOI22_X1 U16982 ( .A1(n15383), .A2(n15385), .B1(n15338), .B2(n15381), .ZN(
        P2_U3433) );
  INV_X1 U16983 ( .A(n15339), .ZN(n15345) );
  NOR2_X1 U16984 ( .A1(n15339), .A2(n15369), .ZN(n15344) );
  OAI211_X1 U16985 ( .C1(n15342), .C2(n15376), .A(n15341), .B(n15340), .ZN(
        n15343) );
  AOI211_X1 U16986 ( .C1(n15362), .C2(n15345), .A(n15344), .B(n15343), .ZN(
        n15386) );
  INV_X1 U16987 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15346) );
  AOI22_X1 U16988 ( .A1(n15383), .A2(n15386), .B1(n15346), .B2(n15381), .ZN(
        P2_U3436) );
  AOI21_X1 U16989 ( .B1(n15366), .B2(n15348), .A(n15347), .ZN(n15350) );
  OAI211_X1 U16990 ( .C1(n15352), .C2(n15351), .A(n15350), .B(n15349), .ZN(
        n15353) );
  INV_X1 U16991 ( .A(n15353), .ZN(n15387) );
  INV_X1 U16992 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15354) );
  AOI22_X1 U16993 ( .A1(n15383), .A2(n15387), .B1(n15354), .B2(n15381), .ZN(
        P2_U3439) );
  INV_X1 U16994 ( .A(n15355), .ZN(n15361) );
  NOR2_X1 U16995 ( .A1(n15355), .A2(n15369), .ZN(n15360) );
  OAI211_X1 U16996 ( .C1(n15358), .C2(n15376), .A(n15357), .B(n15356), .ZN(
        n15359) );
  AOI211_X1 U16997 ( .C1(n15362), .C2(n15361), .A(n15360), .B(n15359), .ZN(
        n15388) );
  INV_X1 U16998 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15363) );
  AOI22_X1 U16999 ( .A1(n15383), .A2(n15388), .B1(n15363), .B2(n15381), .ZN(
        P2_U3442) );
  AOI21_X1 U17000 ( .B1(n15366), .B2(n15365), .A(n15364), .ZN(n15367) );
  OAI211_X1 U17001 ( .C1(n15370), .C2(n15369), .A(n15368), .B(n15367), .ZN(
        n15371) );
  INV_X1 U17002 ( .A(n15371), .ZN(n15389) );
  INV_X1 U17003 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15372) );
  AOI22_X1 U17004 ( .A1(n15383), .A2(n15389), .B1(n15372), .B2(n15381), .ZN(
        P2_U3448) );
  AND2_X1 U17005 ( .A1(n15374), .A2(n15373), .ZN(n15379) );
  OAI21_X1 U17006 ( .B1(n15377), .B2(n15376), .A(n15375), .ZN(n15378) );
  NOR3_X1 U17007 ( .A1(n15380), .A2(n15379), .A3(n15378), .ZN(n15391) );
  INV_X1 U17008 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15382) );
  AOI22_X1 U17009 ( .A1(n15383), .A2(n15391), .B1(n15382), .B2(n15381), .ZN(
        P2_U3463) );
  AOI22_X1 U17010 ( .A1(n15392), .A2(n15384), .B1(n7908), .B2(n15390), .ZN(
        P2_U3499) );
  AOI22_X1 U17011 ( .A1(n15392), .A2(n15385), .B1(n9496), .B2(n15390), .ZN(
        P2_U3500) );
  AOI22_X1 U17012 ( .A1(n15392), .A2(n15386), .B1(n9495), .B2(n15390), .ZN(
        P2_U3501) );
  AOI22_X1 U17013 ( .A1(n15392), .A2(n15387), .B1(n9494), .B2(n15390), .ZN(
        P2_U3502) );
  AOI22_X1 U17014 ( .A1(n15392), .A2(n15388), .B1(n9563), .B2(n15390), .ZN(
        P2_U3503) );
  AOI22_X1 U17015 ( .A1(n15392), .A2(n15389), .B1(n9578), .B2(n15390), .ZN(
        P2_U3505) );
  AOI22_X1 U17016 ( .A1(n15392), .A2(n15391), .B1(n9818), .B2(n15390), .ZN(
        P2_U3510) );
  NOR2_X1 U17017 ( .A1(P3_U3897), .A2(n15535), .ZN(P3_U3150) );
  INV_X1 U17018 ( .A(n15397), .ZN(n15393) );
  OAI21_X1 U17019 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n15394), .A(n15393), .ZN(
        n15395) );
  AOI22_X1 U17020 ( .A1(n15398), .A2(n15396), .B1(n15543), .B2(n15395), .ZN(
        n15405) );
  OAI21_X1 U17021 ( .B1(n15398), .B2(n15562), .A(n15397), .ZN(n15401) );
  AOI22_X1 U17022 ( .A1(n15562), .A2(n15399), .B1(n15535), .B2(
        P3_ADDR_REG_0__SCAN_IN), .ZN(n15400) );
  OAI211_X1 U17023 ( .C1(n15555), .C2(n15402), .A(n15401), .B(n15400), .ZN(
        n15403) );
  INV_X1 U17024 ( .A(n15403), .ZN(n15404) );
  OAI211_X1 U17025 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n10659), .A(n15405), .B(
        n15404), .ZN(P3_U3182) );
  AOI21_X1 U17026 ( .B1(n8820), .B2(n15408), .A(n15407), .ZN(n15424) );
  INV_X1 U17027 ( .A(n15409), .ZN(n15410) );
  OAI21_X1 U17028 ( .B1(n15559), .B2(n7187), .A(n15410), .ZN(n15417) );
  OR3_X1 U17029 ( .A1(n15413), .A2(n15412), .A3(n15411), .ZN(n15414) );
  AOI21_X1 U17030 ( .B1(n15415), .B2(n15414), .A(n15564), .ZN(n15416) );
  AOI211_X1 U17031 ( .C1(n15419), .C2(n15418), .A(n15417), .B(n15416), .ZN(
        n15423) );
  XNOR2_X1 U17032 ( .A(n15420), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n15421) );
  NAND2_X1 U17033 ( .A1(n15562), .A2(n15421), .ZN(n15422) );
  OAI211_X1 U17034 ( .C1(n15424), .C2(n15571), .A(n15423), .B(n15422), .ZN(
        P3_U3185) );
  AOI21_X1 U17035 ( .B1(n15427), .B2(n15426), .A(n15425), .ZN(n15442) );
  OAI21_X1 U17036 ( .B1(n15430), .B2(n15429), .A(n15428), .ZN(n15435) );
  AOI21_X1 U17037 ( .B1(n15535), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n15431), .ZN(
        n15432) );
  OAI21_X1 U17038 ( .B1(n15555), .B2(n15433), .A(n15432), .ZN(n15434) );
  AOI21_X1 U17039 ( .B1(n15435), .B2(n15543), .A(n15434), .ZN(n15441) );
  AND2_X1 U17040 ( .A1(n15437), .A2(n15436), .ZN(n15438) );
  OAI21_X1 U17041 ( .B1(n15439), .B2(n15438), .A(n15562), .ZN(n15440) );
  OAI211_X1 U17042 ( .C1(n15442), .C2(n15571), .A(n15441), .B(n15440), .ZN(
        P3_U3186) );
  AOI21_X1 U17043 ( .B1(n15445), .B2(n15444), .A(n15443), .ZN(n15460) );
  INV_X1 U17044 ( .A(n15446), .ZN(n15447) );
  NOR2_X1 U17045 ( .A1(n15448), .A2(n15447), .ZN(n15449) );
  XNOR2_X1 U17046 ( .A(n15450), .B(n15449), .ZN(n15455) );
  AOI21_X1 U17047 ( .B1(n15535), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n15451), .ZN(
        n15452) );
  OAI21_X1 U17048 ( .B1(n15555), .B2(n15453), .A(n15452), .ZN(n15454) );
  AOI21_X1 U17049 ( .B1(n15455), .B2(n15543), .A(n15454), .ZN(n15459) );
  XOR2_X1 U17050 ( .A(P3_REG1_REG_5__SCAN_IN), .B(n15456), .Z(n15457) );
  NAND2_X1 U17051 ( .A1(n15562), .A2(n15457), .ZN(n15458) );
  OAI211_X1 U17052 ( .C1(n15460), .C2(n15571), .A(n15459), .B(n15458), .ZN(
        P3_U3187) );
  AOI21_X1 U17053 ( .B1(n11359), .B2(n15462), .A(n15461), .ZN(n15476) );
  NAND2_X1 U17054 ( .A1(n15464), .A2(n15463), .ZN(n15465) );
  XNOR2_X1 U17055 ( .A(n15466), .B(n15465), .ZN(n15468) );
  OAI22_X1 U17056 ( .A1(n15468), .A2(n15564), .B1(n15467), .B2(n15555), .ZN(
        n15469) );
  AOI211_X1 U17057 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15535), .A(n15470), .B(
        n15469), .ZN(n15475) );
  OAI21_X1 U17058 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15472), .A(n15471), .ZN(
        n15473) );
  NAND2_X1 U17059 ( .A1(n15473), .A2(n15562), .ZN(n15474) );
  OAI211_X1 U17060 ( .C1(n15476), .C2(n15571), .A(n15475), .B(n15474), .ZN(
        P3_U3191) );
  AOI21_X1 U17061 ( .B1(n15479), .B2(n15478), .A(n15477), .ZN(n15494) );
  OAI21_X1 U17062 ( .B1(n15482), .B2(n15481), .A(n15480), .ZN(n15487) );
  AOI21_X1 U17063 ( .B1(n15535), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n15483), 
        .ZN(n15484) );
  OAI21_X1 U17064 ( .B1(n15555), .B2(n15485), .A(n15484), .ZN(n15486) );
  AOI21_X1 U17065 ( .B1(n15487), .B2(n15562), .A(n15486), .ZN(n15493) );
  OAI21_X1 U17066 ( .B1(n15490), .B2(n15489), .A(n15488), .ZN(n15491) );
  NAND2_X1 U17067 ( .A1(n15491), .A2(n15543), .ZN(n15492) );
  OAI211_X1 U17068 ( .C1(n15494), .C2(n15571), .A(n15493), .B(n15492), .ZN(
        P3_U3192) );
  AOI21_X1 U17069 ( .B1(n11417), .B2(n15496), .A(n15495), .ZN(n15510) );
  OAI21_X1 U17070 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n15498), .A(n15497), 
        .ZN(n15503) );
  AOI21_X1 U17071 ( .B1(n15535), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n15499), 
        .ZN(n15500) );
  OAI21_X1 U17072 ( .B1(n15555), .B2(n15501), .A(n15500), .ZN(n15502) );
  AOI21_X1 U17073 ( .B1(n15503), .B2(n15562), .A(n15502), .ZN(n15509) );
  OAI21_X1 U17074 ( .B1(n15506), .B2(n15505), .A(n15504), .ZN(n15507) );
  NAND2_X1 U17075 ( .A1(n15507), .A2(n15543), .ZN(n15508) );
  OAI211_X1 U17076 ( .C1(n15510), .C2(n15571), .A(n15509), .B(n15508), .ZN(
        P3_U3193) );
  AOI21_X1 U17077 ( .B1(n15513), .B2(n15512), .A(n15511), .ZN(n15528) );
  OAI21_X1 U17078 ( .B1(n15516), .B2(n15515), .A(n15514), .ZN(n15521) );
  AOI21_X1 U17079 ( .B1(n15535), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n15517), 
        .ZN(n15518) );
  OAI21_X1 U17080 ( .B1(n15555), .B2(n15519), .A(n15518), .ZN(n15520) );
  AOI21_X1 U17081 ( .B1(n15521), .B2(n15562), .A(n15520), .ZN(n15527) );
  AOI21_X1 U17082 ( .B1(n15523), .B2(n15522), .A(n15564), .ZN(n15525) );
  NAND2_X1 U17083 ( .A1(n15525), .A2(n15524), .ZN(n15526) );
  OAI211_X1 U17084 ( .C1(n15528), .C2(n15571), .A(n15527), .B(n15526), .ZN(
        P3_U3194) );
  AOI21_X1 U17085 ( .B1(n15531), .B2(n15530), .A(n15529), .ZN(n15547) );
  OAI21_X1 U17086 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n15533), .A(n15532), 
        .ZN(n15539) );
  AOI21_X1 U17087 ( .B1(n15535), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n15534), 
        .ZN(n15536) );
  OAI21_X1 U17088 ( .B1(n15555), .B2(n15537), .A(n15536), .ZN(n15538) );
  AOI21_X1 U17089 ( .B1(n15539), .B2(n15562), .A(n15538), .ZN(n15546) );
  OAI21_X1 U17090 ( .B1(n15542), .B2(n15541), .A(n15540), .ZN(n15544) );
  NAND2_X1 U17091 ( .A1(n15544), .A2(n15543), .ZN(n15545) );
  OAI211_X1 U17092 ( .C1(n15547), .C2(n15571), .A(n15546), .B(n15545), .ZN(
        P3_U3195) );
  AOI21_X1 U17093 ( .B1(n15550), .B2(n15549), .A(n15548), .ZN(n15572) );
  OAI21_X1 U17094 ( .B1(n15553), .B2(n15552), .A(n15551), .ZN(n15563) );
  NOR2_X1 U17095 ( .A1(n15555), .A2(n15554), .ZN(n15561) );
  INV_X1 U17096 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15558) );
  INV_X1 U17097 ( .A(n15556), .ZN(n15557) );
  OAI21_X1 U17098 ( .B1(n15559), .B2(n15558), .A(n15557), .ZN(n15560) );
  AOI211_X1 U17099 ( .C1(n15563), .C2(n15562), .A(n15561), .B(n15560), .ZN(
        n15570) );
  AOI21_X1 U17100 ( .B1(n15566), .B2(n15565), .A(n15564), .ZN(n15568) );
  NAND2_X1 U17101 ( .A1(n15568), .A2(n15567), .ZN(n15569) );
  OAI211_X1 U17102 ( .C1(n15572), .C2(n15571), .A(n15570), .B(n15569), .ZN(
        P3_U3196) );
  INV_X1 U17103 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15574) );
  AOI22_X1 U17104 ( .A1(n15601), .A2(n15574), .B1(n15573), .B2(n15599), .ZN(
        P3_U3393) );
  INV_X1 U17105 ( .A(n15575), .ZN(n15577) );
  AOI211_X1 U17106 ( .C1(n15591), .C2(n15578), .A(n15577), .B(n15576), .ZN(
        n15602) );
  AOI22_X1 U17107 ( .A1(n15601), .A2(n15579), .B1(n15602), .B2(n15599), .ZN(
        P3_U3396) );
  INV_X1 U17108 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15584) );
  INV_X1 U17109 ( .A(n15580), .ZN(n15581) );
  AOI211_X1 U17110 ( .C1(n15583), .C2(n15591), .A(n15582), .B(n15581), .ZN(
        n15603) );
  AOI22_X1 U17111 ( .A1(n15601), .A2(n15584), .B1(n15603), .B2(n15599), .ZN(
        P3_U3405) );
  INV_X1 U17112 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15588) );
  AOI211_X1 U17113 ( .C1(n15591), .C2(n15587), .A(n15586), .B(n15585), .ZN(
        n15605) );
  AOI22_X1 U17114 ( .A1(n15601), .A2(n15588), .B1(n15605), .B2(n15599), .ZN(
        P3_U3414) );
  INV_X1 U17115 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15593) );
  AOI211_X1 U17116 ( .C1(n15592), .C2(n15591), .A(n15590), .B(n15589), .ZN(
        n15607) );
  AOI22_X1 U17117 ( .A1(n15601), .A2(n15593), .B1(n15607), .B2(n15599), .ZN(
        P3_U3417) );
  INV_X1 U17118 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15600) );
  NAND3_X1 U17119 ( .A1(n11409), .A2(n15595), .A3(n15594), .ZN(n15596) );
  AND3_X1 U17120 ( .A1(n15598), .A2(n15597), .A3(n15596), .ZN(n15610) );
  AOI22_X1 U17121 ( .A1(n15601), .A2(n15600), .B1(n15610), .B2(n15599), .ZN(
        P3_U3420) );
  AOI22_X1 U17122 ( .A1(n15611), .A2(n15602), .B1(n10186), .B2(n15608), .ZN(
        P3_U3461) );
  AOI22_X1 U17123 ( .A1(n15611), .A2(n15603), .B1(n10367), .B2(n15608), .ZN(
        P3_U3464) );
  AOI22_X1 U17124 ( .A1(n15611), .A2(n15605), .B1(n15604), .B2(n15608), .ZN(
        P3_U3467) );
  AOI22_X1 U17125 ( .A1(n15611), .A2(n15607), .B1(n15606), .B2(n15608), .ZN(
        P3_U3468) );
  AOI22_X1 U17126 ( .A1(n15611), .A2(n15610), .B1(n15609), .B2(n15608), .ZN(
        P3_U3469) );
  AOI21_X1 U17127 ( .B1(n15614), .B2(n15613), .A(n15612), .ZN(SUB_1596_U59) );
  OAI21_X1 U17128 ( .B1(n15617), .B2(n15616), .A(n15615), .ZN(SUB_1596_U58) );
  XOR2_X1 U17129 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15618), .Z(SUB_1596_U53) );
  AOI21_X1 U17130 ( .B1(n15621), .B2(n15620), .A(n15619), .ZN(SUB_1596_U56) );
  AOI21_X1 U17131 ( .B1(n15624), .B2(n15623), .A(n15622), .ZN(n15625) );
  XOR2_X1 U17132 ( .A(n15625), .B(P2_ADDR_REG_3__SCAN_IN), .Z(SUB_1596_U60) );
  AOI21_X1 U17133 ( .B1(n15628), .B2(n15627), .A(n15626), .ZN(SUB_1596_U5) );
  CLKBUF_X1 U7517 ( .A(n8334), .Z(n9476) );
endmodule

