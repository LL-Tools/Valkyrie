

module b17_C_SARLock_k_64_8 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, U355, U356, U357, U358, 
        U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, 
        U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, 
        U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, 
        U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, 
        U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, 
        U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, 
        U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, 
        U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9605,
         n9606, n9607, n9608, n9609, n9611, n9612, n9613, n9614, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861;

  OR2_X1 U11040 ( .A1(n14839), .A2(n10100), .ZN(n14802) );
  INV_X1 U11041 ( .A(n14921), .ZN(n14909) );
  NAND2_X1 U11042 ( .A1(n17516), .A2(n17631), .ZN(n17764) );
  NAND2_X1 U11043 ( .A1(n11440), .A2(n11439), .ZN(n13964) );
  CLKBUF_X3 U11044 ( .A(n15825), .Z(n9618) );
  CLKBUF_X2 U11045 ( .A(n14425), .Z(n9617) );
  CLKBUF_X2 U11046 ( .A(n11207), .Z(n9603) );
  INV_X2 U11047 ( .A(n17097), .ZN(n17077) );
  AND2_X1 U11049 ( .A1(n12383), .A2(n10259), .ZN(n10572) );
  CLKBUF_X2 U11050 ( .A(n10316), .Z(n12378) );
  CLKBUF_X2 U11051 ( .A(n11694), .Z(n9607) );
  INV_X1 U11052 ( .A(n10165), .ZN(n17039) );
  CLKBUF_X2 U11053 ( .A(n17109), .Z(n9600) );
  AND2_X1 U11054 ( .A1(n11043), .A2(n11038), .ZN(n11073) );
  AND2_X1 U11055 ( .A1(n11043), .A2(n13203), .ZN(n11123) );
  AND2_X1 U11056 ( .A1(n11045), .A2(n13203), .ZN(n11186) );
  AND2_X1 U11057 ( .A1(n11045), .A2(n11038), .ZN(n11138) );
  NAND2_X2 U11060 ( .A1(n9765), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12445) );
  AND2_X1 U11061 ( .A1(n13300), .A2(n13301), .ZN(n9599) );
  AND2_X1 U11062 ( .A1(n13300), .A2(n13301), .ZN(n12383) );
  INV_X4 U11063 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13301) );
  NOR2_X2 U11064 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13324) );
  CLKBUF_X1 U11065 ( .A(n20820), .Z(n9595) );
  NOR2_X1 U11066 ( .A1(n20775), .A2(n20858), .ZN(n20820) );
  OAI22_X1 U11067 ( .A1(n10517), .A2(n12225), .B1(n19558), .B2(n10516), .ZN(
        n10518) );
  NAND3_X1 U11068 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U11069 ( .A1(n9824), .A2(n10416), .ZN(n10437) );
  AND2_X1 U11070 ( .A1(n10364), .A2(n10372), .ZN(n12895) );
  INV_X2 U11071 ( .A(n9777), .ZN(n13874) );
  OR2_X1 U11072 ( .A1(n10666), .A2(n10665), .ZN(n13728) );
  BUF_X1 U11073 ( .A(n12441), .Z(n17106) );
  INV_X1 U11074 ( .A(n12441), .ZN(n16949) );
  INV_X1 U11075 ( .A(n12420), .ZN(n16906) );
  OAI21_X1 U11076 ( .B1(n14458), .B2(n10138), .A(n10137), .ZN(n12323) );
  INV_X2 U11077 ( .A(n19188), .ZN(n10362) );
  AOI21_X1 U11078 ( .B1(n14898), .B2(n14896), .A(n14883), .ZN(n14887) );
  INV_X2 U11079 ( .A(n17005), .ZN(n12486) );
  INV_X2 U11080 ( .A(n17109), .ZN(n17038) );
  INV_X1 U11081 ( .A(n17764), .ZN(n17754) );
  NAND2_X1 U11082 ( .A1(n17556), .A2(n17670), .ZN(n17522) );
  INV_X1 U11083 ( .A(n19958), .ZN(n19925) );
  OAI211_X1 U11084 ( .C1(n9865), .C2(n11891), .A(n9636), .B(n9858), .ZN(n13607) );
  NAND2_X1 U11085 ( .A1(n10394), .A2(n13369), .ZN(n16215) );
  OR2_X1 U11087 ( .A1(n15234), .A2(n9947), .ZN(n14921) );
  NOR2_X1 U11088 ( .A1(n11960), .A2(n16160), .ZN(n11963) );
  NAND2_X1 U11089 ( .A1(n14967), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15234) );
  NAND2_X1 U11090 ( .A1(n16123), .A2(n10674), .ZN(n14837) );
  INV_X1 U11091 ( .A(n16749), .ZN(n16692) );
  INV_X1 U11092 ( .A(n10165), .ZN(n17101) );
  OAI21_X1 U11093 ( .B1(n15603), .B2(n15602), .A(n18771), .ZN(n17152) );
  INV_X1 U11094 ( .A(n17678), .ZN(n17607) );
  INV_X1 U11095 ( .A(n19905), .ZN(n19920) );
  INV_X1 U11096 ( .A(n19961), .ZN(n19948) );
  INV_X1 U11097 ( .A(n16761), .ZN(n16777) );
  INV_X1 U11098 ( .A(n16770), .ZN(n16789) );
  OR2_X1 U11099 ( .A1(n12407), .A2(n12404), .ZN(n9596) );
  CLKBUF_X3 U11100 ( .A(n20157), .Z(n9614) );
  NOR2_X2 U11101 ( .A1(n17195), .A2(n17364), .ZN(n17194) );
  AND2_X1 U11102 ( .A1(n11043), .A2(n12999), .ZN(n11207) );
  NOR2_X2 U11103 ( .A1(n16112), .A2(n10765), .ZN(n14967) );
  OAI21_X1 U11104 ( .B1(n13229), .B2(n13227), .A(n13228), .ZN(n19791) );
  AOI21_X2 U11105 ( .B1(n14929), .B2(n13691), .A(n10794), .ZN(n14919) );
  OAI21_X2 U11106 ( .B1(n9782), .B2(n15548), .A(n12978), .ZN(n13029) );
  OAI21_X2 U11107 ( .B1(n16274), .B2(n17670), .A(n17436), .ZN(n17428) );
  INV_X4 U11109 ( .A(n10388), .ZN(n15359) );
  AND2_X2 U11110 ( .A1(n9913), .A2(n9908), .ZN(n9907) );
  INV_X1 U11111 ( .A(n12445), .ZN(n9597) );
  INV_X1 U11112 ( .A(n12445), .ZN(n9598) );
  NOR2_X1 U11113 ( .A1(n18563), .A2(n18722), .ZN(n17109) );
  NAND2_X2 U11114 ( .A1(n14461), .A2(n12273), .ZN(n12293) );
  AND2_X4 U11115 ( .A1(n11044), .A2(n11043), .ZN(n11329) );
  INV_X4 U11116 ( .A(n12442), .ZN(n17087) );
  NAND2_X2 U11117 ( .A1(n14837), .A2(n13754), .ZN(n14839) );
  CLKBUF_X1 U11118 ( .A(n10491), .Z(n9601) );
  NOR2_X2 U11120 ( .A1(n11982), .A2(n14821), .ZN(n11953) );
  BUF_X4 U11122 ( .A(n11084), .Z(n9605) );
  CLKBUF_X3 U11123 ( .A(n11694), .Z(n9606) );
  AOI211_X2 U11124 ( .C1(n18050), .C2(n16281), .A(n16280), .B(n16279), .ZN(
        n16282) );
  NOR2_X1 U11125 ( .A1(n17276), .A2(n17774), .ZN(n9608) );
  INV_X1 U11126 ( .A(n17664), .ZN(n17682) );
  OR2_X1 U11127 ( .A1(n9948), .A2(n15219), .ZN(n15193) );
  OR2_X1 U11128 ( .A1(n13885), .A2(n11774), .ZN(n14026) );
  OR2_X1 U11129 ( .A1(n14032), .A2(n10084), .ZN(n13891) );
  AND2_X1 U11130 ( .A1(n11918), .A2(n15773), .ZN(n14298) );
  AND2_X1 U11131 ( .A1(n9748), .A2(n9747), .ZN(n10671) );
  NAND2_X1 U11132 ( .A1(n11906), .A2(n9618), .ZN(n15773) );
  AND2_X1 U11133 ( .A1(n9842), .A2(n9683), .ZN(n14321) );
  OR3_X2 U11134 ( .A1(n13964), .A2(n10079), .A3(n10082), .ZN(n9656) );
  OAI21_X1 U11135 ( .B1(n11892), .B2(n13607), .A(n13605), .ZN(n15834) );
  NAND2_X1 U11136 ( .A1(n12523), .A2(n12522), .ZN(n12528) );
  NAND2_X1 U11137 ( .A1(n9861), .A2(n9860), .ZN(n9864) );
  NAND2_X1 U11138 ( .A1(n12684), .A2(n17676), .ZN(n17636) );
  OR2_X1 U11139 ( .A1(n14238), .A2(n14239), .ZN(n9785) );
  INV_X1 U11140 ( .A(n11900), .ZN(n15825) );
  NAND2_X1 U11141 ( .A1(n17975), .A2(n12524), .ZN(n18028) );
  NAND2_X1 U11142 ( .A1(n13712), .A2(n10802), .ZN(n10804) );
  NAND2_X1 U11143 ( .A1(n10483), .A2(n13351), .ZN(n19486) );
  NOR2_X1 U11144 ( .A1(n9657), .A2(n13942), .ZN(n14063) );
  NOR2_X1 U11145 ( .A1(n17152), .A2(n17383), .ZN(n17304) );
  NOR2_X1 U11146 ( .A1(n10478), .A2(n10458), .ZN(n10509) );
  NOR2_X1 U11147 ( .A1(n18559), .A2(n18583), .ZN(n17889) );
  NOR2_X1 U11148 ( .A1(n9893), .A2(n10443), .ZN(n10444) );
  INV_X2 U11149 ( .A(n18585), .ZN(n18559) );
  AND2_X1 U11150 ( .A1(n13596), .A2(n13558), .ZN(n13557) );
  NAND2_X1 U11151 ( .A1(n11252), .A2(n11251), .ZN(n12986) );
  NOR2_X1 U11152 ( .A1(n17348), .A2(n17411), .ZN(n17404) );
  NAND2_X1 U11153 ( .A1(n10410), .A2(n10381), .ZN(n10428) );
  AND2_X2 U11154 ( .A1(n10392), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10432) );
  AND2_X1 U11155 ( .A1(n12641), .A2(n9934), .ZN(n17347) );
  AOI21_X1 U11156 ( .B1(n12973), .B2(n14406), .A(n11160), .ZN(n11163) );
  INV_X1 U11157 ( .A(n18763), .ZN(n18125) );
  AOI211_X2 U11158 ( .C1(n17078), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n12440), .B(n12439), .ZN(n17292) );
  NAND2_X1 U11159 ( .A1(n10382), .A2(n10808), .ZN(n12893) );
  INV_X1 U11160 ( .A(n10808), .ZN(n10698) );
  NAND3_X1 U11161 ( .A1(n9814), .A2(n9808), .A3(n12599), .ZN(n18158) );
  OR2_X1 U11162 ( .A1(n10328), .A2(n10327), .ZN(n10833) );
  AND2_X1 U11163 ( .A1(n11147), .A2(n11154), .ZN(n11159) );
  OR2_X1 U11164 ( .A1(n11107), .A2(n11106), .ZN(n20162) );
  INV_X4 U11165 ( .A(n12405), .ZN(n17073) );
  INV_X4 U11166 ( .A(n10169), .ZN(n17070) );
  CLKBUF_X2 U11167 ( .A(n11186), .Z(n11693) );
  BUF_X2 U11169 ( .A(n11073), .Z(n13772) );
  BUF_X2 U11170 ( .A(n11191), .Z(n13784) );
  CLKBUF_X2 U11171 ( .A(n11123), .Z(n13775) );
  CLKBUF_X2 U11172 ( .A(n11089), .Z(n11708) );
  CLKBUF_X2 U11173 ( .A(n12377), .Z(n12370) );
  AND2_X1 U11174 ( .A1(n11038), .A2(n13186), .ZN(n11100) );
  INV_X4 U11175 ( .A(n16801), .ZN(n17095) );
  INV_X2 U11176 ( .A(n17100), .ZN(n12418) );
  CLKBUF_X2 U11177 ( .A(n11133), .Z(n13774) );
  INV_X2 U11178 ( .A(n13321), .ZN(n10317) );
  NOR2_X2 U11179 ( .A1(n11036), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11043) );
  NOR2_X1 U11180 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10172) );
  INV_X2 U11181 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11268) );
  AND2_X1 U11182 ( .A1(n9891), .A2(n9890), .ZN(n14775) );
  INV_X1 U11183 ( .A(n9866), .ZN(n16264) );
  AOI211_X1 U11184 ( .C1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n13768), .A(
        n13767), .B(n13766), .ZN(n13769) );
  OAI21_X1 U11185 ( .B1(n15982), .B2(n15983), .A(n19000), .ZN(n10027) );
  NAND2_X1 U11186 ( .A1(n9902), .A2(n9900), .ZN(n14786) );
  OAI21_X1 U11187 ( .B1(n15109), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15108), .ZN(n16095) );
  NAND2_X1 U11188 ( .A1(n15094), .A2(n9671), .ZN(n9902) );
  NAND2_X1 U11189 ( .A1(n14845), .A2(n14844), .ZN(n15094) );
  AOI21_X1 U11190 ( .B1(n15623), .B2(n20070), .A(n11835), .ZN(n11917) );
  NAND2_X1 U11191 ( .A1(n9906), .A2(n9904), .ZN(n14845) );
  AND2_X1 U11192 ( .A1(n14173), .A2(n11920), .ZN(n10148) );
  NAND2_X1 U11193 ( .A1(n11908), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11909) );
  XNOR2_X1 U11194 ( .A(n13891), .B(n13809), .ZN(n13817) );
  AND3_X1 U11195 ( .A1(n14300), .A2(n13818), .A3(n9741), .ZN(n14163) );
  AND2_X1 U11196 ( .A1(n9660), .A2(n14033), .ZN(n15763) );
  AND2_X1 U11197 ( .A1(n12534), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16274) );
  AND2_X1 U11198 ( .A1(n14061), .A2(n14047), .ZN(n15787) );
  AND2_X1 U11199 ( .A1(n10653), .A2(n10652), .ZN(n9946) );
  XNOR2_X1 U11200 ( .A(n10743), .B(n15284), .ZN(n15294) );
  NAND3_X1 U11201 ( .A1(n9758), .A2(n15300), .A3(n10582), .ZN(n15304) );
  NOR2_X1 U11202 ( .A1(n17474), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17473) );
  OAI21_X1 U11203 ( .B1(n9874), .B2(n17662), .A(n9871), .ZN(n17503) );
  OR2_X1 U11204 ( .A1(n10108), .A2(n10105), .ZN(n9666) );
  NAND2_X1 U11205 ( .A1(n9874), .A2(n9876), .ZN(n17556) );
  CLKBUF_X1 U11206 ( .A(n17573), .Z(n9613) );
  NOR2_X1 U11207 ( .A1(n9845), .A2(n9844), .ZN(n9843) );
  NAND2_X1 U11208 ( .A1(n9950), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17188) );
  AND2_X1 U11209 ( .A1(n18612), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18717) );
  NAND2_X1 U11210 ( .A1(n17606), .A2(n17636), .ZN(n17955) );
  AND2_X1 U11211 ( .A1(n10553), .A2(n10552), .ZN(n10566) );
  INV_X1 U11212 ( .A(n10615), .ZN(n9609) );
  XOR2_X1 U11213 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11882), .Z(
        n13468) );
  OR2_X1 U11214 ( .A1(n14340), .A2(n14336), .ZN(n9846) );
  NAND2_X1 U11215 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17656), .ZN(n17631) );
  OR3_X1 U11216 ( .A1(n10600), .A2(n10599), .A3(n10598), .ZN(n10613) );
  NOR2_X1 U11217 ( .A1(n14255), .A2(n15957), .ZN(n14254) );
  AND2_X1 U11218 ( .A1(n13252), .A2(n11408), .ZN(n9633) );
  INV_X1 U11219 ( .A(n17770), .ZN(n17757) );
  OAI211_X1 U11220 ( .C1(n13797), .C2(n11384), .A(n11383), .B(n11382), .ZN(
        n13252) );
  AOI21_X1 U11221 ( .B1(n9752), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A(n9751), 
        .ZN(n9750) );
  OR2_X1 U11222 ( .A1(n10475), .A2(n10474), .ZN(n10476) );
  NOR2_X1 U11223 ( .A1(n14954), .A2(n9909), .ZN(n9828) );
  NAND2_X1 U11224 ( .A1(n14042), .A2(n13917), .ZN(n14029) );
  OR2_X1 U11225 ( .A1(n13293), .A2(n10467), .ZN(n19249) );
  NOR2_X1 U11226 ( .A1(n17296), .A2(n17151), .ZN(n17234) );
  AND2_X1 U11227 ( .A1(n10482), .A2(n10461), .ZN(n19551) );
  XNOR2_X1 U11228 ( .A(n11846), .B(n11386), .ZN(n11838) );
  NAND2_X1 U11229 ( .A1(n11846), .A2(n11837), .ZN(n11900) );
  OR2_X1 U11230 ( .A1(n13293), .A2(n10471), .ZN(n10622) );
  NAND2_X1 U11231 ( .A1(n10483), .A2(n19158), .ZN(n10629) );
  AND2_X1 U11232 ( .A1(n10482), .A2(n10459), .ZN(n15381) );
  NAND2_X1 U11233 ( .A1(n11381), .A2(n9787), .ZN(n11846) );
  NAND2_X1 U11234 ( .A1(n12678), .A2(n17700), .ZN(n17689) );
  AND2_X1 U11235 ( .A1(n10482), .A2(n12969), .ZN(n10483) );
  NAND2_X1 U11236 ( .A1(n17684), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17683) );
  NAND2_X1 U11237 ( .A1(n18875), .A2(n18876), .ZN(n18874) );
  XNOR2_X1 U11238 ( .A(n12516), .B(n12515), .ZN(n17684) );
  XNOR2_X1 U11239 ( .A(n11279), .B(n11278), .ZN(n14386) );
  NAND2_X1 U11240 ( .A1(n10773), .A2(n10772), .ZN(n10782) );
  NAND2_X1 U11241 ( .A1(n10017), .A2(n10016), .ZN(n12516) );
  AOI21_X1 U11242 ( .B1(n11858), .B2(n11277), .A(n11239), .ZN(n11299) );
  INV_X1 U11243 ( .A(n14395), .ZN(n14394) );
  INV_X1 U11244 ( .A(n19023), .ZN(n16204) );
  XNOR2_X1 U11245 ( .A(n11238), .B(n11236), .ZN(n11277) );
  AOI21_X1 U11246 ( .B1(n20428), .B2(n20754), .A(n9784), .ZN(n14395) );
  NOR2_X2 U11247 ( .A1(n19091), .A2(n19285), .ZN(n13539) );
  NAND2_X1 U11248 ( .A1(n11230), .A2(n11229), .ZN(n11238) );
  NOR2_X2 U11249 ( .A1(n16089), .A2(n19285), .ZN(n13567) );
  NOR2_X2 U11250 ( .A1(n15340), .A2(n19285), .ZN(n15341) );
  NAND2_X1 U11251 ( .A1(n17730), .A2(n12511), .ZN(n17714) );
  XNOR2_X1 U11252 ( .A(n12986), .B(n20305), .ZN(n20428) );
  OAI21_X1 U11253 ( .B1(n11869), .B2(n11868), .A(n11867), .ZN(n13028) );
  XNOR2_X1 U11254 ( .A(n11286), .B(n11285), .ZN(n11869) );
  NAND2_X1 U11255 ( .A1(n9763), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17730) );
  NAND2_X1 U11256 ( .A1(n11245), .A2(n11244), .ZN(n11252) );
  NAND2_X1 U11257 ( .A1(n12779), .A2(n12833), .ZN(n12812) );
  CLKBUF_X1 U11258 ( .A(n17404), .Z(n17412) );
  XNOR2_X1 U11259 ( .A(n12509), .B(n12508), .ZN(n9763) );
  NOR2_X1 U11260 ( .A1(n9951), .A2(n12646), .ZN(n9914) );
  NAND2_X1 U11261 ( .A1(n20267), .A2(n11185), .ZN(n11245) );
  NAND2_X1 U11262 ( .A1(n17738), .A2(n12506), .ZN(n12509) );
  INV_X2 U11263 ( .A(n10985), .ZN(n13743) );
  OAI211_X1 U11264 ( .C1(n15551), .C2(n20429), .A(n11248), .B(n11247), .ZN(
        n11251) );
  NAND2_X1 U11265 ( .A1(n11303), .A2(n11302), .ZN(n20305) );
  NAND2_X1 U11266 ( .A1(n10413), .A2(n10152), .ZN(n10440) );
  NAND2_X1 U11267 ( .A1(n17739), .A2(n17740), .ZN(n17738) );
  OAI211_X1 U11268 ( .C1(n17750), .C2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n9769), .B(n9767), .ZN(n17739) );
  AOI21_X1 U11269 ( .B1(n10432), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n10421), .ZN(n10424) );
  AND2_X1 U11270 ( .A1(n17698), .A2(n10021), .ZN(n10020) );
  OR2_X1 U11271 ( .A1(n11246), .A2(n11272), .ZN(n11248) );
  OAI21_X1 U11272 ( .B1(n12640), .B2(n12639), .A(n13651), .ZN(n12646) );
  AOI21_X1 U11273 ( .B1(n10432), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10435), .ZN(n10964) );
  AND2_X1 U11274 ( .A1(n9933), .A2(n12632), .ZN(n16399) );
  OR2_X2 U11275 ( .A1(n18611), .A2(n17345), .ZN(n17414) );
  OR2_X1 U11276 ( .A1(n10411), .A2(n19855), .ZN(n10412) );
  AOI21_X1 U11277 ( .B1(n10402), .B2(n9670), .A(n9892), .ZN(n10404) );
  AND2_X1 U11278 ( .A1(n10379), .A2(n10378), .ZN(n10410) );
  NAND2_X1 U11279 ( .A1(n17751), .A2(n17752), .ZN(n17750) );
  AOI21_X1 U11280 ( .B1(n9852), .B2(n9780), .A(n9707), .ZN(n9778) );
  NAND2_X1 U11281 ( .A1(n12513), .A2(n12656), .ZN(n16276) );
  OAI211_X1 U11282 ( .C1(n10097), .C2(n10094), .A(n10096), .B(n10092), .ZN(
        n10379) );
  NAND2_X1 U11283 ( .A1(n17759), .A2(n12500), .ZN(n17751) );
  NOR2_X1 U11284 ( .A1(n12655), .A2(n12512), .ZN(n12513) );
  NAND2_X1 U11285 ( .A1(n11163), .A2(n11180), .ZN(n9852) );
  OAI21_X1 U11286 ( .B1(n13345), .B2(n10400), .A(n9635), .ZN(n9892) );
  AND2_X1 U11287 ( .A1(n10355), .A2(n10354), .ZN(n10356) );
  NAND2_X1 U11288 ( .A1(n10313), .A2(n9756), .ZN(n10363) );
  AND2_X1 U11289 ( .A1(n10312), .A2(n12900), .ZN(n10313) );
  OR2_X1 U11290 ( .A1(n11157), .A2(n11156), .ZN(n12973) );
  AND2_X1 U11291 ( .A1(n12895), .A2(n9746), .ZN(n9745) );
  OR2_X1 U11292 ( .A1(n18088), .A2(n12502), .ZN(n12503) );
  XNOR2_X1 U11293 ( .A(n12502), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17752) );
  INV_X1 U11294 ( .A(n10382), .ZN(n12894) );
  NAND2_X1 U11295 ( .A1(n13874), .A2(n11170), .ZN(n13877) );
  OR2_X1 U11296 ( .A1(n11172), .A2(n13054), .ZN(n11176) );
  AOI211_X2 U11297 ( .C1(n17102), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n12624), .B(n12623), .ZN(n18763) );
  INV_X1 U11298 ( .A(n12667), .ZN(n12501) );
  INV_X4 U11299 ( .A(n10755), .ZN(n19180) );
  AND2_X1 U11300 ( .A1(n11972), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11974) );
  AND2_X1 U11301 ( .A1(n10150), .A2(n10168), .ZN(n9743) );
  OAI211_X1 U11302 ( .C1(n17087), .C2(n17128), .A(n12596), .B(n12595), .ZN(
        n18148) );
  CLKBUF_X3 U11303 ( .A(n10811), .Z(n10755) );
  NAND2_X1 U11304 ( .A1(n11159), .A2(n11158), .ZN(n14406) );
  NOR2_X1 U11305 ( .A1(n11227), .A2(n20754), .ZN(n11836) );
  NAND2_X1 U11306 ( .A1(n12452), .A2(n9770), .ZN(n12667) );
  AND2_X1 U11307 ( .A1(n11148), .A2(n11776), .ZN(n9783) );
  AND2_X1 U11308 ( .A1(n11155), .A2(n11154), .ZN(n11778) );
  INV_X2 U11309 ( .A(n16287), .ZN(n16338) );
  NOR2_X1 U11310 ( .A1(n12906), .A2(n20162), .ZN(n13149) );
  OR2_X1 U11311 ( .A1(n10578), .A2(n10577), .ZN(n10813) );
  AND3_X1 U11312 ( .A1(n12906), .A2(n19976), .A3(n12971), .ZN(n9816) );
  INV_X1 U11313 ( .A(n20162), .ZN(n11776) );
  INV_X1 U11314 ( .A(n11287), .ZN(n20188) );
  OR2_X2 U11315 ( .A1(n11072), .A2(n11071), .ZN(n11154) );
  OR2_X1 U11316 ( .A1(n11213), .A2(n11212), .ZN(n11895) );
  INV_X1 U11317 ( .A(n20182), .ZN(n12971) );
  NAND4_X1 U11318 ( .A1(n11146), .A2(n11145), .A3(n11144), .A4(n11143), .ZN(
        n20157) );
  NOR2_X2 U11319 ( .A1(n11051), .A2(n11050), .ZN(n11287) );
  NOR2_X2 U11320 ( .A1(n20149), .A2(n20147), .ZN(n20148) );
  AND4_X1 U11321 ( .A1(n11137), .A2(n11136), .A3(n11135), .A4(n11134), .ZN(
        n11144) );
  AND4_X1 U11322 ( .A1(n11142), .A2(n11141), .A3(n11140), .A4(n11139), .ZN(
        n11143) );
  AND4_X1 U11323 ( .A1(n11077), .A2(n11076), .A3(n11075), .A4(n11074), .ZN(
        n11083) );
  AND4_X1 U11324 ( .A1(n11081), .A2(n11080), .A3(n11079), .A4(n11078), .ZN(
        n11082) );
  AND4_X1 U11325 ( .A1(n11127), .A2(n11126), .A3(n11125), .A4(n11124), .ZN(
        n11146) );
  AND4_X1 U11326 ( .A1(n11132), .A2(n11131), .A3(n11130), .A4(n11129), .ZN(
        n11145) );
  INV_X2 U11327 ( .A(n9596), .ZN(n17075) );
  INV_X4 U11328 ( .A(n17073), .ZN(n16812) );
  INV_X1 U11329 ( .A(n9596), .ZN(n17092) );
  AND4_X1 U11330 ( .A1(n10237), .A2(n10236), .A3(n10235), .A4(n10234), .ZN(
        n10238) );
  AND4_X1 U11331 ( .A1(n10233), .A2(n10232), .A3(n10231), .A4(n10230), .ZN(
        n10239) );
  AND2_X2 U11332 ( .A1(n12376), .A2(n10259), .ZN(n10523) );
  AND2_X2 U11333 ( .A1(n12382), .A2(n10259), .ZN(n10497) );
  NAND2_X2 U11335 ( .A1(n18758), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18705) );
  INV_X2 U11336 ( .A(n16370), .ZN(U215) );
  NAND2_X2 U11337 ( .A1(n18758), .A2(n18643), .ZN(n18701) );
  CLKBUF_X2 U11338 ( .A(n11100), .Z(n11657) );
  NAND2_X2 U11339 ( .A1(n19867), .A2(n19729), .ZN(n19780) );
  AND2_X2 U11340 ( .A1(n12382), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10496) );
  INV_X2 U11341 ( .A(n17988), .ZN(n9611) );
  AND2_X2 U11342 ( .A1(n12383), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10543) );
  AND2_X2 U11343 ( .A1(n11038), .A2(n13185), .ZN(n11446) );
  AND2_X2 U11344 ( .A1(n11044), .A2(n11045), .ZN(n11191) );
  AND2_X2 U11345 ( .A1(n12381), .A2(n10259), .ZN(n10544) );
  NOR2_X1 U11346 ( .A1(n16775), .A2(n18734), .ZN(n9765) );
  OR2_X2 U11347 ( .A1(n18568), .A2(n12406), .ZN(n10169) );
  OR3_X2 U11348 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n12407), .ZN(n17053) );
  INV_X2 U11349 ( .A(n16374), .ZN(n9612) );
  CLKBUF_X1 U11350 ( .A(n20617), .Z(n20701) );
  NOR2_X1 U11351 ( .A1(n11959), .A2(n13524), .ZN(n11961) );
  AND2_X1 U11352 ( .A1(n10171), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13347) );
  AND2_X1 U11353 ( .A1(n11035), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11038) );
  AND2_X1 U11354 ( .A1(n11037), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11045) );
  AND2_X1 U11355 ( .A1(n13018), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11044) );
  NAND4_X1 U11356 ( .A1(n18722), .A2(n18734), .A3(n18741), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17100) );
  AND2_X2 U11357 ( .A1(n13185), .A2(n12999), .ZN(n11115) );
  NAND2_X1 U11358 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18568) );
  INV_X1 U11359 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13018) );
  INV_X1 U11360 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10170) );
  AND2_X1 U11361 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13300) );
  AND2_X1 U11362 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13186) );
  AND2_X2 U11363 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U11364 ( .A1(n10307), .A2(n15359), .ZN(n9756) );
  AOI21_X1 U11365 ( .B1(n10428), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10417), .ZN(n10425) );
  AND2_X2 U11366 ( .A1(n12381), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10537) );
  NAND4_X1 U11368 ( .A1(n9825), .A2(n10426), .A3(n10427), .A4(n10437), .ZN(
        n10436) );
  NAND2_X2 U11369 ( .A1(n14463), .A2(n14462), .ZN(n14461) );
  XNOR2_X2 U11370 ( .A(n12270), .B(n12271), .ZN(n14463) );
  AND2_X2 U11371 ( .A1(n13249), .A2(n11365), .ZN(n13216) );
  NAND2_X2 U11372 ( .A1(n10131), .A2(n10130), .ZN(n12270) );
  AND2_X1 U11373 ( .A1(n12099), .A2(n19023), .ZN(n10482) );
  OR2_X1 U11374 ( .A1(n12099), .A2(n16204), .ZN(n10478) );
  NAND2_X1 U11375 ( .A1(n12099), .A2(n12098), .ZN(n10136) );
  NAND2_X4 U11376 ( .A1(n10457), .A2(n9893), .ZN(n13351) );
  NAND2_X1 U11378 ( .A1(n10436), .A2(n9759), .ZN(n14425) );
  NOR2_X1 U11379 ( .A1(n14458), .A2(n14457), .ZN(n14456) );
  NAND3_X2 U11380 ( .A1(n11161), .A2(n11122), .A3(n15548), .ZN(n12978) );
  AND2_X2 U11381 ( .A1(n11110), .A2(n11109), .ZN(n11161) );
  NOR2_X2 U11382 ( .A1(n15834), .A2(n15833), .ZN(n15832) );
  AND2_X2 U11383 ( .A1(n14494), .A2(n16073), .ZN(n14484) );
  NOR2_X2 U11384 ( .A1(n14493), .A2(n14495), .ZN(n14494) );
  INV_X2 U11385 ( .A(n13369), .ZN(n13541) );
  AND2_X2 U11386 ( .A1(n13936), .A2(n13939), .ZN(n13937) );
  NOR2_X2 U11387 ( .A1(n14070), .A2(n14071), .ZN(n13936) );
  XNOR2_X2 U11388 ( .A(n11267), .B(n11298), .ZN(n14390) );
  AND3_X1 U11389 ( .A1(n14394), .A2(n11298), .A3(n10074), .ZN(n11381) );
  NOR2_X2 U11390 ( .A1(n14032), .A2(n10086), .ZN(n11772) );
  NAND2_X2 U11391 ( .A1(n13915), .A2(n13916), .ZN(n14032) );
  INV_X1 U11392 ( .A(n14386), .ZN(n9619) );
  INV_X1 U11393 ( .A(n9619), .ZN(n9620) );
  NAND2_X2 U11394 ( .A1(n11253), .A2(n12986), .ZN(n12991) );
  AND2_X1 U11395 ( .A1(n11299), .A2(n10076), .ZN(n10074) );
  OR3_X1 U11396 ( .A1(n10635), .A2(n10634), .A3(n10633), .ZN(n10648) );
  NAND2_X1 U11397 ( .A1(n12081), .A2(n19587), .ZN(n12104) );
  AND2_X1 U11398 ( .A1(n19855), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12098) );
  NOR2_X1 U11399 ( .A1(n18548), .A2(n13658), .ZN(n15397) );
  AND2_X1 U11400 ( .A1(n9955), .A2(n12568), .ZN(n17151) );
  NOR2_X1 U11401 ( .A1(n12569), .A2(n9956), .ZN(n9955) );
  AOI21_X1 U11402 ( .B1(n17074), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(n9927), .ZN(n9926) );
  NOR2_X1 U11403 ( .A1(n17005), .A2(n17063), .ZN(n9927) );
  BUF_X1 U11404 ( .A(n11733), .Z(n11713) );
  NAND2_X1 U11406 ( .A1(n10113), .A2(n9941), .ZN(n10407) );
  AOI21_X1 U11407 ( .B1(n10093), .B2(n10373), .A(n12837), .ZN(n10092) );
  NOR2_X1 U11408 ( .A1(n10809), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U11409 ( .A1(n10075), .A2(n14394), .ZN(n11356) );
  INV_X1 U11410 ( .A(n11324), .ZN(n10075) );
  NAND2_X1 U11411 ( .A1(n9847), .A2(n9843), .ZN(n9842) );
  INV_X1 U11412 ( .A(n10064), .ZN(n9844) );
  OAI21_X1 U11413 ( .B1(n9618), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n14209), .ZN(n9845) );
  AND2_X1 U11414 ( .A1(n11836), .A2(n11887), .ZN(n11837) );
  NAND2_X1 U11415 ( .A1(n13416), .A2(n9777), .ZN(n13857) );
  NAND2_X1 U11416 ( .A1(n13874), .A2(n13894), .ZN(n13867) );
  NAND3_X1 U11417 ( .A1(n19976), .A2(n20176), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11816) );
  AND2_X1 U11418 ( .A1(n11787), .A2(n11819), .ZN(n12840) );
  OR2_X1 U11419 ( .A1(n11820), .A2(n11786), .ZN(n11787) );
  INV_X1 U11420 ( .A(n11816), .ZN(n11824) );
  OR2_X1 U11421 ( .A1(n11820), .A2(n11819), .ZN(n12846) );
  AND2_X1 U11422 ( .A1(n9691), .A2(n9997), .ZN(n9996) );
  NAND2_X1 U11423 ( .A1(n12270), .A2(n12272), .ZN(n12273) );
  AND2_X1 U11424 ( .A1(n10142), .A2(n12145), .ZN(n10141) );
  INV_X1 U11425 ( .A(n14469), .ZN(n10128) );
  NAND2_X1 U11426 ( .A1(n9910), .A2(n9909), .ZN(n9908) );
  NAND2_X1 U11427 ( .A1(n10109), .A2(n9628), .ZN(n14981) );
  AND2_X1 U11428 ( .A1(n14788), .A2(n15048), .ZN(n13671) );
  NOR2_X1 U11429 ( .A1(n9641), .A2(n10061), .ZN(n10060) );
  NOR2_X1 U11430 ( .A1(n10671), .A2(n9940), .ZN(n9938) );
  AND2_X1 U11431 ( .A1(n10656), .A2(n10650), .ZN(n10694) );
  NAND2_X1 U11432 ( .A1(n10436), .A2(n10427), .ZN(n10969) );
  XNOR2_X1 U11433 ( .A(n10966), .B(n10964), .ZN(n10968) );
  NAND2_X1 U11434 ( .A1(n10715), .A2(n10712), .ZN(n10730) );
  NAND2_X1 U11435 ( .A1(n10136), .A2(n12105), .ZN(n12107) );
  NAND3_X1 U11436 ( .A1(n18741), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12401) );
  AOI21_X1 U11437 ( .B1(n17276), .B2(n16276), .A(n17662), .ZN(n12517) );
  XNOR2_X1 U11438 ( .A(n12667), .B(n12653), .ZN(n12502) );
  AND2_X1 U11439 ( .A1(n9875), .A2(n17902), .ZN(n9874) );
  NAND2_X1 U11440 ( .A1(n18140), .A2(n18158), .ZN(n12647) );
  OR2_X1 U11441 ( .A1(n14015), .A2(n11170), .ZN(n13881) );
  NAND2_X1 U11442 ( .A1(n14015), .A2(n13895), .ZN(n13880) );
  OR2_X1 U11443 ( .A1(n13045), .A2(n15553), .ZN(n13404) );
  NAND2_X1 U11444 ( .A1(n15553), .A2(n13152), .ZN(n15585) );
  NAND2_X1 U11445 ( .A1(n10218), .A2(n10217), .ZN(n10334) );
  OR2_X1 U11446 ( .A1(n10216), .A2(n10215), .ZN(n10218) );
  NOR2_X1 U11447 ( .A1(n14713), .A2(n14702), .ZN(n14695) );
  AOI21_X1 U11448 ( .B1(n15399), .B2(n15398), .A(n15397), .ZN(n15601) );
  INV_X1 U11449 ( .A(n16269), .ZN(n12534) );
  NAND2_X1 U11450 ( .A1(n17517), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17497) );
  NAND2_X1 U11451 ( .A1(n15512), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15572) );
  NAND2_X1 U11452 ( .A1(n12528), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9875) );
  OAI21_X1 U11453 ( .B1(n12524), .B2(n9877), .A(n17670), .ZN(n12526) );
  NOR2_X1 U11454 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n9878) );
  INV_X1 U11455 ( .A(n18143), .ZN(n15500) );
  NAND2_X1 U11456 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n9959) );
  OR2_X1 U11457 ( .A1(n12556), .A2(n12557), .ZN(n12550) );
  INV_X1 U11458 ( .A(n12576), .ZN(n9928) );
  NAND2_X1 U11459 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n9925) );
  NOR2_X1 U11460 ( .A1(n11035), .A2(n20754), .ZN(n9780) );
  NAND2_X1 U11461 ( .A1(n20146), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11305) );
  NAND2_X1 U11462 ( .A1(n11305), .A2(n11304), .ZN(n11811) );
  NAND2_X1 U11463 ( .A1(n9666), .A2(n13694), .ZN(n10104) );
  NOR2_X1 U11464 ( .A1(n14993), .A2(n10669), .ZN(n10099) );
  NOR2_X1 U11465 ( .A1(n10583), .A2(n10705), .ZN(n9827) );
  AND2_X1 U11466 ( .A1(n18148), .A2(n18153), .ZN(n12635) );
  INV_X1 U11467 ( .A(n11147), .ZN(n11148) );
  NOR2_X1 U11468 ( .A1(n11642), .A2(n10072), .ZN(n10071) );
  INV_X1 U11469 ( .A(n14060), .ZN(n10072) );
  OR2_X1 U11470 ( .A1(n14048), .A2(n14055), .ZN(n11642) );
  OR2_X1 U11471 ( .A1(n14406), .A2(n20754), .ZN(n13801) );
  INV_X1 U11472 ( .A(n13614), .ZN(n10081) );
  NAND2_X1 U11473 ( .A1(n9704), .A2(n10083), .ZN(n10082) );
  NAND2_X1 U11474 ( .A1(n13963), .A2(n15725), .ZN(n10083) );
  INV_X1 U11475 ( .A(n13929), .ZN(n9978) );
  NOR2_X1 U11476 ( .A1(n14049), .A2(n13852), .ZN(n9979) );
  NAND2_X1 U11477 ( .A1(n13955), .A2(n14082), .ZN(n9970) );
  AND2_X1 U11478 ( .A1(n9975), .A2(n9974), .ZN(n9973) );
  INV_X1 U11479 ( .A(n15730), .ZN(n9974) );
  NOR2_X1 U11480 ( .A1(n13509), .A2(n9976), .ZN(n9975) );
  NAND2_X1 U11481 ( .A1(n10067), .A2(n11899), .ZN(n10066) );
  INV_X1 U11482 ( .A(n11894), .ZN(n10067) );
  NAND2_X1 U11483 ( .A1(n11381), .A2(n11380), .ZN(n9789) );
  NOR2_X1 U11484 ( .A1(n13550), .A2(n9962), .ZN(n9961) );
  INV_X1 U11485 ( .A(n13438), .ZN(n9962) );
  NAND2_X1 U11486 ( .A1(n9854), .A2(n9853), .ZN(n11879) );
  OAI21_X1 U11487 ( .B1(n11870), .B2(n20135), .A(n9855), .ZN(n9854) );
  INV_X1 U11488 ( .A(n14345), .ZN(n14328) );
  INV_X1 U11489 ( .A(n11871), .ZN(n9855) );
  OR2_X1 U11490 ( .A1(n11223), .A2(n11222), .ZN(n11865) );
  AND2_X1 U11491 ( .A1(n11202), .A2(n11200), .ZN(n11185) );
  NAND2_X1 U11492 ( .A1(n13054), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11304) );
  OR2_X1 U11493 ( .A1(n11246), .A2(n11037), .ZN(n11303) );
  NOR2_X1 U11494 ( .A1(n11238), .A2(n11237), .ZN(n11239) );
  OR2_X1 U11495 ( .A1(n10216), .A2(n10217), .ZN(n10703) );
  INV_X1 U11496 ( .A(n10363), .ZN(n10097) );
  NOR2_X1 U11497 ( .A1(n13700), .A2(n13698), .ZN(n13704) );
  NAND2_X1 U11498 ( .A1(n13695), .A2(n13712), .ZN(n13681) );
  AND2_X1 U11499 ( .A1(n10737), .A2(n10709), .ZN(n10749) );
  AND2_X1 U11500 ( .A1(n9989), .A2(n10715), .ZN(n10737) );
  NOR2_X1 U11501 ( .A1(n9990), .A2(n10735), .ZN(n9989) );
  NAND2_X1 U11502 ( .A1(n10415), .A2(n10414), .ZN(n10438) );
  INV_X1 U11503 ( .A(n14478), .ZN(n10132) );
  AOI21_X1 U11504 ( .B1(n10432), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n10409), .ZN(n10413) );
  NAND2_X1 U11505 ( .A1(n12069), .A2(n10170), .ZN(n10402) );
  NAND2_X1 U11506 ( .A1(n10140), .A2(n10139), .ZN(n10138) );
  NAND2_X1 U11507 ( .A1(n12294), .A2(n10140), .ZN(n10137) );
  INV_X1 U11508 ( .A(n14457), .ZN(n10139) );
  AND2_X1 U11509 ( .A1(n12134), .A2(n13290), .ZN(n10142) );
  NAND2_X1 U11510 ( .A1(n12393), .A2(n15359), .ZN(n10393) );
  NOR2_X1 U11511 ( .A1(n14888), .A2(n10032), .ZN(n10031) );
  NOR2_X1 U11512 ( .A1(n9734), .A2(n10118), .ZN(n10117) );
  INV_X1 U11513 ( .A(n16136), .ZN(n10118) );
  NOR2_X1 U11514 ( .A1(n14997), .A2(n10037), .ZN(n10036) );
  INV_X1 U11515 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10037) );
  NOR2_X1 U11516 ( .A1(n10535), .A2(n10534), .ZN(n10818) );
  NOR2_X1 U11517 ( .A1(n14807), .A2(n9901), .ZN(n9900) );
  OR2_X1 U11518 ( .A1(n16046), .A2(n10733), .ZN(n13707) );
  INV_X1 U11519 ( .A(n14954), .ZN(n10107) );
  INV_X1 U11520 ( .A(n14491), .ZN(n10122) );
  NAND2_X1 U11521 ( .A1(n10121), .A2(n14874), .ZN(n10120) );
  INV_X1 U11522 ( .A(n14900), .ZN(n10121) );
  INV_X1 U11523 ( .A(n14853), .ZN(n9836) );
  INV_X1 U11524 ( .A(n13238), .ZN(n10062) );
  INV_X1 U11525 ( .A(n13288), .ZN(n10125) );
  AND2_X1 U11526 ( .A1(n13024), .A2(n13011), .ZN(n10047) );
  INV_X1 U11527 ( .A(n14993), .ZN(n10098) );
  INV_X1 U11528 ( .A(n10099), .ZN(n9945) );
  NOR2_X1 U11529 ( .A1(n10099), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9944) );
  NAND2_X1 U11530 ( .A1(n10667), .A2(n13728), .ZN(n10672) );
  INV_X1 U11531 ( .A(n10656), .ZN(n10667) );
  NAND2_X1 U11532 ( .A1(n15304), .A2(n10155), .ZN(n10653) );
  AND2_X1 U11533 ( .A1(n10694), .A2(n15301), .ZN(n10155) );
  INV_X1 U11534 ( .A(n10694), .ZN(n10088) );
  INV_X1 U11535 ( .A(n13473), .ZN(n9897) );
  NAND2_X1 U11536 ( .A1(n10431), .A2(n10430), .ZN(n10966) );
  NAND2_X1 U11537 ( .A1(n9745), .A2(n12894), .ZN(n9742) );
  AND2_X1 U11538 ( .A1(n14510), .A2(n10362), .ZN(n9746) );
  NOR2_X1 U11539 ( .A1(n10716), .A2(n10726), .ZN(n10715) );
  NOR2_X1 U11540 ( .A1(n10832), .A2(n10831), .ZN(n10837) );
  AND2_X1 U11541 ( .A1(n12959), .A2(n12958), .ZN(n10830) );
  INV_X1 U11542 ( .A(n10465), .ZN(n10451) );
  OAI21_X1 U11543 ( .B1(n10370), .B2(n10308), .A(n9756), .ZN(n10309) );
  AND3_X2 U11544 ( .A1(n10303), .A2(n14510), .A3(n10350), .ZN(n10394) );
  NOR2_X1 U11545 ( .A1(n16801), .A2(n16969), .ZN(n9811) );
  OR2_X1 U11546 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15483), .ZN(
        n12441) );
  INV_X1 U11547 ( .A(n12453), .ZN(n9772) );
  NOR2_X1 U11548 ( .A1(n17503), .A2(n17810), .ZN(n10005) );
  INV_X1 U11549 ( .A(n12528), .ZN(n12533) );
  NOR2_X1 U11550 ( .A1(n15605), .A2(n12631), .ZN(n13654) );
  OR2_X1 U11551 ( .A1(n17713), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10021) );
  NAND2_X1 U11552 ( .A1(n17750), .A2(n12503), .ZN(n12505) );
  INV_X1 U11553 ( .A(n16399), .ZN(n13646) );
  NOR2_X1 U11554 ( .A1(n9922), .A2(n9921), .ZN(n12644) );
  INV_X1 U11555 ( .A(n12573), .ZN(n9921) );
  OR2_X1 U11556 ( .A1(n12995), .A2(n13035), .ZN(n13045) );
  NAND2_X1 U11557 ( .A1(n19931), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13276) );
  OAI22_X1 U11558 ( .A1(n12978), .A2(n12982), .B1(n12981), .B2(n13006), .ZN(
        n13151) );
  AND2_X1 U11559 ( .A1(n13030), .A2(n12980), .ZN(n12981) );
  AND2_X1 U11560 ( .A1(n11268), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13808) );
  NAND2_X1 U11561 ( .A1(n9708), .A2(n10085), .ZN(n10084) );
  INV_X1 U11562 ( .A(n10086), .ZN(n10085) );
  NAND2_X1 U11563 ( .A1(n13937), .A2(n14060), .ZN(n14047) );
  INV_X1 U11564 ( .A(n13952), .ZN(n11556) );
  INV_X1 U11565 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11409) );
  AND3_X1 U11566 ( .A1(n9633), .A2(n13216), .A3(n10077), .ZN(n10164) );
  INV_X1 U11567 ( .A(n11366), .ZN(n11367) );
  NAND2_X1 U11568 ( .A1(n13216), .A2(n13252), .ZN(n13446) );
  NAND2_X1 U11569 ( .A1(n10148), .A2(n14161), .ZN(n9840) );
  NOR2_X1 U11570 ( .A1(n14029), .A2(n9980), .ZN(n14015) );
  OR4_X1 U11571 ( .A1(n13912), .A2(n14028), .A3(n9981), .A4(n9983), .ZN(n9980)
         );
  AND2_X1 U11572 ( .A1(n13845), .A2(n13844), .ZN(n14072) );
  AND3_X1 U11573 ( .A1(n13619), .A2(n13857), .A3(n13618), .ZN(n14097) );
  INV_X1 U11574 ( .A(n14254), .ZN(n10068) );
  OR2_X1 U11575 ( .A1(n15832), .A2(n10066), .ZN(n10065) );
  INV_X1 U11576 ( .A(n20127), .ZN(n15948) );
  INV_X1 U11577 ( .A(n13469), .ZN(n9860) );
  INV_X1 U11578 ( .A(n13468), .ZN(n9861) );
  INV_X1 U11579 ( .A(n11888), .ZN(n10069) );
  INV_X1 U11580 ( .A(n15838), .ZN(n9862) );
  INV_X1 U11581 ( .A(n9864), .ZN(n13467) );
  AND2_X1 U11582 ( .A1(n14329), .A2(n14345), .ZN(n14376) );
  NAND2_X1 U11583 ( .A1(n9855), .A2(n11870), .ZN(n10063) );
  INV_X1 U11584 ( .A(n11870), .ZN(n9856) );
  AND2_X1 U11585 ( .A1(n10063), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9857) );
  NAND2_X1 U11586 ( .A1(n13415), .A2(n13894), .ZN(n13879) );
  AND2_X1 U11587 ( .A1(n14410), .A2(n20754), .ZN(n11833) );
  AOI21_X1 U11588 ( .B1(n13043), .B2(n13152), .A(n13042), .ZN(n13058) );
  NAND4_X1 U11589 ( .A1(n13149), .A2(n11171), .A3(n12971), .A4(n13161), .ZN(
        n13053) );
  INV_X1 U11590 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20689) );
  NOR2_X1 U11591 ( .A1(n20310), .A2(n20483), .ZN(n20647) );
  INV_X1 U11592 ( .A(n19976), .ZN(n20146) );
  NAND2_X1 U11593 ( .A1(n9620), .A2(n20141), .ZN(n20540) );
  AOI21_X1 U11594 ( .B1(n20611), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20310), 
        .ZN(n20699) );
  NAND2_X1 U11595 ( .A1(n9818), .A2(n11829), .ZN(n15553) );
  OAI21_X1 U11596 ( .B1(n11827), .B2(n11826), .A(n9676), .ZN(n9818) );
  AND2_X1 U11597 ( .A1(n20753), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15551) );
  INV_X1 U11598 ( .A(n20157), .ZN(n15548) );
  NAND2_X1 U11599 ( .A1(n13541), .A2(n19852), .ZN(n10382) );
  AND2_X1 U11600 ( .A1(n13340), .A2(n13338), .ZN(n13374) );
  AND2_X1 U11601 ( .A1(n10703), .A2(n10699), .ZN(n10332) );
  AND2_X1 U11602 ( .A1(n13731), .A2(n13666), .ZN(n13722) );
  INV_X1 U11603 ( .A(n12019), .ZN(n13709) );
  OR2_X1 U11604 ( .A1(n13682), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n13695) );
  NAND2_X1 U11605 ( .A1(n10804), .A2(n9691), .ZN(n13672) );
  NAND2_X1 U11606 ( .A1(n9986), .A2(n10795), .ZN(n10802) );
  INV_X1 U11607 ( .A(n10798), .ZN(n9986) );
  NAND2_X1 U11608 ( .A1(n10424), .A2(n10425), .ZN(n10427) );
  AND2_X1 U11609 ( .A1(n10167), .A2(n12113), .ZN(n10146) );
  AND2_X1 U11610 ( .A1(n19071), .A2(n19072), .ZN(n12113) );
  NAND2_X1 U11611 ( .A1(n14695), .A2(n9723), .ZN(n14685) );
  NAND2_X1 U11612 ( .A1(n10851), .A2(n10850), .ZN(n12899) );
  AND2_X1 U11613 ( .A1(n12110), .A2(n12109), .ZN(n12111) );
  INV_X1 U11614 ( .A(n10393), .ZN(n10113) );
  AND2_X1 U11615 ( .A1(n11990), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11949) );
  AND2_X1 U11616 ( .A1(n11953), .A2(n10038), .ZN(n11990) );
  AND2_X1 U11617 ( .A1(n9650), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10038) );
  AOI21_X1 U11618 ( .B1(n9907), .B2(n9911), .A(n9905), .ZN(n9904) );
  INV_X1 U11619 ( .A(n15123), .ZN(n9905) );
  AND2_X1 U11620 ( .A1(n11948), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11980) );
  OR2_X1 U11621 ( .A1(n11019), .A2(n11020), .ZN(n14901) );
  AND2_X1 U11622 ( .A1(n11956), .A2(n9711), .ZN(n11972) );
  NOR2_X1 U11623 ( .A1(n16105), .A2(n13242), .ZN(n14970) );
  AND2_X1 U11624 ( .A1(n10116), .A2(n10978), .ZN(n10115) );
  NAND2_X1 U11625 ( .A1(n13485), .A2(n10116), .ZN(n13125) );
  NAND2_X1 U11626 ( .A1(n14777), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14766) );
  NAND2_X1 U11627 ( .A1(n14695), .A2(n10055), .ZN(n14674) );
  AND2_X1 U11628 ( .A1(n14695), .A2(n9732), .ZN(n14520) );
  INV_X1 U11629 ( .A(n14518), .ZN(n10054) );
  AND2_X1 U11630 ( .A1(n9651), .A2(n14455), .ZN(n10126) );
  OR2_X1 U11631 ( .A1(n14454), .A2(n14449), .ZN(n14451) );
  NOR2_X1 U11632 ( .A1(n14732), .A2(n10043), .ZN(n10042) );
  INV_X1 U11633 ( .A(n14740), .ZN(n10043) );
  AND2_X1 U11634 ( .A1(n15111), .A2(n15110), .ZN(n15112) );
  NOR2_X1 U11635 ( .A1(n15169), .A2(n11995), .ZN(n15142) );
  AND2_X1 U11636 ( .A1(n15142), .A2(n15141), .ZN(n15144) );
  NOR2_X1 U11637 ( .A1(n14850), .A2(n9836), .ZN(n9835) );
  INV_X1 U11638 ( .A(n14871), .ZN(n9834) );
  NAND2_X1 U11639 ( .A1(n14853), .A2(n9839), .ZN(n9837) );
  NAND2_X1 U11640 ( .A1(n9725), .A2(n13164), .ZN(n13221) );
  NAND2_X1 U11641 ( .A1(n9937), .A2(n9936), .ZN(n16112) );
  NOR2_X1 U11642 ( .A1(n9939), .A2(n15245), .ZN(n9936) );
  NAND2_X1 U11643 ( .A1(n10671), .A2(n10670), .ZN(n16123) );
  NAND2_X1 U11644 ( .A1(n9946), .A2(n10651), .ZN(n15283) );
  NAND2_X1 U11645 ( .A1(n15283), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15282) );
  NAND2_X1 U11646 ( .A1(n10742), .A2(n10741), .ZN(n15293) );
  NAND2_X1 U11647 ( .A1(n10048), .A2(n9733), .ZN(n13384) );
  NAND2_X1 U11648 ( .A1(n13476), .A2(n13475), .ZN(n9758) );
  AOI21_X1 U11649 ( .B1(n13451), .B2(n9698), .A(n9899), .ZN(n9898) );
  NOR2_X1 U11650 ( .A1(n13523), .A2(n16195), .ZN(n9899) );
  AOI21_X1 U11651 ( .B1(n13351), .B2(n12098), .A(n12091), .ZN(n12923) );
  XNOR2_X1 U11652 ( .A(n12093), .B(n12094), .ZN(n12922) );
  NAND2_X1 U11653 ( .A1(n10251), .A2(n10224), .ZN(n13334) );
  INV_X1 U11654 ( .A(n19593), .ZN(n19285) );
  AND2_X1 U11655 ( .A1(n16749), .A2(n9888), .ZN(n16538) );
  NAND2_X1 U11656 ( .A1(n17495), .A2(n16591), .ZN(n9888) );
  INV_X1 U11657 ( .A(n18782), .ZN(n18769) );
  AND2_X1 U11658 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16983), .ZN(n16960) );
  INV_X2 U11659 ( .A(n12420), .ZN(n17096) );
  OR2_X2 U11660 ( .A1(n18568), .A2(n12404), .ZN(n10165) );
  NAND2_X1 U11661 ( .A1(n17151), .A2(n18148), .ZN(n15604) );
  INV_X1 U11662 ( .A(n17152), .ZN(n17150) );
  NOR2_X1 U11663 ( .A1(n12642), .A2(n9935), .ZN(n9934) );
  OR2_X1 U11664 ( .A1(n18763), .A2(n18148), .ZN(n9935) );
  AOI21_X1 U11665 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n12648), .A(
        n18493), .ZN(n17612) );
  AOI22_X1 U11666 ( .A1(n17670), .A2(n16259), .B1(n17662), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10014) );
  NOR3_X1 U11667 ( .A1(n17662), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n17436), .ZN(n15511) );
  AND2_X1 U11668 ( .A1(n16274), .A2(n10157), .ZN(n15512) );
  NOR2_X1 U11669 ( .A1(n17473), .A2(n10001), .ZN(n17464) );
  NAND2_X1 U11670 ( .A1(n17503), .A2(n9652), .ZN(n10001) );
  NAND2_X1 U11671 ( .A1(n10002), .A2(n10009), .ZN(n17445) );
  OAI21_X1 U11672 ( .B1(n17474), .B2(n10007), .A(n10006), .ZN(n10009) );
  NOR2_X1 U11673 ( .A1(n10005), .A2(n10003), .ZN(n10002) );
  NAND2_X1 U11674 ( .A1(n9685), .A2(n17825), .ZN(n10007) );
  INV_X1 U11675 ( .A(n12527), .ZN(n9876) );
  OAI21_X1 U11676 ( .B1(n12629), .B2(n12628), .A(n13649), .ZN(n18548) );
  NOR3_X1 U11677 ( .A1(n16399), .A2(n17348), .A3(n9952), .ZN(n9951) );
  INV_X1 U11678 ( .A(n12647), .ZN(n9952) );
  NOR2_X1 U11679 ( .A1(n9775), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9774) );
  INV_X1 U11680 ( .A(n12518), .ZN(n9775) );
  AND2_X1 U11681 ( .A1(n17713), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10022) );
  NAND2_X1 U11682 ( .A1(n17714), .A2(n10021), .ZN(n10019) );
  INV_X1 U11683 ( .A(n10022), .ZN(n10018) );
  INV_X1 U11684 ( .A(n17348), .ZN(n18128) );
  OAI211_X1 U11685 ( .C1(n12454), .C2(n16889), .A(n12586), .B(n12585), .ZN(
        n18143) );
  AOI211_X1 U11686 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n12584), .B(n12583), .ZN(n12585) );
  INV_X1 U11687 ( .A(n18617), .ZN(n18771) );
  AND2_X1 U11688 ( .A1(n19931), .A2(n13260), .ZN(n19905) );
  AND2_X1 U11689 ( .A1(n19972), .A2(n13160), .ZN(n15751) );
  INV_X1 U11690 ( .A(n19972), .ZN(n15760) );
  INV_X1 U11691 ( .A(n14026), .ZN(n15623) );
  AND2_X1 U11692 ( .A1(n11775), .A2(n20701), .ZN(n20070) );
  AND2_X1 U11693 ( .A1(n15800), .A2(n20085), .ZN(n20079) );
  INV_X1 U11694 ( .A(n20089), .ZN(n20071) );
  OR2_X1 U11695 ( .A1(n15541), .A2(n15585), .ZN(n20089) );
  INV_X1 U11696 ( .A(n15800), .ZN(n20086) );
  NAND2_X1 U11697 ( .A1(n9963), .A2(n15570), .ZN(n9822) );
  NAND2_X1 U11698 ( .A1(n15562), .A2(n20131), .ZN(n9963) );
  NOR2_X1 U11699 ( .A1(n14275), .A2(n15566), .ZN(n9823) );
  OAI21_X1 U11700 ( .B1(n11910), .B2(n11919), .A(n11909), .ZN(n11914) );
  NAND2_X1 U11701 ( .A1(n15844), .A2(n20131), .ZN(n9792) );
  XNOR2_X1 U11702 ( .A(n9795), .B(n14289), .ZN(n15845) );
  NAND2_X1 U11703 ( .A1(n9797), .A2(n11912), .ZN(n9796) );
  NOR2_X1 U11704 ( .A1(n15847), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9793) );
  INV_X1 U11705 ( .A(n20120), .ZN(n20130) );
  INV_X1 U11706 ( .A(n20116), .ZN(n20131) );
  INV_X1 U11707 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20611) );
  AND2_X1 U11708 ( .A1(n13374), .A2(n19700), .ZN(n19846) );
  INV_X1 U11709 ( .A(n19826), .ZN(n19036) );
  XNOR2_X1 U11710 ( .A(n12392), .B(n12391), .ZN(n14504) );
  AND2_X1 U11711 ( .A1(n19070), .A2(n12900), .ZN(n19081) );
  XNOR2_X1 U11712 ( .A(n14766), .B(n11950), .ZN(n13765) );
  INV_X1 U11713 ( .A(n16161), .ZN(n16142) );
  OR2_X1 U11714 ( .A1(n18792), .A2(n19852), .ZN(n16152) );
  NAND3_X1 U11715 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19806), .A3(n19593), 
        .ZN(n16138) );
  AOI21_X1 U11716 ( .B1(n14762), .B2(n14763), .A(n13730), .ZN(n13737) );
  XNOR2_X1 U11717 ( .A(n14431), .B(n13738), .ZN(n15020) );
  INV_X1 U11718 ( .A(n19164), .ZN(n16209) );
  INV_X1 U11719 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19830) );
  INV_X1 U11720 ( .A(n16792), .ZN(n16776) );
  NOR2_X1 U11721 ( .A1(n18158), .A2(n16873), .ZN(n16885) );
  INV_X1 U11722 ( .A(n17049), .ZN(n17031) );
  INV_X1 U11723 ( .A(n18158), .ZN(n17199) );
  NOR2_X2 U11724 ( .A1(n17146), .A2(n17199), .ZN(n17147) );
  NAND2_X1 U11725 ( .A1(n17194), .A2(n17199), .ZN(n17187) );
  NOR2_X1 U11726 ( .A1(n15604), .A2(n17152), .ZN(n17283) );
  NOR2_X1 U11727 ( .A1(n17682), .A2(n17857), .ZN(n9916) );
  AOI21_X1 U11728 ( .B1(n17605), .B2(n17496), .A(n9919), .ZN(n9918) );
  NOR2_X1 U11729 ( .A1(n17988), .A2(n18685), .ZN(n9919) );
  NAND2_X1 U11730 ( .A1(n17513), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9917) );
  NAND2_X1 U11731 ( .A1(n17501), .A2(n17500), .ZN(n9920) );
  AND2_X1 U11732 ( .A1(n9931), .A2(n9930), .ZN(n9929) );
  NAND2_X1 U11733 ( .A1(n17497), .A2(n17600), .ZN(n9930) );
  OR2_X1 U11734 ( .A1(n17495), .A2(n17771), .ZN(n9931) );
  AND2_X1 U11735 ( .A1(n11811), .A2(n9815), .ZN(n11797) );
  INV_X1 U11736 ( .A(n10151), .ZN(n10093) );
  INV_X1 U11737 ( .A(n10373), .ZN(n10094) );
  NAND2_X1 U11738 ( .A1(n19976), .A2(n20162), .ZN(n12902) );
  CLKBUF_X1 U11739 ( .A(n11657), .Z(n13781) );
  BUF_X1 U11740 ( .A(n11115), .Z(n13776) );
  OR2_X1 U11741 ( .A1(n11377), .A2(n11376), .ZN(n11839) );
  OR2_X1 U11742 ( .A1(n11345), .A2(n11344), .ZN(n11851) );
  OR2_X1 U11743 ( .A1(n11197), .A2(n11196), .ZN(n11859) );
  INV_X1 U11744 ( .A(n11811), .ZN(n11807) );
  INV_X1 U11745 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10144) );
  INV_X1 U11746 ( .A(n12319), .ZN(n10140) );
  AND2_X1 U11747 ( .A1(n10253), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10257) );
  NOR2_X1 U11748 ( .A1(n13541), .A2(n19855), .ZN(n9942) );
  INV_X1 U11749 ( .A(n10674), .ZN(n9940) );
  NAND2_X1 U11750 ( .A1(n10380), .A2(n10395), .ZN(n10381) );
  INV_X1 U11751 ( .A(n10813), .ZN(n10705) );
  AND4_X1 U11752 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10521) );
  NOR2_X1 U11753 ( .A1(n10508), .A2(n9749), .ZN(n10522) );
  AND2_X1 U11754 ( .A1(n10372), .A2(n19171), .ZN(n10303) );
  OAI211_X1 U11755 ( .C1(n17053), .C2(n16862), .A(n9959), .B(n9958), .ZN(n9957) );
  NAND2_X1 U11756 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n9958) );
  AND2_X1 U11757 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12558), .ZN(
        n12552) );
  NOR2_X1 U11758 ( .A1(n12574), .A2(n9924), .ZN(n9923) );
  AND2_X1 U11759 ( .A1(n11945), .A2(n11944), .ZN(n13807) );
  INV_X1 U11760 ( .A(n11924), .ZN(n11925) );
  NAND2_X1 U11761 ( .A1(n11751), .A2(n10087), .ZN(n10086) );
  INV_X1 U11762 ( .A(n14031), .ZN(n10087) );
  AND2_X1 U11763 ( .A1(n10071), .A2(n13927), .ZN(n10070) );
  NAND2_X1 U11764 ( .A1(n11504), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11536) );
  AND2_X1 U11765 ( .A1(n11489), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11504) );
  INV_X1 U11766 ( .A(n14020), .ZN(n9983) );
  AND2_X1 U11767 ( .A1(n11903), .A2(n11902), .ZN(n11904) );
  INV_X1 U11768 ( .A(n13877), .ZN(n13868) );
  AOI21_X1 U11769 ( .B1(n9623), .B2(n10066), .A(n9675), .ZN(n10064) );
  AND2_X1 U11770 ( .A1(n10068), .A2(n11901), .ZN(n9623) );
  OR2_X1 U11771 ( .A1(n15819), .A2(n15945), .ZN(n11901) );
  NOR2_X1 U11772 ( .A1(n9788), .A2(n9640), .ZN(n9787) );
  INV_X1 U11773 ( .A(n11840), .ZN(n11874) );
  NAND2_X1 U11774 ( .A1(n9779), .A2(n9778), .ZN(n9781) );
  NAND2_X1 U11775 ( .A1(n11166), .A2(n9780), .ZN(n9779) );
  INV_X1 U11776 ( .A(n11859), .ZN(n11232) );
  NAND2_X1 U11777 ( .A1(n12901), .A2(n11170), .ZN(n13048) );
  INV_X1 U11778 ( .A(n12901), .ZN(n11795) );
  INV_X1 U11779 ( .A(n11316), .ZN(n9784) );
  INV_X1 U11780 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20429) );
  NOR2_X1 U11781 ( .A1(n11816), .A2(n11868), .ZN(n11818) );
  NAND2_X1 U11782 ( .A1(n20754), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9819) );
  OR2_X1 U11783 ( .A1(n10209), .A2(n10207), .ZN(n10206) );
  AND2_X1 U11784 ( .A1(n9993), .A2(n12054), .ZN(n9992) );
  AND2_X1 U11785 ( .A1(n14466), .A2(n9994), .ZN(n9993) );
  INV_X1 U11786 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n9994) );
  AND2_X1 U11787 ( .A1(n13704), .A2(n12054), .ZN(n13706) );
  INV_X1 U11788 ( .A(n9724), .ZN(n9998) );
  NOR2_X1 U11789 ( .A1(n13677), .A2(n10000), .ZN(n9999) );
  INV_X1 U11790 ( .A(n10803), .ZN(n10000) );
  NAND2_X1 U11791 ( .A1(n13244), .A2(n10763), .ZN(n10774) );
  AND2_X1 U11792 ( .A1(n10749), .A2(n9637), .ZN(n10763) );
  NAND2_X1 U11793 ( .A1(n13712), .A2(n10774), .ZN(n10773) );
  INV_X1 U11794 ( .A(n10368), .ZN(n12393) );
  INV_X1 U11795 ( .A(n14683), .ZN(n10057) );
  OR2_X1 U11796 ( .A1(n10645), .A2(n10644), .ZN(n10849) );
  NOR2_X1 U11797 ( .A1(n10053), .A2(n10052), .ZN(n10049) );
  NAND2_X1 U11798 ( .A1(n13386), .A2(n15307), .ZN(n10052) );
  INV_X1 U11799 ( .A(n10838), .ZN(n10050) );
  NOR2_X1 U11800 ( .A1(n16014), .A2(n10040), .ZN(n10039) );
  INV_X1 U11801 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10040) );
  NAND2_X1 U11802 ( .A1(n10777), .A2(n10776), .ZN(n9912) );
  NOR2_X1 U11803 ( .A1(n14958), .A2(n10029), .ZN(n10028) );
  INV_X1 U11804 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10029) );
  AND2_X1 U11805 ( .A1(n13116), .A2(n13484), .ZN(n10116) );
  OR2_X1 U11806 ( .A1(n13724), .A2(n13725), .ZN(n13732) );
  AND2_X1 U11807 ( .A1(n9723), .A2(n10056), .ZN(n10055) );
  INV_X1 U11808 ( .A(n14672), .ZN(n10056) );
  INV_X1 U11809 ( .A(n14790), .ZN(n10112) );
  OR2_X1 U11810 ( .A1(n15059), .A2(n10103), .ZN(n10102) );
  NAND2_X1 U11811 ( .A1(n10101), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10100) );
  INV_X1 U11812 ( .A(n10102), .ZN(n10101) );
  INV_X1 U11813 ( .A(n14464), .ZN(n10127) );
  AND2_X1 U11814 ( .A1(n16025), .A2(n13728), .ZN(n13713) );
  OR2_X1 U11815 ( .A1(n16035), .A2(n10733), .ZN(n13717) );
  INV_X1 U11816 ( .A(n13702), .ZN(n9903) );
  NAND2_X1 U11817 ( .A1(n10771), .A2(n9697), .ZN(n9829) );
  INV_X1 U11818 ( .A(n10777), .ZN(n9830) );
  NAND2_X1 U11819 ( .A1(n15293), .A2(n15294), .ZN(n10109) );
  INV_X1 U11820 ( .A(n12069), .ZN(n13739) );
  NAND2_X1 U11821 ( .A1(n10505), .A2(n10504), .ZN(n10567) );
  NAND2_X1 U11822 ( .A1(n10362), .A2(n10114), .ZN(n10368) );
  AND2_X1 U11823 ( .A1(n15345), .A2(n10302), .ZN(n10114) );
  NOR2_X1 U11824 ( .A1(n10550), .A2(n10549), .ZN(n10825) );
  NAND2_X1 U11825 ( .A1(n10447), .A2(n9894), .ZN(n9893) );
  INV_X1 U11826 ( .A(n10456), .ZN(n9894) );
  NAND2_X1 U11827 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18749), .ZN(
        n12407) );
  NAND2_X1 U11828 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18734), .ZN(
        n12406) );
  AOI21_X1 U11829 ( .B1(n12417), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n9766), .ZN(n12489) );
  AND2_X1 U11830 ( .A1(n9765), .A2(n9764), .ZN(n9766) );
  NOR2_X1 U11831 ( .A1(n18722), .A2(n17094), .ZN(n9764) );
  NAND2_X1 U11832 ( .A1(n18722), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12404) );
  NAND2_X1 U11833 ( .A1(n15500), .A2(n17151), .ZN(n12642) );
  NOR2_X1 U11834 ( .A1(n18132), .A2(n12647), .ZN(n12641) );
  INV_X1 U11835 ( .A(n17613), .ZN(n9885) );
  AOI21_X1 U11836 ( .B1(n10020), .B2(n10022), .A(n9673), .ZN(n10016) );
  OAI22_X1 U11837 ( .A1(n17474), .A2(n10004), .B1(n17810), .B2(n9652), .ZN(
        n10003) );
  NAND2_X1 U11838 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17825), .ZN(
        n10004) );
  NAND2_X1 U11839 ( .A1(n9685), .A2(n17662), .ZN(n10006) );
  INV_X1 U11840 ( .A(n15604), .ZN(n18584) );
  INV_X1 U11841 ( .A(n18573), .ZN(n13656) );
  NAND2_X1 U11842 ( .A1(n18762), .A2(n13647), .ZN(n17309) );
  NAND2_X1 U11843 ( .A1(n9816), .A2(n9783), .ZN(n12910) );
  AND2_X1 U11844 ( .A1(n12847), .A2(n12846), .ZN(n12979) );
  INV_X1 U11845 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13989) );
  INV_X1 U11846 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14001) );
  NAND2_X1 U11847 ( .A1(n9852), .A2(n9851), .ZN(n9849) );
  NAND2_X1 U11848 ( .A1(n11166), .A2(n9851), .ZN(n9850) );
  AND2_X1 U11849 ( .A1(n13622), .A2(n13621), .ZN(n13974) );
  AND3_X1 U11850 ( .A1(n13418), .A2(n13857), .A3(n13417), .ZN(n13552) );
  NAND2_X1 U11851 ( .A1(n9968), .A2(n9966), .ZN(n13418) );
  NAND2_X1 U11852 ( .A1(n13415), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n9968) );
  INV_X1 U11853 ( .A(n13807), .ZN(n13888) );
  NOR2_X1 U11854 ( .A1(n11726), .A2(n14184), .ZN(n11727) );
  AOI21_X1 U11855 ( .B1(n11707), .B2(n11706), .A(n11705), .ZN(n13916) );
  AND2_X1 U11856 ( .A1(n13804), .A2(n14186), .ZN(n11705) );
  NOR2_X1 U11857 ( .A1(n11684), .A2(n14193), .ZN(n11685) );
  NAND2_X1 U11858 ( .A1(n11685), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11726) );
  NOR2_X1 U11859 ( .A1(n11639), .A2(n11635), .ZN(n11622) );
  NAND2_X1 U11860 ( .A1(n11622), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11684) );
  AND2_X1 U11861 ( .A1(n11607), .A2(n11606), .ZN(n14060) );
  AND2_X1 U11862 ( .A1(n11589), .A2(n11588), .ZN(n13939) );
  NOR2_X1 U11863 ( .A1(n11571), .A2(n14216), .ZN(n11572) );
  NAND2_X1 U11864 ( .A1(n11572), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11604) );
  NOR2_X1 U11865 ( .A1(n11536), .A2(n14230), .ZN(n11537) );
  NAND2_X1 U11866 ( .A1(n11537), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11571) );
  INV_X1 U11867 ( .A(n13951), .ZN(n14081) );
  OR2_X1 U11868 ( .A1(n10081), .A2(n10080), .ZN(n10079) );
  INV_X1 U11869 ( .A(n13634), .ZN(n10080) );
  NOR3_X1 U11870 ( .A1(n13964), .A2(n10082), .A3(n10081), .ZN(n13635) );
  NOR2_X1 U11871 ( .A1(n11472), .A2(n15717), .ZN(n11489) );
  NOR2_X1 U11872 ( .A1(n13964), .A2(n10082), .ZN(n13967) );
  AND2_X1 U11873 ( .A1(n14093), .A2(n14092), .ZN(n14095) );
  NAND2_X1 U11874 ( .A1(n11443), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11472) );
  NAND2_X1 U11875 ( .A1(n11424), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11442) );
  INV_X1 U11876 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11441) );
  AND2_X1 U11877 ( .A1(n11407), .A2(n11406), .ZN(n13436) );
  INV_X1 U11878 ( .A(n11387), .ZN(n11388) );
  NAND2_X1 U11879 ( .A1(n11388), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11410) );
  NAND2_X1 U11880 ( .A1(n11847), .A2(n11501), .ZN(n11383) );
  AND2_X1 U11881 ( .A1(n13217), .A2(n13250), .ZN(n11365) );
  NAND2_X1 U11882 ( .A1(n11348), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11366) );
  INV_X1 U11883 ( .A(n11357), .ZN(n11348) );
  NAND2_X1 U11884 ( .A1(n11358), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11357) );
  NOR3_X1 U11885 ( .A1(n20078), .A2(n14001), .A3(n13989), .ZN(n11358) );
  INV_X1 U11886 ( .A(n13158), .ZN(n11296) );
  INV_X1 U11887 ( .A(n13399), .ZN(n11295) );
  NOR2_X1 U11888 ( .A1(n9982), .A2(n9983), .ZN(n14023) );
  INV_X1 U11889 ( .A(n14021), .ZN(n9982) );
  NOR2_X1 U11890 ( .A1(n9618), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11911) );
  AND2_X1 U11891 ( .A1(n14065), .A2(n9696), .ZN(n14042) );
  INV_X1 U11892 ( .A(n14039), .ZN(n9977) );
  NAND2_X1 U11893 ( .A1(n14065), .A2(n9687), .ZN(n14040) );
  NAND2_X1 U11894 ( .A1(n14065), .A2(n9979), .ZN(n14051) );
  NAND2_X1 U11895 ( .A1(n14065), .A2(n14056), .ZN(n14058) );
  AND2_X1 U11896 ( .A1(n14063), .A2(n14062), .ZN(n14065) );
  NAND2_X1 U11897 ( .A1(n9842), .A2(n11904), .ZN(n15793) );
  OR3_X1 U11898 ( .A1(n9970), .A2(n13638), .A3(n14072), .ZN(n9969) );
  NOR3_X1 U11899 ( .A1(n13639), .A2(n13638), .A3(n9971), .ZN(n14085) );
  NOR2_X1 U11900 ( .A1(n13639), .A2(n13638), .ZN(n14083) );
  OR2_X1 U11901 ( .A1(n13975), .A2(n13627), .ZN(n13639) );
  OR2_X1 U11902 ( .A1(n11900), .A2(n15916), .ZN(n14359) );
  NAND2_X1 U11903 ( .A1(n14359), .A2(n9786), .ZN(n14239) );
  NAND2_X1 U11904 ( .A1(n11900), .A2(n15916), .ZN(n9786) );
  AND2_X1 U11905 ( .A1(n13557), .A2(n9682), .ZN(n14096) );
  INV_X1 U11906 ( .A(n14097), .ZN(n9972) );
  NOR2_X1 U11907 ( .A1(n13058), .A2(n13045), .ZN(n20092) );
  NAND2_X1 U11908 ( .A1(n13557), .A2(n9973), .ZN(n15733) );
  AND3_X1 U11909 ( .A1(n13508), .A2(n13857), .A3(n13507), .ZN(n13509) );
  NAND2_X1 U11910 ( .A1(n13557), .A2(n9975), .ZN(n15731) );
  NAND2_X1 U11911 ( .A1(n10065), .A2(n9623), .ZN(n15818) );
  AND2_X1 U11912 ( .A1(n13600), .A2(n9960), .ZN(n13596) );
  AND2_X1 U11913 ( .A1(n9961), .A2(n9680), .ZN(n9960) );
  AND2_X1 U11914 ( .A1(n15819), .A2(n11898), .ZN(n14255) );
  NOR2_X1 U11915 ( .A1(n11873), .A2(n20125), .ZN(n14378) );
  NAND2_X1 U11916 ( .A1(n13600), .A2(n9961), .ZN(n13594) );
  NAND2_X1 U11917 ( .A1(n13600), .A2(n13438), .ZN(n13549) );
  NOR2_X1 U11918 ( .A1(n20092), .A2(n14378), .ZN(n14343) );
  OR2_X1 U11919 ( .A1(n13553), .A2(n13552), .ZN(n13602) );
  NOR2_X1 U11920 ( .A1(n13602), .A2(n13601), .ZN(n13600) );
  INV_X1 U11921 ( .A(n11299), .ZN(n11267) );
  INV_X1 U11922 ( .A(n11152), .ZN(n11158) );
  OAI22_X2 U11923 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20832), .B1(n15975), 
        .B2(n20853), .ZN(n20197) );
  AND2_X1 U11924 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20529) );
  INV_X1 U11925 ( .A(n20168), .ZN(n20194) );
  NOR2_X1 U11926 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20617) );
  NAND2_X1 U11927 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20197), .ZN(n20168) );
  NAND2_X1 U11928 ( .A1(n13722), .A2(n13723), .ZN(n13724) );
  NAND2_X1 U11929 ( .A1(n13706), .A2(n14466), .ZN(n13708) );
  NAND2_X1 U11930 ( .A1(n11980), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11982) );
  NAND2_X1 U11931 ( .A1(n13681), .A2(n12018), .ZN(n13700) );
  NAND2_X2 U11932 ( .A1(n10756), .A2(n10811), .ZN(n13712) );
  NAND2_X1 U11933 ( .A1(n9987), .A2(n9702), .ZN(n10798) );
  INV_X1 U11934 ( .A(n9987), .ZN(n10790) );
  NAND2_X1 U11935 ( .A1(n10749), .A2(n9665), .ZN(n10750) );
  NAND2_X1 U11936 ( .A1(n9988), .A2(n10715), .ZN(n10736) );
  INV_X1 U11937 ( .A(n9990), .ZN(n9988) );
  INV_X1 U11938 ( .A(n19028), .ZN(n19006) );
  NAND2_X1 U11939 ( .A1(n12221), .A2(n10133), .ZN(n10130) );
  AND2_X1 U11940 ( .A1(n14970), .A2(n9717), .ZN(n14923) );
  INV_X1 U11941 ( .A(n13464), .ZN(n10123) );
  OR2_X1 U11942 ( .A1(n10892), .A2(n10891), .ZN(n19061) );
  NAND2_X1 U11943 ( .A1(n10442), .A2(n10441), .ZN(n10448) );
  NOR2_X1 U11944 ( .A1(n14456), .A2(n12294), .ZN(n12320) );
  NAND2_X1 U11945 ( .A1(n14695), .A2(n14694), .ZN(n14682) );
  NOR2_X1 U11946 ( .A1(n14479), .A2(n14478), .ZN(n14477) );
  NAND2_X1 U11947 ( .A1(n10059), .A2(n9648), .ZN(n15171) );
  INV_X1 U11948 ( .A(n13221), .ZN(n10059) );
  NOR2_X2 U11949 ( .A1(n10811), .A2(n15345), .ZN(n14510) );
  OAI211_X1 U11950 ( .C1(n10818), .C2(n10955), .A(n10834), .B(n10820), .ZN(
        n12959) );
  NOR2_X1 U11951 ( .A1(n14451), .A2(n14437), .ZN(n14439) );
  NAND2_X1 U11952 ( .A1(n11953), .A2(n9650), .ZN(n11989) );
  NAND2_X1 U11953 ( .A1(n11953), .A2(n10039), .ZN(n11987) );
  NAND2_X1 U11954 ( .A1(n11953), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11985) );
  NAND2_X1 U11955 ( .A1(n15112), .A2(n9722), .ZN(n14471) );
  AND2_X1 U11956 ( .A1(n9643), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10030) );
  NAND2_X1 U11957 ( .A1(n11976), .A2(n9643), .ZN(n11979) );
  NAND2_X1 U11958 ( .A1(n11976), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11977) );
  NOR3_X1 U11959 ( .A1(n14901), .A2(n10122), .A3(n14900), .ZN(n14873) );
  NOR2_X1 U11960 ( .A1(n14901), .A2(n14900), .ZN(n14902) );
  NAND2_X1 U11961 ( .A1(n14970), .A2(n9646), .ZN(n14944) );
  NAND2_X1 U11962 ( .A1(n11956), .A2(n10028), .ZN(n11970) );
  INV_X1 U11963 ( .A(n16102), .ZN(n10119) );
  NOR2_X1 U11964 ( .A1(n9626), .A2(n10035), .ZN(n10034) );
  INV_X1 U11965 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10035) );
  NOR2_X1 U11966 ( .A1(n11962), .A2(n9626), .ZN(n11967) );
  NAND2_X1 U11967 ( .A1(n16137), .A2(n10117), .ZN(n16103) );
  NAND2_X1 U11968 ( .A1(n10033), .A2(n10036), .ZN(n11964) );
  NAND2_X1 U11969 ( .A1(n16137), .A2(n16136), .ZN(n16135) );
  INV_X1 U11970 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14997) );
  NOR2_X1 U11971 ( .A1(n11962), .A2(n14997), .ZN(n11965) );
  NOR2_X1 U11972 ( .A1(n13142), .A2(n13141), .ZN(n16137) );
  NAND2_X1 U11973 ( .A1(n10734), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15301) );
  NAND2_X1 U11974 ( .A1(n10160), .A2(n13729), .ZN(n13730) );
  INV_X1 U11975 ( .A(n14773), .ZN(n13729) );
  NAND2_X1 U11976 ( .A1(n9755), .A2(n9754), .ZN(n9753) );
  INV_X1 U11977 ( .A(n10100), .ZN(n9755) );
  AND3_X1 U11978 ( .A1(n15992), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n13728), .ZN(n14773) );
  NAND2_X1 U11979 ( .A1(n9985), .A2(n9984), .ZN(n14788) );
  NOR2_X1 U11980 ( .A1(n13667), .A2(n10733), .ZN(n9984) );
  OR2_X1 U11981 ( .A1(n14839), .A2(n10102), .ZN(n14809) );
  NAND2_X1 U11982 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10103) );
  AND2_X1 U11983 ( .A1(n13717), .A2(n15073), .ZN(n14813) );
  NAND2_X1 U11984 ( .A1(n9902), .A2(n14826), .ZN(n14816) );
  NAND2_X1 U11985 ( .A1(n15144), .A2(n10041), .ZN(n14713) );
  AND2_X1 U11986 ( .A1(n9726), .A2(n14714), .ZN(n10041) );
  NOR2_X1 U11987 ( .A1(n14839), .A2(n14831), .ZN(n14830) );
  NAND2_X1 U11988 ( .A1(n15112), .A2(n14474), .ZN(n14476) );
  NAND2_X1 U11989 ( .A1(n15109), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15108) );
  INV_X1 U11990 ( .A(n14857), .ZN(n10108) );
  NAND2_X1 U11991 ( .A1(n14855), .A2(n10106), .ZN(n10105) );
  AND2_X1 U11992 ( .A1(n13686), .A2(n10107), .ZN(n10106) );
  NOR3_X1 U11993 ( .A1(n14901), .A2(n9689), .A3(n10120), .ZN(n15111) );
  NAND2_X1 U11994 ( .A1(n9832), .A2(n9831), .ZN(n14872) );
  AOI21_X1 U11995 ( .B1(n14851), .B2(n14850), .A(n9836), .ZN(n9831) );
  OR2_X1 U11996 ( .A1(n15171), .A2(n15172), .ZN(n15169) );
  OAI21_X1 U11997 ( .B1(n14852), .B2(n14851), .A(n14850), .ZN(n14898) );
  INV_X1 U11998 ( .A(n10060), .ZN(n10058) );
  NOR2_X1 U11999 ( .A1(n13221), .A2(n13220), .ZN(n13239) );
  NOR2_X1 U12000 ( .A1(n13221), .A2(n9641), .ZN(n15187) );
  NAND2_X1 U12001 ( .A1(n14970), .A2(n14969), .ZN(n14972) );
  NAND2_X1 U12002 ( .A1(n9829), .A2(n10776), .ZN(n14956) );
  NOR2_X1 U12003 ( .A1(n9642), .A2(n10046), .ZN(n10045) );
  NAND2_X1 U12004 ( .A1(n10771), .A2(n10770), .ZN(n14966) );
  OR3_X1 U12005 ( .A1(n18933), .A2(n10733), .A3(n15245), .ZN(n16106) );
  OR2_X1 U12006 ( .A1(n15264), .A2(n14982), .ZN(n16109) );
  AOI21_X1 U12007 ( .B1(n10655), .B2(n9944), .A(n9943), .ZN(n9747) );
  NOR2_X1 U12008 ( .A1(n10098), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9943) );
  NOR2_X1 U12009 ( .A1(n12948), .A2(n10869), .ZN(n13025) );
  NAND2_X1 U12010 ( .A1(n10854), .A2(n10853), .ZN(n12947) );
  NAND2_X1 U12011 ( .A1(n10109), .A2(n10744), .ZN(n16130) );
  AOI21_X1 U12012 ( .B1(n9688), .B2(n9898), .A(n9897), .ZN(n9896) );
  NOR2_X1 U12013 ( .A1(n12928), .A2(n10051), .ZN(n15306) );
  NAND2_X1 U12014 ( .A1(n9733), .A2(n13386), .ZN(n10051) );
  AOI21_X1 U12015 ( .B1(n10969), .B2(n10968), .A(n10967), .ZN(n13485) );
  AND2_X1 U12016 ( .A1(n13485), .A2(n13484), .ZN(n13482) );
  AND2_X1 U12017 ( .A1(n10095), .A2(n10096), .ZN(n10961) );
  NAND2_X1 U12018 ( .A1(n10374), .A2(n10373), .ZN(n10095) );
  AND2_X1 U12019 ( .A1(n10347), .A2(n19700), .ZN(n11026) );
  XNOR2_X1 U12020 ( .A(n10830), .B(n10829), .ZN(n13066) );
  NOR2_X1 U12021 ( .A1(n12928), .A2(n10838), .ZN(n13231) );
  AND2_X1 U12022 ( .A1(n10367), .A2(n10366), .ZN(n13356) );
  INV_X1 U12023 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U12024 ( .A1(n12096), .A2(n12095), .ZN(n12967) );
  NOR2_X1 U12025 ( .A1(n12106), .A2(n10135), .ZN(n10134) );
  INV_X1 U12026 ( .A(n12105), .ZN(n10135) );
  OR3_X1 U12027 ( .A1(n19200), .A2(n19220), .A3(n19843), .ZN(n19203) );
  INV_X1 U12028 ( .A(n19555), .ZN(n19483) );
  NOR2_X2 U12029 ( .A1(n14507), .A2(n16138), .ZN(n19192) );
  NOR2_X2 U12030 ( .A1(n14505), .A2(n16138), .ZN(n19193) );
  INV_X1 U12031 ( .A(n19192), .ZN(n19184) );
  INV_X1 U12032 ( .A(n19193), .ZN(n19186) );
  AND2_X1 U12033 ( .A1(n10334), .A2(n10228), .ZN(n13338) );
  OR2_X1 U12034 ( .A1(n13650), .A2(n17347), .ZN(n9933) );
  NOR3_X1 U12035 ( .A1(n17347), .A2(n16399), .A3(n18571), .ZN(n18550) );
  NAND2_X1 U12036 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16917), .ZN(n16873) );
  NOR2_X1 U12037 ( .A1(n16930), .A2(n9806), .ZN(n9805) );
  INV_X1 U12038 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n9806) );
  NAND3_X1 U12039 ( .A1(n12604), .A2(n12600), .A3(n9810), .ZN(n9809) );
  AOI21_X1 U12040 ( .B1(n17060), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(n9811), .ZN(n9810) );
  INV_X1 U12041 ( .A(n12602), .ZN(n9812) );
  INV_X1 U12042 ( .A(n12601), .ZN(n9813) );
  INV_X1 U12043 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17112) );
  OAI211_X1 U12044 ( .C1(n17038), .C2(n17124), .A(n12484), .B(n12483), .ZN(
        n12656) );
  AOI211_X1 U12045 ( .C1(n17039), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n12429), .B(n12428), .ZN(n12655) );
  NOR2_X1 U12046 ( .A1(n9772), .A2(n9771), .ZN(n9770) );
  NOR2_X1 U12047 ( .A1(n17038), .A2(n17142), .ZN(n9771) );
  NAND2_X1 U12048 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12496) );
  NOR2_X1 U12049 ( .A1(n17345), .A2(n17309), .ZN(n17326) );
  NAND2_X1 U12050 ( .A1(n16246), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9889) );
  INV_X1 U12051 ( .A(n17782), .ZN(n16235) );
  NOR2_X1 U12052 ( .A1(n17763), .A2(n12649), .ZN(n16246) );
  NAND2_X1 U12053 ( .A1(n17446), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17420) );
  AND2_X1 U12054 ( .A1(n17517), .A2(n9880), .ZN(n17446) );
  AND2_X1 U12055 ( .A1(n9644), .A2(n9881), .ZN(n9880) );
  INV_X1 U12056 ( .A(n17459), .ZN(n9881) );
  NAND2_X1 U12057 ( .A1(n17517), .A2(n9644), .ZN(n17458) );
  NOR2_X1 U12058 ( .A1(n17498), .A2(n9883), .ZN(n9882) );
  INV_X1 U12059 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9883) );
  NOR2_X1 U12060 ( .A1(n17531), .A2(n17532), .ZN(n17517) );
  NOR2_X1 U12061 ( .A1(n17565), .A2(n17566), .ZN(n17551) );
  INV_X1 U12062 ( .A(n17923), .ZN(n17847) );
  NAND2_X1 U12063 ( .A1(n9886), .A2(n9884), .ZN(n17565) );
  AND2_X1 U12064 ( .A1(n9632), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9884) );
  AND2_X1 U12065 ( .A1(n9886), .A2(n9632), .ZN(n17589) );
  INV_X1 U12066 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17638) );
  AND2_X1 U12067 ( .A1(n16607), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9887) );
  NOR2_X1 U12068 ( .A1(n17671), .A2(n17685), .ZN(n17673) );
  NOR2_X1 U12069 ( .A1(n17720), .A2(n17719), .ZN(n17699) );
  INV_X1 U12070 ( .A(n16736), .ZN(n17729) );
  NOR2_X1 U12071 ( .A1(n12643), .A2(n12646), .ZN(n13655) );
  NAND2_X1 U12072 ( .A1(n9622), .A2(n17348), .ZN(n17844) );
  AND2_X1 U12073 ( .A1(n9872), .A2(n17502), .ZN(n9871) );
  INV_X1 U12074 ( .A(n10025), .ZN(n17669) );
  NAND2_X1 U12075 ( .A1(n12520), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17975) );
  NAND2_X1 U12076 ( .A1(n17683), .A2(n12518), .ZN(n12520) );
  NAND2_X1 U12077 ( .A1(n15501), .A2(n13652), .ZN(n18555) );
  INV_X1 U12078 ( .A(n12510), .ZN(n12508) );
  INV_X1 U12079 ( .A(n17889), .ZN(n18077) );
  INV_X1 U12080 ( .A(n17844), .ZN(n18549) );
  NOR2_X1 U12081 ( .A1(n17769), .A2(n18725), .ZN(n17768) );
  NAND2_X1 U12082 ( .A1(n9914), .A2(n9664), .ZN(n18567) );
  AND2_X1 U12083 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18569) );
  NAND2_X1 U12084 ( .A1(n18569), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n18563) );
  NAND3_X1 U12085 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15483) );
  AND2_X1 U12086 ( .A1(n13655), .A2(n13656), .ZN(n18571) );
  OAI211_X1 U12087 ( .C1(n17005), .C2(n15456), .A(n12614), .B(n12613), .ZN(
        n18140) );
  AOI211_X1 U12088 ( .C1(n16949), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n12612), .B(n12611), .ZN(n12613) );
  AOI211_X1 U12089 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n12594), .B(n12593), .ZN(n12595) );
  INV_X1 U12090 ( .A(n17151), .ZN(n18153) );
  INV_X1 U12091 ( .A(n18410), .ZN(n18385) );
  OAI22_X1 U12092 ( .A1(n17844), .A2(n18548), .B1(n18547), .B2(n18555), .ZN(
        n18606) );
  OR2_X1 U12093 ( .A1(n15585), .A2(n9782), .ZN(n13078) );
  AND2_X1 U12094 ( .A1(n12873), .A2(n13078), .ZN(n20848) );
  INV_X1 U12095 ( .A(n19910), .ZN(n19941) );
  AND2_X1 U12096 ( .A1(n19931), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19955) );
  NAND2_X1 U12097 ( .A1(n13270), .A2(n13269), .ZN(n19958) );
  INV_X1 U12098 ( .A(n19937), .ZN(n19950) );
  AND2_X1 U12099 ( .A1(n19920), .A2(n13262), .ZN(n19963) );
  XNOR2_X1 U12100 ( .A(n9965), .B(n9964), .ZN(n15562) );
  INV_X1 U12101 ( .A(n13882), .ZN(n9964) );
  NAND2_X1 U12102 ( .A1(n13881), .A2(n13880), .ZN(n9965) );
  OR2_X1 U12103 ( .A1(n13402), .A2(n9777), .ZN(n13403) );
  INV_X1 U12104 ( .A(n14091), .ZN(n14068) );
  INV_X1 U12105 ( .A(n14068), .ZN(n19970) );
  INV_X1 U12106 ( .A(n19965), .ZN(n14098) );
  OR2_X1 U12107 ( .A1(n13813), .A2(n14158), .ZN(n14133) );
  INV_X1 U12108 ( .A(n15756), .ZN(n14151) );
  OR2_X1 U12109 ( .A1(n15751), .A2(n13162), .ZN(n15759) );
  OR2_X1 U12110 ( .A1(n13151), .A2(n13150), .ZN(n13153) );
  INV_X1 U12111 ( .A(n15759), .ZN(n19974) );
  AND2_X1 U12112 ( .A1(n15587), .A2(n15586), .ZN(n20008) );
  BUF_X1 U12113 ( .A(n20022), .Z(n20035) );
  INV_X1 U12114 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14230) );
  OR2_X1 U12115 ( .A1(n20071), .A2(n11830), .ZN(n15800) );
  INV_X1 U12116 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20078) );
  INV_X1 U12117 ( .A(n20070), .ZN(n20149) );
  NAND2_X1 U12118 ( .A1(n9841), .A2(n9840), .ZN(n14165) );
  NAND2_X1 U12119 ( .A1(n14163), .A2(n14162), .ZN(n9841) );
  NOR4_X1 U12120 ( .A1(n15867), .A2(n14269), .A3(n14272), .A4(n15953), .ZN(
        n15863) );
  OAI21_X1 U12121 ( .B1(n15930), .B2(n14272), .A(n20127), .ZN(n9817) );
  AND2_X1 U12122 ( .A1(n10065), .A2(n10068), .ZN(n15827) );
  NAND2_X1 U12123 ( .A1(n9864), .A2(n9703), .ZN(n9863) );
  OR2_X1 U12124 ( .A1(n13058), .A2(n13057), .ZN(n20116) );
  NOR2_X1 U12125 ( .A1(n13467), .A2(n11888), .ZN(n20068) );
  NAND2_X1 U12126 ( .A1(n14376), .A2(n20109), .ZN(n20127) );
  NAND2_X1 U12127 ( .A1(n11872), .A2(n10063), .ZN(n20077) );
  AND2_X1 U12128 ( .A1(n9857), .A2(n11872), .ZN(n20076) );
  INV_X1 U12129 ( .A(n11277), .ZN(n11279) );
  CLKBUF_X1 U12130 ( .A(n14390), .Z(n20139) );
  NOR2_X1 U12131 ( .A1(n20570), .A2(n13006), .ZN(n13016) );
  NOR2_X1 U12132 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14410) );
  INV_X1 U12133 ( .A(n20225), .ZN(n20228) );
  INV_X1 U12134 ( .A(n20275), .ZN(n20301) );
  OAI21_X1 U12135 ( .B1(n10159), .B2(n20311), .A(n20647), .ZN(n20330) );
  INV_X1 U12136 ( .A(n20325), .ZN(n20329) );
  OR2_X1 U12137 ( .A1(n20403), .A2(n20609), .ZN(n20380) );
  AND2_X1 U12138 ( .A1(n20529), .A2(n20363), .ZN(n20422) );
  INV_X1 U12139 ( .A(n20480), .ZN(n20452) );
  OR2_X1 U12140 ( .A1(n20541), .A2(n20609), .ZN(n20520) );
  INV_X1 U12141 ( .A(n20608), .ZN(n20559) );
  OR2_X1 U12142 ( .A1(n20642), .A2(n20565), .ZN(n20602) );
  INV_X1 U12143 ( .A(n20602), .ZN(n20634) );
  INV_X1 U12144 ( .A(n20493), .ZN(n20692) );
  INV_X1 U12145 ( .A(n20577), .ZN(n20706) );
  INV_X1 U12146 ( .A(n20497), .ZN(n20707) );
  INV_X1 U12147 ( .A(n20581), .ZN(n20712) );
  INV_X1 U12148 ( .A(n20501), .ZN(n20713) );
  INV_X1 U12149 ( .A(n20505), .ZN(n20719) );
  INV_X1 U12150 ( .A(n20588), .ZN(n20724) );
  INV_X1 U12151 ( .A(n20509), .ZN(n20725) );
  INV_X1 U12152 ( .A(n20592), .ZN(n20730) );
  INV_X1 U12153 ( .A(n20514), .ZN(n20731) );
  INV_X1 U12154 ( .A(n20518), .ZN(n20737) );
  INV_X1 U12155 ( .A(n20601), .ZN(n20743) );
  INV_X1 U12156 ( .A(n20525), .ZN(n20744) );
  INV_X1 U12157 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20753) );
  NOR2_X1 U12158 ( .A1(n10374), .A2(n19854), .ZN(n19836) );
  INV_X1 U12159 ( .A(n10027), .ZN(n10026) );
  XOR2_X1 U12160 ( .A(n13725), .B(n13724), .Z(n15992) );
  AND2_X1 U12161 ( .A1(n14674), .A2(n14673), .ZN(n16004) );
  OR2_X1 U12162 ( .A1(n13667), .A2(n13722), .ZN(n16013) );
  NAND2_X1 U12163 ( .A1(n18994), .A2(n10166), .ZN(n18875) );
  INV_X1 U12164 ( .A(n19026), .ZN(n18989) );
  NOR2_X1 U12165 ( .A1(n19587), .A2(n19027), .ZN(n18979) );
  INV_X1 U12166 ( .A(n19004), .ZN(n19027) );
  NAND2_X1 U12167 ( .A1(n9761), .A2(n9760), .ZN(n9759) );
  NAND2_X1 U12168 ( .A1(n10426), .A2(n10427), .ZN(n9760) );
  INV_X1 U12169 ( .A(n18979), .ZN(n18850) );
  AND2_X1 U12170 ( .A1(n19846), .A2(n12017), .ZN(n19008) );
  OR2_X1 U12171 ( .A1(n10929), .A2(n10928), .ZN(n13290) );
  INV_X1 U12172 ( .A(n13245), .ZN(n10145) );
  NAND2_X1 U12173 ( .A1(n19073), .A2(n10146), .ZN(n19063) );
  NAND2_X1 U12174 ( .A1(n19073), .A2(n12113), .ZN(n19060) );
  NAND2_X2 U12175 ( .A1(n10448), .A2(n10447), .ZN(n19023) );
  INV_X1 U12176 ( .A(n19081), .ZN(n19075) );
  XNOR2_X1 U12177 ( .A(n13759), .B(n13758), .ZN(n19086) );
  INV_X1 U12178 ( .A(n19101), .ZN(n19085) );
  AND2_X1 U12179 ( .A1(n14509), .A2(n14508), .ZN(n19087) );
  NAND2_X1 U12180 ( .A1(n12897), .A2(n19700), .ZN(n19102) );
  INV_X1 U12181 ( .A(n16085), .ZN(n19096) );
  INV_X1 U12182 ( .A(n16083), .ZN(n19105) );
  INV_X2 U12183 ( .A(n19117), .ZN(n19147) );
  INV_X1 U12184 ( .A(n14793), .ZN(n16005) );
  NAND2_X1 U12185 ( .A1(n9655), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9947) );
  INV_X1 U12186 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16160) );
  NAND2_X1 U12187 ( .A1(n18792), .A2(n12883), .ZN(n16161) );
  INV_X1 U12188 ( .A(n16154), .ZN(n16146) );
  INV_X1 U12189 ( .A(n16152), .ZN(n16145) );
  OR2_X1 U12190 ( .A1(n14520), .A2(n14519), .ZN(n15993) );
  AND2_X1 U12191 ( .A1(n14451), .A2(n14450), .ZN(n16018) );
  NAND2_X1 U12192 ( .A1(n15094), .A2(n13702), .ZN(n14829) );
  AND2_X1 U12193 ( .A1(n15144), .A2(n10042), .ZN(n14720) );
  XNOR2_X1 U12194 ( .A(n9838), .B(n9693), .ZN(n15155) );
  NOR2_X1 U12195 ( .A1(n9835), .A2(n9834), .ZN(n9833) );
  NAND2_X1 U12196 ( .A1(n15282), .A2(n10655), .ZN(n14995) );
  NAND2_X1 U12197 ( .A1(n9758), .A2(n9757), .ZN(n13493) );
  OAI21_X1 U12198 ( .B1(n10714), .B2(n9688), .A(n9898), .ZN(n13474) );
  INV_X1 U12199 ( .A(n16200), .ZN(n19155) );
  NAND2_X1 U12200 ( .A1(n10714), .A2(n13523), .ZN(n13453) );
  INV_X1 U12201 ( .A(n19152), .ZN(n16184) );
  INV_X1 U12202 ( .A(n16189), .ZN(n19162) );
  INV_X1 U12203 ( .A(n19157), .ZN(n16203) );
  NAND2_X1 U12204 ( .A1(n13560), .A2(n12957), .ZN(n19826) );
  INV_X1 U12205 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19821) );
  INV_X1 U12206 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19813) );
  INV_X1 U12207 ( .A(n15366), .ZN(n19807) );
  INV_X1 U12208 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19805) );
  INV_X1 U12209 ( .A(n12093), .ZN(n13560) );
  XNOR2_X1 U12210 ( .A(n12924), .B(n12923), .ZN(n19808) );
  INV_X1 U12211 ( .A(n12922), .ZN(n12924) );
  XNOR2_X1 U12212 ( .A(n12966), .B(n12968), .ZN(n15366) );
  INV_X1 U12213 ( .A(n12967), .ZN(n12968) );
  AND3_X1 U12214 ( .A1(n12900), .A2(n15359), .A3(n10362), .ZN(n9744) );
  NOR2_X1 U12215 ( .A1(n19442), .A2(n19280), .ZN(n19194) );
  OAI21_X1 U12216 ( .B1(n19292), .B2(n19288), .A(n19287), .ZN(n19315) );
  INV_X1 U12217 ( .A(n19355), .ZN(n19330) );
  OR3_X1 U12218 ( .A1(n15369), .A2(n15371), .A3(n19285), .ZN(n19372) );
  NAND2_X1 U12219 ( .A1(n19414), .A2(n19413), .ZN(n19438) );
  NOR2_X1 U12220 ( .A1(n19510), .A2(n19442), .ZN(n19498) );
  NOR2_X1 U12221 ( .A1(n19555), .A2(n19554), .ZN(n19578) );
  INV_X1 U12222 ( .A(n19524), .ZN(n19595) );
  INV_X1 U12223 ( .A(n19654), .ZN(n19601) );
  INV_X1 U12224 ( .A(n19629), .ZN(n19604) );
  INV_X1 U12225 ( .A(n19578), .ZN(n19622) );
  OAI22_X1 U12226 ( .A1(n16299), .A2(n19186), .B1(n18120), .B2(n19184), .ZN(
        n19521) );
  INV_X1 U12227 ( .A(n19530), .ZN(n19630) );
  NOR2_X2 U12228 ( .A1(n19510), .A2(n19554), .ZN(n19645) );
  OAI22_X1 U12229 ( .A1(n18129), .A2(n19184), .B1(n16297), .B2(n19186), .ZN(
        n19654) );
  INV_X1 U12230 ( .A(n19527), .ZN(n19655) );
  INV_X1 U12231 ( .A(n19536), .ZN(n19673) );
  INV_X1 U12232 ( .A(n19542), .ZN(n19685) );
  NOR2_X2 U12233 ( .A1(n19510), .A2(n19796), .ZN(n19693) );
  AND2_X1 U12234 ( .A1(n12023), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19700) );
  INV_X1 U12235 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19587) );
  INV_X1 U12236 ( .A(n9933), .ZN(n16382) );
  NAND2_X1 U12237 ( .A1(n18771), .A2(n18606), .ZN(n16383) );
  NOR2_X1 U12238 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16596), .ZN(n16585) );
  NOR2_X1 U12239 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16658), .ZN(n16657) );
  NOR2_X2 U12240 ( .A1(n18610), .A2(n16405), .ZN(n16770) );
  OAI211_X1 U12241 ( .C1(n16400), .C2(n18613), .A(n16638), .B(n18769), .ZN(
        n16792) );
  NAND2_X1 U12242 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n9799), .ZN(n9798) );
  NOR2_X1 U12243 ( .A1(n9800), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n9799) );
  INV_X1 U12244 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n9800) );
  NAND2_X1 U12245 ( .A1(n16960), .A2(n9654), .ZN(n16901) );
  NOR2_X1 U12246 ( .A1(n16901), .A2(n16902), .ZN(n16917) );
  NAND2_X1 U12247 ( .A1(n16960), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n16944) );
  NOR2_X1 U12248 ( .A1(n16999), .A2(n17016), .ZN(n16983) );
  NAND3_X1 U12249 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n17031), .ZN(n17016) );
  NOR2_X1 U12250 ( .A1(n17067), .A2(n16407), .ZN(n9807) );
  NAND2_X1 U12251 ( .A1(n17117), .A2(n9653), .ZN(n17049) );
  NAND2_X1 U12252 ( .A1(n17117), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n17090) );
  AND2_X1 U12253 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17121), .ZN(n17117) );
  NOR3_X1 U12254 ( .A1(n16707), .A2(n16728), .A3(n17129), .ZN(n17118) );
  AND2_X1 U12255 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17118), .ZN(n17121) );
  INV_X1 U12256 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17128) );
  NAND2_X1 U12257 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17136), .ZN(n17129) );
  NOR2_X1 U12258 ( .A1(n17132), .A2(n17137), .ZN(n17136) );
  AND2_X1 U12259 ( .A1(n17143), .A2(n9803), .ZN(n17138) );
  INV_X1 U12260 ( .A(n16780), .ZN(n9803) );
  NAND2_X1 U12261 ( .A1(n17138), .A2(P3_EBX_REG_2__SCAN_IN), .ZN(n17137) );
  NOR2_X1 U12262 ( .A1(n15601), .A2(n9804), .ZN(n17143) );
  OR3_X1 U12263 ( .A1(n17348), .A2(n18763), .A3(n18617), .ZN(n9804) );
  INV_X1 U12264 ( .A(n17143), .ZN(n17146) );
  NOR2_X1 U12265 ( .A1(n17372), .A2(n17178), .ZN(n17171) );
  NAND2_X1 U12266 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17182), .ZN(n17178) );
  INV_X1 U12267 ( .A(n17187), .ZN(n9950) );
  NOR2_X1 U12268 ( .A1(n17356), .A2(n17222), .ZN(n17217) );
  NOR2_X1 U12269 ( .A1(n17352), .A2(n17226), .ZN(n17227) );
  NAND2_X1 U12270 ( .A1(n17304), .A2(n9954), .ZN(n17270) );
  AND2_X1 U12271 ( .A1(n17153), .A2(n9735), .ZN(n9954) );
  INV_X1 U12272 ( .A(n12656), .ZN(n17279) );
  INV_X1 U12273 ( .A(n17296), .ZN(n17285) );
  INV_X1 U12274 ( .A(n12653), .ZN(n17297) );
  NOR3_X1 U12275 ( .A1(n15601), .A2(n18125), .A3(n18128), .ZN(n15602) );
  INV_X1 U12276 ( .A(n17300), .ZN(n17306) );
  OAI211_X1 U12277 ( .C1(n17348), .C2(n18773), .A(n17347), .B(n17346), .ZN(
        n17379) );
  BUF_X1 U12278 ( .A(n17379), .Z(n17411) );
  NOR2_X1 U12279 ( .A1(n16254), .A2(n16235), .ZN(n16236) );
  NOR2_X1 U12280 ( .A1(n17420), .A2(n17421), .ZN(n16249) );
  NAND2_X1 U12281 ( .A1(n10008), .A2(n17670), .ZN(n17463) );
  INV_X1 U12282 ( .A(n17473), .ZN(n10008) );
  AOI22_X1 U12283 ( .A1(n17607), .A2(n17847), .B1(n17762), .B2(n17845), .ZN(
        n17573) );
  NAND2_X1 U12284 ( .A1(n9886), .A2(n9887), .ZN(n17640) );
  NOR2_X2 U12285 ( .A1(n17276), .A2(n17774), .ZN(n17664) );
  NAND2_X1 U12286 ( .A1(n17276), .A2(n17717), .ZN(n17678) );
  NOR2_X1 U12287 ( .A1(n17348), .A2(n16383), .ZN(n17717) );
  INV_X1 U12288 ( .A(n18456), .ZN(n18493) );
  NOR2_X2 U12289 ( .A1(n18128), .A2(n16383), .ZN(n17762) );
  NAND2_X1 U12290 ( .A1(n17770), .A2(n17728), .ZN(n17765) );
  INV_X1 U12291 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18726) );
  INV_X1 U12292 ( .A(n17762), .ZN(n17775) );
  INV_X1 U12293 ( .A(n17717), .ZN(n17774) );
  OAI21_X1 U12294 ( .B1(n9869), .B2(n9674), .A(n9867), .ZN(n9866) );
  INV_X1 U12295 ( .A(n16266), .ZN(n10011) );
  OAI21_X1 U12296 ( .B1(n17464), .B2(n17670), .A(n9706), .ZN(n9776) );
  NOR2_X2 U12297 ( .A1(n13655), .A2(n18573), .ZN(n18585) );
  NOR2_X1 U12298 ( .A1(n9873), .A2(n12527), .ZN(n17557) );
  INV_X1 U12299 ( .A(n9875), .ZN(n9873) );
  INV_X1 U12300 ( .A(n12526), .ZN(n17561) );
  OAI21_X2 U12301 ( .B1(n15509), .B2(n15508), .A(n18771), .ZN(n18016) );
  OAI211_X1 U12302 ( .C1(n18547), .C2(n15507), .A(n15506), .B(n15505), .ZN(
        n15508) );
  INV_X1 U12303 ( .A(n18089), .ZN(n18092) );
  NAND2_X1 U12304 ( .A1(n10019), .A2(n10018), .ZN(n17697) );
  OR2_X1 U12305 ( .A1(n17714), .A2(n10022), .ZN(n10015) );
  NOR2_X1 U12306 ( .A1(n18555), .A2(n18016), .ZN(n18050) );
  NAND2_X1 U12307 ( .A1(n17714), .A2(n17713), .ZN(n17712) );
  NAND2_X1 U12308 ( .A1(n18549), .A2(n18101), .ZN(n18110) );
  INV_X1 U12309 ( .A(n18016), .ZN(n18101) );
  INV_X1 U12310 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18589) );
  INV_X1 U12311 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18591) );
  INV_X1 U12312 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18596) );
  INV_X2 U12313 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18749) );
  NOR2_X1 U12314 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18743), .ZN(
        n18745) );
  INV_X1 U12315 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18743) );
  NAND2_X1 U12317 ( .A1(n14288), .A2(n20071), .ZN(n11916) );
  OAI21_X1 U12318 ( .B1(n20075), .B2(n15617), .A(n11834), .ZN(n11835) );
  AOI21_X1 U12319 ( .B1(n15564), .B2(n9823), .A(n9822), .ZN(n9821) );
  NAND2_X1 U12320 ( .A1(n15563), .A2(n20130), .ZN(n9820) );
  NOR2_X1 U12321 ( .A1(n9793), .A2(n9791), .ZN(n9790) );
  NAND2_X1 U12322 ( .A1(n15845), .A2(n20130), .ZN(n9794) );
  NAND2_X1 U12323 ( .A1(n15846), .A2(n9792), .ZN(n9791) );
  OAI21_X1 U12324 ( .B1(n15020), .B2(n19084), .A(n12395), .ZN(n12396) );
  AND2_X1 U12325 ( .A1(n10091), .A2(n10090), .ZN(n13752) );
  AOI21_X1 U12326 ( .B1(n16068), .B2(n16157), .A(n13751), .ZN(n10090) );
  OR2_X1 U12327 ( .A1(n13765), .A2(n16154), .ZN(n10091) );
  NOR2_X1 U12328 ( .A1(n15185), .A2(n10686), .ZN(n11034) );
  OR2_X1 U12329 ( .A1(n16446), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9879) );
  OR2_X1 U12330 ( .A1(n16843), .A2(n16844), .ZN(n9802) );
  AOI21_X1 U12331 ( .B1(n17508), .B2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n9916), .ZN(n9915) );
  NAND2_X1 U12332 ( .A1(n10013), .A2(n10010), .ZN(P3_U2831) );
  AOI211_X1 U12333 ( .C1(n16265), .C2(n18097), .A(n10012), .B(n10011), .ZN(
        n10010) );
  NAND2_X1 U12334 ( .A1(n16264), .A2(n18009), .ZN(n10013) );
  NOR2_X1 U12335 ( .A1(n16267), .A2(n18027), .ZN(n10012) );
  AND4_X1 U12336 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_13__SCAN_IN), .A4(P3_EAX_REG_12__SCAN_IN), .ZN(n9621)
         );
  INV_X1 U12337 ( .A(n11133), .ZN(n13192) );
  INV_X1 U12338 ( .A(n13321), .ZN(n13297) );
  NAND2_X1 U12339 ( .A1(n19976), .A2(n9614), .ZN(n9777) );
  AND2_X2 U12340 ( .A1(n17889), .A2(n9932), .ZN(n9622) );
  INV_X1 U12341 ( .A(n10432), .ZN(n10985) );
  OAI21_X1 U12342 ( .B1(n11166), .B2(n9852), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11246) );
  AND2_X1 U12343 ( .A1(n17770), .A2(n9929), .ZN(n9624) );
  NAND2_X1 U12344 ( .A1(n13937), .A2(n10070), .ZN(n9625) );
  NAND2_X1 U12345 ( .A1(n10036), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9626) );
  AND2_X1 U12346 ( .A1(n11150), .A2(n13053), .ZN(n9627) );
  AND2_X1 U12347 ( .A1(n10744), .A2(n9714), .ZN(n9628) );
  INV_X1 U12348 ( .A(n11891), .ZN(n9859) );
  AND2_X1 U12349 ( .A1(n9668), .A2(n12895), .ZN(n9629) );
  INV_X1 U12350 ( .A(n17662), .ZN(n17670) );
  AND2_X1 U12351 ( .A1(n9817), .A2(n14270), .ZN(n9630) );
  AND2_X1 U12352 ( .A1(n9665), .A2(n10988), .ZN(n9631) );
  AND2_X1 U12353 ( .A1(n9887), .A2(n9885), .ZN(n9632) );
  AND2_X2 U12354 ( .A1(n11045), .A2(n12999), .ZN(n11084) );
  AND2_X1 U12355 ( .A1(n12503), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9634) );
  NAND2_X1 U12356 ( .A1(n10429), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n9635) );
  NAND2_X1 U12357 ( .A1(n15838), .A2(n9859), .ZN(n9636) );
  AND2_X1 U12358 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10315) );
  AND2_X1 U12359 ( .A1(n9631), .A2(n19069), .ZN(n9637) );
  AND2_X1 U12360 ( .A1(n10389), .A2(n12895), .ZN(n9638) );
  AND2_X1 U12361 ( .A1(n12895), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n9639) );
  INV_X1 U12362 ( .A(n10870), .ZN(n11999) );
  INV_X1 U12363 ( .A(n11997), .ZN(n13756) );
  AND2_X1 U12364 ( .A1(n11379), .A2(n11378), .ZN(n9640) );
  OR2_X1 U12365 ( .A1(n10062), .A2(n13220), .ZN(n9641) );
  NAND2_X1 U12366 ( .A1(n10047), .A2(n9710), .ZN(n9642) );
  AND2_X1 U12367 ( .A1(n15144), .A2(n9726), .ZN(n14712) );
  AND2_X1 U12368 ( .A1(n10031), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9643) );
  AND2_X1 U12369 ( .A1(n9882), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9644) );
  AND2_X1 U12370 ( .A1(n14969), .A2(n10125), .ZN(n9645) );
  AND2_X1 U12371 ( .A1(n9645), .A2(n10124), .ZN(n9646) );
  AND3_X1 U12372 ( .A1(n9865), .A2(n9862), .A3(n9863), .ZN(n9647) );
  AND2_X1 U12373 ( .A1(n10060), .A2(n10960), .ZN(n9648) );
  OR2_X1 U12374 ( .A1(n12948), .A2(n9642), .ZN(n9649) );
  AND2_X1 U12375 ( .A1(n10039), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9650) );
  NAND2_X1 U12376 ( .A1(n12947), .A2(n12946), .ZN(n12948) );
  INV_X1 U12377 ( .A(n19249), .ZN(n9752) );
  AND2_X1 U12378 ( .A1(n9722), .A2(n10127), .ZN(n9651) );
  OR2_X1 U12379 ( .A1(n10844), .A2(n10843), .ZN(n13230) );
  AND2_X1 U12380 ( .A1(n17803), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9652) );
  AND2_X1 U12381 ( .A1(n9807), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n9653) );
  AND2_X1 U12382 ( .A1(n9805), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n9654) );
  AND2_X1 U12383 ( .A1(n9949), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9655) );
  NOR2_X2 U12384 ( .A1(n12406), .A2(n16775), .ZN(n12405) );
  INV_X1 U12385 ( .A(n18994), .ZN(n19016) );
  AND2_X2 U12386 ( .A1(n12378), .A2(n10259), .ZN(n10529) );
  OR2_X1 U12387 ( .A1(n13639), .A2(n9969), .ZN(n9657) );
  AND2_X1 U12388 ( .A1(n13759), .A2(n12015), .ZN(n9658) );
  NOR2_X1 U12389 ( .A1(n14839), .A2(n10103), .ZN(n9659) );
  AND2_X2 U12390 ( .A1(n10314), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10601) );
  INV_X1 U12391 ( .A(n10372), .ZN(n10358) );
  AND2_X2 U12392 ( .A1(n10300), .A2(n10299), .ZN(n19188) );
  NOR2_X1 U12393 ( .A1(n12404), .A2(n16775), .ZN(n12494) );
  OR2_X1 U12394 ( .A1(n14032), .A2(n14031), .ZN(n9660) );
  AND2_X1 U12395 ( .A1(n13937), .A2(n10071), .ZN(n9661) );
  OR2_X1 U12396 ( .A1(n14029), .A2(n14028), .ZN(n9662) );
  NOR2_X1 U12397 ( .A1(n12407), .A2(n12406), .ZN(n12417) );
  INV_X1 U12398 ( .A(n12417), .ZN(n12430) );
  OR2_X1 U12399 ( .A1(n11889), .A2(n20100), .ZN(n9663) );
  OR2_X1 U12400 ( .A1(n18153), .A2(n15396), .ZN(n9664) );
  NAND2_X1 U12401 ( .A1(n9847), .A2(n10064), .ZN(n14208) );
  AND2_X1 U12402 ( .A1(n10747), .A2(n10745), .ZN(n9665) );
  OAI21_X1 U12403 ( .B1(n10670), .B2(n9940), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n9939) );
  NAND2_X1 U12404 ( .A1(n17683), .A2(n9774), .ZN(n12524) );
  AND3_X1 U12405 ( .A1(n12690), .A2(n12689), .A3(n10156), .ZN(n9667) );
  AND2_X1 U12406 ( .A1(n15338), .A2(n9942), .ZN(n9668) );
  OAI21_X1 U12407 ( .B1(n14191), .B2(n11919), .A(n9618), .ZN(n14300) );
  INV_X1 U12408 ( .A(n14270), .ZN(n20111) );
  INV_X1 U12409 ( .A(n12648), .ZN(n17516) );
  NOR2_X1 U12410 ( .A1(n17771), .A2(n17757), .ZN(n12648) );
  OR3_X1 U12411 ( .A1(n16857), .A2(n9800), .A3(n9801), .ZN(n9669) );
  AND2_X1 U12412 ( .A1(n10401), .A2(n10698), .ZN(n9670) );
  NOR2_X1 U12413 ( .A1(n14827), .A2(n9903), .ZN(n9671) );
  INV_X1 U12414 ( .A(n9948), .ZN(n14950) );
  INV_X1 U12415 ( .A(n9911), .ZN(n9910) );
  NAND2_X1 U12416 ( .A1(n13694), .A2(n9912), .ZN(n9911) );
  AND2_X1 U12417 ( .A1(n11828), .A2(n9819), .ZN(n9672) );
  AND2_X1 U12418 ( .A1(n10613), .A2(n10612), .ZN(n10615) );
  AND2_X1 U12419 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12514), .ZN(
        n9673) );
  NOR2_X1 U12420 ( .A1(n15572), .A2(n16255), .ZN(n9674) );
  NOR2_X1 U12421 ( .A1(n9618), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9675) );
  AND2_X1 U12422 ( .A1(n11825), .A2(n9672), .ZN(n9676) );
  NAND2_X1 U12423 ( .A1(n12895), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10400) );
  INV_X1 U12424 ( .A(n12837), .ZN(n10375) );
  NAND2_X1 U12425 ( .A1(n10439), .A2(n10440), .ZN(n10447) );
  NOR2_X1 U12426 ( .A1(n15832), .A2(n11894), .ZN(n9677) );
  AND3_X1 U12427 ( .A1(n9920), .A2(n9918), .A3(n9917), .ZN(n9678) );
  OR2_X1 U12428 ( .A1(n16857), .A2(n9798), .ZN(n9679) );
  AND2_X1 U12429 ( .A1(n13500), .A2(n13591), .ZN(n9680) );
  NOR2_X1 U12430 ( .A1(n9957), .A2(n12567), .ZN(n9681) );
  INV_X1 U12431 ( .A(n10110), .ZN(n10350) );
  AND2_X1 U12432 ( .A1(n9973), .A2(n9972), .ZN(n9682) );
  AND2_X1 U12433 ( .A1(n11904), .A2(n15894), .ZN(n9683) );
  INV_X1 U12434 ( .A(n11154), .ZN(n13810) );
  INV_X1 U12435 ( .A(n14329), .ZN(n14344) );
  OR2_X1 U12436 ( .A1(n13058), .A2(n15583), .ZN(n14329) );
  INV_X1 U12437 ( .A(n14785), .ZN(n13720) );
  NAND2_X1 U12438 ( .A1(n10648), .A2(n10647), .ZN(n9684) );
  AND2_X1 U12439 ( .A1(n10812), .A2(n10755), .ZN(n10817) );
  NAND2_X1 U12440 ( .A1(n10097), .A2(n10151), .ZN(n10374) );
  INV_X1 U12441 ( .A(n9782), .ZN(n12849) );
  INV_X1 U12442 ( .A(n12065), .ZN(n13741) );
  OR2_X1 U12443 ( .A1(n17670), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9685) );
  INV_X1 U12444 ( .A(n10823), .ZN(n11998) );
  NAND2_X1 U12445 ( .A1(n13289), .A2(n10142), .ZN(n14498) );
  NAND2_X1 U12446 ( .A1(n11956), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11954) );
  NOR2_X1 U12447 ( .A1(n13221), .A2(n10058), .ZN(n9686) );
  INV_X1 U12448 ( .A(n9848), .ZN(n12839) );
  NAND2_X1 U12449 ( .A1(n11161), .A2(n11122), .ZN(n9848) );
  INV_X1 U12450 ( .A(n11355), .ZN(n10076) );
  AND2_X1 U12451 ( .A1(n9979), .A2(n9978), .ZN(n9687) );
  NOR2_X1 U12452 ( .A1(n13451), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9688) );
  NOR2_X1 U12453 ( .A1(n11966), .A2(n14988), .ZN(n11956) );
  NAND2_X1 U12454 ( .A1(n20169), .A2(n19976), .ZN(n13415) );
  OR2_X1 U12455 ( .A1(n10122), .A2(n14487), .ZN(n9689) );
  INV_X1 U12456 ( .A(n10729), .ZN(n9991) );
  AND2_X1 U12457 ( .A1(n15112), .A2(n9651), .ZN(n9690) );
  AND2_X1 U12458 ( .A1(n9999), .A2(n9998), .ZN(n9691) );
  INV_X1 U12459 ( .A(n10776), .ZN(n9909) );
  OR3_X1 U12460 ( .A1(n13639), .A2(n9970), .A3(n13638), .ZN(n9692) );
  NAND2_X1 U12461 ( .A1(n10044), .A2(n10047), .ZN(n13023) );
  AND2_X1 U12462 ( .A1(n14870), .A2(n14869), .ZN(n9693) );
  INV_X1 U12463 ( .A(n14826), .ZN(n9901) );
  INV_X1 U12464 ( .A(n11796), .ZN(n9815) );
  OR2_X1 U12465 ( .A1(n13964), .A2(n13963), .ZN(n9694) );
  AOI21_X1 U12466 ( .B1(n11838), .B2(n11501), .A(n11391), .ZN(n13447) );
  INV_X1 U12467 ( .A(n13447), .ZN(n10077) );
  NAND2_X1 U12468 ( .A1(n11963), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11962) );
  INV_X1 U12469 ( .A(n11380), .ZN(n9788) );
  OR3_X1 U12470 ( .A1(n14901), .A2(n10120), .A3(n10122), .ZN(n9695) );
  NAND2_X1 U12471 ( .A1(n15144), .A2(n14740), .ZN(n14731) );
  AND2_X1 U12472 ( .A1(n9687), .A2(n9977), .ZN(n9696) );
  AND2_X1 U12473 ( .A1(n10770), .A2(n9830), .ZN(n9697) );
  NAND2_X1 U12474 ( .A1(n13523), .A2(n16195), .ZN(n9698) );
  NOR2_X1 U12475 ( .A1(n20068), .A2(n20067), .ZN(n9699) );
  NAND2_X1 U12476 ( .A1(n17662), .A2(n17572), .ZN(n9700) );
  AND2_X1 U12477 ( .A1(n16960), .A2(n9805), .ZN(n9701) );
  NAND2_X1 U12478 ( .A1(n19180), .A2(n10789), .ZN(n9702) );
  AND2_X1 U12479 ( .A1(n10069), .A2(n9663), .ZN(n9703) );
  AND2_X1 U12480 ( .A1(n13969), .A2(n14092), .ZN(n9704) );
  NOR2_X1 U12481 ( .A1(n14477), .A2(n12221), .ZN(n9705) );
  INV_X1 U12482 ( .A(n14851), .ZN(n9839) );
  INV_X1 U12483 ( .A(n13436), .ZN(n11408) );
  INV_X1 U12484 ( .A(n13230), .ZN(n10053) );
  INV_X1 U12485 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20754) );
  NAND2_X1 U12486 ( .A1(n10749), .A2(n9631), .ZN(n9995) );
  NAND2_X1 U12487 ( .A1(n17662), .A2(n17780), .ZN(n9706) );
  NAND2_X1 U12488 ( .A1(n11165), .A2(n11240), .ZN(n9707) );
  AND2_X1 U12489 ( .A1(n10162), .A2(n11773), .ZN(n9708) );
  AND2_X1 U12490 ( .A1(n13289), .A2(n13290), .ZN(n9709) );
  NOR2_X1 U12491 ( .A1(n9656), .A2(n14079), .ZN(n13951) );
  AND2_X1 U12492 ( .A1(n13026), .A2(n13074), .ZN(n9710) );
  AND2_X1 U12493 ( .A1(n10028), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9711) );
  AND2_X1 U12494 ( .A1(n10117), .A2(n10119), .ZN(n9712) );
  AND2_X1 U12495 ( .A1(n9758), .A2(n10582), .ZN(n9713) );
  AND2_X1 U12496 ( .A1(n16132), .A2(n16127), .ZN(n9714) );
  AND2_X1 U12497 ( .A1(n10070), .A2(n14043), .ZN(n9715) );
  AND2_X1 U12498 ( .A1(n10146), .A2(n10145), .ZN(n9716) );
  AND2_X1 U12499 ( .A1(n9646), .A2(n10123), .ZN(n9717) );
  AND2_X1 U12500 ( .A1(n10050), .A2(n10049), .ZN(n9718) );
  AND2_X1 U12501 ( .A1(n11668), .A2(n11667), .ZN(n13927) );
  NAND2_X1 U12502 ( .A1(n20067), .A2(n9663), .ZN(n9865) );
  NOR2_X1 U12504 ( .A1(n18781), .A2(n13658), .ZN(n18581) );
  INV_X1 U12505 ( .A(n18581), .ZN(n9932) );
  NOR2_X1 U12506 ( .A1(n20428), .A2(n20143), .ZN(n9719) );
  AND2_X1 U12507 ( .A1(n14970), .A2(n9645), .ZN(n9720) );
  AND2_X1 U12508 ( .A1(n13557), .A2(n15939), .ZN(n9721) );
  INV_X1 U12509 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11036) );
  AND2_X1 U12510 ( .A1(n10128), .A2(n14474), .ZN(n9722) );
  NAND2_X1 U12511 ( .A1(n9856), .A2(n11871), .ZN(n11872) );
  INV_X1 U12512 ( .A(n14943), .ZN(n10124) );
  AND2_X1 U12513 ( .A1(n10057), .A2(n14694), .ZN(n9723) );
  AND2_X1 U12514 ( .A1(n19180), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n9724) );
  AND2_X1 U12515 ( .A1(n10044), .A2(n10045), .ZN(n9725) );
  AND2_X1 U12516 ( .A1(n10042), .A2(n14721), .ZN(n9726) );
  INV_X2 U12517 ( .A(n10809), .ZN(n19852) );
  BUF_X4 U12518 ( .A(n10809), .Z(n15338) );
  NAND2_X1 U12519 ( .A1(n10015), .A2(n10020), .ZN(n17696) );
  NAND2_X1 U12520 ( .A1(n19073), .A2(n19072), .ZN(n9727) );
  AND2_X1 U12521 ( .A1(n17117), .A2(n9807), .ZN(n9728) );
  AND2_X1 U12522 ( .A1(n12292), .A2(n12317), .ZN(n9729) );
  NAND2_X1 U12523 ( .A1(n13228), .A2(n12111), .ZN(n13391) );
  AND2_X1 U12524 ( .A1(n11976), .A2(n10031), .ZN(n9730) );
  AND2_X1 U12525 ( .A1(n10133), .A2(n10132), .ZN(n9731) );
  AND2_X1 U12526 ( .A1(n10055), .A2(n10054), .ZN(n9732) );
  AND2_X1 U12527 ( .A1(n10050), .A2(n13230), .ZN(n9733) );
  INV_X1 U12528 ( .A(n13146), .ZN(n10046) );
  INV_X1 U12529 ( .A(n15186), .ZN(n10061) );
  AND2_X1 U12530 ( .A1(n10991), .A2(n10990), .ZN(n9734) );
  AND2_X1 U12531 ( .A1(n13506), .A2(n13505), .ZN(n15939) );
  INV_X1 U12532 ( .A(n15939), .ZN(n9976) );
  INV_X1 U12533 ( .A(n11170), .ZN(n13894) );
  AND2_X1 U12534 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .ZN(n9735) );
  NAND2_X1 U12535 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n9736) );
  INV_X1 U12536 ( .A(n17671), .ZN(n9886) );
  AND2_X1 U12537 ( .A1(n17517), .A2(n9882), .ZN(n9737) );
  OR2_X1 U12538 ( .A1(n18770), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n9738) );
  AND2_X1 U12539 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .ZN(n9739) );
  INV_X1 U12540 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n9997) );
  INV_X1 U12541 ( .A(n15026), .ZN(n9754) );
  INV_X1 U12542 ( .A(n13748), .ZN(n9949) );
  INV_X1 U12543 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n9967) );
  INV_X1 U12544 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10032) );
  INV_X1 U12545 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n9801) );
  OR2_X1 U12546 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9740) );
  AND2_X1 U12547 ( .A1(n14289), .A2(n14290), .ZN(n9741) );
  NAND2_X1 U12548 ( .A1(n17503), .A2(n17803), .ZN(n17480) );
  AOI22_X2 U12549 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20148), .B1(DATAI_29_), 
        .B2(n20199), .ZN(n20672) );
  NOR3_X2 U12550 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19830), .A3(
        n19517), .ZN(n19484) );
  NOR3_X2 U12551 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18124), .A3(n18743), 
        .ZN(n18159) );
  OR2_X1 U12552 ( .A1(n19791), .A2(n19826), .ZN(n19510) );
  OR2_X1 U12553 ( .A1(n19791), .A2(n19036), .ZN(n19555) );
  NAND2_X1 U12554 ( .A1(n19791), .A2(n19826), .ZN(n19280) );
  AOI22_X2 U12555 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20148), .B1(DATAI_25_), 
        .B2(n20199), .ZN(n20656) );
  NOR2_X2 U12556 ( .A1(n19189), .A2(n13541), .ZN(n19586) );
  OR2_X1 U12557 ( .A1(n13562), .A2(n13540), .ZN(n19189) );
  NAND2_X1 U12558 ( .A1(n10391), .A2(n16215), .ZN(n11022) );
  AND2_X2 U12559 ( .A1(n9742), .A2(n15492), .ZN(n10391) );
  NAND2_X2 U12560 ( .A1(n9743), .A2(n9744), .ZN(n15492) );
  NAND4_X1 U12561 ( .A1(n9946), .A2(n10655), .A3(n10651), .A4(n9945), .ZN(
        n9748) );
  INV_X1 U12562 ( .A(n10671), .ZN(n16125) );
  NAND2_X1 U12563 ( .A1(n9750), .A2(n10506), .ZN(n9749) );
  OAI21_X1 U12564 ( .B1(n13534), .B2(n19658), .A(n10809), .ZN(n9751) );
  NOR2_X2 U12565 ( .A1(n14839), .A2(n9753), .ZN(n14777) );
  OR2_X1 U12566 ( .A1(n13476), .A2(n13475), .ZN(n9757) );
  INV_X1 U12567 ( .A(n16095), .ZN(n16096) );
  NOR2_X2 U12568 ( .A1(n14867), .A2(n14860), .ZN(n15109) );
  NAND2_X1 U12569 ( .A1(n14837), .A2(n15129), .ZN(n14867) );
  NAND2_X1 U12570 ( .A1(n9825), .A2(n10437), .ZN(n9761) );
  NAND2_X1 U12571 ( .A1(n17730), .A2(n9762), .ZN(n18062) );
  OR2_X1 U12572 ( .A1(n9763), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9762) );
  NAND2_X1 U12573 ( .A1(n9768), .A2(n18065), .ZN(n9767) );
  INV_X1 U12574 ( .A(n12503), .ZN(n9768) );
  NAND2_X1 U12575 ( .A1(n17750), .A2(n9634), .ZN(n9769) );
  NAND2_X1 U12576 ( .A1(n17768), .A2(n17760), .ZN(n17759) );
  XNOR2_X1 U12577 ( .A(n12667), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17760) );
  NOR3_X2 U12578 ( .A1(n9773), .A2(n12499), .A3(n12498), .ZN(n17769) );
  INV_X1 U12579 ( .A(n12493), .ZN(n9773) );
  OR2_X2 U12580 ( .A1(n17444), .A2(n9776), .ZN(n16269) );
  NOR2_X2 U12581 ( .A1(n17445), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17444) );
  OR2_X4 U12582 ( .A1(n11121), .A2(n11120), .ZN(n19976) );
  NOR2_X2 U12583 ( .A1(n19976), .A2(n9614), .ZN(n11171) );
  NAND2_X2 U12584 ( .A1(n15548), .A2(n19976), .ZN(n11172) );
  NOR2_X1 U12585 ( .A1(n11795), .A2(n19976), .ZN(n11122) );
  XNOR2_X2 U12586 ( .A(n9781), .B(n11241), .ZN(n20267) );
  NAND2_X1 U12587 ( .A1(n11166), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11241) );
  NAND3_X1 U12588 ( .A1(n9816), .A2(n11154), .A3(n9783), .ZN(n9782) );
  NOR2_X2 U12589 ( .A1(n14237), .A2(n9785), .ZN(n14356) );
  NAND2_X1 U12590 ( .A1(n9789), .A2(n9640), .ZN(n11847) );
  NAND2_X1 U12591 ( .A1(n9794), .A2(n9790), .ZN(P1_U3004) );
  NAND2_X1 U12592 ( .A1(n14172), .A2(n9796), .ZN(n9795) );
  INV_X1 U12593 ( .A(n14173), .ZN(n9797) );
  NOR2_X1 U12594 ( .A1(n16857), .A2(n9801), .ZN(n16851) );
  INV_X1 U12595 ( .A(n16857), .ZN(n16847) );
  NAND3_X1 U12596 ( .A1(n9802), .A2(n16842), .A3(n9679), .ZN(P3_U2677) );
  NAND4_X2 U12597 ( .A1(n18741), .A2(n18734), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n17005) );
  NOR3_X1 U12598 ( .A1(n9813), .A2(n9812), .A3(n9809), .ZN(n9808) );
  INV_X1 U12599 ( .A(n12603), .ZN(n9814) );
  NAND3_X1 U12600 ( .A1(n15569), .A2(n9821), .A3(n9820), .ZN(P1_U3000) );
  NAND3_X1 U12601 ( .A1(n10390), .A2(n12893), .A3(n10389), .ZN(n13345) );
  NAND3_X1 U12602 ( .A1(n10390), .A2(n12893), .A3(n9638), .ZN(n11023) );
  INV_X1 U12603 ( .A(n10415), .ZN(n9824) );
  NAND3_X1 U12604 ( .A1(n10438), .A2(n10440), .A3(n10439), .ZN(n9825) );
  NAND2_X1 U12605 ( .A1(n9827), .A2(n10615), .ZN(n10649) );
  NAND2_X1 U12606 ( .A1(n9827), .A2(n9826), .ZN(n10656) );
  NOR2_X1 U12607 ( .A1(n9609), .A2(n9684), .ZN(n9826) );
  NOR2_X1 U12608 ( .A1(n10583), .A2(n10705), .ZN(n10616) );
  NAND2_X1 U12609 ( .A1(n9829), .A2(n9828), .ZN(n10780) );
  NAND2_X1 U12610 ( .A1(n14852), .A2(n14850), .ZN(n9832) );
  OAI21_X1 U12611 ( .B1(n14852), .B2(n9837), .A(n9833), .ZN(n9838) );
  NAND2_X1 U12612 ( .A1(n14300), .A2(n13818), .ZN(n14173) );
  NAND2_X1 U12613 ( .A1(n15832), .A2(n9623), .ZN(n9847) );
  AOI21_X2 U12614 ( .B1(n14223), .B2(n14338), .A(n9846), .ZN(n14209) );
  NAND3_X1 U12615 ( .A1(n9850), .A2(n11168), .A3(n9849), .ZN(n11202) );
  NOR2_X1 U12616 ( .A1(n13018), .A2(n20754), .ZN(n9851) );
  XNOR2_X2 U12617 ( .A(n11202), .B(n11201), .ZN(n11289) );
  NAND2_X2 U12618 ( .A1(n11151), .A2(n9627), .ZN(n11166) );
  NAND2_X1 U12619 ( .A1(n11870), .A2(n20135), .ZN(n9853) );
  NAND3_X1 U12620 ( .A1(n9703), .A2(n9864), .A3(n9859), .ZN(n9858) );
  NAND2_X1 U12621 ( .A1(n9863), .A2(n9865), .ZN(n15839) );
  NAND2_X1 U12622 ( .A1(n9868), .A2(n12537), .ZN(n9867) );
  NAND2_X1 U12623 ( .A1(n12536), .A2(n9870), .ZN(n9868) );
  NAND2_X1 U12624 ( .A1(n9870), .A2(n10014), .ZN(n9869) );
  NAND2_X1 U12625 ( .A1(n15571), .A2(n17670), .ZN(n9870) );
  NAND2_X1 U12626 ( .A1(n12527), .A2(n17670), .ZN(n9872) );
  NAND3_X1 U12627 ( .A1(n12525), .A2(n9878), .A3(n17910), .ZN(n9877) );
  NAND3_X1 U12628 ( .A1(n16438), .A2(n16437), .A3(n9879), .ZN(P3_U2641) );
  XNOR2_X2 U12629 ( .A(n9889), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16749) );
  AND2_X1 U12630 ( .A1(n9639), .A2(n9668), .ZN(n9941) );
  NAND2_X1 U12631 ( .A1(n14981), .A2(n10766), .ZN(n10771) );
  NOR2_X2 U12632 ( .A1(n14775), .A2(n14774), .ZN(n14762) );
  AOI21_X1 U12633 ( .B1(n13721), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14785), .ZN(n9890) );
  OAI21_X1 U12634 ( .B1(n13721), .B2(n9740), .A(n10112), .ZN(n9891) );
  NAND2_X1 U12635 ( .A1(n9895), .A2(n9896), .ZN(n10732) );
  NAND2_X1 U12636 ( .A1(n10714), .A2(n9898), .ZN(n9895) );
  NAND2_X1 U12637 ( .A1(n14966), .A2(n9907), .ZN(n9906) );
  AND2_X1 U12638 ( .A1(n10104), .A2(n15122), .ZN(n9913) );
  OAI21_X2 U12639 ( .B1(n18573), .B2(n15396), .A(n9914), .ZN(n18583) );
  OAI21_X2 U12640 ( .B1(n18567), .B2(n18148), .A(n13646), .ZN(n18573) );
  NAND3_X1 U12641 ( .A1(n9678), .A2(n17499), .A3(n9915), .ZN(P3_U2808) );
  NAND3_X1 U12642 ( .A1(n12571), .A2(n12572), .A3(n9923), .ZN(n9922) );
  NAND4_X1 U12643 ( .A1(n9928), .A2(n9926), .A3(n12575), .A4(n9925), .ZN(n9924) );
  NAND2_X2 U12644 ( .A1(n16383), .A2(n9738), .ZN(n17770) );
  NOR2_X1 U12645 ( .A1(n9938), .A2(n9939), .ZN(n16113) );
  INV_X1 U12646 ( .A(n9938), .ZN(n9937) );
  NAND2_X4 U12647 ( .A1(n10113), .A2(n9629), .ZN(n12069) );
  NAND2_X2 U12648 ( .A1(n15338), .A2(n13369), .ZN(n10808) );
  OR2_X1 U12649 ( .A1(n15234), .A2(n10675), .ZN(n9948) );
  NOR2_X2 U12650 ( .A1(n17188), .A2(n17368), .ZN(n17182) );
  INV_X2 U12651 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18741) );
  INV_X2 U12652 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18734) );
  NOR2_X2 U12653 ( .A1(n17270), .A2(n9953), .ZN(n17245) );
  NAND3_X1 U12654 ( .A1(n9621), .A2(P3_EAX_REG_11__SCAN_IN), .A3(n9739), .ZN(
        n9953) );
  NAND4_X1 U12655 ( .A1(n12565), .A2(n12566), .A3(n12564), .A4(n9681), .ZN(
        n9956) );
  AND2_X4 U12656 ( .A1(n11044), .A2(n13186), .ZN(n11128) );
  NAND2_X1 U12657 ( .A1(n13877), .A2(n9967), .ZN(n9966) );
  INV_X1 U12658 ( .A(n14082), .ZN(n9971) );
  NOR3_X1 U12659 ( .A1(n14029), .A2(n13912), .A3(n14028), .ZN(n14021) );
  INV_X1 U12660 ( .A(n14017), .ZN(n9981) );
  NOR2_X2 U12661 ( .A1(n10808), .A2(n19855), .ZN(n10395) );
  INV_X1 U12662 ( .A(n13722), .ZN(n9985) );
  NOR2_X2 U12663 ( .A1(n10782), .A2(n10781), .ZN(n9987) );
  NAND2_X1 U12664 ( .A1(n9991), .A2(n10712), .ZN(n9990) );
  NAND2_X1 U12665 ( .A1(n13704), .A2(n9992), .ZN(n12019) );
  AND2_X1 U12666 ( .A1(n10749), .A2(n10747), .ZN(n10756) );
  INV_X1 U12667 ( .A(n9995), .ZN(n10762) );
  AND2_X1 U12668 ( .A1(n10804), .A2(n9999), .ZN(n13676) );
  NAND2_X1 U12669 ( .A1(n10804), .A2(n9996), .ZN(n13682) );
  NAND2_X1 U12670 ( .A1(n10804), .A2(n10803), .ZN(n13679) );
  NAND2_X1 U12671 ( .A1(n17714), .A2(n10020), .ZN(n10017) );
  INV_X1 U12672 ( .A(n18028), .ZN(n10023) );
  NAND2_X1 U12673 ( .A1(n10023), .A2(n17662), .ZN(n10025) );
  INV_X1 U12674 ( .A(n17579), .ZN(n12523) );
  NAND2_X1 U12675 ( .A1(n10024), .A2(n10025), .ZN(n17579) );
  NOR2_X1 U12676 ( .A1(n12521), .A2(n9736), .ZN(n10024) );
  NOR2_X1 U12677 ( .A1(n17669), .A2(n12521), .ZN(n17609) );
  NAND2_X2 U12678 ( .A1(n18749), .A2(n18741), .ZN(n16775) );
  NAND2_X1 U12679 ( .A1(n11991), .A2(n10026), .ZN(n12080) );
  NAND2_X1 U12680 ( .A1(n15996), .A2(n18994), .ZN(n15982) );
  AND2_X2 U12681 ( .A1(n11976), .A2(n10030), .ZN(n11978) );
  INV_X1 U12682 ( .A(n11962), .ZN(n10033) );
  NAND2_X1 U12683 ( .A1(n10033), .A2(n10034), .ZN(n11966) );
  INV_X1 U12684 ( .A(n12948), .ZN(n10044) );
  INV_X1 U12685 ( .A(n12928), .ZN(n10048) );
  NAND2_X1 U12686 ( .A1(n9718), .A2(n10048), .ZN(n10851) );
  AND2_X2 U12687 ( .A1(n13937), .A2(n9715), .ZN(n13915) );
  INV_X1 U12688 ( .A(n14043), .ZN(n10073) );
  NAND2_X1 U12689 ( .A1(n11298), .A2(n11299), .ZN(n11324) );
  NAND4_X1 U12690 ( .A1(n9633), .A2(n10077), .A3(n13442), .A4(n13216), .ZN(
        n13441) );
  NAND3_X1 U12691 ( .A1(n10077), .A2(n13216), .A3(n13252), .ZN(n10078) );
  INV_X1 U12692 ( .A(n10078), .ZN(n13435) );
  AND2_X2 U12693 ( .A1(n11772), .A2(n11773), .ZN(n13885) );
  NAND2_X1 U12694 ( .A1(n10089), .A2(n10088), .ZN(n10651) );
  INV_X1 U12695 ( .A(n15304), .ZN(n10089) );
  INV_X1 U12696 ( .A(n10394), .ZN(n10096) );
  OAI21_X1 U12697 ( .B1(n9666), .B2(n14956), .A(n13694), .ZN(n15124) );
  INV_X2 U12698 ( .A(n15345), .ZN(n12900) );
  NAND2_X1 U12699 ( .A1(n15359), .A2(n19188), .ZN(n10110) );
  INV_X1 U12700 ( .A(n10302), .ZN(n10111) );
  NAND3_X1 U12701 ( .A1(n10113), .A2(n12894), .A3(n12895), .ZN(n12896) );
  AND2_X2 U12702 ( .A1(n10276), .A2(n10277), .ZN(n15345) );
  NAND2_X1 U12703 ( .A1(n10115), .A2(n13485), .ZN(n13142) );
  NAND2_X1 U12704 ( .A1(n16137), .A2(n9712), .ZN(n16105) );
  NAND2_X1 U12705 ( .A1(n15112), .A2(n10126), .ZN(n14454) );
  NAND2_X1 U12706 ( .A1(n10129), .A2(n9731), .ZN(n10131) );
  INV_X1 U12707 ( .A(n14479), .ZN(n10129) );
  INV_X1 U12708 ( .A(n14468), .ZN(n10133) );
  NAND2_X1 U12709 ( .A1(n10136), .A2(n10134), .ZN(n12108) );
  XNOR2_X2 U12710 ( .A(n10969), .B(n10968), .ZN(n12099) );
  XNOR2_X2 U12711 ( .A(n12293), .B(n9729), .ZN(n14458) );
  NAND2_X1 U12712 ( .A1(n13289), .A2(n10141), .ZN(n14493) );
  INV_X1 U12713 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10143) );
  INV_X2 U12714 ( .A(n12199), .ZN(n12376) );
  NAND3_X2 U12715 ( .A1(n10144), .A2(n10143), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12199) );
  AND2_X2 U12716 ( .A1(n19073), .A2(n9716), .ZN(n19054) );
  AND2_X1 U12717 ( .A1(n11159), .A2(n11169), .ZN(n11110) );
  XNOR2_X1 U12718 ( .A(n14165), .B(n14164), .ZN(n14267) );
  NAND2_X1 U12719 ( .A1(n11918), .A2(n15773), .ZN(n14191) );
  NAND4_X1 U12720 ( .A1(n11176), .A2(n13048), .A3(n12906), .A4(n12902), .ZN(
        n11160) );
  OAI22_X1 U12721 ( .A1(n14172), .A2(n14294), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13820), .ZN(n13821) );
  NAND2_X1 U12722 ( .A1(n13819), .A2(n15819), .ZN(n14172) );
  NAND2_X1 U12723 ( .A1(n14281), .A2(n20071), .ZN(n11947) );
  NAND2_X1 U12724 ( .A1(n11250), .A2(n11249), .ZN(n11253) );
  INV_X1 U12725 ( .A(n13441), .ZN(n11440) );
  CLKBUF_X1 U12726 ( .A(n13441), .Z(n13497) );
  NAND2_X1 U12727 ( .A1(n10649), .A2(n9684), .ZN(n10650) );
  INV_X1 U12728 ( .A(n10566), .ZN(n10554) );
  OAI22_X1 U12729 ( .A1(n10204), .A2(n10203), .B1(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n19813), .ZN(n10209) );
  INV_X1 U12730 ( .A(n10697), .ZN(n10716) );
  OAI211_X2 U12731 ( .C1(n14298), .C2(n14273), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14180), .ZN(n13818) );
  XNOR2_X1 U12732 ( .A(n10567), .B(n10554), .ZN(n13449) );
  NAND2_X1 U12733 ( .A1(n13951), .A2(n11556), .ZN(n14070) );
  INV_X1 U12734 ( .A(n12218), .ZN(n14729) );
  NAND2_X1 U12735 ( .A1(n13747), .A2(n19855), .ZN(n11952) );
  AOI211_X1 U12736 ( .C1(n9600), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n17108), .B(n17107), .ZN(n17110) );
  AOI211_X1 U12737 ( .C1(n9600), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n17025), .B(n17024), .ZN(n17026) );
  AOI211_X1 U12738 ( .C1(n9600), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n15406), .B(n15405), .ZN(n15407) );
  AOI22_X1 U12739 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12487) );
  NOR2_X1 U12740 ( .A1(n10478), .A2(n9617), .ZN(n10479) );
  NAND2_X1 U12741 ( .A1(n10450), .A2(n9617), .ZN(n10465) );
  NOR2_X1 U12742 ( .A1(n10445), .A2(n9617), .ZN(n10466) );
  NOR2_X2 U12743 ( .A1(n11881), .A2(n11880), .ZN(n11882) );
  NAND2_X1 U12744 ( .A1(n13227), .A2(n13229), .ZN(n13228) );
  AND3_X1 U12745 ( .A1(n10260), .A2(n10259), .A3(n10258), .ZN(n10263) );
  CLKBUF_X1 U12746 ( .A(n14493), .Z(n16077) );
  INV_X1 U12747 ( .A(n19975), .ZN(n15753) );
  NAND2_X1 U12748 ( .A1(n19972), .A2(n13155), .ZN(n19975) );
  INV_X1 U12749 ( .A(n13133), .ZN(n13428) );
  INV_X1 U12750 ( .A(n18998), .ZN(n19022) );
  AND2_X1 U12751 ( .A1(n12802), .A2(n19797), .ZN(n18998) );
  AND3_X1 U12752 ( .A1(n11905), .A2(n15884), .A3(n15596), .ZN(n10147) );
  AND2_X1 U12753 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10149) );
  AND2_X1 U12754 ( .A1(n10364), .A2(n10811), .ZN(n10150) );
  AND3_X1 U12755 ( .A1(n10372), .A2(n19171), .A3(n10362), .ZN(n10151) );
  AND2_X1 U12756 ( .A1(n10410), .A2(n10412), .ZN(n10152) );
  NOR2_X1 U12757 ( .A1(n11957), .A2(n11956), .ZN(n10153) );
  INV_X1 U12758 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20156) );
  INV_X1 U12759 ( .A(n16401), .ZN(n16783) );
  INV_X1 U12760 ( .A(n16783), .ZN(n16758) );
  OR2_X1 U12761 ( .A1(n17053), .A2(n17099), .ZN(n10154) );
  INV_X1 U12762 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11873) );
  OR2_X1 U12763 ( .A1(n17678), .A2(n16267), .ZN(n10156) );
  AND2_X1 U12764 ( .A1(n17662), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10157) );
  OR3_X1 U12765 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17492), .ZN(n10158) );
  INV_X1 U12766 ( .A(n11269), .ZN(n11553) );
  NOR2_X1 U12767 ( .A1(n11154), .A2(n11268), .ZN(n11269) );
  NOR2_X1 U12768 ( .A1(n20564), .A2(n20333), .ZN(n10159) );
  OR2_X1 U12769 ( .A1(n13727), .A2(n13726), .ZN(n10160) );
  INV_X1 U12770 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11033) );
  INV_X1 U12771 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11905) );
  INV_X2 U12772 ( .A(n17147), .ZN(n17139) );
  INV_X1 U12773 ( .A(n14078), .ZN(n19966) );
  NOR2_X1 U12774 ( .A1(n20564), .A2(n20485), .ZN(n10161) );
  AND2_X1 U12775 ( .A1(n13886), .A2(n13807), .ZN(n10162) );
  NAND2_X1 U12776 ( .A1(n15744), .A2(n20070), .ZN(n10163) );
  OR2_X1 U12777 ( .A1(n18882), .A2(n18884), .ZN(n10166) );
  AND2_X1 U12778 ( .A1(n19062), .A2(n19061), .ZN(n10167) );
  NOR2_X1 U12779 ( .A1(n13369), .A2(n10372), .ZN(n10168) );
  INV_X1 U12780 ( .A(n10810), .ZN(n11997) );
  OR2_X1 U12781 ( .A1(n18788), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18966) );
  INV_X1 U12782 ( .A(n15819), .ZN(n11912) );
  AND2_X2 U12783 ( .A1(n12999), .A2(n13186), .ZN(n11133) );
  NAND2_X1 U12784 ( .A1(n11793), .A2(n11792), .ZN(n11800) );
  OR2_X1 U12785 ( .A1(n11800), .A2(n15548), .ZN(n11821) );
  INV_X1 U12786 ( .A(n11794), .ZN(n11790) );
  INV_X1 U12787 ( .A(n11821), .ZN(n11822) );
  INV_X1 U12788 ( .A(n11778), .ZN(n11156) );
  INV_X2 U12789 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10259) );
  NOR2_X1 U12790 ( .A1(n15352), .A2(n10507), .ZN(n10508) );
  NAND2_X1 U12791 ( .A1(n10353), .A2(n10358), .ZN(n10354) );
  AOI22_X1 U12792 ( .A1(n11811), .A2(n11855), .B1(n11824), .B2(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11355) );
  INV_X1 U12793 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11272) );
  OAI21_X1 U12794 ( .B1(n18734), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n12550), .ZN(n12551) );
  AND2_X1 U12795 ( .A1(n11186), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11066) );
  AOI22_X1 U12796 ( .A1(n11329), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11186), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11118) );
  OR2_X1 U12797 ( .A1(n11263), .A2(n11262), .ZN(n11840) );
  OR2_X1 U12798 ( .A1(n11335), .A2(n11334), .ZN(n11855) );
  INV_X1 U12799 ( .A(n12271), .ZN(n12272) );
  OR2_X1 U12800 ( .A1(n13671), .A2(n14813), .ZN(n13716) );
  AOI21_X1 U12801 ( .B1(n12642), .B2(n15504), .A(n13654), .ZN(n12639) );
  AOI21_X1 U12802 ( .B1(n11329), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n11066), .ZN(n11069) );
  INV_X1 U12803 ( .A(n13498), .ZN(n11439) );
  INV_X1 U12804 ( .A(n14357), .ZN(n14224) );
  OR2_X1 U12805 ( .A1(n11315), .A2(n11314), .ZN(n11884) );
  NAND2_X1 U12806 ( .A1(n10206), .A2(n10205), .ZN(n10216) );
  NOR2_X1 U12807 ( .A1(n10611), .A2(n10610), .ZN(n10845) );
  INV_X1 U12808 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14988) );
  OR2_X1 U12809 ( .A1(n18941), .A2(n10733), .ZN(n10767) );
  INV_X1 U12810 ( .A(n19171), .ZN(n10364) );
  INV_X1 U12811 ( .A(n18140), .ZN(n12640) );
  INV_X1 U12812 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16985) );
  INV_X1 U12813 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17076) );
  NOR2_X1 U12814 ( .A1(n17974), .A2(n17910), .ZN(n12522) );
  NOR2_X1 U12815 ( .A1(n17292), .A2(n12504), .ZN(n12507) );
  INV_X1 U12816 ( .A(n12401), .ZN(n12402) );
  AND2_X1 U12817 ( .A1(n13626), .A2(n13625), .ZN(n13627) );
  AND2_X1 U12818 ( .A1(n13806), .A2(n13805), .ZN(n13886) );
  NOR2_X1 U12819 ( .A1(n11768), .A2(n14174), .ZN(n11769) );
  AOI21_X1 U12820 ( .B1(n9618), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n14225), .ZN(n14338) );
  OR2_X1 U12821 ( .A1(n9620), .A2(n20693), .ZN(n14387) );
  INV_X1 U12822 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20234) );
  OR2_X1 U12823 ( .A1(n10865), .A2(n10864), .ZN(n19071) );
  AND2_X1 U12824 ( .A1(n12293), .A2(n9729), .ZN(n12294) );
  AND2_X1 U12825 ( .A1(n14729), .A2(n12220), .ZN(n12221) );
  INV_X1 U12826 ( .A(n10447), .ZN(n10455) );
  OR3_X1 U12827 ( .A1(n18826), .A2(n10733), .A3(n14866), .ZN(n14869) );
  AND4_X1 U12828 ( .A1(n10344), .A2(n13316), .A3(n12879), .A4(n10343), .ZN(
        n10345) );
  AND2_X1 U12829 ( .A1(n10348), .A2(n10305), .ZN(n10371) );
  INV_X1 U12830 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17105) );
  INV_X1 U12831 ( .A(n16274), .ZN(n17435) );
  NAND2_X1 U12832 ( .A1(n12524), .A2(n12519), .ZN(n12521) );
  NOR2_X1 U12833 ( .A1(n17690), .A2(n17689), .ZN(n17688) );
  AOI21_X1 U12834 ( .B1(n12562), .B2(n12626), .A(n12561), .ZN(n13649) );
  INV_X1 U12835 ( .A(n13281), .ZN(n13270) );
  INV_X1 U12836 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15717) );
  NAND2_X1 U12837 ( .A1(n20848), .A2(n13257), .ZN(n19931) );
  AND2_X1 U12838 ( .A1(n11771), .A2(n11770), .ZN(n11773) );
  INV_X1 U12839 ( .A(n13154), .ZN(n13161) );
  NAND2_X1 U12840 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n11925), .ZN(
        n13803) );
  NOR2_X1 U12841 ( .A1(n11410), .A2(n11409), .ZN(n11424) );
  BUF_X4 U12842 ( .A(n11900), .Z(n15819) );
  INV_X1 U12843 ( .A(n20128), .ZN(n20114) );
  INV_X1 U12844 ( .A(n15553), .ZN(n13006) );
  OR2_X1 U12845 ( .A1(n20403), .A2(n20641), .ZN(n20391) );
  INV_X1 U12846 ( .A(n20232), .ZN(n20490) );
  INV_X1 U12847 ( .A(n20696), .ZN(n20538) );
  INV_X1 U12848 ( .A(n11869), .ZN(n20141) );
  OR2_X1 U12849 ( .A1(n19846), .A2(n12024), .ZN(n19004) );
  NAND2_X1 U12850 ( .A1(n14923), .A2(n14922), .ZN(n11019) );
  OR2_X1 U12851 ( .A1(n10917), .A2(n10916), .ZN(n19053) );
  INV_X1 U12852 ( .A(n13757), .ZN(n13758) );
  OR2_X1 U12853 ( .A1(n19102), .A2(n14511), .ZN(n19090) );
  INV_X1 U12854 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13524) );
  NOR2_X1 U12855 ( .A1(n12877), .A2(n15321), .ZN(n13540) );
  AOI211_X1 U12856 ( .C1(n9658), .C2(n19152), .A(n15018), .B(n15017), .ZN(
        n15019) );
  INV_X1 U12857 ( .A(n15112), .ZN(n15113) );
  AND2_X1 U12858 ( .A1(n10682), .A2(n10681), .ZN(n15257) );
  AND2_X1 U12859 ( .A1(n10371), .A2(n10370), .ZN(n13336) );
  INV_X1 U12860 ( .A(n18992), .ZN(n18974) );
  AND2_X1 U12861 ( .A1(n15366), .A2(n19808), .ZN(n19588) );
  AND2_X1 U12862 ( .A1(n19377), .A2(n19376), .ZN(n19380) );
  NAND2_X1 U12863 ( .A1(n19807), .A2(n19808), .ZN(n19442) );
  NOR2_X1 U12864 ( .A1(n18125), .A2(n17348), .ZN(n12632) );
  NOR2_X1 U12865 ( .A1(n13649), .A2(n13648), .ZN(n16381) );
  NOR2_X1 U12866 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16626), .ZN(n16611) );
  INV_X1 U12867 ( .A(n16790), .ZN(n16782) );
  INV_X1 U12868 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16986) );
  INV_X1 U12869 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16918) );
  INV_X1 U12870 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17063) );
  INV_X1 U12871 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17072) );
  NOR2_X1 U12872 ( .A1(n18617), .A2(n16381), .ZN(n17346) );
  INV_X1 U12873 ( .A(n12517), .ZN(n12515) );
  NAND2_X1 U12874 ( .A1(n12531), .A2(n10158), .ZN(n12532) );
  NOR2_X1 U12875 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18124), .ZN(n18410) );
  NAND2_X1 U12876 ( .A1(n11605), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11639) );
  NOR2_X1 U12877 ( .A1(n11604), .A2(n14202), .ZN(n11605) );
  NAND2_X1 U12878 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n11367), .ZN(
        n11387) );
  AND2_X1 U12879 ( .A1(n19931), .A2(n13282), .ZN(n19961) );
  AND2_X1 U12880 ( .A1(n19970), .A2(n13810), .ZN(n19965) );
  INV_X1 U12881 ( .A(n14133), .ZN(n15752) );
  INV_X1 U12882 ( .A(n19870), .ZN(n13152) );
  INV_X1 U12883 ( .A(n13139), .ZN(n20052) );
  NAND2_X1 U12884 ( .A1(n11727), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11768) );
  NOR2_X1 U12885 ( .A1(n11442), .A2(n11441), .ZN(n11443) );
  NOR2_X1 U12886 ( .A1(n20091), .A2(n14343), .ZN(n20103) );
  INV_X1 U12887 ( .A(n14376), .ZN(n20113) );
  INV_X1 U12888 ( .A(n13016), .ZN(n20832) );
  INV_X1 U12889 ( .A(n20751), .ZN(n20170) );
  INV_X1 U12890 ( .A(n20260), .ZN(n20222) );
  OR2_X1 U12891 ( .A1(n9620), .A2(n11869), .ZN(n20609) );
  INV_X1 U12892 ( .A(n20291), .ZN(n20300) );
  OR2_X1 U12893 ( .A1(n20140), .A2(n20139), .ZN(n20276) );
  INV_X1 U12894 ( .A(n20380), .ZN(n20393) );
  INV_X1 U12895 ( .A(n20391), .ZN(n20424) );
  OAI211_X1 U12896 ( .C1(n10161), .C2(n20570), .A(n20490), .B(n20436), .ZN(
        n20453) );
  OR2_X1 U12897 ( .A1(n9620), .A2(n20141), .ZN(n20565) );
  INV_X1 U12898 ( .A(n20520), .ZN(n20511) );
  INV_X1 U12899 ( .A(n20563), .ZN(n20546) );
  NAND2_X1 U12900 ( .A1(n9620), .A2(n11869), .ZN(n20641) );
  NAND2_X1 U12901 ( .A1(n14396), .A2(n20140), .ZN(n20541) );
  OAI211_X1 U12902 ( .C1(n20677), .C2(n20648), .A(n20647), .B(n20646), .ZN(
        n20680) );
  INV_X1 U12903 ( .A(n20596), .ZN(n20736) );
  NAND2_X1 U12904 ( .A1(n20139), .A2(n14394), .ZN(n20642) );
  INV_X1 U12905 ( .A(n20818), .ZN(n20819) );
  NAND2_X1 U12906 ( .A1(n12076), .A2(n18998), .ZN(n12077) );
  NAND2_X1 U12907 ( .A1(n15997), .A2(n15998), .ZN(n15996) );
  OR2_X1 U12908 ( .A1(n15986), .A2(n12027), .ZN(n19028) );
  AND2_X1 U12909 ( .A1(n15984), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n19026) );
  INV_X1 U12910 ( .A(n18850), .ZN(n19038) );
  OR2_X1 U12911 ( .A1(n10880), .A2(n10879), .ZN(n19062) );
  INV_X1 U12912 ( .A(n14425), .ZN(n12969) );
  INV_X1 U12913 ( .A(n19090), .ZN(n14755) );
  INV_X1 U12914 ( .A(n12812), .ZN(n12829) );
  INV_X1 U12915 ( .A(n12833), .ZN(n12809) );
  NOR2_X1 U12916 ( .A1(n12718), .A2(n12075), .ZN(n12802) );
  AND2_X1 U12917 ( .A1(n16161), .A2(n15005), .ZN(n16151) );
  NOR2_X2 U12918 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13540), .ZN(n19593) );
  OAI21_X1 U12919 ( .B1(n11030), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11029), .ZN(n11031) );
  AND2_X1 U12920 ( .A1(n11026), .A2(n19838), .ZN(n16200) );
  AND2_X1 U12921 ( .A1(n11026), .A2(n13336), .ZN(n13479) );
  AND2_X1 U12922 ( .A1(n11026), .A2(n10963), .ZN(n19152) );
  AND2_X1 U12923 ( .A1(n13334), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15321) );
  OAI21_X1 U12924 ( .B1(n15328), .B2(n15331), .A(n15327), .ZN(n19195) );
  INV_X1 U12925 ( .A(n19274), .ZN(n19255) );
  OAI21_X1 U12926 ( .B1(n19292), .B2(n19291), .A(n19290), .ZN(n19314) );
  INV_X1 U12927 ( .A(n19588), .ZN(n19554) );
  NOR2_X1 U12928 ( .A1(n19796), .A2(n19280), .ZN(n19401) );
  NAND2_X1 U12929 ( .A1(n15366), .A2(n19817), .ZN(n19796) );
  NOR2_X1 U12930 ( .A1(n15366), .A2(n19808), .ZN(n19482) );
  INV_X1 U12931 ( .A(n19501), .ZN(n19545) );
  INV_X1 U12932 ( .A(n19482), .ZN(n19518) );
  AND2_X1 U12933 ( .A1(n19592), .A2(n19585), .ZN(n19618) );
  OAI21_X1 U12934 ( .B1(n15380), .B2(n15383), .A(n15379), .ZN(n19646) );
  NOR2_X2 U12935 ( .A1(n19555), .A2(n19796), .ZN(n19695) );
  INV_X1 U12936 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19717) );
  INV_X1 U12937 ( .A(n12632), .ZN(n12645) );
  NOR2_X1 U12938 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16578), .ZN(n16563) );
  NOR2_X1 U12939 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16653), .ZN(n16632) );
  NOR2_X2 U12940 ( .A1(n18743), .A2(n16776), .ZN(n16761) );
  INV_X1 U12941 ( .A(n17166), .ZN(n17163) );
  NOR2_X1 U12942 ( .A1(n17401), .A2(n17265), .ZN(n17261) );
  NOR2_X1 U12943 ( .A1(n17199), .A2(n18584), .ZN(n15605) );
  INV_X1 U12944 ( .A(n17346), .ZN(n17345) );
  NAND2_X1 U12945 ( .A1(n17588), .A2(n12686), .ZN(n17923) );
  INV_X1 U12946 ( .A(n17631), .ZN(n17605) );
  INV_X1 U12947 ( .A(n17765), .ZN(n17656) );
  INV_X1 U12948 ( .A(n17845), .ZN(n17920) );
  NOR2_X1 U12949 ( .A1(n17975), .A2(n17595), .ZN(n17588) );
  INV_X1 U12950 ( .A(n18110), .ZN(n18097) );
  INV_X1 U12951 ( .A(n18259), .ZN(n18267) );
  INV_X1 U12952 ( .A(n18277), .ZN(n18291) );
  INV_X1 U12953 ( .A(n18445), .ZN(n18452) );
  INV_X1 U12954 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18629) );
  INV_X1 U12955 ( .A(n14158), .ZN(n20147) );
  INV_X1 U12956 ( .A(n19955), .ZN(n19913) );
  INV_X1 U12957 ( .A(n19926), .ZN(n19952) );
  AOI21_X1 U12958 ( .B1(n13404), .B2(n13403), .A(n19870), .ZN(n14091) );
  OR2_X1 U12959 ( .A1(n13813), .A2(n20147), .ZN(n15756) );
  AND2_X1 U12960 ( .A1(n13153), .A2(n13152), .ZN(n19972) );
  NOR2_X1 U12961 ( .A1(n20008), .A2(n20036), .ZN(n20022) );
  INV_X1 U12962 ( .A(n20008), .ZN(n20038) );
  NOR2_X1 U12963 ( .A1(n13078), .A2(n13077), .ZN(n13138) );
  NAND2_X1 U12964 ( .A1(n13891), .A2(n13890), .ZN(n14171) );
  OAI21_X1 U12965 ( .B1(n14095), .B2(n13969), .A(n13968), .ZN(n14246) );
  INV_X1 U12966 ( .A(n20079), .ZN(n20075) );
  NAND2_X1 U12967 ( .A1(n13610), .A2(n20103), .ZN(n15953) );
  OR2_X1 U12968 ( .A1(n13044), .A2(n13058), .ZN(n20120) );
  INV_X1 U12969 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20138) );
  INV_X1 U12970 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12990) );
  AOI211_X2 U12971 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20307), .A(n20232), 
        .B(n20145), .ZN(n20204) );
  OR2_X1 U12972 ( .A1(n20276), .A2(n20565), .ZN(n20225) );
  OR2_X1 U12973 ( .A1(n20276), .A2(n20609), .ZN(n20260) );
  OR2_X1 U12974 ( .A1(n20276), .A2(n20641), .ZN(n20291) );
  OR2_X1 U12975 ( .A1(n20276), .A2(n20540), .ZN(n20325) );
  OR2_X1 U12976 ( .A1(n20403), .A2(n20565), .ZN(n20358) );
  AOI22_X1 U12977 ( .A1(n20366), .A2(n20364), .B1(n20362), .B2(n20361), .ZN(
        n20397) );
  NAND2_X1 U12978 ( .A1(n20399), .A2(n20398), .ZN(n20456) );
  OR2_X1 U12979 ( .A1(n20541), .A2(n20565), .ZN(n20480) );
  AOI22_X1 U12980 ( .A1(n20488), .A2(n20486), .B1(n20484), .B2(n20483), .ZN(
        n20526) );
  OR2_X1 U12981 ( .A1(n20541), .A2(n20641), .ZN(n20563) );
  OR2_X1 U12982 ( .A1(n20541), .A2(n20540), .ZN(n20608) );
  NAND2_X1 U12983 ( .A1(n20694), .A2(n20610), .ZN(n20683) );
  OR2_X1 U12984 ( .A1(n20642), .A2(n20540), .ZN(n20751) );
  INV_X1 U12985 ( .A(n20830), .ZN(n20759) );
  INV_X1 U12986 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19855) );
  AND2_X1 U12987 ( .A1(n12078), .A2(n12077), .ZN(n12079) );
  INV_X1 U12988 ( .A(n19008), .ZN(n19032) );
  INV_X1 U12989 ( .A(n12396), .ZN(n12397) );
  AND2_X2 U12990 ( .A1(n12394), .A2(n19700), .ZN(n19070) );
  INV_X1 U12991 ( .A(n19102), .ZN(n14687) );
  AND2_X1 U12992 ( .A1(n16083), .A2(n16085), .ZN(n19111) );
  OR2_X1 U12993 ( .A1(n10349), .A2(n19102), .ZN(n16083) );
  NAND2_X1 U12994 ( .A1(n12836), .A2(n19856), .ZN(n19150) );
  OR2_X1 U12995 ( .A1(n12718), .A2(n15338), .ZN(n12833) );
  INV_X1 U12996 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16122) );
  INV_X1 U12997 ( .A(n16151), .ZN(n16150) );
  OR2_X1 U12998 ( .A1(n18792), .A2(n15338), .ZN(n16154) );
  INV_X1 U12999 ( .A(n11031), .ZN(n11032) );
  NAND2_X1 U13000 ( .A1(n11026), .A2(n19836), .ZN(n16189) );
  AND2_X1 U13001 ( .A1(n10690), .A2(n10689), .ZN(n16196) );
  AOI211_X2 U13002 ( .C1(n15332), .C2(n15331), .A(n15330), .B(n19285), .ZN(
        n19199) );
  INV_X1 U13003 ( .A(n19194), .ZN(n19225) );
  NOR2_X1 U13004 ( .A1(n15356), .A2(n19285), .ZN(n19243) );
  OR2_X1 U13005 ( .A1(n19280), .A2(n19518), .ZN(n19274) );
  OR2_X1 U13006 ( .A1(n19375), .A2(n19518), .ZN(n19318) );
  OR2_X1 U13007 ( .A1(n19280), .A2(n19554), .ZN(n19355) );
  OR2_X1 U13008 ( .A1(n19375), .A2(n19554), .ZN(n19368) );
  INV_X1 U13009 ( .A(n19401), .ZN(n19397) );
  OR2_X1 U13010 ( .A1(n19375), .A2(n19796), .ZN(n19436) );
  NAND2_X1 U13011 ( .A1(n19483), .A2(n19444), .ZN(n19473) );
  INV_X1 U13012 ( .A(n19498), .ZN(n19509) );
  OR2_X1 U13013 ( .A1(n19510), .A2(n19518), .ZN(n19582) );
  INV_X1 U13014 ( .A(n19521), .ZN(n19598) );
  INV_X1 U13015 ( .A(n19684), .ZN(n19616) );
  AOI21_X1 U13016 ( .B1(n13536), .B2(n15378), .A(n13535), .ZN(n19699) );
  NOR2_X1 U13017 ( .A1(n18550), .A2(n17345), .ZN(n18782) );
  OR2_X1 U13018 ( .A1(n18629), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18777) );
  INV_X1 U13019 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17685) );
  INV_X1 U13020 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17720) );
  INV_X1 U13021 ( .A(n17283), .ZN(n17308) );
  NAND2_X1 U13022 ( .A1(n17326), .A2(n18125), .ZN(n17325) );
  INV_X1 U13023 ( .A(n17326), .ZN(n17344) );
  INV_X1 U13024 ( .A(n18009), .ZN(n18021) );
  NAND2_X1 U13025 ( .A1(n17988), .A2(n18016), .ZN(n18089) );
  INV_X1 U13026 ( .A(n18050), .ZN(n18108) );
  INV_X1 U13027 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18600) );
  AOI21_X1 U13028 ( .B1(n18771), .B2(n18582), .A(n13661), .ZN(n18748) );
  INV_X1 U13029 ( .A(n18481), .ZN(n18473) );
  CLKBUF_X1 U13030 ( .A(n16373), .Z(n16374) );
  NAND2_X1 U13031 ( .A1(n11917), .A2(n11916), .ZN(P1_U2971) );
  OAI21_X1 U13032 ( .B1(n11034), .B2(n11033), .A(n11032), .ZN(P2_U3029) );
  AND2_X4 U13033 ( .A1(n13324), .A2(n10170), .ZN(n10314) );
  INV_X2 U13034 ( .A(n12199), .ZN(n10293) );
  AOI22_X1 U13035 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12376), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10176) );
  AND2_X4 U13036 ( .A1(n13347), .A2(n13301), .ZN(n12377) );
  AOI22_X1 U13037 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10175) );
  AND2_X2 U13038 ( .A1(n10143), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13346) );
  AND2_X4 U13039 ( .A1(n13346), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12382) );
  AND2_X4 U13040 ( .A1(n10172), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12381) );
  AOI22_X1 U13041 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10174) );
  AND2_X4 U13042 ( .A1(n10315), .A2(n10170), .ZN(n10316) );
  AOI22_X1 U13043 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10173) );
  NAND4_X1 U13044 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10182) );
  AOI22_X1 U13045 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U13046 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U13047 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U13048 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10177) );
  NAND4_X1 U13049 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(
        n10181) );
  MUX2_X2 U13050 ( .A(n10182), .B(n10181), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13369) );
  AOI22_X1 U13051 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12376), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U13052 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U13053 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U13054 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10183) );
  NAND4_X1 U13055 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n10187) );
  NAND2_X1 U13056 ( .A1(n10187), .A2(n10259), .ZN(n10194) );
  AOI22_X1 U13057 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10314), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U13058 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13059 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U13060 ( .A1(n12376), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10188) );
  NAND4_X1 U13061 ( .A1(n10191), .A2(n10190), .A3(n10189), .A4(n10188), .ZN(
        n10192) );
  NAND2_X1 U13062 ( .A1(n10192), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10193) );
  NAND2_X2 U13063 ( .A1(n10194), .A2(n10193), .ZN(n10809) );
  XNOR2_X1 U13064 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U13065 ( .A1(n19830), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10199) );
  INV_X1 U13066 ( .A(n10199), .ZN(n10195) );
  NAND2_X1 U13067 ( .A1(n10200), .A2(n10195), .ZN(n10197) );
  NAND2_X1 U13068 ( .A1(n19821), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10196) );
  NAND2_X1 U13069 ( .A1(n10197), .A2(n10196), .ZN(n10204) );
  XNOR2_X1 U13070 ( .A(n13301), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10198) );
  XNOR2_X1 U13071 ( .A(n10204), .B(n10198), .ZN(n10225) );
  INV_X1 U13072 ( .A(n10225), .ZN(n10210) );
  OAI21_X1 U13073 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19830), .A(
        n10199), .ZN(n10337) );
  INV_X1 U13074 ( .A(n10337), .ZN(n10720) );
  XNOR2_X1 U13075 ( .A(n10200), .B(n10199), .ZN(n10227) );
  OAI211_X1 U13076 ( .C1(n15338), .C2(n10720), .A(n13541), .B(n10227), .ZN(
        n10202) );
  INV_X1 U13077 ( .A(n10200), .ZN(n10331) );
  OAI21_X1 U13078 ( .B1(n10331), .B2(n10337), .A(n10698), .ZN(n10201) );
  OAI211_X1 U13079 ( .C1(n10382), .C2(n10210), .A(n10202), .B(n10201), .ZN(
        n10214) );
  NOR2_X1 U13080 ( .A1(n13301), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10203) );
  XNOR2_X1 U13081 ( .A(n10259), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10207) );
  NAND2_X1 U13082 ( .A1(n19805), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10205) );
  INV_X1 U13083 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15494) );
  NAND2_X1 U13084 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15494), .ZN(
        n10217) );
  INV_X1 U13085 ( .A(n10207), .ZN(n10208) );
  XNOR2_X1 U13086 ( .A(n10209), .B(n10208), .ZN(n10699) );
  NAND2_X1 U13087 ( .A1(n13369), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U13088 ( .A1(n12837), .A2(n15338), .ZN(n10211) );
  NAND2_X1 U13089 ( .A1(n10211), .A2(n10210), .ZN(n10212) );
  NAND2_X1 U13090 ( .A1(n10808), .A2(n10225), .ZN(n10329) );
  NAND2_X1 U13091 ( .A1(n10212), .A2(n10329), .ZN(n10213) );
  NAND3_X1 U13092 ( .A1(n10214), .A2(n10332), .A3(n10213), .ZN(n10221) );
  INV_X1 U13093 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15600) );
  AND2_X1 U13094 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15600), .ZN(
        n10215) );
  OAI21_X1 U13095 ( .B1(n10332), .B2(n10808), .A(n10334), .ZN(n10219) );
  INV_X1 U13096 ( .A(n10219), .ZN(n10220) );
  NAND2_X1 U13097 ( .A1(n10221), .A2(n10220), .ZN(n10222) );
  MUX2_X1 U13098 ( .A(n10222), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19855), .Z(n10251) );
  INV_X1 U13099 ( .A(n10334), .ZN(n10223) );
  NAND2_X1 U13100 ( .A1(n10375), .A2(n10223), .ZN(n10224) );
  NAND2_X1 U13101 ( .A1(n13334), .A2(n15338), .ZN(n13312) );
  NAND2_X1 U13102 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19850) );
  INV_X1 U13103 ( .A(n19850), .ZN(n19845) );
  NAND2_X1 U13104 ( .A1(n19717), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19864) );
  INV_X2 U13105 ( .A(n19864), .ZN(n19867) );
  NAND2_X2 U13106 ( .A1(n19867), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19776) );
  NOR2_X1 U13107 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19713) );
  INV_X1 U13108 ( .A(n19713), .ZN(n19723) );
  NAND3_X1 U13109 ( .A1(n19717), .A2(n19776), .A3(n19723), .ZN(n12835) );
  NOR2_X1 U13110 ( .A1(n19845), .A2(n12835), .ZN(n13371) );
  INV_X1 U13111 ( .A(n13371), .ZN(n13313) );
  NAND2_X1 U13112 ( .A1(n10332), .A2(n10225), .ZN(n10336) );
  INV_X1 U13113 ( .A(n10336), .ZN(n10226) );
  NAND2_X1 U13114 ( .A1(n10227), .A2(n10226), .ZN(n10228) );
  NAND2_X1 U13115 ( .A1(n13338), .A2(n19850), .ZN(n10229) );
  OAI22_X1 U13116 ( .A1(n13312), .A2(n13313), .B1(n10229), .B2(n15338), .ZN(
        n10240) );
  AOI22_X1 U13117 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U13118 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10232) );
  AOI22_X1 U13119 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U13120 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10230) );
  AOI22_X1 U13121 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10314), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U13122 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U13123 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10235) );
  AOI22_X1 U13124 ( .A1(n12376), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10234) );
  MUX2_X2 U13125 ( .A(n10239), .B(n10238), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10372) );
  NAND2_X1 U13126 ( .A1(n10240), .A2(n10358), .ZN(n10346) );
  AOI22_X1 U13127 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U13128 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U13129 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U13130 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10241) );
  NAND4_X1 U13131 ( .A1(n10244), .A2(n10243), .A3(n10242), .A4(n10241), .ZN(
        n10250) );
  AOI22_X1 U13132 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12376), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10248) );
  AOI22_X1 U13133 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10247) );
  AOI22_X1 U13134 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U13135 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10245) );
  NAND4_X1 U13136 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        n10249) );
  MUX2_X2 U13137 ( .A(n10250), .B(n10249), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10388) );
  AOI21_X1 U13138 ( .B1(n10251), .B2(n13541), .A(n15359), .ZN(n10252) );
  NAND2_X1 U13139 ( .A1(n13312), .A2(n10252), .ZN(n10344) );
  AOI22_X1 U13140 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U13141 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U13142 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__5__SCAN_IN), .B2(n10293), .ZN(n10255) );
  AOI22_X1 U13143 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10254) );
  NAND4_X1 U13144 ( .A1(n10257), .A2(n10256), .A3(n10255), .A4(n10254), .ZN(
        n10265) );
  AOI22_X1 U13145 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U13146 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U13147 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U13148 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12376), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10261) );
  NAND3_X1 U13149 ( .A1(n10263), .A2(n10262), .A3(n10261), .ZN(n10264) );
  NAND2_X2 U13150 ( .A1(n10265), .A2(n10264), .ZN(n10302) );
  AOI22_X1 U13151 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10269) );
  AOI22_X1 U13152 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10268) );
  AOI22_X1 U13153 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U13154 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10266) );
  NAND4_X1 U13155 ( .A1(n10269), .A2(n10268), .A3(n10267), .A4(n10266), .ZN(
        n10270) );
  NAND2_X1 U13156 ( .A1(n10270), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10277) );
  AOI22_X1 U13157 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10314), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10274) );
  AOI22_X1 U13158 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n12381), .ZN(n10273) );
  AOI22_X1 U13159 ( .A1(n12376), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U13160 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10316), .B1(
        n10317), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10271) );
  NAND4_X1 U13161 ( .A1(n10274), .A2(n10273), .A3(n10272), .A4(n10271), .ZN(
        n10275) );
  NAND2_X1 U13162 ( .A1(n10275), .A2(n10259), .ZN(n10276) );
  AOI22_X1 U13163 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12376), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U13164 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U13165 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U13166 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10278) );
  NAND4_X1 U13167 ( .A1(n10281), .A2(n10280), .A3(n10279), .A4(n10278), .ZN(
        n10287) );
  AOI22_X1 U13168 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U13169 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U13170 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U13171 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10282) );
  NAND4_X1 U13172 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10286) );
  MUX2_X2 U13173 ( .A(n10287), .B(n10286), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19171) );
  AOI22_X1 U13174 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12376), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U13175 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10290) );
  AOI22_X1 U13176 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12383), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13177 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10288) );
  NAND4_X1 U13178 ( .A1(n10291), .A2(n10290), .A3(n10289), .A4(n10288), .ZN(
        n10292) );
  NAND2_X1 U13179 ( .A1(n10292), .A2(n10259), .ZN(n10300) );
  AOI22_X1 U13180 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13181 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U13182 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10295) );
  AOI22_X1 U13183 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10316), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10294) );
  NAND4_X1 U13184 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10298) );
  NAND2_X1 U13185 ( .A1(n10298), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10299) );
  NAND3_X1 U13186 ( .A1(n10394), .A2(n13338), .A3(n19850), .ZN(n10341) );
  NAND2_X2 U13187 ( .A1(n10111), .A2(n19188), .ZN(n10349) );
  NAND2_X1 U13188 ( .A1(n10302), .A2(n10362), .ZN(n10301) );
  NAND2_X1 U13189 ( .A1(n10349), .A2(n10301), .ZN(n10307) );
  AND2_X1 U13190 ( .A1(n19852), .A2(n13369), .ZN(n12016) );
  OAI21_X1 U13191 ( .B1(n10307), .B2(n15345), .A(n12016), .ZN(n10348) );
  INV_X2 U13192 ( .A(n10302), .ZN(n10811) );
  NAND2_X1 U13193 ( .A1(n10349), .A2(n10388), .ZN(n10312) );
  NAND2_X1 U13194 ( .A1(n10312), .A2(n10303), .ZN(n10304) );
  NAND2_X1 U13195 ( .A1(n15492), .A2(n10304), .ZN(n10305) );
  AND3_X1 U13196 ( .A1(n12900), .A2(n10388), .A3(n19852), .ZN(n10370) );
  NAND2_X1 U13197 ( .A1(n13369), .A2(n12900), .ZN(n10306) );
  NAND2_X1 U13198 ( .A1(n10306), .A2(n10372), .ZN(n10308) );
  INV_X1 U13199 ( .A(n10309), .ZN(n10310) );
  OAI211_X1 U13200 ( .C1(n10341), .C2(n12835), .A(n10371), .B(n10310), .ZN(
        n10311) );
  INV_X1 U13201 ( .A(n10311), .ZN(n13316) );
  INV_X1 U13202 ( .A(n12016), .ZN(n19854) );
  AND2_X2 U13203 ( .A1(n12370), .A2(n10259), .ZN(n10490) );
  AND2_X1 U13204 ( .A1(n10314), .A2(n10259), .ZN(n10491) );
  AOI22_X1 U13205 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9601), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10321) );
  AND2_X2 U13206 ( .A1(n12376), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10524) );
  AOI22_X1 U13207 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10523), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10320) );
  AND2_X2 U13208 ( .A1(n12370), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10536) );
  INV_X1 U13209 ( .A(n10315), .ZN(n13325) );
  NOR2_X1 U13210 ( .A1(n13325), .A2(n10259), .ZN(n13304) );
  AND2_X2 U13211 ( .A1(n13304), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12186) );
  AOI22_X1 U13212 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n12186), .ZN(n10319) );
  AND2_X2 U13213 ( .A1(n10317), .A2(n10259), .ZN(n13295) );
  AOI22_X1 U13214 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10529), .B1(
        n13295), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10318) );
  NAND4_X1 U13215 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n10318), .ZN(
        n10328) );
  AND2_X1 U13216 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10322) );
  AND2_X1 U13217 ( .A1(n13347), .A2(n10322), .ZN(n10542) );
  AOI22_X1 U13218 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n10542), .ZN(n10326) );
  AOI22_X1 U13219 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__2__SCAN_IN), .B2(n10544), .ZN(n10325) );
  AOI22_X1 U13220 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13221 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10572), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10323) );
  NAND4_X1 U13222 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10327) );
  NAND2_X1 U13223 ( .A1(n10698), .A2(n10833), .ZN(n10330) );
  NAND2_X1 U13224 ( .A1(n10330), .A2(n10329), .ZN(n10696) );
  NOR2_X1 U13225 ( .A1(n10331), .A2(n10337), .ZN(n10333) );
  OAI21_X1 U13226 ( .B1(n10696), .B2(n10333), .A(n10332), .ZN(n10335) );
  AND2_X1 U13227 ( .A1(n10335), .A2(n10334), .ZN(n19834) );
  NAND2_X1 U13228 ( .A1(n19836), .A2(n19834), .ZN(n12879) );
  OAI21_X1 U13229 ( .B1(n10337), .B2(n10336), .A(n13338), .ZN(n10338) );
  INV_X1 U13230 ( .A(n10338), .ZN(n10340) );
  OR2_X1 U13231 ( .A1(n13304), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n15490) );
  INV_X1 U13232 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n10339) );
  OAI21_X1 U13233 ( .B1(n10496), .B2(n15490), .A(n10339), .ZN(n19823) );
  MUX2_X1 U13234 ( .A(n10340), .B(n19823), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n16220) );
  INV_X1 U13235 ( .A(n16220), .ZN(n19837) );
  OAI21_X1 U13236 ( .B1(n10374), .B2(n19837), .A(n10341), .ZN(n10342) );
  NAND2_X1 U13237 ( .A1(n10342), .A2(n15338), .ZN(n10343) );
  NAND2_X1 U13238 ( .A1(n10346), .A2(n10345), .ZN(n10347) );
  AND2_X1 U13239 ( .A1(n19844), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12023) );
  NAND2_X1 U13240 ( .A1(n10363), .A2(n15338), .ZN(n13344) );
  AOI21_X1 U13241 ( .B1(n13344), .B2(n10348), .A(n10364), .ZN(n10361) );
  NAND2_X1 U13242 ( .A1(n10349), .A2(n19171), .ZN(n10351) );
  AND3_X1 U13243 ( .A1(n10351), .A2(n12900), .A3(n10110), .ZN(n10357) );
  AND2_X1 U13244 ( .A1(n10755), .A2(n10362), .ZN(n10352) );
  NAND2_X1 U13245 ( .A1(n10352), .A2(n10372), .ZN(n10355) );
  NAND2_X1 U13246 ( .A1(n15359), .A2(n10755), .ZN(n10353) );
  NAND2_X1 U13247 ( .A1(n10357), .A2(n10356), .ZN(n10377) );
  MUX2_X1 U13248 ( .A(n10358), .B(n10377), .S(n13541), .Z(n10360) );
  NOR2_X1 U13249 ( .A1(n12893), .A2(n15359), .ZN(n10359) );
  NOR3_X1 U13250 ( .A1(n10361), .A2(n10360), .A3(n10359), .ZN(n10367) );
  MUX2_X1 U13251 ( .A(n10393), .B(n10363), .S(n19171), .Z(n10380) );
  NAND2_X1 U13252 ( .A1(n10349), .A2(n19852), .ZN(n10376) );
  NAND2_X1 U13253 ( .A1(n10380), .A2(n10376), .ZN(n10411) );
  NAND2_X1 U13254 ( .A1(n10411), .A2(n12893), .ZN(n10365) );
  NAND2_X1 U13255 ( .A1(n10365), .A2(n12895), .ZN(n10366) );
  NAND2_X1 U13256 ( .A1(n13356), .A2(n10368), .ZN(n10369) );
  NAND2_X1 U13257 ( .A1(n11026), .A2(n10369), .ZN(n10688) );
  INV_X1 U13258 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12275) );
  AND2_X1 U13259 ( .A1(n10372), .A2(n15338), .ZN(n10373) );
  NOR2_X1 U13260 ( .A1(n13369), .A2(n19855), .ZN(n19851) );
  OAI21_X1 U13261 ( .B1(n10377), .B2(n10376), .A(n19851), .ZN(n10378) );
  NAND2_X1 U13262 ( .A1(n19855), .A2(n19844), .ZN(n10406) );
  NAND2_X1 U13263 ( .A1(n11022), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10383) );
  OAI21_X1 U13264 ( .B1(n19821), .B2(n10406), .A(n10383), .ZN(n10384) );
  AOI21_X2 U13265 ( .B1(n10428), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10384), .ZN(n10414) );
  INV_X1 U13266 ( .A(n16215), .ZN(n10385) );
  NAND2_X1 U13267 ( .A1(n10385), .A2(n19852), .ZN(n13381) );
  OAI21_X1 U13268 ( .B1(n19171), .B2(n13369), .A(n10302), .ZN(n10386) );
  INV_X1 U13269 ( .A(n10386), .ZN(n10387) );
  NOR2_X1 U13270 ( .A1(n10387), .A2(n10150), .ZN(n10390) );
  AND3_X1 U13271 ( .A1(n19188), .A2(n10388), .A3(n12900), .ZN(n10389) );
  NAND3_X1 U13272 ( .A1(n13381), .A2(n10391), .A3(n11023), .ZN(n10392) );
  INV_X1 U13273 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10398) );
  AND2_X4 U13274 ( .A1(n10395), .A2(n10394), .ZN(n12065) );
  NAND2_X1 U13275 ( .A1(n12065), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U13276 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10396) );
  OAI211_X1 U13277 ( .C1(n12069), .C2(n10398), .A(n10397), .B(n10396), .ZN(
        n10399) );
  AOI21_X2 U13278 ( .B1(n10432), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10399), .ZN(n10415) );
  INV_X1 U13279 ( .A(n10400), .ZN(n10401) );
  INV_X1 U13280 ( .A(n10406), .ZN(n10429) );
  NAND2_X1 U13281 ( .A1(n10428), .A2(n10402), .ZN(n10403) );
  NAND2_X1 U13282 ( .A1(n10404), .A2(n10403), .ZN(n10439) );
  NAND2_X1 U13283 ( .A1(n12065), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U13284 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10405) );
  NAND4_X1 U13285 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10409) );
  INV_X1 U13286 ( .A(n10414), .ZN(n10416) );
  OAI21_X1 U13287 ( .B1(n19813), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n19844), 
        .ZN(n10417) );
  INV_X1 U13288 ( .A(n10425), .ZN(n10423) );
  INV_X1 U13289 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10420) );
  NAND2_X1 U13290 ( .A1(n12065), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10419) );
  NAND2_X1 U13291 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10418) );
  OAI211_X1 U13292 ( .C1(n12069), .C2(n10420), .A(n10419), .B(n10418), .ZN(
        n10421) );
  INV_X1 U13293 ( .A(n10424), .ZN(n10422) );
  NAND2_X1 U13294 ( .A1(n10423), .A2(n10422), .ZN(n10426) );
  NAND2_X1 U13295 ( .A1(n10428), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10431) );
  NAND2_X1 U13296 ( .A1(n10429), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10430) );
  INV_X1 U13297 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13663) );
  NAND2_X1 U13298 ( .A1(n12065), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10434) );
  NAND2_X1 U13299 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10433) );
  OAI211_X1 U13300 ( .C1(n12069), .C2(n13663), .A(n10434), .B(n10433), .ZN(
        n10435) );
  NAND2_X1 U13301 ( .A1(n10438), .A2(n10437), .ZN(n10456) );
  INV_X1 U13302 ( .A(n10439), .ZN(n10442) );
  INV_X1 U13303 ( .A(n10440), .ZN(n10441) );
  INV_X1 U13304 ( .A(n10448), .ZN(n10443) );
  NAND2_X1 U13305 ( .A1(n9617), .A2(n10444), .ZN(n10472) );
  OR2_X1 U13306 ( .A1(n12099), .A2(n10472), .ZN(n19377) );
  BUF_X4 U13307 ( .A(n12099), .Z(n13293) );
  INV_X1 U13308 ( .A(n10444), .ZN(n10445) );
  NAND2_X1 U13309 ( .A1(n13293), .A2(n10466), .ZN(n19515) );
  INV_X1 U13310 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10446) );
  OAI22_X1 U13311 ( .A1(n12275), .A2(n19377), .B1(n19515), .B2(n10446), .ZN(
        n10454) );
  INV_X1 U13312 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12283) );
  NAND2_X1 U13313 ( .A1(n16204), .A2(n10456), .ZN(n10449) );
  NOR2_X1 U13314 ( .A1(n9617), .A2(n10449), .ZN(n10470) );
  NAND2_X1 U13315 ( .A1(n13293), .A2(n10470), .ZN(n19443) );
  INV_X1 U13316 ( .A(n10449), .ZN(n10450) );
  NAND2_X1 U13317 ( .A1(n13293), .A2(n10451), .ZN(n19584) );
  INV_X1 U13318 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10452) );
  OAI22_X1 U13319 ( .A1(n12283), .A2(n19443), .B1(n19584), .B2(n10452), .ZN(
        n10453) );
  NOR2_X1 U13320 ( .A1(n10454), .A2(n10453), .ZN(n10464) );
  NAND2_X1 U13321 ( .A1(n10456), .A2(n10455), .ZN(n10457) );
  NAND2_X1 U13322 ( .A1(n14425), .A2(n13351), .ZN(n10458) );
  INV_X1 U13323 ( .A(n10458), .ZN(n10459) );
  AOI22_X1 U13324 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10509), .B1(
        n15381), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10463) );
  INV_X2 U13325 ( .A(n13351), .ZN(n19158) );
  NAND2_X1 U13326 ( .A1(n9617), .A2(n19158), .ZN(n10460) );
  NOR2_X2 U13327 ( .A1(n10478), .A2(n10460), .ZN(n19289) );
  INV_X1 U13328 ( .A(n10460), .ZN(n10461) );
  AOI22_X1 U13329 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19289), .B1(
        n19551), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10462) );
  NAND3_X1 U13330 ( .A1(n10464), .A2(n10463), .A3(n10462), .ZN(n10477) );
  INV_X1 U13331 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10469) );
  OR2_X1 U13332 ( .A1(n12099), .A2(n10465), .ZN(n19319) );
  INV_X1 U13333 ( .A(n10466), .ZN(n10467) );
  INV_X1 U13334 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10468) );
  OAI22_X1 U13335 ( .A1(n10469), .A2(n19319), .B1(n19249), .B2(n10468), .ZN(
        n10475) );
  INV_X1 U13336 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12274) );
  INV_X1 U13337 ( .A(n10470), .ZN(n10471) );
  INV_X1 U13338 ( .A(n10472), .ZN(n10473) );
  NAND2_X1 U13339 ( .A1(n13293), .A2(n10473), .ZN(n13534) );
  OAI22_X1 U13340 ( .A1(n12274), .A2(n10622), .B1(n13534), .B2(n19668), .ZN(
        n10474) );
  NOR2_X1 U13341 ( .A1(n10477), .A2(n10476), .ZN(n10488) );
  INV_X1 U13342 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10480) );
  NAND2_X1 U13343 ( .A1(n10479), .A2(n13351), .ZN(n15352) );
  NAND2_X1 U13344 ( .A1(n10479), .A2(n19158), .ZN(n10630) );
  INV_X1 U13345 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19176) );
  OAI22_X1 U13346 ( .A1(n10480), .A2(n15352), .B1(n10630), .B2(n19176), .ZN(
        n10481) );
  INV_X1 U13347 ( .A(n10481), .ZN(n10487) );
  INV_X1 U13348 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10484) );
  INV_X1 U13349 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12282) );
  OAI22_X1 U13350 ( .A1(n10484), .A2(n19486), .B1(n10629), .B2(n12282), .ZN(
        n10485) );
  INV_X1 U13351 ( .A(n10485), .ZN(n10486) );
  NAND3_X1 U13352 ( .A1(n10488), .A2(n10487), .A3(n10486), .ZN(n10489) );
  NAND2_X1 U13353 ( .A1(n10489), .A2(n15338), .ZN(n10505) );
  AOI22_X1 U13354 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10524), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U13355 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10494) );
  AOI22_X1 U13356 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12186), .ZN(n10493) );
  AOI22_X1 U13357 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10529), .B1(
        n13295), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10492) );
  NAND4_X1 U13358 ( .A1(n10495), .A2(n10494), .A3(n10493), .A4(n10492), .ZN(
        n10503) );
  AOI22_X1 U13359 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__3__SCAN_IN), .B2(n10537), .ZN(n10501) );
  AOI22_X1 U13360 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13361 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13362 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10498) );
  NAND4_X1 U13363 ( .A1(n10501), .A2(n10500), .A3(n10499), .A4(n10498), .ZN(
        n10502) );
  NOR2_X1 U13364 ( .A1(n10503), .A2(n10502), .ZN(n10702) );
  INV_X1 U13365 ( .A(n10702), .ZN(n10839) );
  NAND2_X1 U13366 ( .A1(n10839), .A2(n19852), .ZN(n10504) );
  INV_X1 U13367 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n19658) );
  NAND2_X1 U13368 ( .A1(n15381), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10506) );
  INV_X1 U13369 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10507) );
  INV_X1 U13370 ( .A(n10622), .ZN(n19200) );
  INV_X1 U13371 ( .A(n19515), .ZN(n19512) );
  AOI22_X1 U13372 ( .A1(n19200), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n19512), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10515) );
  NAND2_X1 U13373 ( .A1(n10509), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10514) );
  INV_X1 U13374 ( .A(n19319), .ZN(n19324) );
  INV_X1 U13375 ( .A(n19443), .ZN(n19448) );
  AOI22_X1 U13376 ( .A1(n19324), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n19448), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10513) );
  INV_X1 U13377 ( .A(n19377), .ZN(n10511) );
  INV_X1 U13378 ( .A(n19584), .ZN(n10510) );
  AOI22_X1 U13379 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10510), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10512) );
  INV_X1 U13380 ( .A(n19486), .ZN(n19479) );
  INV_X1 U13381 ( .A(n10629), .ZN(n19412) );
  AOI22_X1 U13382 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19479), .B1(
        n19412), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10520) );
  INV_X1 U13383 ( .A(n10630), .ZN(n15329) );
  INV_X1 U13384 ( .A(n19289), .ZN(n10517) );
  INV_X1 U13385 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12225) );
  INV_X1 U13386 ( .A(n19551), .ZN(n19558) );
  INV_X1 U13387 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10516) );
  AOI21_X1 U13388 ( .B1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n15329), .A(
        n10518), .ZN(n10519) );
  NAND4_X1 U13389 ( .A1(n10522), .A2(n10521), .A3(n10520), .A4(n10519), .ZN(
        n10553) );
  AOI22_X1 U13390 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13391 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U13392 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13393 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10525) );
  NAND4_X1 U13394 ( .A1(n10528), .A2(n10527), .A3(n10526), .A4(n10525), .ZN(
        n10535) );
  AOI22_X1 U13395 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13396 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13397 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13398 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12186), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10530) );
  NAND4_X1 U13399 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n10534) );
  AOI22_X1 U13400 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13401 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12186), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13402 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13403 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10538) );
  NAND4_X1 U13404 ( .A1(n10541), .A2(n10540), .A3(n10539), .A4(n10538), .ZN(
        n10550) );
  AOI22_X1 U13405 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13406 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13407 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13408 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10545) );
  NAND4_X1 U13409 ( .A1(n10548), .A2(n10547), .A3(n10546), .A4(n10545), .ZN(
        n10549) );
  NOR2_X1 U13410 ( .A1(n10818), .A2(n10825), .ZN(n10551) );
  NAND2_X1 U13411 ( .A1(n19852), .A2(n10551), .ZN(n10559) );
  INV_X1 U13412 ( .A(n10833), .ZN(n10558) );
  NAND2_X1 U13413 ( .A1(n10559), .A2(n10558), .ZN(n10552) );
  INV_X1 U13414 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10728) );
  INV_X1 U13415 ( .A(n10818), .ZN(n15004) );
  INV_X1 U13416 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15003) );
  NOR2_X1 U13417 ( .A1(n15004), .A2(n15003), .ZN(n15002) );
  INV_X1 U13418 ( .A(n10825), .ZN(n10555) );
  NAND2_X1 U13419 ( .A1(n15002), .A2(n10555), .ZN(n10557) );
  NOR2_X1 U13420 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15004), .ZN(
        n10556) );
  XOR2_X1 U13421 ( .A(n10825), .B(n10556), .Z(n12887) );
  NAND2_X1 U13422 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12887), .ZN(
        n12886) );
  NAND2_X1 U13423 ( .A1(n10557), .A2(n12886), .ZN(n10560) );
  XNOR2_X1 U13424 ( .A(n10728), .B(n10560), .ZN(n12934) );
  XNOR2_X1 U13425 ( .A(n10559), .B(n10558), .ZN(n12933) );
  NAND2_X1 U13426 ( .A1(n12934), .A2(n12933), .ZN(n10562) );
  NAND2_X1 U13427 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10560), .ZN(
        n10561) );
  NAND2_X1 U13428 ( .A1(n10562), .A2(n10561), .ZN(n10563) );
  INV_X1 U13429 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16195) );
  XNOR2_X1 U13430 ( .A(n10563), .B(n16195), .ZN(n13450) );
  NAND2_X1 U13431 ( .A1(n13449), .A2(n13450), .ZN(n10565) );
  NAND2_X1 U13432 ( .A1(n10563), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10564) );
  NAND2_X1 U13433 ( .A1(n10565), .A2(n10564), .ZN(n10579) );
  NAND2_X1 U13434 ( .A1(n10567), .A2(n10566), .ZN(n10583) );
  AOI22_X1 U13435 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10524), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13436 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13437 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n12186), .ZN(n10569) );
  AOI22_X1 U13438 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10529), .B1(
        n13295), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10568) );
  NAND4_X1 U13439 ( .A1(n10571), .A2(n10570), .A3(n10569), .A4(n10568), .ZN(
        n10578) );
  AOI22_X1 U13440 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .B2(n10537), .ZN(n10576) );
  AOI22_X1 U13441 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10575) );
  AOI22_X1 U13442 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13443 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10573) );
  NAND4_X1 U13444 ( .A1(n10576), .A2(n10575), .A3(n10574), .A4(n10573), .ZN(
        n10577) );
  XNOR2_X1 U13445 ( .A(n10583), .B(n10705), .ZN(n10580) );
  XNOR2_X1 U13446 ( .A(n10579), .B(n10580), .ZN(n13476) );
  INV_X1 U13447 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13475) );
  INV_X1 U13448 ( .A(n10579), .ZN(n10581) );
  NAND2_X1 U13449 ( .A1(n10581), .A2(n10580), .ZN(n10582) );
  AOI22_X1 U13450 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n10509), .B1(
        n19551), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13451 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19289), .B1(
        n15381), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10594) );
  INV_X1 U13452 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10585) );
  INV_X1 U13453 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10584) );
  OAI22_X1 U13454 ( .A1(n10585), .A2(n19249), .B1(n19584), .B2(n10584), .ZN(
        n10587) );
  INV_X1 U13455 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12333) );
  INV_X1 U13456 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12334) );
  OAI22_X1 U13457 ( .A1(n12333), .A2(n19443), .B1(n13534), .B2(n12334), .ZN(
        n10586) );
  NOR2_X1 U13458 ( .A1(n10587), .A2(n10586), .ZN(n10593) );
  INV_X1 U13459 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10588) );
  INV_X1 U13460 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12325) );
  OAI22_X1 U13461 ( .A1(n10588), .A2(n19319), .B1(n19377), .B2(n12325), .ZN(
        n10591) );
  INV_X1 U13462 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12324) );
  INV_X1 U13463 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10589) );
  OAI22_X1 U13464 ( .A1(n12324), .A2(n10622), .B1(n19515), .B2(n10589), .ZN(
        n10590) );
  NOR2_X1 U13465 ( .A1(n10591), .A2(n10590), .ZN(n10592) );
  NAND4_X1 U13466 ( .A1(n10595), .A2(n10594), .A3(n10593), .A4(n10592), .ZN(
        n10600) );
  INV_X1 U13467 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10596) );
  INV_X1 U13468 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12332) );
  OAI22_X1 U13469 ( .A1(n10596), .A2(n15352), .B1(n10629), .B2(n12332), .ZN(
        n10599) );
  INV_X1 U13470 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13121) );
  INV_X1 U13471 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10597) );
  OAI22_X1 U13472 ( .A1(n13121), .A2(n10630), .B1(n19486), .B2(n10597), .ZN(
        n10598) );
  AOI22_X1 U13473 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13474 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U13475 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12186), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13476 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10602) );
  NAND4_X1 U13477 ( .A1(n10605), .A2(n10604), .A3(n10603), .A4(n10602), .ZN(
        n10611) );
  AOI22_X1 U13478 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U13479 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13480 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13481 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10606) );
  NAND4_X1 U13482 ( .A1(n10609), .A2(n10608), .A3(n10607), .A4(n10606), .ZN(
        n10610) );
  NAND2_X1 U13483 ( .A1(n10845), .A2(n19852), .ZN(n10612) );
  XNOR2_X1 U13484 ( .A(n10616), .B(n9609), .ZN(n10734) );
  INV_X1 U13485 ( .A(n10734), .ZN(n10614) );
  INV_X1 U13486 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15308) );
  NAND2_X1 U13487 ( .A1(n10614), .A2(n15308), .ZN(n15300) );
  AOI22_X1 U13488 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19289), .B1(
        n15381), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10628) );
  AOI22_X1 U13489 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10509), .B1(
        n19551), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10627) );
  INV_X1 U13490 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12344) );
  INV_X1 U13491 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12353) );
  OAI22_X1 U13492 ( .A1(n12344), .A2(n19377), .B1(n19443), .B2(n12353), .ZN(
        n10619) );
  INV_X1 U13493 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12345) );
  INV_X1 U13494 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10617) );
  OAI22_X1 U13495 ( .A1(n12345), .A2(n19319), .B1(n19584), .B2(n10617), .ZN(
        n10618) );
  NOR2_X1 U13496 ( .A1(n10619), .A2(n10618), .ZN(n10626) );
  INV_X1 U13497 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10621) );
  INV_X1 U13498 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10620) );
  OAI22_X1 U13499 ( .A1(n10621), .A2(n19249), .B1(n19515), .B2(n10620), .ZN(
        n10624) );
  INV_X1 U13500 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12343) );
  INV_X1 U13501 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12355) );
  OAI22_X1 U13502 ( .A1(n12343), .A2(n10622), .B1(n13534), .B2(n12355), .ZN(
        n10623) );
  NOR2_X1 U13503 ( .A1(n10624), .A2(n10623), .ZN(n10625) );
  NAND4_X1 U13504 ( .A1(n10628), .A2(n10627), .A3(n10626), .A4(n10625), .ZN(
        n10635) );
  INV_X1 U13505 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19198) );
  INV_X1 U13506 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12351) );
  OAI22_X1 U13507 ( .A1(n19198), .A2(n10630), .B1(n10629), .B2(n12351), .ZN(
        n10634) );
  INV_X1 U13508 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10632) );
  INV_X1 U13509 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10631) );
  OAI22_X1 U13510 ( .A1(n10632), .A2(n15352), .B1(n19486), .B2(n10631), .ZN(
        n10633) );
  AOI22_X1 U13511 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10524), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10639) );
  AOI22_X1 U13512 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13513 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n12186), .ZN(n10637) );
  AOI22_X1 U13514 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10529), .B1(
        n13295), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10636) );
  NAND4_X1 U13515 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10636), .ZN(
        n10645) );
  AOI22_X1 U13516 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n10537), .ZN(n10643) );
  AOI22_X1 U13517 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U13518 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10641) );
  AOI22_X1 U13519 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10640) );
  NAND4_X1 U13520 ( .A1(n10643), .A2(n10642), .A3(n10641), .A4(n10640), .ZN(
        n10644) );
  INV_X1 U13521 ( .A(n10849), .ZN(n10646) );
  NAND2_X1 U13522 ( .A1(n10646), .A2(n19852), .ZN(n10647) );
  INV_X1 U13523 ( .A(n15301), .ZN(n15303) );
  NAND2_X1 U13524 ( .A1(n15303), .A2(n9684), .ZN(n10652) );
  NAND2_X1 U13525 ( .A1(n15304), .A2(n15301), .ZN(n10654) );
  NAND2_X1 U13526 ( .A1(n10654), .A2(n10694), .ZN(n10655) );
  AOI22_X1 U13527 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10523), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U13528 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U13529 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n12186), .ZN(n10658) );
  AOI22_X1 U13530 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10529), .B1(
        n13295), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10657) );
  NAND4_X1 U13531 ( .A1(n10660), .A2(n10659), .A3(n10658), .A4(n10657), .ZN(
        n10666) );
  AOI22_X1 U13532 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n10537), .ZN(n10664) );
  AOI22_X1 U13533 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U13534 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13535 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10661) );
  NAND4_X1 U13536 ( .A1(n10664), .A2(n10663), .A3(n10662), .A4(n10661), .ZN(
        n10665) );
  NAND2_X1 U13537 ( .A1(n10656), .A2(n10733), .ZN(n10668) );
  NAND2_X1 U13538 ( .A1(n10672), .A2(n10668), .ZN(n14993) );
  INV_X1 U13539 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10669) );
  INV_X1 U13540 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16176) );
  XNOR2_X1 U13541 ( .A(n10672), .B(n16176), .ZN(n16126) );
  INV_X1 U13542 ( .A(n16126), .ZN(n10670) );
  INV_X1 U13543 ( .A(n10672), .ZN(n10673) );
  NAND2_X1 U13544 ( .A1(n10673), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10674) );
  INV_X1 U13545 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10765) );
  INV_X1 U13546 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10675) );
  NAND2_X1 U13547 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13748) );
  OAI21_X1 U13548 ( .B1(n19162), .B2(n13479), .A(n14921), .ZN(n10685) );
  INV_X1 U13549 ( .A(n13479), .ZN(n10676) );
  NAND2_X1 U13550 ( .A1(n10676), .A2(n10688), .ZN(n19164) );
  NAND2_X1 U13551 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19163) );
  NAND2_X1 U13552 ( .A1(n10728), .A2(n19163), .ZN(n12930) );
  NAND3_X1 U13553 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n12930), .ZN(n10677) );
  NAND2_X1 U13554 ( .A1(n19164), .A2(n10677), .ZN(n10682) );
  INV_X1 U13555 ( .A(n19163), .ZN(n10678) );
  OR2_X1 U13556 ( .A1(n10688), .A2(n10678), .ZN(n10680) );
  INV_X1 U13557 ( .A(n11026), .ZN(n10679) );
  NOR2_X2 U13558 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19806) );
  NAND2_X1 U13559 ( .A1(n19806), .A2(n19844), .ZN(n18788) );
  NAND2_X1 U13560 ( .A1(n10679), .A2(n18966), .ZN(n16197) );
  AND2_X1 U13561 ( .A1(n10680), .A2(n16197), .ZN(n13480) );
  OR2_X1 U13562 ( .A1(n10688), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12932) );
  NAND2_X1 U13563 ( .A1(n13480), .A2(n12932), .ZN(n13477) );
  NOR3_X1 U13564 ( .A1(n13475), .A2(n16195), .A3(n15308), .ZN(n15285) );
  NAND2_X1 U13565 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15285), .ZN(
        n10691) );
  AND2_X1 U13566 ( .A1(n10691), .A2(n19164), .ZN(n15273) );
  NOR2_X1 U13567 ( .A1(n13477), .A2(n15273), .ZN(n10681) );
  NAND2_X1 U13568 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15213) );
  NAND3_X1 U13569 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15210) );
  INV_X1 U13570 ( .A(n15210), .ZN(n15211) );
  NAND2_X1 U13571 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15211), .ZN(
        n10683) );
  NOR2_X1 U13572 ( .A1(n15213), .A2(n10683), .ZN(n13749) );
  INV_X1 U13573 ( .A(n13749), .ZN(n10693) );
  NAND2_X1 U13574 ( .A1(n19164), .A2(n10693), .ZN(n10684) );
  NAND2_X1 U13575 ( .A1(n15257), .A2(n10684), .ZN(n15148) );
  INV_X1 U13576 ( .A(n15148), .ZN(n15201) );
  OAI211_X1 U13577 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n10688), .A(
        n10685), .B(n15201), .ZN(n15185) );
  NOR2_X1 U13578 ( .A1(n16209), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10686) );
  NOR2_X1 U13579 ( .A1(n10728), .A2(n19163), .ZN(n12931) );
  INV_X1 U13580 ( .A(n12931), .ZN(n10687) );
  OR2_X1 U13581 ( .A1(n10688), .A2(n10687), .ZN(n10690) );
  NAND2_X1 U13582 ( .A1(n13479), .A2(n12930), .ZN(n10689) );
  NOR2_X1 U13583 ( .A1(n16196), .A2(n10691), .ZN(n16172) );
  AND2_X1 U13584 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10692) );
  NAND2_X1 U13585 ( .A1(n16172), .A2(n10692), .ZN(n15261) );
  NOR2_X1 U13586 ( .A1(n15261), .A2(n10693), .ZN(n15204) );
  AOI22_X1 U13587 ( .A1(n14909), .A2(n19162), .B1(n9949), .B2(n15204), .ZN(
        n11030) );
  NAND2_X1 U13588 ( .A1(n10694), .A2(n10733), .ZN(n10711) );
  OR2_X1 U13589 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(
        n10695) );
  MUX2_X1 U13590 ( .A(n10825), .B(n10695), .S(n19180), .Z(n10726) );
  MUX2_X1 U13591 ( .A(n10696), .B(n10420), .S(n19180), .Z(n10697) );
  NAND2_X1 U13592 ( .A1(n10755), .A2(n10698), .ZN(n10719) );
  NOR2_X1 U13593 ( .A1(n10698), .A2(n19180), .ZN(n10721) );
  NAND2_X1 U13594 ( .A1(n10721), .A2(n10699), .ZN(n10701) );
  NAND2_X1 U13595 ( .A1(n19180), .A2(n13663), .ZN(n10700) );
  OAI211_X1 U13596 ( .C1(n10702), .C2(n10719), .A(n10701), .B(n10700), .ZN(
        n10712) );
  INV_X1 U13597 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19005) );
  INV_X1 U13598 ( .A(n10703), .ZN(n10704) );
  NAND2_X1 U13599 ( .A1(n10721), .A2(n10704), .ZN(n10708) );
  INV_X1 U13600 ( .A(n10719), .ZN(n10706) );
  NAND2_X1 U13601 ( .A1(n10706), .A2(n10705), .ZN(n10707) );
  OAI211_X1 U13602 ( .C1(n19005), .C2(n10755), .A(n10708), .B(n10707), .ZN(
        n10729) );
  MUX2_X1 U13603 ( .A(n10845), .B(P2_EBX_REG_5__SCAN_IN), .S(n19180), .Z(
        n10735) );
  INV_X1 U13604 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18976) );
  MUX2_X1 U13605 ( .A(n10849), .B(n18976), .S(n19180), .Z(n10709) );
  NOR2_X1 U13606 ( .A1(n10737), .A2(n10709), .ZN(n10710) );
  OR2_X1 U13607 ( .A1(n10749), .A2(n10710), .ZN(n18975) );
  NAND2_X1 U13608 ( .A1(n10711), .A2(n18975), .ZN(n10743) );
  INV_X1 U13609 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15284) );
  INV_X1 U13610 ( .A(n13728), .ZN(n10733) );
  NAND2_X1 U13611 ( .A1(n13449), .A2(n10733), .ZN(n10714) );
  OR2_X1 U13612 ( .A1(n10715), .A2(n10712), .ZN(n10713) );
  NAND2_X1 U13613 ( .A1(n10730), .A2(n10713), .ZN(n13523) );
  INV_X1 U13614 ( .A(n10715), .ZN(n10718) );
  NAND2_X1 U13615 ( .A1(n10726), .A2(n10716), .ZN(n10717) );
  NAND2_X1 U13616 ( .A1(n10718), .A2(n10717), .ZN(n14421) );
  OR2_X1 U13617 ( .A1(n10818), .A2(n10719), .ZN(n10723) );
  AND2_X1 U13618 ( .A1(n19180), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10724) );
  AOI21_X1 U13619 ( .B1(n10721), .B2(n10720), .A(n10724), .ZN(n10722) );
  NAND2_X1 U13620 ( .A1(n10723), .A2(n10722), .ZN(n19025) );
  NAND2_X1 U13621 ( .A1(n19025), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15009) );
  NAND2_X1 U13622 ( .A1(n10724), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10725) );
  NAND2_X1 U13623 ( .A1(n10726), .A2(n10725), .ZN(n13582) );
  NOR2_X1 U13624 ( .A1(n15009), .A2(n13582), .ZN(n10727) );
  NAND2_X1 U13625 ( .A1(n15009), .A2(n13582), .ZN(n12881) );
  OAI21_X1 U13626 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10727), .A(
        n12881), .ZN(n12938) );
  XNOR2_X1 U13627 ( .A(n14421), .B(n10728), .ZN(n12937) );
  OR2_X1 U13628 ( .A1(n12938), .A2(n12937), .ZN(n12935) );
  OAI21_X1 U13629 ( .B1(n14421), .B2(n10728), .A(n12935), .ZN(n13451) );
  XNOR2_X1 U13630 ( .A(n10730), .B(n9991), .ZN(n19003) );
  XNOR2_X1 U13631 ( .A(n19003), .B(n13475), .ZN(n13473) );
  NAND2_X1 U13632 ( .A1(n19003), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10731) );
  NAND2_X1 U13633 ( .A1(n10732), .A2(n10731), .ZN(n15299) );
  NAND2_X1 U13634 ( .A1(n10734), .A2(n10733), .ZN(n10739) );
  AND2_X1 U13635 ( .A1(n10736), .A2(n10735), .ZN(n10738) );
  OR2_X1 U13636 ( .A1(n10738), .A2(n10737), .ZN(n18990) );
  NAND2_X1 U13637 ( .A1(n10739), .A2(n18990), .ZN(n10740) );
  XNOR2_X1 U13638 ( .A(n10740), .B(n15308), .ZN(n15298) );
  NAND2_X1 U13639 ( .A1(n15299), .A2(n15298), .ZN(n10742) );
  NAND2_X1 U13640 ( .A1(n10740), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10741) );
  NAND2_X1 U13641 ( .A1(n10743), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10744) );
  INV_X1 U13642 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10981) );
  MUX2_X1 U13643 ( .A(n13728), .B(n10981), .S(n19180), .Z(n10747) );
  NAND2_X1 U13644 ( .A1(n19180), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10745) );
  OR2_X1 U13645 ( .A1(n10756), .A2(n10745), .ZN(n10746) );
  NAND2_X1 U13646 ( .A1(n10750), .A2(n10746), .ZN(n18953) );
  NOR2_X1 U13647 ( .A1(n18953), .A2(n10733), .ZN(n10753) );
  NAND2_X1 U13648 ( .A1(n10753), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16132) );
  INV_X1 U13649 ( .A(n10747), .ZN(n10748) );
  XNOR2_X1 U13650 ( .A(n10749), .B(n10748), .ZN(n18965) );
  NAND2_X1 U13651 ( .A1(n18965), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16127) );
  NAND2_X1 U13652 ( .A1(n19180), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10751) );
  MUX2_X1 U13653 ( .A(n19180), .B(n10751), .S(n10750), .Z(n10752) );
  NAND2_X1 U13654 ( .A1(n9995), .A2(n10752), .ZN(n18941) );
  NAND2_X1 U13655 ( .A1(n10767), .A2(n14587), .ZN(n15262) );
  INV_X1 U13656 ( .A(n10753), .ZN(n10754) );
  NAND2_X1 U13657 ( .A1(n10754), .A2(n16176), .ZN(n16131) );
  OR2_X1 U13658 ( .A1(n18965), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16129) );
  AND2_X1 U13659 ( .A1(n16131), .A2(n16129), .ZN(n14980) );
  INV_X1 U13660 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19069) );
  NAND2_X1 U13661 ( .A1(n10762), .A2(n19069), .ZN(n10760) );
  NOR2_X1 U13662 ( .A1(n10762), .A2(n19069), .ZN(n10757) );
  NAND2_X1 U13663 ( .A1(n19180), .A2(n10757), .ZN(n10758) );
  AND2_X1 U13664 ( .A1(n13712), .A2(n10758), .ZN(n10759) );
  NAND2_X1 U13665 ( .A1(n10760), .A2(n10759), .ZN(n18933) );
  OR2_X1 U13666 ( .A1(n18933), .A2(n10733), .ZN(n10761) );
  INV_X1 U13667 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15245) );
  NAND2_X1 U13668 ( .A1(n10761), .A2(n15245), .ZN(n16107) );
  INV_X1 U13669 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13244) );
  AND3_X1 U13670 ( .A1(n19180), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10760), .ZN(
        n10764) );
  OR2_X1 U13671 ( .A1(n10773), .A2(n10764), .ZN(n18921) );
  OAI21_X1 U13672 ( .B1(n18921), .B2(n10733), .A(n10765), .ZN(n14985) );
  AND4_X1 U13673 ( .A1(n15262), .A2(n14980), .A3(n16107), .A4(n14985), .ZN(
        n10766) );
  INV_X1 U13674 ( .A(n10767), .ZN(n10768) );
  NAND2_X1 U13675 ( .A1(n10768), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16108) );
  NAND2_X1 U13676 ( .A1(n13728), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10769) );
  OR2_X1 U13677 ( .A1(n18921), .A2(n10769), .ZN(n14984) );
  AND3_X1 U13678 ( .A1(n16108), .A2(n14984), .A3(n16106), .ZN(n10770) );
  NAND2_X1 U13679 ( .A1(n19180), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10772) );
  NAND3_X1 U13680 ( .A1(n19180), .A2(n10774), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n10775) );
  AND2_X1 U13681 ( .A1(n10782), .A2(n10775), .ZN(n18912) );
  NAND2_X1 U13682 ( .A1(n18912), .A2(n13728), .ZN(n14964) );
  INV_X1 U13683 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14968) );
  NOR2_X1 U13684 ( .A1(n14964), .A2(n14968), .ZN(n10777) );
  NAND2_X1 U13685 ( .A1(n14964), .A2(n14968), .ZN(n10776) );
  AND2_X1 U13686 ( .A1(n19180), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10781) );
  INV_X1 U13687 ( .A(n10781), .ZN(n10778) );
  XNOR2_X1 U13688 ( .A(n10782), .B(n10778), .ZN(n18904) );
  AOI21_X1 U13689 ( .B1(n18904), .B2(n13728), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14954) );
  AND2_X1 U13690 ( .A1(n13728), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10779) );
  NAND2_X1 U13691 ( .A1(n18904), .A2(n10779), .ZN(n14952) );
  NAND2_X1 U13692 ( .A1(n10780), .A2(n14952), .ZN(n14942) );
  NAND2_X1 U13693 ( .A1(n19180), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10783) );
  MUX2_X1 U13694 ( .A(n19180), .B(n10783), .S(n10790), .Z(n10784) );
  OR2_X1 U13695 ( .A1(n10790), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10788) );
  NAND2_X1 U13696 ( .A1(n10784), .A2(n10788), .ZN(n18891) );
  INV_X1 U13697 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15219) );
  OAI21_X1 U13698 ( .B1(n18891), .B2(n10733), .A(n15219), .ZN(n14940) );
  NAND2_X1 U13699 ( .A1(n14942), .A2(n14940), .ZN(n14929) );
  INV_X1 U13700 ( .A(n18891), .ZN(n10786) );
  AND2_X1 U13701 ( .A1(n13728), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10785) );
  NAND2_X1 U13702 ( .A1(n10786), .A2(n10785), .ZN(n14939) );
  AND2_X1 U13703 ( .A1(n19180), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10787) );
  NAND2_X1 U13704 ( .A1(n10788), .A2(n10787), .ZN(n10791) );
  INV_X1 U13705 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11006) );
  INV_X1 U13706 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11010) );
  NAND2_X1 U13707 ( .A1(n11006), .A2(n11010), .ZN(n10789) );
  NAND2_X1 U13708 ( .A1(n10791), .A2(n10798), .ZN(n18879) );
  INV_X1 U13709 ( .A(n18879), .ZN(n10793) );
  AND2_X1 U13710 ( .A1(n13728), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10792) );
  NAND2_X1 U13711 ( .A1(n10793), .A2(n10792), .ZN(n14930) );
  AND2_X1 U13712 ( .A1(n14939), .A2(n14930), .ZN(n13691) );
  INV_X1 U13713 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15203) );
  OAI21_X1 U13714 ( .B1(n18879), .B2(n10733), .A(n15203), .ZN(n14931) );
  INV_X1 U13715 ( .A(n14931), .ZN(n10794) );
  INV_X1 U13716 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10795) );
  AND2_X1 U13717 ( .A1(n19180), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10797) );
  INV_X1 U13718 ( .A(n13712), .ZN(n10796) );
  AOI21_X1 U13719 ( .B1(n10798), .B2(n10797), .A(n10796), .ZN(n10799) );
  NAND2_X1 U13720 ( .A1(n10802), .A2(n10799), .ZN(n18872) );
  OR2_X1 U13721 ( .A1(n18872), .A2(n10733), .ZN(n10800) );
  XNOR2_X1 U13722 ( .A(n10800), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14918) );
  NAND2_X1 U13723 ( .A1(n14919), .A2(n14918), .ZN(n14917) );
  NAND2_X1 U13724 ( .A1(n13728), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10801) );
  OR2_X1 U13725 ( .A1(n18872), .A2(n10801), .ZN(n13690) );
  NAND2_X1 U13726 ( .A1(n14917), .A2(n13690), .ZN(n14852) );
  NAND2_X1 U13727 ( .A1(n19180), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10803) );
  OR2_X1 U13728 ( .A1(n10804), .A2(n10803), .ZN(n10805) );
  NAND2_X1 U13729 ( .A1(n10805), .A2(n13679), .ZN(n18861) );
  OAI21_X1 U13730 ( .B1(n18861), .B2(n10733), .A(n11033), .ZN(n14850) );
  INV_X1 U13731 ( .A(n18861), .ZN(n10807) );
  AND2_X1 U13732 ( .A1(n13728), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10806) );
  NAND2_X1 U13733 ( .A1(n10807), .A2(n10806), .ZN(n13692) );
  NAND2_X1 U13734 ( .A1(n14850), .A2(n13692), .ZN(n14851) );
  XNOR2_X1 U13735 ( .A(n14852), .B(n14851), .ZN(n14914) );
  NOR2_X1 U13736 ( .A1(n10374), .A2(n10808), .ZN(n19838) );
  NAND2_X2 U13737 ( .A1(n14510), .A2(n10812), .ZN(n10870) );
  INV_X1 U13738 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10972) );
  NOR2_X1 U13739 ( .A1(n12900), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10810) );
  AND2_X2 U13740 ( .A1(n15338), .A2(n19587), .ZN(n10823) );
  AOI22_X1 U13741 ( .A1(n13756), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n10823), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10815) );
  NAND2_X1 U13742 ( .A1(n10817), .A2(n10813), .ZN(n10814) );
  OAI211_X1 U13743 ( .C1(n10870), .C2(n10972), .A(n10815), .B(n10814), .ZN(
        n13386) );
  INV_X1 U13744 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19733) );
  AOI22_X1 U13745 ( .A1(n13756), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10823), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10816) );
  OAI21_X1 U13746 ( .B1(n10870), .B2(n19733), .A(n10816), .ZN(n12926) );
  INV_X1 U13747 ( .A(n10817), .ZN(n10955) );
  MUX2_X1 U13748 ( .A(n12900), .B(n19830), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10820) );
  INV_X1 U13749 ( .A(n10349), .ZN(n10819) );
  NAND2_X1 U13750 ( .A1(n10819), .A2(n10823), .ZN(n10834) );
  INV_X1 U13751 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19024) );
  AOI21_X1 U13752 ( .B1(n15338), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10822) );
  NAND2_X1 U13753 ( .A1(n15345), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10821) );
  OAI211_X1 U13754 ( .C1(n10870), .C2(n19024), .A(n10822), .B(n10821), .ZN(
        n12958) );
  INV_X1 U13755 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19731) );
  AOI22_X1 U13756 ( .A1(n10810), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10823), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10824) );
  OAI21_X1 U13757 ( .B1(n10870), .B2(n19731), .A(n10824), .ZN(n10829) );
  OR2_X1 U13758 ( .A1(n10825), .A2(n10955), .ZN(n10828) );
  NAND2_X1 U13759 ( .A1(n10349), .A2(n12900), .ZN(n10826) );
  MUX2_X1 U13760 ( .A(n10826), .B(n19821), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10827) );
  NAND2_X1 U13761 ( .A1(n10828), .A2(n10827), .ZN(n13065) );
  NOR2_X1 U13762 ( .A1(n13066), .A2(n13065), .ZN(n10832) );
  NOR2_X1 U13763 ( .A1(n10830), .A2(n10829), .ZN(n10831) );
  NAND2_X1 U13764 ( .A1(n10817), .A2(n10833), .ZN(n10835) );
  OAI211_X1 U13765 ( .C1(n19587), .C2(n19813), .A(n10835), .B(n10834), .ZN(
        n10836) );
  XNOR2_X1 U13766 ( .A(n10837), .B(n10836), .ZN(n12927) );
  NOR2_X1 U13767 ( .A1(n12926), .A2(n12927), .ZN(n12928) );
  NOR2_X1 U13768 ( .A1(n10837), .A2(n10836), .ZN(n10838) );
  NAND2_X1 U13769 ( .A1(n10817), .A2(n10839), .ZN(n10841) );
  NAND2_X1 U13770 ( .A1(n13756), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10840) );
  NAND2_X1 U13771 ( .A1(n10841), .A2(n10840), .ZN(n10844) );
  INV_X1 U13772 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13454) );
  AOI22_X1 U13773 ( .A1(n10823), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10842) );
  OAI21_X1 U13774 ( .B1(n10870), .B2(n13454), .A(n10842), .ZN(n10843) );
  INV_X1 U13775 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n15310) );
  AOI22_X1 U13776 ( .A1(n13756), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n10823), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10848) );
  INV_X1 U13777 ( .A(n10845), .ZN(n10846) );
  NAND2_X1 U13778 ( .A1(n10817), .A2(n10846), .ZN(n10847) );
  OAI211_X1 U13779 ( .C1(n10870), .C2(n15310), .A(n10848), .B(n10847), .ZN(
        n15307) );
  NAND2_X1 U13780 ( .A1(n10817), .A2(n10849), .ZN(n10850) );
  INV_X1 U13781 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19737) );
  AOI22_X1 U13782 ( .A1(n13756), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n10823), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10852) );
  OAI21_X1 U13783 ( .B1(n10870), .B2(n19737), .A(n10852), .ZN(n12898) );
  NAND2_X1 U13784 ( .A1(n12899), .A2(n12898), .ZN(n10854) );
  NAND2_X1 U13785 ( .A1(n10817), .A2(n13728), .ZN(n10853) );
  INV_X1 U13786 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19739) );
  AOI22_X1 U13787 ( .A1(n13756), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n10823), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10855) );
  OAI21_X1 U13788 ( .B1(n10870), .B2(n19739), .A(n10855), .ZN(n12946) );
  INV_X1 U13789 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U13790 ( .A1(n13756), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10823), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13791 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10536), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U13792 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13793 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12186), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13794 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10856) );
  NAND4_X1 U13795 ( .A1(n10859), .A2(n10858), .A3(n10857), .A4(n10856), .ZN(
        n10865) );
  AOI22_X1 U13796 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U13797 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U13798 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10861) );
  AOI22_X1 U13799 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10860) );
  NAND4_X1 U13800 ( .A1(n10863), .A2(n10862), .A3(n10861), .A4(n10860), .ZN(
        n10864) );
  NAND2_X1 U13801 ( .A1(n10817), .A2(n19071), .ZN(n10866) );
  OAI211_X1 U13802 ( .C1(n10870), .C2(n10868), .A(n10867), .B(n10866), .ZN(
        n13011) );
  INV_X1 U13803 ( .A(n13011), .ZN(n10869) );
  AOI22_X1 U13804 ( .A1(n11999), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10882) );
  AOI22_X1 U13805 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10874) );
  AOI22_X1 U13806 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U13807 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12186), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U13808 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10871) );
  NAND4_X1 U13809 ( .A1(n10874), .A2(n10873), .A3(n10872), .A4(n10871), .ZN(
        n10880) );
  AOI22_X1 U13810 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U13811 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U13812 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U13813 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10875) );
  NAND4_X1 U13814 ( .A1(n10878), .A2(n10877), .A3(n10876), .A4(n10875), .ZN(
        n10879) );
  AOI22_X1 U13815 ( .A1(n10817), .A2(n19062), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n13756), .ZN(n10881) );
  NAND2_X1 U13816 ( .A1(n10882), .A2(n10881), .ZN(n13024) );
  INV_X1 U13817 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13818 ( .A1(n13756), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U13819 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10523), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U13820 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U13821 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n12186), .ZN(n10884) );
  AOI22_X1 U13822 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10529), .B1(
        n13295), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10883) );
  NAND4_X1 U13823 ( .A1(n10886), .A2(n10885), .A3(n10884), .A4(n10883), .ZN(
        n10892) );
  AOI22_X1 U13824 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n10542), .ZN(n10890) );
  AOI22_X1 U13825 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10544), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U13826 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10888) );
  AOI22_X1 U13827 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10543), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10887) );
  NAND4_X1 U13828 ( .A1(n10890), .A2(n10889), .A3(n10888), .A4(n10887), .ZN(
        n10891) );
  NAND2_X1 U13829 ( .A1(n10817), .A2(n19061), .ZN(n10893) );
  OAI211_X1 U13830 ( .C1(n10870), .C2(n10895), .A(n10894), .B(n10893), .ZN(
        n13026) );
  INV_X1 U13831 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19745) );
  AOI22_X1 U13832 ( .A1(n13756), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U13833 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10524), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U13834 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U13835 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n12186), .ZN(n10897) );
  AOI22_X1 U13836 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10529), .B1(
        n13295), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10896) );
  NAND4_X1 U13837 ( .A1(n10899), .A2(n10898), .A3(n10897), .A4(n10896), .ZN(
        n10905) );
  AOI22_X1 U13838 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__3__SCAN_IN), .B2(n10537), .ZN(n10903) );
  AOI22_X1 U13839 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U13840 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U13841 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10900) );
  NAND4_X1 U13842 ( .A1(n10903), .A2(n10902), .A3(n10901), .A4(n10900), .ZN(
        n10904) );
  NOR2_X1 U13843 ( .A1(n10905), .A2(n10904), .ZN(n13245) );
  OR2_X1 U13844 ( .A1(n10955), .A2(n13245), .ZN(n10906) );
  OAI211_X1 U13845 ( .C1(n10870), .C2(n19745), .A(n10907), .B(n10906), .ZN(
        n13074) );
  INV_X1 U13846 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n14973) );
  AOI22_X1 U13847 ( .A1(n13756), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10919) );
  AOI22_X1 U13848 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13849 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13850 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12186), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13851 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10529), .B1(
        n13295), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10908) );
  NAND4_X1 U13852 ( .A1(n10911), .A2(n10910), .A3(n10909), .A4(n10908), .ZN(
        n10917) );
  AOI22_X1 U13853 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n10542), .ZN(n10915) );
  AOI22_X1 U13854 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U13855 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U13856 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10544), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10912) );
  NAND4_X1 U13857 ( .A1(n10915), .A2(n10914), .A3(n10913), .A4(n10912), .ZN(
        n10916) );
  NAND2_X1 U13858 ( .A1(n10817), .A2(n19053), .ZN(n10918) );
  OAI211_X1 U13859 ( .C1(n10870), .C2(n14973), .A(n10919), .B(n10918), .ZN(
        n13146) );
  INV_X1 U13860 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n14957) );
  AOI22_X1 U13861 ( .A1(n13756), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10931) );
  AOI22_X1 U13862 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U13863 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U13864 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12186), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U13865 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10920) );
  NAND4_X1 U13866 ( .A1(n10923), .A2(n10922), .A3(n10921), .A4(n10920), .ZN(
        n10929) );
  AOI22_X1 U13867 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U13868 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U13869 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U13870 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10924) );
  NAND4_X1 U13871 ( .A1(n10927), .A2(n10926), .A3(n10925), .A4(n10924), .ZN(
        n10928) );
  NAND2_X1 U13872 ( .A1(n10817), .A2(n13290), .ZN(n10930) );
  OAI211_X1 U13873 ( .C1(n10870), .C2(n14957), .A(n10931), .B(n10930), .ZN(
        n13164) );
  INV_X1 U13874 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n14945) );
  AOI22_X1 U13875 ( .A1(n13756), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U13876 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U13877 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U13878 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12186), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U13879 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10529), .B1(
        n13295), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10932) );
  NAND4_X1 U13880 ( .A1(n10935), .A2(n10934), .A3(n10933), .A4(n10932), .ZN(
        n10941) );
  AOI22_X1 U13881 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n10544), .ZN(n10939) );
  AOI22_X1 U13882 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13883 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13884 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10936) );
  NAND4_X1 U13885 ( .A1(n10939), .A2(n10938), .A3(n10937), .A4(n10936), .ZN(
        n10940) );
  NOR2_X1 U13886 ( .A1(n10941), .A2(n10940), .ZN(n19049) );
  OR2_X1 U13887 ( .A1(n10955), .A2(n19049), .ZN(n10942) );
  OAI211_X1 U13888 ( .C1(n10870), .C2(n14945), .A(n10943), .B(n10942), .ZN(
        n10944) );
  INV_X1 U13889 ( .A(n10944), .ZN(n13220) );
  INV_X1 U13890 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19750) );
  AOI22_X1 U13891 ( .A1(n13756), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U13892 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n10524), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U13893 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13894 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12186), .ZN(n10946) );
  AOI22_X1 U13895 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10529), .B1(
        n13295), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10945) );
  NAND4_X1 U13896 ( .A1(n10948), .A2(n10947), .A3(n10946), .A4(n10945), .ZN(
        n10954) );
  AOI22_X1 U13897 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n10537), .ZN(n10952) );
  AOI22_X1 U13898 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U13899 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U13900 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10949) );
  NAND4_X1 U13901 ( .A1(n10952), .A2(n10951), .A3(n10950), .A4(n10949), .ZN(
        n10953) );
  NOR2_X1 U13902 ( .A1(n10954), .A2(n10953), .ZN(n13460) );
  OR2_X1 U13903 ( .A1(n10955), .A2(n13460), .ZN(n10956) );
  OAI211_X1 U13904 ( .C1(n10870), .C2(n19750), .A(n10957), .B(n10956), .ZN(
        n13238) );
  INV_X1 U13905 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U13906 ( .A1(n13756), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10958) );
  OAI21_X1 U13907 ( .B1(n10870), .B2(n11014), .A(n10958), .ZN(n15186) );
  INV_X1 U13908 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19753) );
  AOI22_X1 U13909 ( .A1(n13756), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10959) );
  OAI21_X1 U13910 ( .B1(n10870), .B2(n19753), .A(n10959), .ZN(n10960) );
  OAI21_X1 U13911 ( .B1(n9686), .B2(n10960), .A(n15171), .ZN(n18869) );
  NAND2_X1 U13912 ( .A1(n16215), .A2(n15492), .ZN(n13340) );
  INV_X1 U13913 ( .A(n13340), .ZN(n10962) );
  OR2_X1 U13914 ( .A1(n10961), .A2(n13345), .ZN(n13299) );
  OAI21_X1 U13915 ( .B1(n19852), .B2(n10962), .A(n13299), .ZN(n10963) );
  INV_X1 U13916 ( .A(n10964), .ZN(n10965) );
  NOR2_X1 U13917 ( .A1(n10966), .A2(n10965), .ZN(n10967) );
  NAND2_X1 U13918 ( .A1(n13743), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10971) );
  AOI22_X1 U13919 ( .A1(n13739), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10970) );
  OAI211_X1 U13920 ( .C1(n13741), .C2(n10972), .A(n10971), .B(n10970), .ZN(
        n13484) );
  NAND2_X1 U13921 ( .A1(n13743), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10974) );
  AOI22_X1 U13922 ( .A1(n13739), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10973) );
  OAI211_X1 U13923 ( .C1(n13741), .C2(n15310), .A(n10974), .B(n10973), .ZN(
        n13116) );
  NAND2_X1 U13924 ( .A1(n12065), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U13925 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10975) );
  OAI211_X1 U13926 ( .C1(n12069), .C2(n18976), .A(n10976), .B(n10975), .ZN(
        n10977) );
  AOI21_X1 U13927 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10977), .ZN(n13124) );
  INV_X1 U13928 ( .A(n13124), .ZN(n10978) );
  NAND2_X1 U13929 ( .A1(n12065), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10980) );
  NAND2_X1 U13930 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10979) );
  OAI211_X1 U13931 ( .C1(n10981), .C2(n12069), .A(n10980), .B(n10979), .ZN(
        n10982) );
  AOI21_X1 U13932 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10982), .ZN(n13141) );
  AOI22_X1 U13933 ( .A1(n13739), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10984) );
  NAND2_X1 U13934 ( .A1(n12065), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10983) );
  OAI211_X1 U13935 ( .C1(n10985), .C2(n16176), .A(n10984), .B(n10983), .ZN(
        n16136) );
  NAND2_X1 U13936 ( .A1(n13743), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10991) );
  INV_X1 U13937 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10988) );
  NAND2_X1 U13938 ( .A1(n12065), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10987) );
  NAND2_X1 U13939 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10986) );
  OAI211_X1 U13940 ( .C1(n12069), .C2(n10988), .A(n10987), .B(n10986), .ZN(
        n10989) );
  INV_X1 U13941 ( .A(n10989), .ZN(n10990) );
  NAND2_X1 U13942 ( .A1(n12065), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10993) );
  NAND2_X1 U13943 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10992) );
  OAI211_X1 U13944 ( .C1(n12069), .C2(n19069), .A(n10993), .B(n10992), .ZN(
        n10994) );
  AOI21_X1 U13945 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n10994), .ZN(n16102) );
  NAND2_X1 U13946 ( .A1(n12065), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10996) );
  NAND2_X1 U13947 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10995) );
  OAI211_X1 U13948 ( .C1(n12069), .C2(n13244), .A(n10996), .B(n10995), .ZN(
        n10997) );
  AOI21_X1 U13949 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10997), .ZN(n13242) );
  NAND2_X1 U13950 ( .A1(n13743), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10999) );
  AOI22_X1 U13951 ( .A1(n13739), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10998) );
  OAI211_X1 U13952 ( .C1(n13741), .C2(n14973), .A(n10999), .B(n10998), .ZN(
        n14969) );
  INV_X1 U13953 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11002) );
  NAND2_X1 U13954 ( .A1(n12065), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11001) );
  NAND2_X1 U13955 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11000) );
  OAI211_X1 U13956 ( .C1(n12069), .C2(n11002), .A(n11001), .B(n11000), .ZN(
        n11003) );
  AOI21_X1 U13957 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11003), .ZN(n13288) );
  NAND2_X1 U13958 ( .A1(n12065), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11005) );
  NAND2_X1 U13959 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11004) );
  OAI211_X1 U13960 ( .C1(n11006), .C2(n12069), .A(n11005), .B(n11004), .ZN(
        n11007) );
  AOI21_X1 U13961 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11007), .ZN(n14943) );
  NAND2_X1 U13962 ( .A1(n12065), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11009) );
  NAND2_X1 U13963 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11008) );
  OAI211_X1 U13964 ( .C1(n12069), .C2(n11010), .A(n11009), .B(n11008), .ZN(
        n11011) );
  AOI21_X1 U13965 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11011), .ZN(n13464) );
  NAND2_X1 U13966 ( .A1(n13743), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11013) );
  AOI22_X1 U13967 ( .A1(n13739), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11012) );
  OAI211_X1 U13968 ( .C1(n13741), .C2(n11014), .A(n11013), .B(n11012), .ZN(
        n14922) );
  INV_X1 U13969 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11017) );
  NAND2_X1 U13970 ( .A1(n12065), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11016) );
  NAND2_X1 U13971 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11015) );
  OAI211_X1 U13972 ( .C1(n12069), .C2(n11017), .A(n11016), .B(n11015), .ZN(
        n11018) );
  AOI21_X1 U13973 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11018), .ZN(n11020) );
  NAND2_X1 U13974 ( .A1(n11019), .A2(n11020), .ZN(n11021) );
  AND2_X1 U13975 ( .A1(n14901), .A2(n11021), .ZN(n18863) );
  NAND2_X1 U13976 ( .A1(n11022), .A2(n19852), .ZN(n11024) );
  NAND2_X1 U13977 ( .A1(n11024), .A2(n11023), .ZN(n11025) );
  NAND2_X1 U13978 ( .A1(n11026), .A2(n11025), .ZN(n19157) );
  NOR2_X1 U13979 ( .A1(n18966), .A2(n19753), .ZN(n14910) );
  AOI21_X1 U13980 ( .B1(n18863), .B2(n16203), .A(n14910), .ZN(n11027) );
  OAI21_X1 U13981 ( .B1(n18869), .B2(n16184), .A(n11027), .ZN(n11028) );
  AOI21_X1 U13982 ( .B1(n14914), .B2(n16200), .A(n11028), .ZN(n11029) );
  INV_X1 U13983 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11035) );
  NOR2_X4 U13984 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13185) );
  AOI22_X1 U13985 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U13986 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11329), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11041) );
  INV_X1 U13987 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U13988 ( .A1(n11138), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11040) );
  AND2_X2 U13989 ( .A1(n11044), .A2(n13185), .ZN(n11089) );
  AOI22_X1 U13990 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11039) );
  NAND4_X1 U13991 ( .A1(n11042), .A2(n11041), .A3(n11040), .A4(n11039), .ZN(
        n11051) );
  NOR2_X4 U13992 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13203) );
  AOI22_X1 U13993 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11191), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11049) );
  AND2_X4 U13994 ( .A1(n13186), .A2(n13203), .ZN(n11733) );
  AOI22_X1 U13995 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11048) );
  AND2_X4 U13996 ( .A1(n13203), .A2(n13185), .ZN(n11694) );
  AOI22_X1 U13997 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U13998 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11186), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11046) );
  NAND4_X1 U13999 ( .A1(n11049), .A2(n11048), .A3(n11047), .A4(n11046), .ZN(
        n11050) );
  AOI22_X1 U14000 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14001 ( .A1(n11329), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11186), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14002 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11138), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14003 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11052) );
  NAND4_X1 U14004 ( .A1(n11055), .A2(n11054), .A3(n11053), .A4(n11052), .ZN(
        n11061) );
  AOI22_X1 U14005 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U14006 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14007 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U14008 ( .A1(n11191), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11056) );
  NAND4_X1 U14009 ( .A1(n11059), .A2(n11058), .A3(n11057), .A4(n11056), .ZN(
        n11060) );
  NOR2_X1 U14010 ( .A1(n11061), .A2(n11060), .ZN(n11153) );
  NAND2_X1 U14011 ( .A1(n11287), .A2(n11153), .ZN(n11147) );
  AOI22_X1 U14012 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U14013 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U14014 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U14015 ( .A1(n11191), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11062) );
  NAND4_X1 U14016 ( .A1(n11065), .A2(n11064), .A3(n11063), .A4(n11062), .ZN(
        n11072) );
  AOI22_X1 U14017 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11138), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14018 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U14019 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11067) );
  NAND4_X1 U14020 ( .A1(n11070), .A2(n11069), .A3(n11068), .A4(n11067), .ZN(
        n11071) );
  AOI22_X1 U14021 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11138), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U14022 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U14023 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11075) );
  AOI22_X1 U14024 ( .A1(n11329), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11186), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U14025 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11081) );
  AOI22_X1 U14026 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U14027 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11079) );
  AOI22_X1 U14028 ( .A1(n11191), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11078) );
  NAND2_X2 U14029 ( .A1(n11083), .A2(n11082), .ZN(n20182) );
  NAND2_X2 U14030 ( .A1(n11287), .A2(n20182), .ZN(n11152) );
  AOI22_X1 U14031 ( .A1(n11186), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U14032 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11138), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U14033 ( .A1(n11191), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U14034 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11085) );
  NAND4_X1 U14035 ( .A1(n11088), .A2(n11087), .A3(n11086), .A4(n11085), .ZN(
        n11095) );
  AOI22_X1 U14036 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11093) );
  AOI22_X1 U14037 ( .A1(n11329), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11089), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11092) );
  AOI22_X1 U14038 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11207), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U14039 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11090) );
  NAND4_X1 U14040 ( .A1(n11093), .A2(n11092), .A3(n11091), .A4(n11090), .ZN(
        n11094) );
  OR2_X2 U14041 ( .A1(n11095), .A2(n11094), .ZN(n12906) );
  NAND2_X1 U14042 ( .A1(n11152), .A2(n12906), .ZN(n11169) );
  NAND2_X1 U14043 ( .A1(n11152), .A2(n20182), .ZN(n11108) );
  AND2_X2 U14044 ( .A1(n20182), .A2(n11153), .ZN(n12901) );
  AOI22_X1 U14045 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11138), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14046 ( .A1(n11329), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11186), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14047 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14048 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11096) );
  NAND4_X1 U14049 ( .A1(n11099), .A2(n11098), .A3(n11097), .A4(n11096), .ZN(
        n11107) );
  AOI22_X1 U14050 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11105) );
  AOI22_X1 U14051 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U14052 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11103) );
  AND2_X1 U14053 ( .A1(n11694), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11101) );
  AOI21_X1 U14054 ( .B1(n11191), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n11101), .ZN(n11102) );
  NAND4_X1 U14055 ( .A1(n11105), .A2(n11104), .A3(n11103), .A4(n11102), .ZN(
        n11106) );
  MUX2_X1 U14056 ( .A(n11108), .B(n12901), .S(n20162), .Z(n11109) );
  AOI22_X1 U14057 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U14058 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U14059 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14060 ( .A1(n11191), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11111) );
  NAND4_X1 U14061 ( .A1(n11114), .A2(n11113), .A3(n11112), .A4(n11111), .ZN(
        n11121) );
  AOI22_X1 U14062 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11138), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U14063 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11117) );
  AOI22_X1 U14064 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11116) );
  NAND4_X1 U14065 ( .A1(n11119), .A2(n11118), .A3(n11117), .A4(n11116), .ZN(
        n11120) );
  NAND2_X1 U14066 ( .A1(n11123), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11127) );
  NAND2_X1 U14067 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11126) );
  NAND2_X1 U14068 ( .A1(n11191), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11125) );
  NAND2_X1 U14069 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11124) );
  NAND2_X1 U14070 ( .A1(n11186), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11132) );
  NAND2_X1 U14071 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11131) );
  NAND2_X1 U14072 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11130) );
  NAND2_X1 U14073 ( .A1(n11084), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11129) );
  NAND2_X1 U14074 ( .A1(n11100), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11137) );
  NAND2_X1 U14075 ( .A1(n11329), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11136) );
  NAND2_X1 U14076 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11135) );
  NAND2_X1 U14077 ( .A1(n11133), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14078 ( .A1(n11138), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11142) );
  NAND2_X1 U14079 ( .A1(n11207), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11141) );
  NAND2_X1 U14080 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11140) );
  NAND2_X1 U14081 ( .A1(n11115), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11139) );
  INV_X1 U14082 ( .A(n13029), .ZN(n11151) );
  NAND2_X1 U14083 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20765) );
  OAI21_X1 U14084 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20765), .ZN(n12915) );
  INV_X1 U14085 ( .A(n12915), .ZN(n11149) );
  NAND2_X1 U14086 ( .A1(n12849), .A2(n11149), .ZN(n11150) );
  NAND2_X1 U14087 ( .A1(n11154), .A2(n20188), .ZN(n13154) );
  NAND2_X1 U14088 ( .A1(n11152), .A2(n13054), .ZN(n11157) );
  NAND2_X1 U14089 ( .A1(n12971), .A2(n20188), .ZN(n11155) );
  AND2_X2 U14090 ( .A1(n12906), .A2(n9614), .ZN(n11170) );
  NAND2_X1 U14091 ( .A1(n11161), .A2(n15548), .ZN(n11162) );
  NAND2_X1 U14092 ( .A1(n11162), .A2(n20146), .ZN(n11180) );
  INV_X1 U14093 ( .A(n20529), .ZN(n20685) );
  NAND2_X1 U14094 ( .A1(n20689), .A2(n20611), .ZN(n20564) );
  AND2_X1 U14095 ( .A1(n20685), .A2(n20564), .ZN(n20482) );
  NAND2_X1 U14096 ( .A1(n20482), .A2(n11833), .ZN(n11165) );
  INV_X1 U14097 ( .A(n15551), .ZN(n11164) );
  NAND2_X1 U14098 ( .A1(n11164), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11240) );
  INV_X1 U14099 ( .A(n20267), .ZN(n11184) );
  INV_X1 U14100 ( .A(n11833), .ZN(n11167) );
  MUX2_X1 U14101 ( .A(n15551), .B(n11167), .S(n20611), .Z(n11168) );
  INV_X1 U14102 ( .A(n14406), .ZN(n11182) );
  NAND2_X1 U14103 ( .A1(n12973), .A2(n9614), .ZN(n11181) );
  INV_X1 U14104 ( .A(n11169), .ZN(n11173) );
  OR2_X1 U14105 ( .A1(n11170), .A2(n11171), .ZN(n12872) );
  OAI22_X1 U14106 ( .A1(n11173), .A2(n12872), .B1(n11778), .B2(n11172), .ZN(
        n11178) );
  NAND2_X1 U14107 ( .A1(n13149), .A2(n11287), .ZN(n13046) );
  NAND2_X1 U14108 ( .A1(n14410), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19872) );
  INV_X1 U14109 ( .A(n19872), .ZN(n11174) );
  AND2_X1 U14110 ( .A1(n12902), .A2(n11174), .ZN(n11175) );
  NAND4_X1 U14111 ( .A1(n13048), .A2(n11176), .A3(n13046), .A4(n11175), .ZN(
        n11177) );
  NOR2_X1 U14112 ( .A1(n11178), .A2(n11177), .ZN(n11179) );
  OAI211_X1 U14113 ( .C1(n11182), .C2(n11181), .A(n11180), .B(n11179), .ZN(
        n11200) );
  INV_X1 U14114 ( .A(n11185), .ZN(n11183) );
  NAND2_X1 U14115 ( .A1(n11184), .A2(n11183), .ZN(n20205) );
  NAND2_X1 U14116 ( .A1(n20205), .A2(n11245), .ZN(n14385) );
  AOI22_X1 U14117 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U14118 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11128), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U14119 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U14120 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n9603), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11187) );
  NAND4_X1 U14121 ( .A1(n11190), .A2(n11189), .A3(n11188), .A4(n11187), .ZN(
        n11197) );
  AOI22_X1 U14122 ( .A1(n11329), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U14123 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n9605), .B1(n9606), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11194) );
  AOI22_X1 U14124 ( .A1(n13771), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11193) );
  AOI22_X1 U14125 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11192) );
  NAND4_X1 U14126 ( .A1(n11195), .A2(n11194), .A3(n11193), .A4(n11192), .ZN(
        n11196) );
  OR2_X1 U14127 ( .A1(n11304), .A2(n11232), .ZN(n11198) );
  OAI21_X1 U14128 ( .B1(n14385), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11198), 
        .ZN(n11199) );
  INV_X1 U14129 ( .A(n11199), .ZN(n11858) );
  INV_X1 U14130 ( .A(n11200), .ZN(n11201) );
  NAND2_X1 U14131 ( .A1(n11289), .A2(n20754), .ZN(n11226) );
  AOI22_X1 U14132 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11206) );
  AOI22_X1 U14133 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14134 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U14135 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11203) );
  NAND4_X1 U14136 ( .A1(n11206), .A2(n11205), .A3(n11204), .A4(n11203), .ZN(
        n11213) );
  AOI22_X1 U14137 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14138 ( .A1(n11329), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14139 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11209) );
  AOI22_X1 U14140 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11208) );
  NAND4_X1 U14141 ( .A1(n11211), .A2(n11210), .A3(n11209), .A4(n11208), .ZN(
        n11212) );
  NAND2_X1 U14142 ( .A1(n13054), .A2(n11895), .ZN(n11227) );
  NOR2_X1 U14143 ( .A1(n11304), .A2(n11895), .ZN(n11231) );
  AOI22_X1 U14144 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14145 ( .A1(n11073), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13773), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14146 ( .A1(n13771), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9603), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14147 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11214) );
  NAND4_X1 U14148 ( .A1(n11217), .A2(n11216), .A3(n11215), .A4(n11214), .ZN(
        n11223) );
  AOI22_X1 U14149 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13784), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14150 ( .A1(n11089), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11220) );
  AOI22_X1 U14151 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11219) );
  AOI22_X1 U14152 ( .A1(n11713), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11218) );
  NAND4_X1 U14153 ( .A1(n11221), .A2(n11220), .A3(n11219), .A4(n11218), .ZN(
        n11222) );
  MUX2_X1 U14154 ( .A(n11836), .B(n11231), .S(n11865), .Z(n11224) );
  INV_X1 U14155 ( .A(n11224), .ZN(n11225) );
  NAND2_X1 U14156 ( .A1(n11226), .A2(n11225), .ZN(n11286) );
  INV_X1 U14157 ( .A(n13054), .ZN(n20176) );
  AOI21_X1 U14158 ( .B1(n20146), .B2(n11865), .A(n20754), .ZN(n11228) );
  OAI211_X1 U14159 ( .C1(n11816), .C2(n20156), .A(n11228), .B(n11227), .ZN(
        n11285) );
  NAND2_X1 U14160 ( .A1(n11286), .A2(n11285), .ZN(n11230) );
  INV_X1 U14161 ( .A(n11836), .ZN(n11229) );
  INV_X1 U14162 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11235) );
  INV_X1 U14163 ( .A(n11231), .ZN(n11234) );
  OR2_X1 U14164 ( .A1(n11305), .A2(n11232), .ZN(n11233) );
  OAI211_X1 U14165 ( .C1(n11816), .C2(n11235), .A(n11234), .B(n11233), .ZN(
        n11237) );
  INV_X1 U14166 ( .A(n11237), .ZN(n11236) );
  INV_X1 U14167 ( .A(n11240), .ZN(n11243) );
  INV_X1 U14168 ( .A(n11241), .ZN(n11242) );
  OAI21_X1 U14169 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11243), .A(
        n11242), .ZN(n11244) );
  INV_X1 U14170 ( .A(n11252), .ZN(n11250) );
  XNOR2_X1 U14171 ( .A(n20529), .B(n20429), .ZN(n20151) );
  NAND2_X1 U14172 ( .A1(n20151), .A2(n11833), .ZN(n11247) );
  INV_X1 U14173 ( .A(n11251), .ZN(n11249) );
  AOI22_X1 U14174 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14175 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14176 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U14177 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11254) );
  NAND4_X1 U14178 ( .A1(n11257), .A2(n11256), .A3(n11255), .A4(n11254), .ZN(
        n11263) );
  AOI22_X1 U14179 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11261) );
  AOI22_X1 U14180 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11260) );
  AOI22_X1 U14181 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11259) );
  AOI22_X1 U14182 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11258) );
  NAND4_X1 U14183 ( .A1(n11261), .A2(n11260), .A3(n11259), .A4(n11258), .ZN(
        n11262) );
  OAI22_X2 U14184 ( .A1(n12991), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11874), 
        .B2(n11304), .ZN(n11266) );
  INV_X1 U14185 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20167) );
  OAI22_X1 U14186 ( .A1(n11305), .A2(n11874), .B1(n11816), .B2(n20167), .ZN(
        n11264) );
  INV_X1 U14187 ( .A(n11264), .ZN(n11265) );
  XNOR2_X2 U14188 ( .A(n11266), .B(n11265), .ZN(n11298) );
  NOR2_X2 U14189 ( .A1(n20188), .A2(n11268), .ZN(n11501) );
  NAND2_X1 U14190 ( .A1(n14390), .A2(n11501), .ZN(n11275) );
  NAND2_X1 U14191 ( .A1(n13161), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11361) );
  NOR2_X2 U14192 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13804) );
  XNOR2_X1 U14193 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14000) );
  AOI21_X1 U14194 ( .B1(n13804), .B2(n14000), .A(n13808), .ZN(n11271) );
  NAND2_X1 U14195 ( .A1(n11269), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11270) );
  OAI211_X1 U14196 ( .C1(n11361), .C2(n11272), .A(n11271), .B(n11270), .ZN(
        n11273) );
  INV_X1 U14197 ( .A(n11273), .ZN(n11274) );
  NAND2_X1 U14198 ( .A1(n11275), .A2(n11274), .ZN(n11276) );
  NAND2_X1 U14199 ( .A1(n13808), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11297) );
  NAND2_X1 U14200 ( .A1(n11276), .A2(n11297), .ZN(n13158) );
  INV_X1 U14201 ( .A(n11858), .ZN(n11278) );
  NAND2_X1 U14202 ( .A1(n14386), .A2(n11501), .ZN(n11284) );
  NAND2_X1 U14203 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n11268), .ZN(
        n11281) );
  NAND2_X1 U14204 ( .A1(n11269), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n11280) );
  OAI211_X1 U14205 ( .C1(n11361), .C2(n11035), .A(n11281), .B(n11280), .ZN(
        n11282) );
  INV_X1 U14206 ( .A(n11282), .ZN(n11283) );
  NAND2_X1 U14207 ( .A1(n11284), .A2(n11283), .ZN(n13401) );
  NAND2_X1 U14208 ( .A1(n11869), .A2(n11287), .ZN(n11288) );
  NAND2_X1 U14209 ( .A1(n11288), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13263) );
  AOI22_X1 U14210 ( .A1(n11269), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n11268), .ZN(n11292) );
  INV_X1 U14211 ( .A(n11361), .ZN(n11290) );
  NAND2_X1 U14212 ( .A1(n11290), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11291) );
  NAND2_X1 U14213 ( .A1(n11292), .A2(n11291), .ZN(n11293) );
  AOI21_X1 U14214 ( .B1(n11289), .B2(n11501), .A(n11293), .ZN(n13264) );
  OR2_X1 U14215 ( .A1(n13263), .A2(n13264), .ZN(n13265) );
  NAND2_X1 U14216 ( .A1(n13264), .A2(n13804), .ZN(n11294) );
  NAND2_X1 U14217 ( .A1(n13265), .A2(n11294), .ZN(n13400) );
  NAND2_X1 U14218 ( .A1(n13401), .A2(n13400), .ZN(n13399) );
  NAND2_X1 U14219 ( .A1(n11296), .A2(n11295), .ZN(n13156) );
  NAND2_X1 U14220 ( .A1(n13156), .A2(n11297), .ZN(n13183) );
  NAND2_X1 U14221 ( .A1(n20234), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20333) );
  INV_X1 U14222 ( .A(n20333), .ZN(n20363) );
  INV_X1 U14223 ( .A(n20422), .ZN(n20400) );
  OAI21_X1 U14224 ( .B1(n20685), .B2(n20429), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11300) );
  NAND2_X1 U14225 ( .A1(n20400), .A2(n11300), .ZN(n20431) );
  NOR2_X1 U14226 ( .A1(n15551), .A2(n20234), .ZN(n11301) );
  AOI21_X1 U14227 ( .B1(n20431), .B2(n11833), .A(n11301), .ZN(n11302) );
  AOI22_X1 U14228 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14229 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14230 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11307) );
  AOI22_X1 U14231 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11306) );
  NAND4_X1 U14232 ( .A1(n11309), .A2(n11308), .A3(n11307), .A4(n11306), .ZN(
        n11315) );
  AOI22_X1 U14233 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14234 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14235 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14236 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11310) );
  NAND4_X1 U14237 ( .A1(n11313), .A2(n11312), .A3(n11311), .A4(n11310), .ZN(
        n11314) );
  AOI22_X1 U14238 ( .A1(n11811), .A2(n11884), .B1(n11824), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11316) );
  XNOR2_X1 U14239 ( .A(n11324), .B(n14394), .ZN(n20140) );
  NAND2_X1 U14240 ( .A1(n20140), .A2(n11501), .ZN(n11323) );
  AND2_X1 U14241 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11318) );
  INV_X1 U14242 ( .A(n11358), .ZN(n11317) );
  OAI21_X1 U14243 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11318), .A(
        n11317), .ZN(n13990) );
  AOI22_X1 U14244 ( .A1(n13804), .A2(n13990), .B1(n13808), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11320) );
  NAND2_X1 U14245 ( .A1(n13799), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11319) );
  OAI211_X1 U14246 ( .C1(n11361), .C2(n11036), .A(n11320), .B(n11319), .ZN(
        n11321) );
  INV_X1 U14247 ( .A(n11321), .ZN(n11322) );
  NAND2_X1 U14248 ( .A1(n11323), .A2(n11322), .ZN(n13182) );
  AND2_X2 U14249 ( .A1(n13183), .A2(n13182), .ZN(n13249) );
  AOI22_X1 U14250 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14251 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14252 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14253 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11325) );
  NAND4_X1 U14254 ( .A1(n11328), .A2(n11327), .A3(n11326), .A4(n11325), .ZN(
        n11335) );
  AOI22_X1 U14255 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14256 ( .A1(n11329), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14257 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14258 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11330) );
  NAND4_X1 U14259 ( .A1(n11333), .A2(n11332), .A3(n11331), .A4(n11330), .ZN(
        n11334) );
  AOI22_X1 U14260 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14261 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14262 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14263 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11336) );
  NAND4_X1 U14264 ( .A1(n11339), .A2(n11338), .A3(n11337), .A4(n11336), .ZN(
        n11345) );
  AOI22_X1 U14265 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14266 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14267 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14268 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11340) );
  NAND4_X1 U14269 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(
        n11344) );
  NAND2_X1 U14270 ( .A1(n11811), .A2(n11851), .ZN(n11347) );
  NAND2_X1 U14271 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11346) );
  NAND2_X1 U14272 ( .A1(n11347), .A2(n11346), .ZN(n11380) );
  XNOR2_X1 U14273 ( .A(n11381), .B(n9788), .ZN(n11853) );
  NAND2_X1 U14274 ( .A1(n11853), .A2(n11501), .ZN(n11354) );
  INV_X2 U14275 ( .A(n11553), .ZN(n13799) );
  INV_X1 U14276 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11351) );
  INV_X1 U14277 ( .A(n13808), .ZN(n11473) );
  NAND2_X1 U14278 ( .A1(n11357), .A2(n11351), .ZN(n11349) );
  NAND2_X1 U14279 ( .A1(n11349), .A2(n11366), .ZN(n19936) );
  NAND2_X1 U14280 ( .A1(n19936), .A2(n13804), .ZN(n11350) );
  OAI21_X1 U14281 ( .B1(n11351), .B2(n11473), .A(n11350), .ZN(n11352) );
  AOI21_X1 U14282 ( .B1(n13799), .B2(P1_EAX_REG_5__SCAN_IN), .A(n11352), .ZN(
        n11353) );
  NAND2_X1 U14283 ( .A1(n11354), .A2(n11353), .ZN(n13217) );
  XNOR2_X1 U14284 ( .A(n11356), .B(n10076), .ZN(n11857) );
  NAND2_X1 U14285 ( .A1(n11857), .A2(n11501), .ZN(n11364) );
  OAI21_X1 U14286 ( .B1(n11358), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11357), .ZN(n20074) );
  INV_X2 U14287 ( .A(n13804), .ZN(n13797) );
  OAI21_X1 U14288 ( .B1(n14399), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11268), .ZN(n11360) );
  NAND2_X1 U14289 ( .A1(n13799), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11359) );
  OAI211_X1 U14290 ( .C1(n11361), .C2(n12990), .A(n11360), .B(n11359), .ZN(
        n11362) );
  OAI21_X1 U14291 ( .B1(n20074), .B2(n13797), .A(n11362), .ZN(n11363) );
  NAND2_X1 U14292 ( .A1(n11364), .A2(n11363), .ZN(n13250) );
  OAI21_X1 U14293 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11367), .A(
        n11387), .ZN(n19924) );
  INV_X1 U14294 ( .A(n19924), .ZN(n11384) );
  AOI22_X1 U14295 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14296 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11370) );
  INV_X1 U14297 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20193) );
  AOI22_X1 U14298 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14299 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11368) );
  NAND4_X1 U14300 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n11377) );
  AOI22_X1 U14301 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14302 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14303 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14304 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11372) );
  NAND4_X1 U14305 ( .A1(n11375), .A2(n11374), .A3(n11373), .A4(n11372), .ZN(
        n11376) );
  NAND2_X1 U14306 ( .A1(n11811), .A2(n11839), .ZN(n11379) );
  NAND2_X1 U14307 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11378) );
  AOI22_X1 U14308 ( .A1(n13799), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n13808), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11382) );
  INV_X1 U14309 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20203) );
  NAND2_X1 U14310 ( .A1(n11811), .A2(n11895), .ZN(n11385) );
  OAI21_X1 U14311 ( .B1(n20203), .B2(n11816), .A(n11385), .ZN(n11386) );
  OAI21_X1 U14312 ( .B1(n11388), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n11410), .ZN(n19909) );
  NAND2_X1 U14313 ( .A1(n19909), .A2(n13804), .ZN(n11390) );
  AOI22_X1 U14314 ( .A1(n13799), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n13808), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11389) );
  NAND2_X1 U14315 ( .A1(n11390), .A2(n11389), .ZN(n11391) );
  XNOR2_X1 U14316 ( .A(n11410), .B(n11409), .ZN(n14258) );
  NAND2_X1 U14317 ( .A1(n14258), .A2(n13804), .ZN(n11407) );
  INV_X1 U14318 ( .A(n11501), .ZN(n11518) );
  AOI22_X1 U14319 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11128), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14320 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14321 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14322 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11392) );
  NAND4_X1 U14323 ( .A1(n11395), .A2(n11394), .A3(n11393), .A4(n11392), .ZN(
        n11401) );
  AOI22_X1 U14324 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14325 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14326 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14327 ( .A1(n13771), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11396) );
  NAND4_X1 U14328 ( .A1(n11399), .A2(n11398), .A3(n11397), .A4(n11396), .ZN(
        n11400) );
  NOR2_X1 U14329 ( .A1(n11401), .A2(n11400), .ZN(n11404) );
  NAND2_X1 U14330 ( .A1(n13799), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11403) );
  NAND2_X1 U14331 ( .A1(n13808), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11402) );
  OAI211_X1 U14332 ( .C1(n11518), .C2(n11404), .A(n11403), .B(n11402), .ZN(
        n11405) );
  INV_X1 U14333 ( .A(n11405), .ZN(n11406) );
  XOR2_X1 U14334 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11424), .Z(n19892) );
  AOI22_X1 U14335 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13784), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14336 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11128), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14337 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14338 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n9603), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11411) );
  NAND4_X1 U14339 ( .A1(n11414), .A2(n11413), .A3(n11412), .A4(n11411), .ZN(
        n11420) );
  AOI22_X1 U14340 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14341 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11708), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14342 ( .A1(n9605), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n9606), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14343 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11415) );
  NAND4_X1 U14344 ( .A1(n11418), .A2(n11417), .A3(n11416), .A4(n11415), .ZN(
        n11419) );
  OR2_X1 U14345 ( .A1(n11420), .A2(n11419), .ZN(n11421) );
  AOI22_X1 U14346 ( .A1(n11501), .A2(n11421), .B1(n13808), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11423) );
  NAND2_X1 U14347 ( .A1(n13799), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11422) );
  OAI211_X1 U14348 ( .C1(n19892), .C2(n13797), .A(n11423), .B(n11422), .ZN(
        n13442) );
  XNOR2_X1 U14349 ( .A(n11442), .B(n11441), .ZN(n14249) );
  AOI22_X1 U14350 ( .A1(n11446), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14351 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14352 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14353 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11425) );
  NAND4_X1 U14354 ( .A1(n11428), .A2(n11427), .A3(n11426), .A4(n11425), .ZN(
        n11434) );
  AOI22_X1 U14355 ( .A1(n11693), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14356 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14357 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14358 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11429) );
  NAND4_X1 U14359 ( .A1(n11432), .A2(n11431), .A3(n11430), .A4(n11429), .ZN(
        n11433) );
  NOR2_X1 U14360 ( .A1(n11434), .A2(n11433), .ZN(n11437) );
  NAND2_X1 U14361 ( .A1(n13799), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11436) );
  NAND2_X1 U14362 ( .A1(n13808), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11435) );
  OAI211_X1 U14363 ( .C1(n11518), .C2(n11437), .A(n11436), .B(n11435), .ZN(
        n11438) );
  AOI21_X1 U14364 ( .B1(n14249), .B2(n13804), .A(n11438), .ZN(n13498) );
  INV_X1 U14365 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15735) );
  OAI21_X1 U14366 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11443), .A(
        n11472), .ZN(n15824) );
  NAND2_X1 U14367 ( .A1(n15824), .A2(n13804), .ZN(n11444) );
  OAI21_X1 U14368 ( .B1(n11473), .B2(n15735), .A(n11444), .ZN(n11445) );
  AOI21_X1 U14369 ( .B1(n13799), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11445), .ZN(
        n13963) );
  BUF_X1 U14370 ( .A(n11446), .Z(n13782) );
  AOI22_X1 U14371 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13784), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14372 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13773), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14373 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9603), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U14374 ( .A1(n11693), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11447) );
  NAND4_X1 U14375 ( .A1(n11450), .A2(n11449), .A3(n11448), .A4(n11447), .ZN(
        n11456) );
  AOI22_X1 U14376 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14377 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14378 ( .A1(n9605), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14379 ( .A1(n11713), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11451) );
  NAND4_X1 U14380 ( .A1(n11454), .A2(n11453), .A3(n11452), .A4(n11451), .ZN(
        n11455) );
  OR2_X1 U14381 ( .A1(n11456), .A2(n11455), .ZN(n11457) );
  NAND2_X1 U14382 ( .A1(n11501), .A2(n11457), .ZN(n15725) );
  INV_X1 U14383 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14159) );
  AOI22_X1 U14384 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13784), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U14385 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14386 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14387 ( .A1(n11713), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11458) );
  NAND4_X1 U14388 ( .A1(n11461), .A2(n11460), .A3(n11459), .A4(n11458), .ZN(
        n11467) );
  AOI22_X1 U14389 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14390 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9603), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14391 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14392 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11462) );
  NAND4_X1 U14393 ( .A1(n11465), .A2(n11464), .A3(n11463), .A4(n11462), .ZN(
        n11466) );
  OAI21_X1 U14394 ( .B1(n11467), .B2(n11466), .A(n11501), .ZN(n11471) );
  INV_X1 U14395 ( .A(n11489), .ZN(n11468) );
  XNOR2_X1 U14396 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11468), .ZN(
        n14244) );
  INV_X1 U14397 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14242) );
  OAI22_X1 U14398 ( .A1(n14244), .A2(n13797), .B1(n11473), .B2(n14242), .ZN(
        n11469) );
  INV_X1 U14399 ( .A(n11469), .ZN(n11470) );
  OAI211_X1 U14400 ( .C1(n11553), .C2(n14159), .A(n11471), .B(n11470), .ZN(
        n13969) );
  INV_X1 U14401 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n11488) );
  XNOR2_X1 U14402 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11472), .ZN(
        n15814) );
  OAI22_X1 U14403 ( .A1(n15814), .A2(n13797), .B1(n11473), .B2(n15717), .ZN(
        n11474) );
  INV_X1 U14404 ( .A(n11474), .ZN(n11487) );
  AOI22_X1 U14405 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13784), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U14406 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14407 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9603), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14408 ( .A1(n11693), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11475) );
  NAND4_X1 U14409 ( .A1(n11478), .A2(n11477), .A3(n11476), .A4(n11475), .ZN(
        n11484) );
  AOI22_X1 U14410 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14411 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14412 ( .A1(n9605), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14413 ( .A1(n11713), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11479) );
  NAND4_X1 U14414 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n11483) );
  OR2_X1 U14415 ( .A1(n11484), .A2(n11483), .ZN(n11485) );
  NAND2_X1 U14416 ( .A1(n11501), .A2(n11485), .ZN(n11486) );
  OAI211_X1 U14417 ( .C1(n11553), .C2(n11488), .A(n11487), .B(n11486), .ZN(
        n14092) );
  XOR2_X1 U14418 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11504), .Z(
        n15711) );
  AOI22_X1 U14419 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14420 ( .A1(n13771), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9603), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11492) );
  AOI22_X1 U14421 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14422 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11490) );
  NAND4_X1 U14423 ( .A1(n11493), .A2(n11492), .A3(n11491), .A4(n11490), .ZN(
        n11499) );
  AOI22_X1 U14424 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11497) );
  AOI22_X1 U14425 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11128), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11496) );
  AOI22_X1 U14426 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14427 ( .A1(n11713), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11494) );
  NAND4_X1 U14428 ( .A1(n11497), .A2(n11496), .A3(n11495), .A4(n11494), .ZN(
        n11498) );
  OR2_X1 U14429 ( .A1(n11499), .A2(n11498), .ZN(n11500) );
  AOI22_X1 U14430 ( .A1(n11501), .A2(n11500), .B1(n13808), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11503) );
  NAND2_X1 U14431 ( .A1(n13799), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11502) );
  OAI211_X1 U14432 ( .C1(n15711), .C2(n13797), .A(n11503), .B(n11502), .ZN(
        n13614) );
  XNOR2_X1 U14433 ( .A(n11536), .B(n14230), .ZN(n14228) );
  NAND2_X1 U14434 ( .A1(n14228), .A2(n13804), .ZN(n11521) );
  AOI22_X1 U14435 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14436 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14437 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14438 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11505) );
  NAND4_X1 U14439 ( .A1(n11508), .A2(n11507), .A3(n11506), .A4(n11505), .ZN(
        n11514) );
  AOI22_X1 U14440 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14441 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14442 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14443 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11509) );
  NAND4_X1 U14444 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11513) );
  NOR2_X1 U14445 ( .A1(n11514), .A2(n11513), .ZN(n11517) );
  NAND2_X1 U14446 ( .A1(n13799), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11516) );
  NAND2_X1 U14447 ( .A1(n13808), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11515) );
  OAI211_X1 U14448 ( .C1(n11518), .C2(n11517), .A(n11516), .B(n11515), .ZN(
        n11519) );
  INV_X1 U14449 ( .A(n11519), .ZN(n11520) );
  NAND2_X1 U14450 ( .A1(n11521), .A2(n11520), .ZN(n13634) );
  AOI22_X1 U14451 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14452 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14453 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14454 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11522) );
  NAND4_X1 U14455 ( .A1(n11525), .A2(n11524), .A3(n11523), .A4(n11522), .ZN(
        n11531) );
  AOI22_X1 U14456 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13782), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14457 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U14458 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14459 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11526) );
  NAND4_X1 U14460 ( .A1(n11529), .A2(n11528), .A3(n11527), .A4(n11526), .ZN(
        n11530) );
  NOR2_X1 U14461 ( .A1(n11531), .A2(n11530), .ZN(n11535) );
  OAI21_X1 U14462 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n14399), .A(
        n11268), .ZN(n11532) );
  INV_X1 U14463 ( .A(n11532), .ZN(n11533) );
  AOI21_X1 U14464 ( .B1(n13799), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11533), .ZN(
        n11534) );
  OAI21_X1 U14465 ( .B1(n13801), .B2(n11535), .A(n11534), .ZN(n11539) );
  OAI21_X1 U14466 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11537), .A(
        n11571), .ZN(n15806) );
  OR2_X1 U14467 ( .A1(n13797), .A2(n15806), .ZN(n11538) );
  NAND2_X1 U14468 ( .A1(n11539), .A2(n11538), .ZN(n14079) );
  INV_X1 U14469 ( .A(n13801), .ZN(n11744) );
  AOI22_X1 U14470 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14471 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14472 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14473 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n9603), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11540) );
  NAND4_X1 U14474 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(
        n11549) );
  AOI22_X1 U14475 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n13773), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14476 ( .A1(n9605), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14477 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11128), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14478 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11544) );
  NAND4_X1 U14479 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11548) );
  OR2_X1 U14480 ( .A1(n11549), .A2(n11548), .ZN(n11555) );
  INV_X1 U14481 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n11552) );
  INV_X1 U14482 ( .A(n11571), .ZN(n11550) );
  XNOR2_X1 U14483 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11550), .ZN(
        n14215) );
  AOI22_X1 U14484 ( .A1(n13804), .A2(n14215), .B1(n13808), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11551) );
  OAI21_X1 U14485 ( .B1(n11553), .B2(n11552), .A(n11551), .ZN(n11554) );
  AOI21_X1 U14486 ( .B1(n11744), .B2(n11555), .A(n11554), .ZN(n13952) );
  AOI22_X1 U14487 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U14488 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U14489 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14490 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11557) );
  NAND4_X1 U14491 ( .A1(n11560), .A2(n11559), .A3(n11558), .A4(n11557), .ZN(
        n11566) );
  AOI22_X1 U14492 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14493 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14494 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14495 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11561) );
  NAND4_X1 U14496 ( .A1(n11564), .A2(n11563), .A3(n11562), .A4(n11561), .ZN(
        n11565) );
  NOR2_X1 U14497 ( .A1(n11566), .A2(n11565), .ZN(n11570) );
  NAND2_X1 U14498 ( .A1(n11268), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11567) );
  NAND2_X1 U14499 ( .A1(n13797), .A2(n11567), .ZN(n11568) );
  AOI21_X1 U14500 ( .B1(n13799), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11568), .ZN(
        n11569) );
  OAI21_X1 U14501 ( .B1(n13801), .B2(n11570), .A(n11569), .ZN(n11574) );
  INV_X1 U14502 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14216) );
  OAI21_X1 U14503 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11572), .A(
        n11604), .ZN(n15795) );
  OR2_X1 U14504 ( .A1(n13797), .A2(n15795), .ZN(n11573) );
  NAND2_X1 U14505 ( .A1(n11574), .A2(n11573), .ZN(n14071) );
  AOI22_X1 U14506 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13782), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14507 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11128), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14508 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U14509 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11575) );
  NAND4_X1 U14510 ( .A1(n11578), .A2(n11577), .A3(n11576), .A4(n11575), .ZN(
        n11584) );
  AOI22_X1 U14511 ( .A1(n13771), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9603), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14512 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14513 ( .A1(n13781), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14514 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11579) );
  NAND4_X1 U14515 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n11583) );
  NOR2_X1 U14516 ( .A1(n11584), .A2(n11583), .ZN(n11587) );
  INV_X1 U14517 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14202) );
  OAI21_X1 U14518 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14202), .A(n13797), 
        .ZN(n11585) );
  AOI21_X1 U14519 ( .B1(n13799), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11585), .ZN(
        n11586) );
  OAI21_X1 U14520 ( .B1(n13801), .B2(n11587), .A(n11586), .ZN(n11589) );
  XNOR2_X1 U14521 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n11604), .ZN(
        n14204) );
  NAND2_X1 U14522 ( .A1(n13804), .A2(n14204), .ZN(n11588) );
  AOI22_X1 U14523 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14524 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11128), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U14525 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U14526 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11590) );
  NAND4_X1 U14527 ( .A1(n11593), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n11599) );
  AOI22_X1 U14528 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14529 ( .A1(n13771), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14530 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14531 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11594) );
  NAND4_X1 U14532 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n11598) );
  NOR2_X1 U14533 ( .A1(n11599), .A2(n11598), .ZN(n11603) );
  NAND2_X1 U14534 ( .A1(n11268), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11600) );
  NAND2_X1 U14535 ( .A1(n13797), .A2(n11600), .ZN(n11601) );
  AOI21_X1 U14536 ( .B1(n13799), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11601), .ZN(
        n11602) );
  OAI21_X1 U14537 ( .B1(n13801), .B2(n11603), .A(n11602), .ZN(n11607) );
  OAI21_X1 U14538 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11605), .A(
        n11639), .ZN(n15786) );
  OR2_X1 U14539 ( .A1(n13797), .A2(n15786), .ZN(n11606) );
  AOI22_X1 U14540 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13782), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14541 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14542 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9603), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14543 ( .A1(n11694), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11608) );
  NAND4_X1 U14544 ( .A1(n11611), .A2(n11610), .A3(n11609), .A4(n11608), .ZN(
        n11617) );
  AOI22_X1 U14545 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14546 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11329), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14547 ( .A1(n11693), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14548 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11612) );
  NAND4_X1 U14549 ( .A1(n11615), .A2(n11614), .A3(n11613), .A4(n11612), .ZN(
        n11616) );
  NOR2_X1 U14550 ( .A1(n11617), .A2(n11616), .ZN(n11621) );
  NAND2_X1 U14551 ( .A1(n11268), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11618) );
  NAND2_X1 U14552 ( .A1(n13797), .A2(n11618), .ZN(n11619) );
  AOI21_X1 U14553 ( .B1(n13799), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11619), .ZN(
        n11620) );
  OAI21_X1 U14554 ( .B1(n13801), .B2(n11621), .A(n11620), .ZN(n11624) );
  INV_X1 U14555 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11635) );
  OAI21_X1 U14556 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11622), .A(
        n11684), .ZN(n15779) );
  OR2_X1 U14557 ( .A1(n13797), .A2(n15779), .ZN(n11623) );
  NAND2_X1 U14558 ( .A1(n11624), .A2(n11623), .ZN(n14048) );
  AOI22_X1 U14559 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U14560 ( .A1(n11128), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U14561 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14562 ( .A1(n11693), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11625) );
  NAND4_X1 U14563 ( .A1(n11628), .A2(n11627), .A3(n11626), .A4(n11625), .ZN(
        n11634) );
  AOI22_X1 U14564 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14565 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U14566 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14567 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11629) );
  NAND4_X1 U14568 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n11633) );
  NOR2_X1 U14569 ( .A1(n11634), .A2(n11633), .ZN(n11638) );
  OAI21_X1 U14570 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n11635), .A(n13797), 
        .ZN(n11636) );
  AOI21_X1 U14571 ( .B1(n13799), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11636), .ZN(
        n11637) );
  OAI21_X1 U14572 ( .B1(n13801), .B2(n11638), .A(n11637), .ZN(n11641) );
  XNOR2_X1 U14573 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n11639), .ZN(
        n15780) );
  NAND2_X1 U14574 ( .A1(n15780), .A2(n13804), .ZN(n11640) );
  NAND2_X1 U14575 ( .A1(n11641), .A2(n11640), .ZN(n14055) );
  AOI22_X1 U14576 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14577 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11329), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14578 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14579 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11643) );
  NAND4_X1 U14580 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n11652) );
  AOI22_X1 U14581 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14582 ( .A1(n13771), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14583 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14584 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11647) );
  NAND4_X1 U14585 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(
        n11651) );
  NOR2_X1 U14586 ( .A1(n11652), .A2(n11651), .ZN(n11669) );
  AOI22_X1 U14587 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11329), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14588 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11133), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14589 ( .A1(n11693), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14590 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11653) );
  NAND4_X1 U14591 ( .A1(n11656), .A2(n11655), .A3(n11654), .A4(n11653), .ZN(
        n11663) );
  AOI22_X1 U14592 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14593 ( .A1(n13771), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14594 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14595 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11658) );
  NAND4_X1 U14596 ( .A1(n11661), .A2(n11660), .A3(n11659), .A4(n11658), .ZN(
        n11662) );
  NOR2_X1 U14597 ( .A1(n11663), .A2(n11662), .ZN(n11670) );
  XNOR2_X1 U14598 ( .A(n11669), .B(n11670), .ZN(n11666) );
  INV_X1 U14599 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14193) );
  OAI21_X1 U14600 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14193), .A(n13797), 
        .ZN(n11664) );
  AOI21_X1 U14601 ( .B1(n13799), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11664), .ZN(
        n11665) );
  OAI21_X1 U14602 ( .B1(n13801), .B2(n11666), .A(n11665), .ZN(n11668) );
  XNOR2_X1 U14603 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n11684), .ZN(
        n14195) );
  NAND2_X1 U14604 ( .A1(n13804), .A2(n14195), .ZN(n11667) );
  NOR2_X1 U14605 ( .A1(n11670), .A2(n11669), .ZN(n11702) );
  AOI22_X1 U14606 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14607 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11708), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14608 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14609 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11671) );
  NAND4_X1 U14610 ( .A1(n11674), .A2(n11673), .A3(n11672), .A4(n11671), .ZN(
        n11680) );
  INV_X1 U14611 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14606) );
  AOI22_X1 U14612 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14613 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n13773), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14614 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14615 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n9603), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11675) );
  NAND4_X1 U14616 ( .A1(n11678), .A2(n11677), .A3(n11676), .A4(n11675), .ZN(
        n11679) );
  OR2_X1 U14617 ( .A1(n11680), .A2(n11679), .ZN(n11701) );
  INV_X1 U14618 ( .A(n11701), .ZN(n11681) );
  XNOR2_X1 U14619 ( .A(n11702), .B(n11681), .ZN(n11682) );
  NAND2_X1 U14620 ( .A1(n11682), .A2(n11744), .ZN(n11688) );
  INV_X1 U14621 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15649) );
  AOI21_X1 U14622 ( .B1(n15649), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11683) );
  AOI21_X1 U14623 ( .B1(n13799), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11683), .ZN(
        n11687) );
  OAI21_X1 U14624 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n11685), .A(
        n11726), .ZN(n15772) );
  NOR2_X1 U14625 ( .A1(n15772), .A2(n13797), .ZN(n11686) );
  AOI21_X1 U14626 ( .B1(n11688), .B2(n11687), .A(n11686), .ZN(n14043) );
  AOI22_X1 U14627 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14628 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11329), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14629 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14630 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11689) );
  NAND4_X1 U14631 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n11700) );
  AOI22_X1 U14632 ( .A1(n13771), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14633 ( .A1(n9605), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14634 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14635 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11695) );
  NAND4_X1 U14636 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n11699) );
  NOR2_X1 U14637 ( .A1(n11700), .A2(n11699), .ZN(n11721) );
  NAND2_X1 U14638 ( .A1(n11702), .A2(n11701), .ZN(n11720) );
  XOR2_X1 U14639 ( .A(n11721), .B(n11720), .Z(n11703) );
  NAND2_X1 U14640 ( .A1(n11703), .A2(n11744), .ZN(n11707) );
  INV_X1 U14641 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14184) );
  OAI21_X1 U14642 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14184), .A(n13797), 
        .ZN(n11704) );
  AOI21_X1 U14643 ( .B1(n13799), .B2(P1_EAX_REG_25__SCAN_IN), .A(n11704), .ZN(
        n11706) );
  XNOR2_X1 U14644 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B(n11726), .ZN(
        n14186) );
  AOI22_X1 U14645 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11329), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14646 ( .A1(n13771), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11128), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14647 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14648 ( .A1(n9606), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11709) );
  NAND4_X1 U14649 ( .A1(n11712), .A2(n11711), .A3(n11710), .A4(n11709), .ZN(
        n11719) );
  AOI22_X1 U14650 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14651 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13775), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14652 ( .A1(n9605), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11713), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14653 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11714) );
  NAND4_X1 U14654 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11714), .ZN(
        n11718) );
  NOR2_X1 U14655 ( .A1(n11719), .A2(n11718), .ZN(n11731) );
  OR2_X1 U14656 ( .A1(n11721), .A2(n11720), .ZN(n11730) );
  XNOR2_X1 U14657 ( .A(n11731), .B(n11730), .ZN(n11725) );
  NAND2_X1 U14658 ( .A1(n11268), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11722) );
  NAND2_X1 U14659 ( .A1(n13797), .A2(n11722), .ZN(n11723) );
  AOI21_X1 U14660 ( .B1(n13799), .B2(P1_EAX_REG_26__SCAN_IN), .A(n11723), .ZN(
        n11724) );
  OAI21_X1 U14661 ( .B1(n11725), .B2(n13801), .A(n11724), .ZN(n11729) );
  OAI21_X1 U14662 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n11727), .A(
        n11768), .ZN(n15767) );
  OR2_X1 U14663 ( .A1(n13797), .A2(n15767), .ZN(n11728) );
  NAND2_X1 U14664 ( .A1(n11729), .A2(n11728), .ZN(n14031) );
  OR2_X1 U14665 ( .A1(n11731), .A2(n11730), .ZN(n11762) );
  AOI22_X1 U14666 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11708), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14667 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14668 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14669 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11734) );
  NAND4_X1 U14670 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n11743) );
  AOI22_X1 U14671 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14672 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11329), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U14673 ( .A1(n13771), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9603), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14674 ( .A1(n11693), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9606), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11738) );
  NAND4_X1 U14675 ( .A1(n11741), .A2(n11740), .A3(n11739), .A4(n11738), .ZN(
        n11742) );
  NOR2_X1 U14676 ( .A1(n11743), .A2(n11742), .ZN(n11763) );
  XOR2_X1 U14677 ( .A(n11762), .B(n11763), .Z(n11745) );
  NAND2_X1 U14678 ( .A1(n11745), .A2(n11744), .ZN(n11748) );
  INV_X1 U14679 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14174) );
  OAI21_X1 U14680 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14174), .A(n13797), 
        .ZN(n11746) );
  AOI21_X1 U14681 ( .B1(n13799), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11746), .ZN(
        n11747) );
  NAND2_X1 U14682 ( .A1(n11748), .A2(n11747), .ZN(n11750) );
  XNOR2_X1 U14683 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B(n11768), .ZN(
        n14176) );
  NAND2_X1 U14684 ( .A1(n13804), .A2(n14176), .ZN(n11749) );
  NAND2_X1 U14685 ( .A1(n11750), .A2(n11749), .ZN(n13904) );
  INV_X1 U14686 ( .A(n13904), .ZN(n11751) );
  AOI22_X1 U14687 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U14688 ( .A1(n13771), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U14689 ( .A1(n13781), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U14690 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11752) );
  NAND4_X1 U14691 ( .A1(n11755), .A2(n11754), .A3(n11753), .A4(n11752), .ZN(
        n11761) );
  AOI22_X1 U14692 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13773), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14693 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13782), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14694 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14695 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11756) );
  NAND4_X1 U14696 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11760) );
  NOR2_X1 U14697 ( .A1(n11761), .A2(n11760), .ZN(n11939) );
  OR2_X1 U14698 ( .A1(n11763), .A2(n11762), .ZN(n11938) );
  XNOR2_X1 U14699 ( .A(n11939), .B(n11938), .ZN(n11767) );
  NAND2_X1 U14700 ( .A1(n11268), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11764) );
  NAND2_X1 U14701 ( .A1(n13797), .A2(n11764), .ZN(n11765) );
  AOI21_X1 U14702 ( .B1(n13799), .B2(P1_EAX_REG_28__SCAN_IN), .A(n11765), .ZN(
        n11766) );
  OAI21_X1 U14703 ( .B1(n11767), .B2(n13801), .A(n11766), .ZN(n11771) );
  NAND2_X1 U14704 ( .A1(n11769), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11924) );
  OAI21_X1 U14705 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11769), .A(
        n11924), .ZN(n15617) );
  OR2_X1 U14706 ( .A1(n13797), .A2(n15617), .ZN(n11770) );
  NOR2_X1 U14707 ( .A1(n11772), .A2(n11773), .ZN(n11774) );
  NAND3_X1 U14708 ( .A1(n20754), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15973) );
  INV_X1 U14709 ( .A(n15973), .ZN(n11775) );
  AND2_X1 U14710 ( .A1(n11776), .A2(n12906), .ZN(n11777) );
  OAI211_X1 U14711 ( .C1(n11795), .C2(n20188), .A(n11778), .B(n11777), .ZN(
        n12907) );
  AND2_X1 U14712 ( .A1(n11152), .A2(n20146), .ZN(n11779) );
  NOR2_X1 U14713 ( .A1(n12907), .A2(n11779), .ZN(n12974) );
  NAND2_X1 U14714 ( .A1(n12974), .A2(n12901), .ZN(n15541) );
  NAND2_X1 U14715 ( .A1(n20182), .A2(n9614), .ZN(n11868) );
  XNOR2_X1 U14716 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11791) );
  NAND2_X1 U14717 ( .A1(n20611), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11794) );
  NAND2_X1 U14718 ( .A1(n11791), .A2(n11790), .ZN(n11781) );
  NAND2_X1 U14719 ( .A1(n20689), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11780) );
  NAND2_X1 U14720 ( .A1(n11781), .A2(n11780), .ZN(n11804) );
  XNOR2_X1 U14721 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11803) );
  NAND2_X1 U14722 ( .A1(n11804), .A2(n11803), .ZN(n11783) );
  NAND2_X1 U14723 ( .A1(n20429), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11782) );
  NAND2_X1 U14724 ( .A1(n11783), .A2(n11782), .ZN(n11789) );
  XNOR2_X1 U14725 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11788) );
  NAND2_X1 U14726 ( .A1(n11789), .A2(n11788), .ZN(n11785) );
  NAND2_X1 U14727 ( .A1(n20234), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11784) );
  NAND2_X1 U14728 ( .A1(n11785), .A2(n11784), .ZN(n11820) );
  AND2_X1 U14729 ( .A1(n20138), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11786) );
  NAND2_X1 U14730 ( .A1(n12990), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11819) );
  NAND2_X1 U14731 ( .A1(n11818), .A2(n12840), .ZN(n11829) );
  NAND2_X1 U14732 ( .A1(n12840), .A2(n11811), .ZN(n11828) );
  XNOR2_X1 U14733 ( .A(n11789), .B(n11788), .ZN(n12843) );
  XNOR2_X1 U14734 ( .A(n11791), .B(n11790), .ZN(n12842) );
  NAND2_X1 U14735 ( .A1(n11811), .A2(n9614), .ZN(n11793) );
  NAND2_X1 U14736 ( .A1(n12971), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11792) );
  NOR2_X1 U14737 ( .A1(n12842), .A2(n11800), .ZN(n11799) );
  AOI21_X1 U14738 ( .B1(n12971), .B2(n19976), .A(n9614), .ZN(n11813) );
  OAI21_X1 U14739 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20611), .A(
        n11794), .ZN(n11796) );
  OAI21_X1 U14740 ( .B1(n20146), .B2(n11795), .A(n9815), .ZN(n11798) );
  OAI22_X1 U14741 ( .A1(n11813), .A2(n11798), .B1(n11818), .B2(n11797), .ZN(
        n11801) );
  NAND2_X1 U14742 ( .A1(n11799), .A2(n11801), .ZN(n11810) );
  INV_X1 U14743 ( .A(n11800), .ZN(n11802) );
  OAI211_X1 U14744 ( .C1(n11802), .C2(n11801), .A(n12842), .B(n11821), .ZN(
        n11809) );
  XNOR2_X1 U14745 ( .A(n11804), .B(n11803), .ZN(n12841) );
  NAND2_X1 U14746 ( .A1(n11824), .A2(n12841), .ZN(n11806) );
  INV_X1 U14747 ( .A(n11813), .ZN(n11805) );
  OAI211_X1 U14748 ( .C1(n11807), .C2(n12841), .A(n11806), .B(n11805), .ZN(
        n11808) );
  NAND3_X1 U14749 ( .A1(n11810), .A2(n11809), .A3(n11808), .ZN(n11815) );
  INV_X1 U14750 ( .A(n12841), .ZN(n11812) );
  NAND3_X1 U14751 ( .A1(n11813), .A2(n11812), .A3(n11811), .ZN(n11814) );
  AOI22_X1 U14752 ( .A1(n11816), .A2(n12843), .B1(n11815), .B2(n11814), .ZN(
        n11817) );
  AOI21_X1 U14753 ( .B1(n11818), .B2(n12843), .A(n11817), .ZN(n11827) );
  NOR2_X1 U14754 ( .A1(n11824), .A2(n12846), .ZN(n11826) );
  INV_X1 U14755 ( .A(n12846), .ZN(n11823) );
  NAND3_X1 U14756 ( .A1(n11824), .A2(n11823), .A3(n11822), .ZN(n11825) );
  NAND2_X1 U14757 ( .A1(n15551), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19870) );
  NOR2_X1 U14758 ( .A1(n11833), .A2(n20701), .ZN(n20849) );
  NOR2_X1 U14759 ( .A1(n20849), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11830) );
  NAND2_X1 U14760 ( .A1(n20754), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11832) );
  INV_X1 U14761 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n14399) );
  NAND2_X1 U14762 ( .A1(n14399), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11831) );
  NAND2_X1 U14763 ( .A1(n11832), .A2(n11831), .ZN(n20085) );
  AND2_X2 U14764 ( .A1(n11833), .A2(n11268), .ZN(n20128) );
  AOI22_X1 U14765 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_28__SCAN_IN), .ZN(n11834) );
  INV_X1 U14766 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14290) );
  INV_X1 U14767 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14303) );
  INV_X1 U14768 ( .A(n11868), .ZN(n11887) );
  AND2_X1 U14769 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14313) );
  NAND2_X1 U14770 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n14313), .ZN(
        n14299) );
  INV_X1 U14771 ( .A(n14299), .ZN(n14273) );
  INV_X1 U14772 ( .A(n11838), .ZN(n11843) );
  INV_X1 U14773 ( .A(n11839), .ZN(n11844) );
  INV_X1 U14774 ( .A(n11855), .ZN(n11841) );
  AND2_X1 U14775 ( .A1(n11865), .A2(n11859), .ZN(n11875) );
  OR2_X1 U14776 ( .A1(n11840), .A2(n11875), .ZN(n11883) );
  NAND2_X1 U14777 ( .A1(n11884), .A2(n11883), .ZN(n11854) );
  NOR2_X1 U14778 ( .A1(n11841), .A2(n11854), .ZN(n11850) );
  NAND2_X1 U14779 ( .A1(n11850), .A2(n11851), .ZN(n11845) );
  NOR2_X1 U14780 ( .A1(n11844), .A2(n11845), .ZN(n11896) );
  XNOR2_X1 U14781 ( .A(n11895), .B(n11896), .ZN(n11842) );
  OAI22_X1 U14782 ( .A1(n11843), .A2(n11868), .B1(n11842), .B2(n11172), .ZN(
        n11893) );
  NOR2_X1 U14783 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n11893), .ZN(
        n11894) );
  XNOR2_X1 U14784 ( .A(n11845), .B(n11844), .ZN(n11849) );
  NAND3_X1 U14785 ( .A1(n11847), .A2(n11846), .A3(n11887), .ZN(n11848) );
  OAI21_X1 U14786 ( .B1(n11849), .B2(n11172), .A(n11848), .ZN(n13606) );
  NOR2_X1 U14787 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13606), .ZN(
        n11892) );
  INV_X1 U14788 ( .A(n11172), .ZN(n11897) );
  XOR2_X1 U14789 ( .A(n11851), .B(n11850), .Z(n11852) );
  AOI22_X1 U14790 ( .A1(n11853), .A2(n11887), .B1(n11897), .B2(n11852), .ZN(
        n11890) );
  INV_X1 U14791 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15970) );
  NOR2_X1 U14792 ( .A1(n11890), .A2(n15970), .ZN(n11891) );
  XNOR2_X1 U14793 ( .A(n11855), .B(n11854), .ZN(n11856) );
  AOI22_X1 U14794 ( .A1(n11857), .A2(n11887), .B1(n11897), .B2(n11856), .ZN(
        n11889) );
  INV_X1 U14795 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20100) );
  NAND2_X1 U14796 ( .A1(n11858), .A2(n9614), .ZN(n11864) );
  NOR2_X1 U14797 ( .A1(n11865), .A2(n11859), .ZN(n11860) );
  NOR2_X1 U14798 ( .A1(n11860), .A2(n11875), .ZN(n11862) );
  NAND2_X1 U14799 ( .A1(n11776), .A2(n20182), .ZN(n11861) );
  AOI21_X1 U14800 ( .B1(n11862), .B2(n11897), .A(n11861), .ZN(n11863) );
  NAND2_X1 U14801 ( .A1(n11864), .A2(n11863), .ZN(n11871) );
  NAND2_X1 U14802 ( .A1(n20146), .A2(n12906), .ZN(n11876) );
  OAI21_X1 U14803 ( .B1(n11172), .B2(n11865), .A(n11876), .ZN(n11866) );
  INV_X1 U14804 ( .A(n11866), .ZN(n11867) );
  NAND2_X1 U14805 ( .A1(n13028), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11870) );
  INV_X1 U14806 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20135) );
  XNOR2_X1 U14807 ( .A(n11879), .B(n11873), .ZN(n13175) );
  XNOR2_X1 U14808 ( .A(n11875), .B(n11874), .ZN(n11877) );
  OAI21_X1 U14809 ( .B1(n11877), .B2(n11172), .A(n11876), .ZN(n11878) );
  AOI21_X1 U14810 ( .B1(n14390), .B2(n11887), .A(n11878), .ZN(n13176) );
  NOR2_X1 U14811 ( .A1(n13175), .A2(n13176), .ZN(n11881) );
  NOR2_X1 U14812 ( .A1(n11879), .A2(n11873), .ZN(n11880) );
  INV_X1 U14813 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20107) );
  NOR2_X1 U14814 ( .A1(n11882), .A2(n20107), .ZN(n11888) );
  XNOR2_X1 U14815 ( .A(n11884), .B(n11883), .ZN(n11885) );
  NOR2_X1 U14816 ( .A1(n11885), .A2(n11172), .ZN(n11886) );
  AOI21_X1 U14817 ( .B1(n20140), .B2(n11887), .A(n11886), .ZN(n13469) );
  XOR2_X1 U14818 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11889), .Z(
        n20067) );
  XOR2_X1 U14819 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11890), .Z(
        n15838) );
  NAND2_X1 U14820 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13606), .ZN(
        n13605) );
  XNOR2_X1 U14821 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n11893), .ZN(
        n15833) );
  NAND3_X1 U14822 ( .A1(n11897), .A2(n11896), .A3(n11895), .ZN(n11898) );
  INV_X1 U14823 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15957) );
  NAND2_X1 U14824 ( .A1(n14255), .A2(n15957), .ZN(n11899) );
  INV_X1 U14825 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15945) );
  INV_X1 U14826 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15895) );
  INV_X1 U14827 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15916) );
  AOI21_X1 U14828 ( .B1(n15895), .B2(n15916), .A(n15819), .ZN(n14225) );
  INV_X1 U14829 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14268) );
  NAND2_X1 U14830 ( .A1(n15819), .A2(n14268), .ZN(n14234) );
  INV_X1 U14831 ( .A(n14234), .ZN(n14238) );
  AOI21_X1 U14832 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n9618), .ZN(n14237) );
  OAI21_X1 U14833 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n9618), .A(
        n14356), .ZN(n14223) );
  INV_X1 U14834 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15896) );
  AOI22_X1 U14835 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15819), .B1(
        n15825), .B2(n15896), .ZN(n14340) );
  NOR2_X1 U14836 ( .A1(n15825), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14336) );
  NAND2_X1 U14837 ( .A1(n9618), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14235) );
  OAI21_X1 U14838 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n9618), .ZN(n14236) );
  NAND2_X1 U14839 ( .A1(n14235), .A2(n14236), .ZN(n14357) );
  NAND2_X1 U14840 ( .A1(n14224), .A2(n14338), .ZN(n14210) );
  INV_X1 U14841 ( .A(n14210), .ZN(n11903) );
  OAI21_X1 U14842 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(n9618), .ZN(n11902) );
  INV_X1 U14843 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15894) );
  AOI22_X1 U14844 ( .A1(n9618), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n15894), .B2(n15819), .ZN(n15794) );
  NAND2_X1 U14845 ( .A1(n15793), .A2(n15794), .ZN(n14199) );
  NAND3_X1 U14846 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14269) );
  OAI21_X1 U14847 ( .B1(n14199), .B2(n14269), .A(n15819), .ZN(n15774) );
  NAND2_X1 U14848 ( .A1(n15774), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11918) );
  INV_X1 U14849 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15884) );
  INV_X1 U14850 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15596) );
  NAND2_X1 U14851 ( .A1(n14321), .A2(n10147), .ZN(n11906) );
  OAI21_X1 U14852 ( .B1(n9618), .B2(n14273), .A(n14191), .ZN(n11907) );
  NAND2_X1 U14853 ( .A1(n14303), .A2(n11907), .ZN(n11910) );
  NOR2_X1 U14854 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14312) );
  INV_X1 U14855 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15853) );
  NAND2_X1 U14856 ( .A1(n14312), .A2(n15853), .ZN(n11919) );
  INV_X1 U14857 ( .A(n11907), .ZN(n11908) );
  INV_X1 U14858 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14289) );
  AOI21_X1 U14859 ( .B1(n11912), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11911), .ZN(n11913) );
  NAND2_X1 U14860 ( .A1(n11914), .A2(n11913), .ZN(n11915) );
  XOR2_X1 U14861 ( .A(n14290), .B(n11915), .Z(n14288) );
  NAND2_X1 U14862 ( .A1(n11918), .A2(n15819), .ZN(n14180) );
  NAND2_X1 U14863 ( .A1(n11912), .A2(n14163), .ZN(n11922) );
  NAND2_X1 U14864 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14294) );
  INV_X1 U14865 ( .A(n14294), .ZN(n11920) );
  NAND2_X1 U14866 ( .A1(n10148), .A2(n15819), .ZN(n11921) );
  NAND2_X1 U14867 ( .A1(n11922), .A2(n11921), .ZN(n11923) );
  INV_X1 U14868 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14285) );
  XNOR2_X1 U14869 ( .A(n11923), .B(n14285), .ZN(n14281) );
  OAI21_X1 U14870 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n11925), .A(
        n13803), .ZN(n15607) );
  AOI22_X1 U14871 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(n20128), .ZN(n11926) );
  OAI21_X1 U14872 ( .B1(n20075), .B2(n15607), .A(n11926), .ZN(n11927) );
  INV_X1 U14873 ( .A(n11927), .ZN(n11946) );
  AOI22_X1 U14874 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U14875 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U14876 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U14877 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11928) );
  NAND4_X1 U14878 ( .A1(n11931), .A2(n11930), .A3(n11929), .A4(n11928), .ZN(
        n11937) );
  AOI22_X1 U14879 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U14880 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U14881 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U14882 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11932) );
  NAND4_X1 U14883 ( .A1(n11935), .A2(n11934), .A3(n11933), .A4(n11932), .ZN(
        n11936) );
  NOR2_X1 U14884 ( .A1(n11937), .A2(n11936), .ZN(n13793) );
  OR2_X1 U14885 ( .A1(n11939), .A2(n11938), .ZN(n13792) );
  XNOR2_X1 U14886 ( .A(n13793), .B(n13792), .ZN(n11943) );
  NAND2_X1 U14887 ( .A1(n11268), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11940) );
  NAND2_X1 U14888 ( .A1(n13797), .A2(n11940), .ZN(n11941) );
  AOI21_X1 U14889 ( .B1(n13799), .B2(P1_EAX_REG_29__SCAN_IN), .A(n11941), .ZN(
        n11942) );
  OAI21_X1 U14890 ( .B1(n11943), .B2(n13801), .A(n11942), .ZN(n11945) );
  OR2_X1 U14891 ( .A1(n15607), .A2(n13797), .ZN(n11944) );
  XNOR2_X2 U14892 ( .A(n13885), .B(n13888), .ZN(n15744) );
  NAND3_X1 U14893 ( .A1(n11947), .A2(n11946), .A3(n10163), .ZN(P1_U2970) );
  NAND2_X1 U14894 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11959) );
  NAND2_X1 U14895 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11961), .ZN(
        n11960) );
  INV_X1 U14896 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14958) );
  INV_X1 U14897 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11969) );
  AND2_X2 U14898 ( .A1(n11974), .A2(n10149), .ZN(n11976) );
  INV_X1 U14899 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14888) );
  INV_X1 U14900 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18813) );
  NAND2_X1 U14901 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n11978), .ZN(
        n11981) );
  INV_X1 U14902 ( .A(n11981), .ZN(n11948) );
  INV_X1 U14903 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14821) );
  INV_X1 U14904 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16014) );
  INV_X1 U14905 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11986) );
  INV_X1 U14906 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14779) );
  XNOR2_X1 U14907 ( .A(n11949), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13747) );
  INV_X1 U14908 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11950) );
  NAND2_X1 U14909 ( .A1(n11950), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11951) );
  AND2_X4 U14910 ( .A1(n11952), .A2(n11951), .ZN(n18994) );
  OAI21_X1 U14911 ( .B1(n11953), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n11985), .ZN(n16030) );
  OAI21_X1 U14912 ( .B1(n11980), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n11982), .ZN(n16053) );
  OAI21_X1 U14913 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11978), .A(
        n11981), .ZN(n16101) );
  OAI21_X1 U14914 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9730), .A(
        n11979), .ZN(n18832) );
  OAI21_X1 U14915 ( .B1(n11976), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n11977), .ZN(n18855) );
  NAND2_X1 U14916 ( .A1(n11954), .A2(n14958), .ZN(n11955) );
  AND2_X1 U14917 ( .A1(n11970), .A2(n11955), .ZN(n18906) );
  AND2_X1 U14918 ( .A1(n11966), .A2(n14988), .ZN(n11957) );
  AOI21_X1 U14919 ( .B1(n16122), .B2(n11964), .A(n11967), .ZN(n18946) );
  AOI21_X1 U14920 ( .B1(n14997), .B2(n11962), .A(n11965), .ZN(n18963) );
  AOI21_X1 U14921 ( .B1(n16160), .B2(n11960), .A(n11963), .ZN(n18996) );
  AOI21_X1 U14922 ( .B1(n13524), .B2(n11959), .A(n11961), .ZN(n13522) );
  OAI22_X1 U14923 ( .A1(n19855), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19042) );
  INV_X1 U14924 ( .A(n19042), .ZN(n13575) );
  INV_X1 U14925 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U14926 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n11958), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19855), .ZN(n13574) );
  NOR2_X1 U14927 ( .A1(n13575), .A2(n13574), .ZN(n14416) );
  OAI21_X1 U14928 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n11959), .ZN(n14417) );
  NAND2_X1 U14929 ( .A1(n14416), .A2(n14417), .ZN(n13520) );
  NOR2_X1 U14930 ( .A1(n13522), .A2(n13520), .ZN(n19015) );
  OAI21_X1 U14931 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11961), .A(
        n11960), .ZN(n19014) );
  NAND2_X1 U14932 ( .A1(n19015), .A2(n19014), .ZN(n18993) );
  NOR2_X1 U14933 ( .A1(n18996), .A2(n18993), .ZN(n18980) );
  OAI21_X1 U14934 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11963), .A(
        n11962), .ZN(n18981) );
  NAND2_X1 U14935 ( .A1(n18980), .A2(n18981), .ZN(n18962) );
  NOR2_X1 U14936 ( .A1(n18963), .A2(n18962), .ZN(n18955) );
  OAI21_X1 U14937 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n11965), .A(
        n11964), .ZN(n18956) );
  NAND2_X1 U14938 ( .A1(n18955), .A2(n18956), .ZN(n18944) );
  NOR2_X1 U14939 ( .A1(n18946), .A2(n18944), .ZN(n18930) );
  OAI21_X1 U14940 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n11967), .A(
        n11966), .ZN(n18932) );
  NAND2_X1 U14941 ( .A1(n18930), .A2(n18932), .ZN(n18925) );
  NOR2_X1 U14942 ( .A1(n10153), .A2(n18925), .ZN(n18910) );
  OR2_X1 U14943 ( .A1(n11956), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11968) );
  NAND2_X1 U14944 ( .A1(n11954), .A2(n11968), .ZN(n18911) );
  NAND2_X1 U14945 ( .A1(n18910), .A2(n18911), .ZN(n18900) );
  NOR2_X1 U14946 ( .A1(n18906), .A2(n18900), .ZN(n18899) );
  AND2_X1 U14947 ( .A1(n11970), .A2(n11969), .ZN(n11971) );
  OR2_X1 U14948 ( .A1(n11971), .A2(n11972), .ZN(n18893) );
  NAND2_X1 U14949 ( .A1(n18899), .A2(n18893), .ZN(n18882) );
  NOR2_X1 U14950 ( .A1(n11972), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11973) );
  OR2_X1 U14951 ( .A1(n11974), .A2(n11973), .ZN(n14936) );
  INV_X1 U14952 ( .A(n14936), .ZN(n18884) );
  XNOR2_X1 U14953 ( .A(n11974), .B(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n18876) );
  NAND2_X1 U14954 ( .A1(n18994), .A2(n18874), .ZN(n18865) );
  AOI21_X1 U14955 ( .B1(n11974), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11975) );
  OR2_X1 U14956 ( .A1(n11976), .A2(n11975), .ZN(n18866) );
  NAND2_X1 U14957 ( .A1(n18865), .A2(n18866), .ZN(n18864) );
  NAND2_X1 U14958 ( .A1(n18994), .A2(n18864), .ZN(n18854) );
  NAND2_X1 U14959 ( .A1(n18855), .A2(n18854), .ZN(n18853) );
  NAND2_X1 U14960 ( .A1(n18853), .A2(n18994), .ZN(n18842) );
  AOI21_X1 U14961 ( .B1(n14888), .B2(n11977), .A(n9730), .ZN(n14890) );
  INV_X1 U14962 ( .A(n14890), .ZN(n18843) );
  NAND2_X1 U14963 ( .A1(n18842), .A2(n18843), .ZN(n18841) );
  NAND2_X1 U14964 ( .A1(n18994), .A2(n18841), .ZN(n18831) );
  NAND2_X1 U14965 ( .A1(n18832), .A2(n18831), .ZN(n18830) );
  NAND2_X1 U14966 ( .A1(n18830), .A2(n18994), .ZN(n18819) );
  AOI21_X1 U14967 ( .B1(n18813), .B2(n11979), .A(n11978), .ZN(n14862) );
  INV_X1 U14968 ( .A(n14862), .ZN(n18820) );
  NAND2_X1 U14969 ( .A1(n18819), .A2(n18820), .ZN(n18818) );
  NAND2_X1 U14970 ( .A1(n18994), .A2(n18818), .ZN(n15521) );
  NAND2_X1 U14971 ( .A1(n16101), .A2(n15521), .ZN(n15520) );
  NAND2_X1 U14972 ( .A1(n15520), .A2(n18994), .ZN(n16062) );
  INV_X1 U14973 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14841) );
  AOI21_X1 U14974 ( .B1(n14841), .B2(n11981), .A(n11980), .ZN(n14843) );
  INV_X1 U14975 ( .A(n14843), .ZN(n16063) );
  NAND2_X1 U14976 ( .A1(n16062), .A2(n16063), .ZN(n16061) );
  NAND2_X1 U14977 ( .A1(n18994), .A2(n16061), .ZN(n16052) );
  NAND2_X1 U14978 ( .A1(n16053), .A2(n16052), .ZN(n16051) );
  NAND2_X1 U14979 ( .A1(n16051), .A2(n18994), .ZN(n16040) );
  AND2_X1 U14980 ( .A1(n11982), .A2(n14821), .ZN(n11983) );
  NOR2_X1 U14981 ( .A1(n11953), .A2(n11983), .ZN(n14819) );
  INV_X1 U14982 ( .A(n14819), .ZN(n16041) );
  NAND2_X1 U14983 ( .A1(n16040), .A2(n16041), .ZN(n16039) );
  NAND2_X1 U14984 ( .A1(n18994), .A2(n16039), .ZN(n16029) );
  NAND2_X1 U14985 ( .A1(n16030), .A2(n16029), .ZN(n16028) );
  NAND2_X1 U14986 ( .A1(n16028), .A2(n18994), .ZN(n16020) );
  INV_X1 U14987 ( .A(n11987), .ZN(n11984) );
  AOI21_X1 U14988 ( .B1(n16014), .B2(n11985), .A(n11984), .ZN(n14799) );
  INV_X1 U14989 ( .A(n14799), .ZN(n16021) );
  NAND2_X1 U14990 ( .A1(n16020), .A2(n16021), .ZN(n16019) );
  NAND2_X1 U14991 ( .A1(n18994), .A2(n16019), .ZN(n16007) );
  NAND2_X1 U14992 ( .A1(n11987), .A2(n11986), .ZN(n11988) );
  NAND2_X1 U14993 ( .A1(n11989), .A2(n11988), .ZN(n16008) );
  NAND2_X1 U14994 ( .A1(n16007), .A2(n16008), .ZN(n16006) );
  NAND2_X1 U14995 ( .A1(n16006), .A2(n18994), .ZN(n15997) );
  AOI21_X1 U14996 ( .B1(n14779), .B2(n11989), .A(n11990), .ZN(n14781) );
  INV_X1 U14997 ( .A(n14781), .ZN(n15998) );
  XNOR2_X1 U14998 ( .A(n11990), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15983) );
  NAND2_X1 U14999 ( .A1(n15982), .A2(n15983), .ZN(n11991) );
  INV_X1 U15000 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19844) );
  NOR4_X1 U15001 ( .A1(n19844), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATEBS16_REG_SCAN_IN), .A4(P2_STATE2_REG_2__SCAN_IN), .ZN(n14419)
         );
  INV_X1 U15002 ( .A(n14419), .ZN(n19705) );
  INV_X1 U15003 ( .A(n19705), .ZN(n19000) );
  INV_X1 U15004 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n14904) );
  AOI22_X1 U15005 ( .A1(n13756), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11992) );
  OAI21_X1 U15006 ( .B1(n10870), .B2(n14904), .A(n11992), .ZN(n11993) );
  INV_X1 U15007 ( .A(n11993), .ZN(n15172) );
  INV_X1 U15008 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19756) );
  AOI22_X1 U15009 ( .A1(n13756), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11994) );
  OAI21_X1 U15010 ( .B1(n10870), .B2(n19756), .A(n11994), .ZN(n14745) );
  INV_X1 U15011 ( .A(n14745), .ZN(n11995) );
  INV_X1 U15012 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19758) );
  AOI22_X1 U15013 ( .A1(n13756), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11996) );
  OAI21_X1 U15014 ( .B1(n10870), .B2(n19758), .A(n11996), .ZN(n15141) );
  INV_X1 U15015 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14860) );
  INV_X1 U15016 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n12871) );
  INV_X1 U15017 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19760) );
  OAI222_X1 U15018 ( .A1(n14860), .A2(n11998), .B1(n11997), .B2(n12871), .C1(
        n10870), .C2(n19760), .ZN(n14740) );
  NAND2_X1 U15019 ( .A1(n11999), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15020 ( .A1(n13756), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12000) );
  AND2_X1 U15021 ( .A1(n12001), .A2(n12000), .ZN(n14732) );
  INV_X1 U15022 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19763) );
  AOI22_X1 U15023 ( .A1(n13756), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12002) );
  OAI21_X1 U15024 ( .B1(n10870), .B2(n19763), .A(n12002), .ZN(n14721) );
  INV_X1 U15025 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n14832) );
  AOI22_X1 U15026 ( .A1(n13756), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12003) );
  OAI21_X1 U15027 ( .B1(n10870), .B2(n14832), .A(n12003), .ZN(n14714) );
  NAND2_X1 U15028 ( .A1(n11999), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U15029 ( .A1(n10810), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12004) );
  AND2_X1 U15030 ( .A1(n12005), .A2(n12004), .ZN(n14702) );
  INV_X1 U15031 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19768) );
  AOI22_X1 U15032 ( .A1(n10810), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12006) );
  OAI21_X1 U15033 ( .B1(n10870), .B2(n19768), .A(n12006), .ZN(n14694) );
  NAND2_X1 U15034 ( .A1(n11999), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U15035 ( .A1(n13756), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12007) );
  AND2_X1 U15036 ( .A1(n12008), .A2(n12007), .ZN(n14683) );
  NAND2_X1 U15037 ( .A1(n11999), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15038 ( .A1(n10810), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12009) );
  AND2_X1 U15039 ( .A1(n12010), .A2(n12009), .ZN(n14672) );
  NAND2_X1 U15040 ( .A1(n11999), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15041 ( .A1(n10810), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12011) );
  AND2_X1 U15042 ( .A1(n12012), .A2(n12011), .ZN(n14518) );
  INV_X1 U15043 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19777) );
  AOI22_X1 U15044 ( .A1(n10810), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n10823), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12013) );
  OAI21_X1 U15045 ( .B1(n10870), .B2(n19777), .A(n12013), .ZN(n12014) );
  NAND2_X1 U15046 ( .A1(n14520), .A2(n12014), .ZN(n13759) );
  OR2_X1 U15047 ( .A1(n14520), .A2(n12014), .ZN(n12015) );
  INV_X1 U15048 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19797) );
  NAND2_X1 U15049 ( .A1(n13371), .A2(n19797), .ZN(n13382) );
  INV_X1 U15050 ( .A(n13382), .ZN(n16213) );
  AND2_X1 U15051 ( .A1(n12016), .A2(n16213), .ZN(n12017) );
  AND2_X1 U15052 ( .A1(n19180), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13677) );
  NAND2_X1 U15053 ( .A1(n19180), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12018) );
  AND2_X1 U15054 ( .A1(n19180), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n13698) );
  INV_X1 U15055 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n12054) );
  INV_X1 U15056 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14466) );
  NAND2_X1 U15057 ( .A1(n13712), .A2(n12019), .ZN(n13731) );
  NAND2_X1 U15058 ( .A1(n19180), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13666) );
  NAND2_X1 U15059 ( .A1(n19180), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n13723) );
  AND2_X1 U15060 ( .A1(n19180), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13725) );
  AND2_X1 U15061 ( .A1(n19180), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12020) );
  XNOR2_X1 U15062 ( .A(n13732), .B(n12020), .ZN(n13727) );
  NAND2_X1 U15063 ( .A1(n13338), .A2(n19700), .ZN(n12021) );
  OR2_X1 U15064 ( .A1(n16215), .A2(n12021), .ZN(n12718) );
  AND2_X1 U15065 ( .A1(n19850), .A2(n19797), .ZN(n12022) );
  NOR2_X1 U15066 ( .A1(n12718), .A2(n12022), .ZN(n12026) );
  AND2_X1 U15067 ( .A1(n12026), .A2(n15338), .ZN(n15984) );
  NOR2_X1 U15068 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19587), .ZN(n19378) );
  NAND2_X1 U15069 ( .A1(n12023), .A2(n19378), .ZN(n16222) );
  NAND3_X1 U15070 ( .A1(n18966), .A2(n16222), .A3(n19705), .ZN(n12024) );
  OAI22_X1 U15071 ( .A1(n13727), .A2(n18989), .B1(n19777), .B2(n19004), .ZN(
        n12030) );
  AND2_X1 U15072 ( .A1(n12809), .A2(n13382), .ZN(n15986) );
  INV_X1 U15073 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12025) );
  AND2_X1 U15074 ( .A1(n12026), .A2(n12025), .ZN(n12027) );
  AOI22_X1 U15075 ( .A1(n19028), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19038), .ZN(n12028) );
  INV_X1 U15076 ( .A(n12028), .ZN(n12029) );
  AOI211_X1 U15077 ( .C1(n9658), .C2(n19008), .A(n12030), .B(n12029), .ZN(
        n12078) );
  INV_X1 U15078 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n12033) );
  NAND2_X1 U15079 ( .A1(n12065), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12032) );
  NAND2_X1 U15080 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12031) );
  OAI211_X1 U15081 ( .C1(n12033), .C2(n12069), .A(n12032), .B(n12031), .ZN(
        n12034) );
  AOI21_X1 U15082 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n12034), .ZN(n14900) );
  NAND2_X1 U15083 ( .A1(n13743), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12036) );
  AOI22_X1 U15084 ( .A1(n13739), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n12035) );
  OAI211_X1 U15085 ( .C1(n13741), .C2(n19756), .A(n12036), .B(n12035), .ZN(
        n14491) );
  NAND2_X1 U15086 ( .A1(n13743), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12038) );
  AOI22_X1 U15087 ( .A1(n13739), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12037) );
  OAI211_X1 U15088 ( .C1(n13741), .C2(n19758), .A(n12038), .B(n12037), .ZN(
        n14874) );
  INV_X1 U15089 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12041) );
  NAND2_X1 U15090 ( .A1(n12065), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12040) );
  NAND2_X1 U15091 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12039) );
  OAI211_X1 U15092 ( .C1(n12069), .C2(n12041), .A(n12040), .B(n12039), .ZN(
        n12042) );
  AOI21_X1 U15093 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12042), .ZN(n14487) );
  INV_X1 U15094 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12045) );
  NAND2_X1 U15095 ( .A1(n13743), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12044) );
  AOI22_X1 U15096 ( .A1(n13739), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n12043) );
  OAI211_X1 U15097 ( .C1(n13741), .C2(n12045), .A(n12044), .B(n12043), .ZN(
        n15110) );
  NAND2_X1 U15098 ( .A1(n13743), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12051) );
  INV_X1 U15099 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12048) );
  NAND2_X1 U15100 ( .A1(n12065), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12047) );
  NAND2_X1 U15101 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12046) );
  OAI211_X1 U15102 ( .C1(n12069), .C2(n12048), .A(n12047), .B(n12046), .ZN(
        n12049) );
  INV_X1 U15103 ( .A(n12049), .ZN(n12050) );
  NAND2_X1 U15104 ( .A1(n12051), .A2(n12050), .ZN(n14474) );
  NAND2_X1 U15105 ( .A1(n12065), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12053) );
  NAND2_X1 U15106 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12052) );
  OAI211_X1 U15107 ( .C1(n12069), .C2(n12054), .A(n12053), .B(n12052), .ZN(
        n12055) );
  AOI21_X1 U15108 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12055), .ZN(n14469) );
  NAND2_X1 U15109 ( .A1(n12065), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12057) );
  NAND2_X1 U15110 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12056) );
  OAI211_X1 U15111 ( .C1(n12069), .C2(n14466), .A(n12057), .B(n12056), .ZN(
        n12058) );
  AOI21_X1 U15112 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12058), .ZN(n14464) );
  NAND2_X1 U15113 ( .A1(n13743), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12060) );
  AOI22_X1 U15114 ( .A1(n13739), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12059) );
  OAI211_X1 U15115 ( .C1(n13741), .C2(n19768), .A(n12060), .B(n12059), .ZN(
        n14455) );
  INV_X1 U15116 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12063) );
  NAND2_X1 U15117 ( .A1(n12065), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12062) );
  NAND2_X1 U15118 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12061) );
  OAI211_X1 U15119 ( .C1(n12069), .C2(n12063), .A(n12062), .B(n12061), .ZN(
        n12064) );
  AOI21_X1 U15120 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12064), .ZN(n14449) );
  INV_X1 U15121 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12068) );
  NAND2_X1 U15122 ( .A1(n12065), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12067) );
  NAND2_X1 U15123 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12066) );
  OAI211_X1 U15124 ( .C1(n12069), .C2(n12068), .A(n12067), .B(n12066), .ZN(
        n12070) );
  AOI21_X1 U15125 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12070), .ZN(n14437) );
  INV_X1 U15126 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19774) );
  NAND2_X1 U15127 ( .A1(n13743), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12072) );
  AOI22_X1 U15128 ( .A1(n13739), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12071) );
  OAI211_X1 U15129 ( .C1(n13741), .C2(n19774), .A(n12072), .B(n12071), .ZN(
        n14429) );
  NAND2_X1 U15130 ( .A1(n14439), .A2(n14429), .ZN(n14431) );
  AOI22_X1 U15131 ( .A1(n13739), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12073) );
  OAI21_X1 U15132 ( .B1(n13741), .B2(n19777), .A(n12073), .ZN(n12074) );
  AOI21_X1 U15133 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12074), .ZN(n13738) );
  INV_X1 U15134 ( .A(n15020), .ZN(n12076) );
  NAND2_X1 U15135 ( .A1(n15338), .A2(n19850), .ZN(n12075) );
  NAND2_X1 U15136 ( .A1(n12080), .A2(n12079), .ZN(P2_U2825) );
  NAND2_X1 U15137 ( .A1(n14425), .A2(n12098), .ZN(n12085) );
  NAND2_X1 U15138 ( .A1(n10362), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12081) );
  NAND2_X1 U15139 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19511) );
  NAND2_X1 U15140 ( .A1(n19511), .A2(n19813), .ZN(n12083) );
  NAND2_X1 U15141 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15367) );
  INV_X1 U15142 ( .A(n15367), .ZN(n12082) );
  NAND2_X1 U15143 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12082), .ZN(
        n12100) );
  AND2_X1 U15144 ( .A1(n12083), .A2(n12100), .ZN(n19284) );
  AOI22_X1 U15145 ( .A1(n12104), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19806), .B2(n19284), .ZN(n12084) );
  NAND2_X1 U15146 ( .A1(n12085), .A2(n12084), .ZN(n12087) );
  NAND3_X1 U15147 ( .A1(n19188), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n15338), 
        .ZN(n12112) );
  INV_X1 U15148 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19170) );
  NOR2_X1 U15149 ( .A1(n12112), .A2(n19170), .ZN(n12086) );
  OR2_X1 U15150 ( .A1(n12087), .A2(n12086), .ZN(n12088) );
  NAND2_X1 U15151 ( .A1(n12087), .A2(n12086), .ZN(n12097) );
  NAND2_X1 U15152 ( .A1(n12088), .A2(n12097), .ZN(n12966) );
  NAND2_X1 U15153 ( .A1(n12104), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12090) );
  NAND2_X1 U15154 ( .A1(n19821), .A2(n19830), .ZN(n19405) );
  NAND2_X1 U15155 ( .A1(n19511), .A2(n19405), .ZN(n19283) );
  INV_X1 U15156 ( .A(n19283), .ZN(n12089) );
  NAND2_X1 U15157 ( .A1(n12089), .A2(n19806), .ZN(n19481) );
  NAND2_X1 U15158 ( .A1(n12090), .A2(n19481), .ZN(n12091) );
  INV_X1 U15159 ( .A(n12098), .ZN(n12885) );
  AOI22_X1 U15160 ( .A1(n12104), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19806), .B2(n19830), .ZN(n12092) );
  OAI21_X2 U15161 ( .B1(n19023), .B2(n12885), .A(n12092), .ZN(n12093) );
  INV_X1 U15162 ( .A(n12112), .ZN(n12317) );
  NAND2_X1 U15163 ( .A1(n12317), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12094) );
  NAND2_X1 U15164 ( .A1(n12923), .A2(n12922), .ZN(n12096) );
  NAND2_X1 U15165 ( .A1(n13560), .A2(n12094), .ZN(n12095) );
  OAI21_X2 U15166 ( .B1(n12966), .B2(n12967), .A(n12097), .ZN(n13227) );
  INV_X1 U15167 ( .A(n12100), .ZN(n12101) );
  NAND2_X1 U15168 ( .A1(n12101), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19660) );
  OAI211_X1 U15169 ( .C1(n12101), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19660), .B(n19806), .ZN(n12102) );
  INV_X1 U15170 ( .A(n12102), .ZN(n12103) );
  AOI21_X1 U15171 ( .B1(n12104), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12103), .ZN(n12105) );
  NOR2_X1 U15172 ( .A1(n12112), .A2(n19176), .ZN(n12106) );
  NAND2_X1 U15173 ( .A1(n12107), .A2(n12106), .ZN(n12110) );
  AND2_X2 U15174 ( .A1(n12108), .A2(n12110), .ZN(n13229) );
  NAND2_X1 U15175 ( .A1(n10362), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12109) );
  INV_X1 U15176 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19179) );
  NOR2_X1 U15177 ( .A1(n12112), .A2(n19179), .ZN(n13392) );
  AND2_X2 U15178 ( .A1(n13391), .A2(n13392), .ZN(n19073) );
  INV_X1 U15179 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15351) );
  NAND2_X1 U15180 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13122) );
  NOR2_X1 U15181 ( .A1(n15351), .A2(n13122), .ZN(n19072) );
  AND2_X2 U15182 ( .A1(n19054), .A2(n19053), .ZN(n13289) );
  AOI22_X1 U15183 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15184 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U15185 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12186), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15186 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12114) );
  NAND4_X1 U15187 ( .A1(n12117), .A2(n12116), .A3(n12115), .A4(n12114), .ZN(
        n12123) );
  AOI22_X1 U15188 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15189 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U15190 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15191 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12118) );
  NAND4_X1 U15192 ( .A1(n12121), .A2(n12120), .A3(n12119), .A4(n12118), .ZN(
        n12122) );
  OR2_X1 U15193 ( .A1(n12123), .A2(n12122), .ZN(n14500) );
  AOI22_X1 U15194 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15195 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12126) );
  AOI22_X1 U15196 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12186), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15197 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12124) );
  NAND4_X1 U15198 ( .A1(n12127), .A2(n12126), .A3(n12125), .A4(n12124), .ZN(
        n12133) );
  AOI22_X1 U15199 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15200 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15201 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15202 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12128) );
  NAND4_X1 U15203 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12132) );
  NOR2_X1 U15204 ( .A1(n12133), .A2(n12132), .ZN(n19045) );
  OR2_X1 U15205 ( .A1(n13460), .A2(n19049), .ZN(n13461) );
  NOR2_X1 U15206 ( .A1(n19045), .A2(n13461), .ZN(n14499) );
  AND2_X1 U15207 ( .A1(n14500), .A2(n14499), .ZN(n12134) );
  AOI22_X1 U15208 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10524), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15209 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15210 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n12186), .ZN(n12136) );
  AOI22_X1 U15211 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n13295), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12135) );
  NAND4_X1 U15212 ( .A1(n12138), .A2(n12137), .A3(n12136), .A4(n12135), .ZN(
        n12144) );
  AOI22_X1 U15213 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n10537), .ZN(n12142) );
  AOI22_X1 U15214 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15215 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15216 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12139) );
  NAND4_X1 U15217 ( .A1(n12142), .A2(n12141), .A3(n12140), .A4(n12139), .ZN(
        n12143) );
  NOR2_X1 U15218 ( .A1(n12144), .A2(n12143), .ZN(n16079) );
  INV_X1 U15219 ( .A(n16079), .ZN(n12145) );
  AOI22_X1 U15220 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10601), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15221 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15222 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n12186), .ZN(n12147) );
  AOI22_X1 U15223 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n13295), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12146) );
  NAND4_X1 U15224 ( .A1(n12149), .A2(n12148), .A3(n12147), .A4(n12146), .ZN(
        n12155) );
  AOI22_X1 U15225 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .B2(n10537), .ZN(n12153) );
  AOI22_X1 U15226 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15227 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15228 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12150) );
  NAND4_X1 U15229 ( .A1(n12153), .A2(n12152), .A3(n12151), .A4(n12150), .ZN(
        n12154) );
  NOR2_X1 U15230 ( .A1(n12155), .A2(n12154), .ZN(n14495) );
  AOI22_X1 U15231 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10601), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15232 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15233 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n12186), .ZN(n12157) );
  AOI22_X1 U15234 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13295), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12156) );
  NAND4_X1 U15235 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n12156), .ZN(
        n12165) );
  AOI22_X1 U15236 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n10537), .ZN(n12163) );
  AOI22_X1 U15237 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15238 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15239 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12160) );
  NAND4_X1 U15240 ( .A1(n12163), .A2(n12162), .A3(n12161), .A4(n12160), .ZN(
        n12164) );
  OR2_X1 U15241 ( .A1(n12165), .A2(n12164), .ZN(n16073) );
  AOI22_X1 U15242 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15243 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15244 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12186), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15245 ( .A1(n13295), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12166) );
  NAND4_X1 U15246 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n12175) );
  AOI22_X1 U15247 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10537), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15248 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15249 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15250 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12170) );
  NAND4_X1 U15251 ( .A1(n12173), .A2(n12172), .A3(n12171), .A4(n12170), .ZN(
        n12174) );
  OR2_X1 U15252 ( .A1(n12175), .A2(n12174), .ZN(n14485) );
  NAND2_X1 U15253 ( .A1(n14484), .A2(n14485), .ZN(n14483) );
  AOI22_X1 U15254 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10601), .B1(
        n10524), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15255 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15256 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n12186), .ZN(n12177) );
  AOI22_X1 U15257 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n13295), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12176) );
  NAND4_X1 U15258 ( .A1(n12179), .A2(n12178), .A3(n12177), .A4(n12176), .ZN(
        n12185) );
  AOI22_X1 U15259 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__6__SCAN_IN), .B2(n10537), .ZN(n12183) );
  AOI22_X1 U15260 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15261 ( .A1(n10523), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15262 ( .A1(n10544), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12180) );
  NAND4_X1 U15263 ( .A1(n12183), .A2(n12182), .A3(n12181), .A4(n12180), .ZN(
        n12184) );
  NOR2_X1 U15264 ( .A1(n12185), .A2(n12184), .ZN(n14730) );
  OR2_X2 U15265 ( .A1(n14483), .A2(n14730), .ZN(n12218) );
  AOI22_X1 U15266 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10523), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15267 ( .A1(n10490), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15268 ( .A1(n10536), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n12186), .ZN(n12188) );
  AOI22_X1 U15269 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n13295), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12187) );
  NAND4_X1 U15270 ( .A1(n12190), .A2(n12189), .A3(n12188), .A4(n12187), .ZN(
        n12196) );
  AOI22_X1 U15271 ( .A1(n10496), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n10544), .ZN(n12194) );
  AOI22_X1 U15272 ( .A1(n10497), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15273 ( .A1(n10524), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15274 ( .A1(n10537), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12191) );
  NAND4_X1 U15275 ( .A1(n12194), .A2(n12193), .A3(n12192), .A4(n12191), .ZN(
        n12195) );
  NOR2_X1 U15276 ( .A1(n12196), .A2(n12195), .ZN(n12242) );
  INV_X1 U15277 ( .A(n12382), .ZN(n12354) );
  INV_X1 U15278 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12198) );
  INV_X1 U15279 ( .A(n12381), .ZN(n12352) );
  INV_X1 U15280 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12197) );
  OAI22_X1 U15281 ( .A1(n12354), .A2(n12198), .B1(n12352), .B2(n12197), .ZN(
        n12203) );
  INV_X1 U15282 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12201) );
  INV_X1 U15283 ( .A(n12383), .ZN(n12356) );
  INV_X1 U15284 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12200) );
  OAI22_X1 U15285 ( .A1(n12199), .A2(n12201), .B1(n12356), .B2(n12200), .ZN(
        n12202) );
  NOR2_X1 U15286 ( .A1(n12203), .A2(n12202), .ZN(n12206) );
  AOI22_X1 U15287 ( .A1(n12370), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10314), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12205) );
  INV_X1 U15288 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n19228) );
  AOI22_X1 U15289 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12204) );
  XNOR2_X1 U15290 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12373) );
  NAND4_X1 U15291 ( .A1(n12206), .A2(n12205), .A3(n12204), .A4(n12373), .ZN(
        n12216) );
  INV_X1 U15292 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12208) );
  INV_X1 U15293 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12207) );
  OAI22_X1 U15294 ( .A1(n12354), .A2(n12208), .B1(n12352), .B2(n12207), .ZN(
        n12211) );
  INV_X1 U15295 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12209) );
  INV_X1 U15296 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13547) );
  OAI22_X1 U15297 ( .A1(n12199), .A2(n12209), .B1(n12356), .B2(n13547), .ZN(
        n12210) );
  NOR2_X1 U15298 ( .A1(n12211), .A2(n12210), .ZN(n12214) );
  INV_X1 U15299 ( .A(n12373), .ZN(n12384) );
  AOI22_X1 U15300 ( .A1(n12370), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10314), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15301 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12212) );
  NAND4_X1 U15302 ( .A1(n12214), .A2(n12384), .A3(n12213), .A4(n12212), .ZN(
        n12215) );
  NAND2_X1 U15303 ( .A1(n12216), .A2(n12215), .ZN(n12217) );
  NOR2_X1 U15304 ( .A1(n19852), .A2(n12217), .ZN(n12222) );
  XOR2_X1 U15305 ( .A(n12242), .B(n12222), .Z(n12219) );
  XNOR2_X2 U15306 ( .A(n12218), .B(n12219), .ZN(n14479) );
  INV_X1 U15307 ( .A(n12217), .ZN(n12244) );
  NAND2_X1 U15308 ( .A1(n19852), .A2(n12244), .ZN(n14478) );
  INV_X1 U15309 ( .A(n12219), .ZN(n12220) );
  INV_X1 U15310 ( .A(n12222), .ZN(n12241) );
  INV_X1 U15311 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12223) );
  INV_X1 U15312 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15344) );
  OAI22_X1 U15313 ( .A1(n12354), .A2(n12223), .B1(n12352), .B2(n15344), .ZN(
        n12227) );
  INV_X1 U15314 ( .A(n10314), .ZN(n12358) );
  INV_X1 U15315 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12224) );
  OAI22_X1 U15316 ( .A1(n12358), .A2(n12225), .B1(n12356), .B2(n12224), .ZN(
        n12226) );
  NOR2_X1 U15317 ( .A1(n12227), .A2(n12226), .ZN(n12230) );
  AOI22_X1 U15318 ( .A1(n12370), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15319 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12228) );
  NAND4_X1 U15320 ( .A1(n12230), .A2(n12229), .A3(n12228), .A4(n12373), .ZN(
        n12240) );
  INV_X1 U15321 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12232) );
  INV_X1 U15322 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12231) );
  OAI22_X1 U15323 ( .A1(n12354), .A2(n12232), .B1(n12352), .B2(n12231), .ZN(
        n12235) );
  INV_X1 U15324 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12233) );
  OAI22_X1 U15325 ( .A1(n12199), .A2(n12233), .B1(n12356), .B2(n19658), .ZN(
        n12234) );
  NOR2_X1 U15326 ( .A1(n12235), .A2(n12234), .ZN(n12238) );
  INV_X1 U15327 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n19627) );
  AOI22_X1 U15328 ( .A1(n12370), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10314), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15329 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12236) );
  NAND4_X1 U15330 ( .A1(n12238), .A2(n12384), .A3(n12237), .A4(n12236), .ZN(
        n12239) );
  NAND2_X1 U15331 ( .A1(n12240), .A2(n12239), .ZN(n12243) );
  OAI21_X1 U15332 ( .B1(n12242), .B2(n12241), .A(n12243), .ZN(n12247) );
  INV_X1 U15333 ( .A(n12242), .ZN(n12245) );
  INV_X1 U15334 ( .A(n12243), .ZN(n12246) );
  NAND3_X1 U15335 ( .A1(n12245), .A2(n12246), .A3(n12244), .ZN(n12248) );
  AOI22_X1 U15336 ( .A1(n12247), .A2(n12248), .B1(n12246), .B2(n19852), .ZN(
        n14468) );
  INV_X1 U15337 ( .A(n12248), .ZN(n12267) );
  INV_X1 U15338 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12249) );
  OAI22_X1 U15339 ( .A1(n12354), .A2(n12249), .B1(n12352), .B2(n19170), .ZN(
        n12253) );
  INV_X1 U15340 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12251) );
  INV_X1 U15341 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12250) );
  OAI22_X1 U15342 ( .A1(n12358), .A2(n12251), .B1(n12356), .B2(n12250), .ZN(
        n12252) );
  NOR2_X1 U15343 ( .A1(n12253), .A2(n12252), .ZN(n12256) );
  AOI22_X1 U15344 ( .A1(n12370), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15345 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12254) );
  NAND4_X1 U15346 ( .A1(n12256), .A2(n12255), .A3(n12254), .A4(n12373), .ZN(
        n12266) );
  INV_X1 U15347 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12258) );
  INV_X1 U15348 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12257) );
  OAI22_X1 U15349 ( .A1(n12354), .A2(n12258), .B1(n12352), .B2(n12257), .ZN(
        n12261) );
  INV_X1 U15350 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12259) );
  INV_X1 U15351 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13573) );
  OAI22_X1 U15352 ( .A1(n12199), .A2(n12259), .B1(n12356), .B2(n13573), .ZN(
        n12260) );
  NOR2_X1 U15353 ( .A1(n12261), .A2(n12260), .ZN(n12264) );
  INV_X1 U15354 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19633) );
  AOI22_X1 U15355 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10314), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15356 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12262) );
  NAND4_X1 U15357 ( .A1(n12264), .A2(n12384), .A3(n12263), .A4(n12262), .ZN(
        n12265) );
  AND2_X1 U15358 ( .A1(n12266), .A2(n12265), .ZN(n12268) );
  NAND2_X1 U15359 ( .A1(n12267), .A2(n12268), .ZN(n12297) );
  OAI211_X1 U15360 ( .C1(n12267), .C2(n12268), .A(n12317), .B(n12297), .ZN(
        n12271) );
  INV_X1 U15361 ( .A(n12268), .ZN(n12269) );
  NOR2_X1 U15362 ( .A1(n15338), .A2(n12269), .ZN(n14462) );
  INV_X1 U15363 ( .A(n12270), .ZN(n14711) );
  OAI22_X1 U15364 ( .A1(n12354), .A2(n12274), .B1(n12352), .B2(n19176), .ZN(
        n12278) );
  INV_X1 U15365 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12276) );
  OAI22_X1 U15366 ( .A1(n12358), .A2(n12276), .B1(n12356), .B2(n12275), .ZN(
        n12277) );
  NOR2_X1 U15367 ( .A1(n12278), .A2(n12277), .ZN(n12281) );
  AOI22_X1 U15368 ( .A1(n12370), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15369 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12279) );
  NAND4_X1 U15370 ( .A1(n12281), .A2(n12280), .A3(n12279), .A4(n12373), .ZN(
        n12291) );
  OAI22_X1 U15371 ( .A1(n12354), .A2(n12283), .B1(n12352), .B2(n12282), .ZN(
        n12286) );
  INV_X1 U15372 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12284) );
  OAI22_X1 U15373 ( .A1(n12358), .A2(n12284), .B1(n12356), .B2(n19668), .ZN(
        n12285) );
  NOR2_X1 U15374 ( .A1(n12286), .A2(n12285), .ZN(n12289) );
  AOI22_X1 U15375 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12376), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15376 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12287) );
  NAND4_X1 U15377 ( .A1(n12289), .A2(n12384), .A3(n12288), .A4(n12287), .ZN(
        n12290) );
  AND2_X1 U15378 ( .A1(n12291), .A2(n12290), .ZN(n12295) );
  XNOR2_X1 U15379 ( .A(n12297), .B(n12295), .ZN(n12292) );
  NAND2_X1 U15380 ( .A1(n19852), .A2(n12295), .ZN(n14457) );
  INV_X1 U15381 ( .A(n12295), .ZN(n12296) );
  NOR2_X1 U15382 ( .A1(n12297), .A2(n12296), .ZN(n12318) );
  INV_X1 U15383 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12298) );
  OAI22_X1 U15384 ( .A1(n12354), .A2(n12298), .B1(n12352), .B2(n19179), .ZN(
        n12302) );
  INV_X1 U15385 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12300) );
  INV_X1 U15386 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12299) );
  OAI22_X1 U15387 ( .A1(n12358), .A2(n12300), .B1(n12356), .B2(n12299), .ZN(
        n12301) );
  NOR2_X1 U15388 ( .A1(n12302), .A2(n12301), .ZN(n12305) );
  AOI22_X1 U15389 ( .A1(n12370), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12376), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15390 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12303) );
  NAND4_X1 U15391 ( .A1(n12305), .A2(n12304), .A3(n12303), .A4(n12373), .ZN(
        n12316) );
  INV_X1 U15392 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12307) );
  INV_X1 U15393 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12306) );
  OAI22_X1 U15394 ( .A1(n12354), .A2(n12307), .B1(n12352), .B2(n12306), .ZN(
        n12311) );
  INV_X1 U15395 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12309) );
  INV_X1 U15396 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12308) );
  OAI22_X1 U15397 ( .A1(n12358), .A2(n12309), .B1(n12356), .B2(n12308), .ZN(
        n12310) );
  NOR2_X1 U15398 ( .A1(n12311), .A2(n12310), .ZN(n12314) );
  AOI22_X1 U15399 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15400 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12312) );
  NAND4_X1 U15401 ( .A1(n12314), .A2(n12384), .A3(n12313), .A4(n12312), .ZN(
        n12315) );
  AND2_X1 U15402 ( .A1(n12316), .A2(n12315), .ZN(n12321) );
  NAND2_X1 U15403 ( .A1(n12318), .A2(n12321), .ZN(n14440) );
  OAI211_X1 U15404 ( .C1(n12318), .C2(n12321), .A(n14440), .B(n12317), .ZN(
        n12319) );
  AOI21_X2 U15405 ( .B1(n12320), .B2(n12319), .A(n12323), .ZN(n14448) );
  INV_X1 U15406 ( .A(n12321), .ZN(n12322) );
  NOR2_X1 U15407 ( .A1(n15338), .A2(n12322), .ZN(n14447) );
  NAND2_X1 U15408 ( .A1(n14448), .A2(n14447), .ZN(n14446) );
  INV_X1 U15409 ( .A(n12323), .ZN(n14441) );
  OAI22_X1 U15410 ( .A1(n12354), .A2(n12324), .B1(n12352), .B2(n13121), .ZN(
        n12328) );
  INV_X1 U15411 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12326) );
  OAI22_X1 U15412 ( .A1(n12358), .A2(n12326), .B1(n12356), .B2(n12325), .ZN(
        n12327) );
  NOR2_X1 U15413 ( .A1(n12328), .A2(n12327), .ZN(n12331) );
  AOI22_X1 U15414 ( .A1(n12370), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12376), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15415 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12329) );
  NAND4_X1 U15416 ( .A1(n12331), .A2(n12330), .A3(n12329), .A4(n12373), .ZN(
        n12342) );
  OAI22_X1 U15417 ( .A1(n12354), .A2(n12333), .B1(n12352), .B2(n12332), .ZN(
        n12337) );
  INV_X1 U15418 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12335) );
  OAI22_X1 U15419 ( .A1(n12358), .A2(n12335), .B1(n12356), .B2(n12334), .ZN(
        n12336) );
  NOR2_X1 U15420 ( .A1(n12337), .A2(n12336), .ZN(n12340) );
  AOI22_X1 U15421 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15422 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12338) );
  NAND4_X1 U15423 ( .A1(n12340), .A2(n12384), .A3(n12339), .A4(n12338), .ZN(
        n12341) );
  NAND2_X1 U15424 ( .A1(n12342), .A2(n12341), .ZN(n14442) );
  AOI21_X2 U15425 ( .B1(n14446), .B2(n14441), .A(n14442), .ZN(n14433) );
  OAI22_X1 U15426 ( .A1(n12354), .A2(n12343), .B1(n12352), .B2(n19198), .ZN(
        n12347) );
  OAI22_X1 U15427 ( .A1(n12199), .A2(n12345), .B1(n12356), .B2(n12344), .ZN(
        n12346) );
  NOR2_X1 U15428 ( .A1(n12347), .A2(n12346), .ZN(n12350) );
  AOI22_X1 U15429 ( .A1(n12370), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10314), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15430 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12348) );
  NAND4_X1 U15431 ( .A1(n12350), .A2(n12349), .A3(n12348), .A4(n12373), .ZN(
        n12365) );
  OAI22_X1 U15432 ( .A1(n12354), .A2(n12353), .B1(n12352), .B2(n12351), .ZN(
        n12360) );
  INV_X1 U15433 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12357) );
  OAI22_X1 U15434 ( .A1(n12358), .A2(n12357), .B1(n12356), .B2(n12355), .ZN(
        n12359) );
  NOR2_X1 U15435 ( .A1(n12360), .A2(n12359), .ZN(n12363) );
  AOI22_X1 U15436 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15437 ( .A1(n10317), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12361) );
  NAND4_X1 U15438 ( .A1(n12363), .A2(n12384), .A3(n12362), .A4(n12361), .ZN(
        n12364) );
  NAND2_X1 U15439 ( .A1(n12365), .A2(n12364), .ZN(n12367) );
  OR3_X1 U15440 ( .A1(n14440), .A2(n19852), .A3(n14442), .ZN(n12366) );
  NOR2_X1 U15441 ( .A1(n12366), .A2(n12367), .ZN(n12368) );
  AOI21_X1 U15442 ( .B1(n12367), .B2(n12366), .A(n12368), .ZN(n14432) );
  NAND2_X1 U15443 ( .A1(n14433), .A2(n14432), .ZN(n14434) );
  INV_X1 U15444 ( .A(n12368), .ZN(n12369) );
  NAND2_X1 U15445 ( .A1(n14434), .A2(n12369), .ZN(n12392) );
  AOI22_X1 U15446 ( .A1(n12370), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10314), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15447 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12371) );
  NAND2_X1 U15448 ( .A1(n12372), .A2(n12371), .ZN(n12390) );
  AOI22_X1 U15449 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15450 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12374) );
  NAND3_X1 U15451 ( .A1(n12375), .A2(n12374), .A3(n12373), .ZN(n12389) );
  AOI22_X1 U15452 ( .A1(n12377), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12376), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15453 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12378), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12379) );
  NAND2_X1 U15454 ( .A1(n12380), .A2(n12379), .ZN(n12388) );
  AOI22_X1 U15455 ( .A1(n12382), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12381), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15456 ( .A1(n10314), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9599), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12385) );
  NAND3_X1 U15457 ( .A1(n12386), .A2(n12385), .A3(n12384), .ZN(n12387) );
  OAI22_X1 U15458 ( .A1(n12390), .A2(n12389), .B1(n12388), .B2(n12387), .ZN(
        n12391) );
  NAND2_X1 U15459 ( .A1(n13356), .A2(n12393), .ZN(n13294) );
  INV_X1 U15460 ( .A(n13299), .ZN(n13335) );
  INV_X1 U15461 ( .A(n13334), .ZN(n13337) );
  NAND2_X1 U15462 ( .A1(n13335), .A2(n13337), .ZN(n13319) );
  NAND2_X1 U15463 ( .A1(n13294), .A2(n13319), .ZN(n12394) );
  NAND2_X1 U15464 ( .A1(n14504), .A2(n19081), .ZN(n12398) );
  INV_X2 U15465 ( .A(n19070), .ZN(n19084) );
  NAND2_X1 U15466 ( .A1(n19084), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12395) );
  NAND2_X1 U15467 ( .A1(n12398), .A2(n12397), .ZN(P2_U2857) );
  INV_X4 U15468 ( .A(n17053), .ZN(n17102) );
  INV_X2 U15469 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18722) );
  NAND2_X1 U15470 ( .A1(n18722), .A2(n18734), .ZN(n12399) );
  NOR2_X2 U15471 ( .A1(n12399), .A2(n16775), .ZN(n12442) );
  INV_X1 U15472 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16968) );
  AOI22_X1 U15473 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12400) );
  OAI21_X1 U15474 ( .B1(n17087), .B2(n16968), .A(n12400), .ZN(n12415) );
  INV_X1 U15475 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14637) );
  NOR2_X4 U15476 ( .A1(n18722), .A2(n12401), .ZN(n17097) );
  AOI22_X1 U15477 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12413) );
  INV_X1 U15478 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15435) );
  NAND2_X2 U15479 ( .A1(n18722), .A2(n12402), .ZN(n12454) );
  AOI22_X1 U15480 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12403) );
  OAI21_X1 U15481 ( .B1(n17005), .B2(n15435), .A(n12403), .ZN(n12411) );
  INV_X1 U15482 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17119) );
  INV_X2 U15483 ( .A(n12494), .ZN(n12420) );
  AOI22_X1 U15484 ( .A1(n17096), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12409) );
  INV_X4 U15485 ( .A(n12430), .ZN(n17078) );
  OR3_X2 U15486 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18568), .ZN(n16801) );
  AOI22_X1 U15487 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12408) );
  OAI211_X1 U15488 ( .C1(n17119), .C2(n17038), .A(n12409), .B(n12408), .ZN(
        n12410) );
  AOI211_X1 U15489 ( .C1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .C2(n16949), .A(
        n12411), .B(n12410), .ZN(n12412) );
  OAI211_X1 U15490 ( .C1(n14637), .C2(n17077), .A(n12413), .B(n12412), .ZN(
        n12414) );
  AOI211_X4 U15491 ( .C1(n17102), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n12415), .B(n12414), .ZN(n17276) );
  AOI22_X1 U15492 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16972), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12416) );
  INV_X1 U15493 ( .A(n12416), .ZN(n12429) );
  AOI22_X1 U15494 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U15495 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12426) );
  BUF_X4 U15496 ( .A(n12418), .Z(n17060) );
  INV_X1 U15497 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U15498 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12419) );
  OAI21_X1 U15499 ( .B1(n17005), .B2(n17003), .A(n12419), .ZN(n12424) );
  INV_X4 U15500 ( .A(n17087), .ZN(n17115) );
  AOI22_X1 U15501 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15502 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16906), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12421) );
  OAI211_X1 U15503 ( .C1(n17038), .C2(n17128), .A(n12422), .B(n12421), .ZN(
        n12423) );
  AOI211_X1 U15504 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n12424), .B(n12423), .ZN(n12425) );
  NAND3_X1 U15505 ( .A1(n12427), .A2(n12426), .A3(n12425), .ZN(n12428) );
  INV_X1 U15506 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U15507 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17101), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12431) );
  OAI21_X1 U15508 ( .B1(n17087), .B2(n17037), .A(n12431), .ZN(n12440) );
  INV_X1 U15509 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15459) );
  AOI22_X1 U15510 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16906), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12438) );
  INV_X1 U15511 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17035) );
  INV_X1 U15512 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17134) );
  OAI22_X1 U15513 ( .A1(n17100), .A2(n17035), .B1(n17038), .B2(n17134), .ZN(
        n12436) );
  AOI22_X1 U15514 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15515 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15516 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12432) );
  NAND3_X1 U15517 ( .A1(n12434), .A2(n12433), .A3(n12432), .ZN(n12435) );
  AOI211_X1 U15518 ( .C1(n17097), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n12436), .B(n12435), .ZN(n12437) );
  OAI211_X1 U15519 ( .C1(n12445), .C2(n15459), .A(n12438), .B(n12437), .ZN(
        n12439) );
  INV_X1 U15520 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U15521 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12486), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U15522 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12442), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15523 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12443) );
  OAI211_X1 U15524 ( .C1(n17106), .C2(n17076), .A(n12444), .B(n12443), .ZN(
        n12451) );
  AOI22_X1 U15525 ( .A1(n12405), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12417), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U15526 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9597), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U15527 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16906), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12447) );
  NAND2_X1 U15528 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12446) );
  NAND4_X1 U15529 ( .A1(n12449), .A2(n12448), .A3(n12447), .A4(n12446), .ZN(
        n12450) );
  AOI211_X1 U15530 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n12451), .B(n12450), .ZN(n12452) );
  INV_X1 U15531 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14558) );
  AOI22_X1 U15532 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12464) );
  INV_X1 U15533 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U15534 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U15535 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16906), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12455) );
  OAI211_X1 U15536 ( .C1(n17106), .C2(n17054), .A(n12456), .B(n12455), .ZN(
        n12462) );
  AOI22_X1 U15537 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15538 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n17102), .B1(
        n12405), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U15539 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12486), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12458) );
  NAND2_X1 U15540 ( .A1(n9600), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12457) );
  NAND4_X1 U15541 ( .A1(n12460), .A2(n12459), .A3(n12458), .A4(n12457), .ZN(
        n12461) );
  AOI211_X1 U15542 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n12462), .B(n12461), .ZN(n12463) );
  OAI211_X1 U15543 ( .C1(n14558), .C2(n12454), .A(n12464), .B(n12463), .ZN(
        n12653) );
  NAND2_X1 U15544 ( .A1(n12667), .A2(n12653), .ZN(n12504) );
  INV_X1 U15545 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17018) );
  AOI22_X1 U15546 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17070), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12474) );
  INV_X1 U15547 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U15548 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U15549 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12465) );
  OAI211_X1 U15550 ( .C1(n17038), .C2(n17131), .A(n12466), .B(n12465), .ZN(
        n12472) );
  AOI22_X1 U15551 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16972), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U15552 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16906), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U15553 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12468) );
  NAND2_X1 U15554 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12467) );
  NAND4_X1 U15555 ( .A1(n12470), .A2(n12469), .A3(n12468), .A4(n12467), .ZN(
        n12471) );
  AOI211_X1 U15556 ( .C1(n12486), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n12472), .B(n12471), .ZN(n12473) );
  OAI211_X1 U15557 ( .C1(n17077), .C2(n17018), .A(n12474), .B(n12473), .ZN(
        n12654) );
  NAND2_X1 U15558 ( .A1(n12507), .A2(n12654), .ZN(n12512) );
  INV_X1 U15559 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17124) );
  AOI22_X1 U15560 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12484) );
  INV_X1 U15561 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16992) );
  AOI22_X1 U15562 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16972), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15563 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n17075), .B1(
        n16906), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12475) );
  OAI211_X1 U15564 ( .C1(n17106), .C2(n16992), .A(n12476), .B(n12475), .ZN(
        n12482) );
  AOI22_X1 U15565 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U15566 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U15567 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12478) );
  NAND2_X1 U15568 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12477) );
  NAND4_X1 U15569 ( .A1(n12480), .A2(n12479), .A3(n12478), .A4(n12477), .ZN(
        n12481) );
  AOI211_X1 U15570 ( .C1(n12486), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n12482), .B(n12481), .ZN(n12483) );
  NOR2_X4 U15571 ( .A1(n17276), .A2(n16276), .ZN(n17662) );
  NAND2_X1 U15572 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17662), .ZN(
        n12485) );
  INV_X1 U15573 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16255) );
  OAI22_X1 U15574 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17662), .B1(
        n12485), .B2(n16255), .ZN(n12537) );
  NAND2_X1 U15575 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17780) );
  INV_X1 U15576 ( .A(n12487), .ZN(n12492) );
  AOI22_X1 U15577 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12405), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U15578 ( .A1(n12418), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12488) );
  NAND3_X1 U15579 ( .A1(n12490), .A2(n12489), .A3(n12488), .ZN(n12491) );
  AOI211_X1 U15580 ( .C1(n17097), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n12492), .B(n12491), .ZN(n12493) );
  INV_X1 U15581 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15423) );
  AOI22_X1 U15582 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12495) );
  OAI21_X1 U15583 ( .B1(n12420), .B2(n15423), .A(n12495), .ZN(n12499) );
  AOI22_X1 U15584 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12497) );
  INV_X1 U15585 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17099) );
  NAND3_X1 U15586 ( .A1(n12497), .A2(n10154), .A3(n12496), .ZN(n12498) );
  INV_X1 U15587 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18725) );
  INV_X1 U15588 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18728) );
  NAND2_X1 U15589 ( .A1(n12501), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12500) );
  INV_X1 U15590 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18088) );
  INV_X1 U15591 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18065) );
  XOR2_X1 U15592 ( .A(n12504), .B(n17292), .Z(n17740) );
  NAND2_X1 U15593 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12505), .ZN(
        n12506) );
  INV_X1 U15594 ( .A(n12654), .ZN(n17288) );
  XNOR2_X1 U15595 ( .A(n12507), .B(n17288), .ZN(n12510) );
  NAND2_X1 U15596 ( .A1(n12510), .A2(n12509), .ZN(n12511) );
  INV_X1 U15597 ( .A(n12655), .ZN(n17282) );
  XNOR2_X1 U15598 ( .A(n12512), .B(n17282), .ZN(n17713) );
  INV_X1 U15599 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17715) );
  XNOR2_X1 U15600 ( .A(n12513), .B(n17279), .ZN(n12514) );
  XOR2_X1 U15601 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12514), .Z(
        n17698) );
  NAND2_X1 U15602 ( .A1(n12517), .A2(n12516), .ZN(n12518) );
  NAND2_X1 U15603 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17982) );
  INV_X1 U15604 ( .A(n17982), .ZN(n17952) );
  NAND2_X1 U15605 ( .A1(n17952), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17968) );
  INV_X1 U15606 ( .A(n17968), .ZN(n12519) );
  INV_X1 U15607 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17974) );
  INV_X1 U15608 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17910) );
  NOR4_X1 U15609 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12525) );
  INV_X1 U15610 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17572) );
  NAND2_X1 U15611 ( .A1(n12526), .A2(n9700), .ZN(n12527) );
  INV_X1 U15612 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17902) );
  NOR2_X1 U15613 ( .A1(n17572), .A2(n17902), .ZN(n17898) );
  NAND2_X1 U15614 ( .A1(n17898), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17862) );
  INV_X1 U15615 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17523) );
  INV_X1 U15616 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17525) );
  NOR2_X1 U15617 ( .A1(n17523), .A2(n17525), .ZN(n17860) );
  NAND2_X1 U15618 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17860), .ZN(
        n17849) );
  NOR2_X1 U15619 ( .A1(n17862), .A2(n17849), .ZN(n17851) );
  NAND2_X1 U15620 ( .A1(n17851), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15495) );
  INV_X1 U15621 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17489) );
  NOR2_X1 U15622 ( .A1(n15495), .A2(n17489), .ZN(n17801) );
  NAND2_X1 U15623 ( .A1(n12533), .A2(n17801), .ZN(n12531) );
  NOR2_X1 U15624 ( .A1(n17662), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17545) );
  NAND2_X1 U15625 ( .A1(n17545), .A2(n17523), .ZN(n12529) );
  NOR2_X1 U15626 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12529), .ZN(
        n17504) );
  INV_X1 U15627 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12530) );
  NAND2_X1 U15628 ( .A1(n17504), .A2(n12530), .ZN(n17492) );
  NAND2_X2 U15629 ( .A1(n17522), .A2(n12532), .ZN(n17474) );
  INV_X1 U15630 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17897) );
  INV_X1 U15631 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17500) );
  NOR3_X1 U15632 ( .A1(n17897), .A2(n17849), .A3(n17500), .ZN(n17803) );
  NAND2_X1 U15633 ( .A1(n17898), .A2(n12533), .ZN(n17502) );
  INV_X1 U15634 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17810) );
  INV_X1 U15635 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17792) );
  OAI21_X1 U15636 ( .B1(n16255), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n15572), .ZN(n12535) );
  INV_X1 U15637 ( .A(n12535), .ZN(n12536) );
  NAND2_X1 U15638 ( .A1(n17792), .A2(n16269), .ZN(n17436) );
  INV_X1 U15639 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16242) );
  NAND2_X1 U15640 ( .A1(n15511), .A2(n16242), .ZN(n15571) );
  NAND2_X1 U15641 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16255), .ZN(
        n16259) );
  INV_X1 U15642 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16935) );
  AOI22_X1 U15643 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12538) );
  OAI21_X1 U15644 ( .B1(n12445), .B2(n16935), .A(n12538), .ZN(n12547) );
  AOI22_X1 U15645 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12545) );
  INV_X1 U15646 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15445) );
  OAI22_X1 U15647 ( .A1(n17005), .A2(n15445), .B1(n17038), .B2(n17076), .ZN(
        n12543) );
  AOI22_X1 U15648 ( .A1(n17096), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12405), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12541) );
  AOI22_X1 U15649 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17115), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12540) );
  AOI22_X1 U15650 ( .A1(n12418), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12539) );
  NAND3_X1 U15651 ( .A1(n12541), .A2(n12540), .A3(n12539), .ZN(n12542) );
  AOI211_X1 U15652 ( .C1(n17097), .C2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n12543), .B(n12542), .ZN(n12544) );
  OAI211_X1 U15653 ( .C1(n12430), .C2(n17072), .A(n12545), .B(n12544), .ZN(
        n12546) );
  AOI211_X4 U15654 ( .C1(n17102), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n12547), .B(n12546), .ZN(n17348) );
  NAND3_X1 U15655 ( .A1(n18726), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18617) );
  OAI22_X1 U15656 ( .A1(n18741), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18591), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12548) );
  INV_X1 U15657 ( .A(n12548), .ZN(n12627) );
  NAND2_X1 U15658 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18589), .ZN(
        n12555) );
  INV_X1 U15659 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18607) );
  NOR2_X1 U15660 ( .A1(n12548), .A2(n12555), .ZN(n12549) );
  AOI21_X1 U15661 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18591), .A(
        n12549), .ZN(n12556) );
  AOI22_X1 U15662 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18596), .B2(n18734), .ZN(
        n12557) );
  OAI22_X1 U15663 ( .A1(n18600), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(
        n12551), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12560) );
  NAND2_X1 U15664 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12551), .ZN(
        n12558) );
  OAI22_X1 U15665 ( .A1(n18607), .A2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n12560), .B2(n12552), .ZN(n12561) );
  INV_X1 U15666 ( .A(n12561), .ZN(n12553) );
  OAI21_X1 U15667 ( .B1(n12627), .B2(n12555), .A(n12553), .ZN(n12554) );
  AOI21_X1 U15668 ( .B1(n12627), .B2(n12555), .A(n12554), .ZN(n13648) );
  OAI21_X1 U15669 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18589), .A(
        n12555), .ZN(n12629) );
  XOR2_X1 U15670 ( .A(n12557), .B(n12556), .Z(n12562) );
  NOR2_X1 U15671 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18600), .ZN(
        n12559) );
  AOI22_X1 U15672 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12560), .B1(
        n12559), .B2(n12558), .ZN(n12626) );
  AOI21_X1 U15673 ( .B1(n13648), .B2(n12629), .A(n13649), .ZN(n18547) );
  AOI22_X1 U15674 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12563) );
  OAI21_X1 U15675 ( .B1(n16986), .B2(n10165), .A(n12563), .ZN(n12569) );
  INV_X1 U15676 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16862) );
  AOI22_X1 U15677 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12568) );
  INV_X1 U15678 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16800) );
  OAI22_X1 U15679 ( .A1(n17100), .A2(n16985), .B1(n17005), .B2(n16800), .ZN(
        n12567) );
  AOI22_X1 U15680 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U15681 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17096), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U15682 ( .A1(n16949), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12564) );
  INV_X1 U15683 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17052) );
  INV_X1 U15684 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16919) );
  OAI22_X1 U15685 ( .A1(n12420), .A2(n17052), .B1(n17073), .B2(n16919), .ZN(
        n12576) );
  AOI22_X1 U15686 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U15687 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12570) );
  OAI21_X1 U15688 ( .B1(n16918), .B2(n16801), .A(n12570), .ZN(n12574) );
  AOI22_X1 U15689 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n17075), .B1(
        n16972), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12573) );
  AOI22_X1 U15690 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12572) );
  AOI22_X1 U15691 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12571) );
  NAND2_X1 U15692 ( .A1(n12644), .A2(n18128), .ZN(n15502) );
  NOR2_X1 U15693 ( .A1(n17151), .A2(n15502), .ZN(n15501) );
  INV_X1 U15694 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U15695 ( .A1(n12405), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12586) );
  INV_X1 U15696 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17019) );
  AOI22_X1 U15697 ( .A1(n17096), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U15698 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16972), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12577) );
  OAI211_X1 U15699 ( .C1(n17038), .C2(n17019), .A(n12578), .B(n12577), .ZN(
        n12584) );
  AOI22_X1 U15700 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U15701 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15702 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12486), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12580) );
  NAND2_X1 U15703 ( .A1(n16949), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12579) );
  NAND4_X1 U15704 ( .A1(n12582), .A2(n12581), .A3(n12580), .A4(n12579), .ZN(
        n12583) );
  AOI22_X1 U15705 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12596) );
  INV_X1 U15706 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U15707 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17096), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12588) );
  AOI22_X1 U15708 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12587) );
  OAI211_X1 U15709 ( .C1(n17038), .C2(n17013), .A(n12588), .B(n12587), .ZN(
        n12594) );
  AOI22_X1 U15710 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16972), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U15711 ( .A1(n16812), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15712 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12590) );
  NAND2_X1 U15713 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12589) );
  NAND4_X1 U15714 ( .A1(n12592), .A2(n12591), .A3(n12590), .A4(n12589), .ZN(
        n12593) );
  NOR2_X1 U15715 ( .A1(n17151), .A2(n18148), .ZN(n15399) );
  INV_X1 U15716 ( .A(n12644), .ZN(n18132) );
  INV_X1 U15717 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16969) );
  AOI22_X1 U15718 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U15719 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n12405), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15720 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17115), .B1(
        n17096), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12597) );
  OAI211_X1 U15721 ( .C1(n14637), .C2(n17106), .A(n12598), .B(n12597), .ZN(
        n12603) );
  AOI22_X1 U15722 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n16972), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U15723 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17078), .ZN(n12601) );
  AOI22_X1 U15724 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n9600), .ZN(n12600) );
  NAND2_X1 U15725 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12599) );
  INV_X1 U15726 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15456) );
  AOI22_X1 U15727 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12614) );
  INV_X1 U15728 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17046) );
  AOI22_X1 U15729 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16906), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U15730 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12605) );
  OAI211_X1 U15731 ( .C1(n17038), .C2(n17046), .A(n12606), .B(n12605), .ZN(
        n12612) );
  AOI22_X1 U15732 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12610) );
  AOI22_X1 U15733 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U15734 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12608) );
  NAND2_X1 U15735 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12607) );
  NAND4_X1 U15736 ( .A1(n12610), .A2(n12609), .A3(n12608), .A4(n12607), .ZN(
        n12611) );
  AOI22_X1 U15737 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12615) );
  OAI21_X1 U15738 ( .B1(n17087), .B2(n17105), .A(n12615), .ZN(n12624) );
  AOI22_X1 U15739 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12622) );
  INV_X1 U15740 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17094) );
  AOI22_X1 U15741 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12616) );
  OAI21_X1 U15742 ( .B1(n17077), .B2(n17094), .A(n12616), .ZN(n12620) );
  INV_X1 U15743 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14657) );
  AOI22_X1 U15744 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15745 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17096), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12617) );
  OAI211_X1 U15746 ( .C1(n14657), .C2(n17005), .A(n12618), .B(n12617), .ZN(
        n12619) );
  AOI211_X1 U15747 ( .C1(n9600), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n12620), .B(n12619), .ZN(n12621) );
  OAI211_X1 U15748 ( .C1(n10165), .C2(n17112), .A(n12622), .B(n12621), .ZN(
        n12623) );
  NAND2_X1 U15749 ( .A1(n12641), .A2(n12645), .ZN(n12625) );
  AOI211_X1 U15750 ( .C1(n18143), .C2(n15604), .A(n15399), .B(n12625), .ZN(
        n13652) );
  NAND2_X1 U15751 ( .A1(n12627), .A2(n12626), .ZN(n12628) );
  NAND2_X1 U15752 ( .A1(n17348), .A2(n18125), .ZN(n12631) );
  NAND2_X1 U15753 ( .A1(n12645), .A2(n12631), .ZN(n18781) );
  NAND3_X1 U15754 ( .A1(n12641), .A2(n18584), .A3(n18143), .ZN(n13658) );
  NAND2_X1 U15755 ( .A1(n18158), .A2(n18763), .ZN(n12638) );
  INV_X1 U15756 ( .A(n12638), .ZN(n12630) );
  NAND4_X1 U15757 ( .A1(n12640), .A2(n15500), .A3(n12630), .A4(n12635), .ZN(
        n12643) );
  NAND2_X1 U15758 ( .A1(n12644), .A2(n18148), .ZN(n15504) );
  OR2_X1 U15759 ( .A1(n15504), .A2(n17151), .ZN(n15499) );
  AOI21_X1 U15760 ( .B1(n12642), .B2(n15499), .A(n18125), .ZN(n12637) );
  AOI211_X1 U15761 ( .C1(n15500), .C2(n18148), .A(n12632), .B(n18132), .ZN(
        n12634) );
  OAI21_X1 U15762 ( .B1(n12635), .B2(n17199), .A(n18143), .ZN(n12633) );
  OAI21_X1 U15763 ( .B1(n12635), .B2(n12634), .A(n12633), .ZN(n12636) );
  AOI211_X2 U15764 ( .C1(n12640), .C2(n12638), .A(n12637), .B(n12636), .ZN(
        n13651) );
  NAND2_X1 U15765 ( .A1(n12644), .A2(n12640), .ZN(n15396) );
  NOR2_X1 U15766 ( .A1(n12644), .A2(n12643), .ZN(n13650) );
  NAND2_X1 U15767 ( .A1(n16264), .A2(n17664), .ZN(n12691) );
  NAND2_X1 U15768 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18112) );
  NAND2_X1 U15769 ( .A1(n18743), .A2(n18112), .ZN(n18770) );
  NAND2_X1 U15770 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17728) );
  INV_X1 U15771 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16428) );
  INV_X1 U15772 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17763) );
  NAND2_X1 U15773 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16736) );
  NAND2_X1 U15774 ( .A1(n17729), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17719) );
  NAND2_X1 U15775 ( .A1(n17699), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17671) );
  NAND3_X1 U15776 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16647) );
  NOR2_X1 U15777 ( .A1(n16647), .A2(n17638), .ZN(n16607) );
  NAND2_X1 U15778 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17613) );
  NAND2_X1 U15779 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17566) );
  NAND2_X1 U15780 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17551), .ZN(
        n17531) );
  NAND2_X1 U15781 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17532) );
  NAND2_X1 U15782 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17498) );
  NAND2_X1 U15783 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17459) );
  NAND2_X1 U15784 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17421) );
  NAND2_X1 U15785 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16249), .ZN(
        n12649) );
  INV_X1 U15786 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18702) );
  NAND2_X1 U15787 ( .A1(n18726), .A2(n18743), .ZN(n18729) );
  OR3_X2 U15788 ( .A1(n18729), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n17988) );
  NOR2_X1 U15789 ( .A1(n18702), .A2(n17988), .ZN(n16262) );
  INV_X1 U15790 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18767) );
  NAND2_X1 U15791 ( .A1(n18767), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17771) );
  NOR2_X1 U15792 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18626) );
  INV_X1 U15793 ( .A(n18626), .ZN(n18766) );
  AOI21_X1 U15794 ( .B1(n18112), .B2(n18766), .A(n18745), .ZN(n18124) );
  INV_X1 U15795 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18779) );
  NAND3_X1 U15796 ( .A1(n18779), .A2(n18743), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18408) );
  OR2_X2 U15797 ( .A1(n18385), .A2(n18408), .ZN(n18456) );
  OR2_X1 U15798 ( .A1(n12649), .A2(n17612), .ZN(n16227) );
  XNOR2_X1 U15799 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12651) );
  NOR2_X1 U15800 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17516), .ZN(
        n16247) );
  INV_X1 U15801 ( .A(n17771), .ZN(n17602) );
  NOR2_X1 U15802 ( .A1(n17763), .A2(n17420), .ZN(n16411) );
  NAND3_X1 U15803 ( .A1(n16411), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16408) );
  AOI22_X1 U15804 ( .A1(n17602), .A2(n16408), .B1(n18493), .B2(n12649), .ZN(
        n12650) );
  NAND2_X1 U15805 ( .A1(n12650), .A2(n17770), .ZN(n16248) );
  NOR2_X1 U15806 ( .A1(n16247), .A2(n16248), .ZN(n16226) );
  OAI22_X1 U15807 ( .A1(n16227), .A2(n12651), .B1(n16226), .B2(n16428), .ZN(
        n12652) );
  AOI211_X1 U15808 ( .C1(n17605), .C2(n16749), .A(n16262), .B(n12652), .ZN(
        n12690) );
  INV_X1 U15809 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18727) );
  NAND2_X1 U15810 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16238) );
  NOR2_X1 U15811 ( .A1(n16238), .A2(n16242), .ZN(n12687) );
  INV_X1 U15812 ( .A(n12687), .ZN(n16254) );
  INV_X1 U15813 ( .A(n15495), .ZN(n17833) );
  INV_X1 U15814 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17825) );
  NOR2_X1 U15815 ( .A1(n17489), .A2(n17825), .ZN(n17779) );
  INV_X1 U15816 ( .A(n17779), .ZN(n17805) );
  NOR2_X1 U15817 ( .A1(n17805), .A2(n17780), .ZN(n16268) );
  NAND2_X1 U15818 ( .A1(n17833), .A2(n16268), .ZN(n16229) );
  NOR2_X1 U15819 ( .A1(n17968), .A2(n17974), .ZN(n17606) );
  NOR2_X1 U15820 ( .A1(n12501), .A2(n17769), .ZN(n12664) );
  NOR2_X1 U15821 ( .A1(n12664), .A2(n12653), .ZN(n12662) );
  NOR2_X1 U15822 ( .A1(n17292), .A2(n12662), .ZN(n12661) );
  NAND2_X1 U15823 ( .A1(n12661), .A2(n12654), .ZN(n12659) );
  NOR2_X1 U15824 ( .A1(n12655), .A2(n12659), .ZN(n12658) );
  NAND2_X1 U15825 ( .A1(n12658), .A2(n12656), .ZN(n12657) );
  NOR2_X1 U15826 ( .A1(n17276), .A2(n12657), .ZN(n12683) );
  XOR2_X1 U15827 ( .A(n17276), .B(n12657), .Z(n17690) );
  XNOR2_X1 U15828 ( .A(n17279), .B(n12658), .ZN(n12676) );
  XNOR2_X1 U15829 ( .A(n17282), .B(n12659), .ZN(n12660) );
  NAND2_X1 U15830 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12660), .ZN(
        n12675) );
  XOR2_X1 U15831 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12660), .Z(
        n17711) );
  XNOR2_X1 U15832 ( .A(n17288), .B(n12661), .ZN(n12673) );
  XOR2_X1 U15833 ( .A(n12662), .B(n17292), .Z(n12663) );
  NAND2_X1 U15834 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12663), .ZN(
        n12671) );
  XOR2_X1 U15835 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n12663), .Z(
        n17737) );
  XNOR2_X1 U15836 ( .A(n17297), .B(n12664), .ZN(n12669) );
  OR2_X1 U15837 ( .A1(n18088), .A2(n12669), .ZN(n12670) );
  INV_X1 U15838 ( .A(n17769), .ZN(n12668) );
  AOI21_X1 U15839 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12667), .A(
        n12668), .ZN(n12666) );
  NOR2_X1 U15840 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12667), .ZN(
        n12665) );
  AOI221_X1 U15841 ( .B1(n12668), .B2(n12667), .C1(n12666), .C2(n18725), .A(
        n12665), .ZN(n17748) );
  XOR2_X1 U15842 ( .A(n18088), .B(n12669), .Z(n17747) );
  NAND2_X1 U15843 ( .A1(n17748), .A2(n17747), .ZN(n17746) );
  NAND2_X1 U15844 ( .A1(n12670), .A2(n17746), .ZN(n17736) );
  NAND2_X1 U15845 ( .A1(n17737), .A2(n17736), .ZN(n17735) );
  NAND2_X1 U15846 ( .A1(n12671), .A2(n17735), .ZN(n12672) );
  NAND2_X1 U15847 ( .A1(n12673), .A2(n12672), .ZN(n12674) );
  XOR2_X1 U15848 ( .A(n12673), .B(n12672), .Z(n17726) );
  NAND2_X1 U15849 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17726), .ZN(
        n17725) );
  NAND2_X1 U15850 ( .A1(n12674), .A2(n17725), .ZN(n17710) );
  NAND2_X1 U15851 ( .A1(n17711), .A2(n17710), .ZN(n17709) );
  NAND2_X1 U15852 ( .A1(n12675), .A2(n17709), .ZN(n12677) );
  NAND2_X1 U15853 ( .A1(n12676), .A2(n12677), .ZN(n12678) );
  XOR2_X1 U15854 ( .A(n12677), .B(n12676), .Z(n17701) );
  NAND2_X1 U15855 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17701), .ZN(
        n17700) );
  INV_X1 U15856 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17691) );
  NOR2_X2 U15857 ( .A1(n17688), .A2(n17691), .ZN(n12679) );
  NAND2_X1 U15858 ( .A1(n12683), .A2(n12679), .ZN(n12684) );
  INV_X1 U15859 ( .A(n12679), .ZN(n12682) );
  NAND2_X1 U15860 ( .A1(n17690), .A2(n17689), .ZN(n12681) );
  NAND2_X1 U15861 ( .A1(n12683), .A2(n12682), .ZN(n12680) );
  OAI211_X1 U15862 ( .C1(n12683), .C2(n12682), .A(n12681), .B(n12680), .ZN(
        n17677) );
  NAND2_X1 U15863 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17677), .ZN(
        n17676) );
  NAND2_X1 U15864 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17895) );
  INV_X1 U15865 ( .A(n17895), .ZN(n12686) );
  NAND2_X1 U15866 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12686), .ZN(
        n15496) );
  NOR2_X4 U15867 ( .A1(n17955), .A2(n15496), .ZN(n17845) );
  NOR2_X2 U15868 ( .A1(n16229), .A2(n17920), .ZN(n17782) );
  NAND2_X1 U15869 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16236), .ZN(
        n12685) );
  XOR2_X1 U15870 ( .A(n18727), .B(n12685), .Z(n16265) );
  NAND2_X1 U15871 ( .A1(n16265), .A2(n17762), .ZN(n12689) );
  INV_X1 U15872 ( .A(n17606), .ZN(n17936) );
  INV_X1 U15873 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17960) );
  NOR2_X1 U15874 ( .A1(n17936), .A2(n17960), .ZN(n17894) );
  INV_X1 U15875 ( .A(n17894), .ZN(n17595) );
  INV_X1 U15876 ( .A(n16229), .ZN(n16257) );
  NAND2_X1 U15877 ( .A1(n17847), .A2(n16257), .ZN(n16239) );
  INV_X1 U15878 ( .A(n16239), .ZN(n17783) );
  NAND3_X1 U15879 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n12687), .A3(
        n17783), .ZN(n12688) );
  XNOR2_X1 U15880 ( .A(n18727), .B(n12688), .ZN(n16267) );
  NAND2_X1 U15881 ( .A1(n12691), .A2(n9667), .ZN(P3_U2799) );
  NOR2_X1 U15882 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12693) );
  NOR4_X1 U15883 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12692) );
  NAND4_X1 U15884 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12693), .A4(n12692), .ZN(n12717) );
  NOR2_X1 U15885 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12717), .ZN(n16362)
         );
  NOR4_X1 U15886 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n12697) );
  NOR4_X1 U15887 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12696) );
  NOR4_X1 U15888 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12695) );
  NOR4_X1 U15889 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12694) );
  AND4_X1 U15890 ( .A1(n12697), .A2(n12696), .A3(n12695), .A4(n12694), .ZN(
        n12703) );
  NOR4_X1 U15891 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_8__SCAN_IN), .A3(P1_ADDRESS_REG_1__SCAN_IN), .A4(
        P1_ADDRESS_REG_0__SCAN_IN), .ZN(n12701) );
  NOR4_X1 U15892 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12700) );
  NOR4_X1 U15893 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12699) );
  INV_X1 U15894 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n12698) );
  AND4_X1 U15895 ( .A1(n12701), .A2(n12700), .A3(n12699), .A4(n12698), .ZN(
        n12702) );
  NAND2_X1 U15896 ( .A1(n12703), .A2(n12702), .ZN(n12704) );
  AND2_X2 U15897 ( .A1(n12704), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14158)
         );
  INV_X1 U15898 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n20859) );
  NOR3_X1 U15899 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20859), .ZN(n12706) );
  NOR4_X1 U15900 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12705) );
  NAND4_X1 U15901 ( .A1(n14158), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n12706), .A4(
        n12705), .ZN(U214) );
  NOR4_X1 U15902 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12710) );
  NOR4_X1 U15903 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n12709) );
  NOR4_X1 U15904 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12708) );
  NOR4_X1 U15905 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12707) );
  AND4_X1 U15906 ( .A1(n12710), .A2(n12709), .A3(n12708), .A4(n12707), .ZN(
        n12715) );
  NOR4_X1 U15907 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_11__SCAN_IN), .A4(
        P2_ADDRESS_REG_22__SCAN_IN), .ZN(n12713) );
  NOR4_X1 U15908 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_23__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n12712) );
  NOR4_X1 U15909 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_28__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n12711) );
  INV_X1 U15910 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19730) );
  AND4_X1 U15911 ( .A1(n12713), .A2(n12712), .A3(n12711), .A4(n19730), .ZN(
        n12714) );
  NAND2_X1 U15912 ( .A1(n12715), .A2(n12714), .ZN(n12716) );
  NAND2_X2 U15913 ( .A1(n12716), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n14505)
         );
  NOR2_X1 U15914 ( .A1(n14505), .A2(n12717), .ZN(n16285) );
  NAND2_X1 U15915 ( .A1(n16285), .A2(U214), .ZN(U212) );
  INV_X1 U15916 ( .A(n19700), .ZN(n19849) );
  NOR2_X1 U15917 ( .A1(n15492), .A2(n19849), .ZN(n12832) );
  NAND2_X1 U15918 ( .A1(n12832), .A2(n13338), .ZN(n19012) );
  INV_X1 U15919 ( .A(n19012), .ZN(n19035) );
  INV_X1 U15920 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19866) );
  OAI211_X1 U15921 ( .C1(n19035), .C2(n19866), .A(n18788), .B(n12718), .ZN(
        P2_U2814) );
  NOR2_X1 U15922 ( .A1(n19846), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n12720)
         );
  INV_X1 U15923 ( .A(n12893), .ZN(n12719) );
  AOI22_X1 U15924 ( .A1(n12720), .A2(n18788), .B1(n12719), .B2(n19846), .ZN(
        P2_U3612) );
  INV_X1 U15925 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12723) );
  INV_X1 U15926 ( .A(n12802), .ZN(n12779) );
  INV_X1 U15927 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13136) );
  NOR2_X1 U15928 ( .A1(n14505), .A2(n13136), .ZN(n12721) );
  AOI21_X1 U15929 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n14505), .A(n12721), .ZN(
        n13241) );
  INV_X1 U15930 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12722) );
  OAI222_X1 U15931 ( .A1(n12723), .A2(n12812), .B1(n12779), .B2(n13241), .C1(
        n12722), .C2(n12833), .ZN(P2_U2982) );
  INV_X1 U15932 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n12728) );
  INV_X1 U15933 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n12724) );
  OR2_X1 U15934 ( .A1(n14505), .A2(n12724), .ZN(n12726) );
  NAND2_X1 U15935 ( .A1(n14505), .A2(BUF2_REG_5__SCAN_IN), .ZN(n12725) );
  AND2_X1 U15936 ( .A1(n12726), .A2(n12725), .ZN(n19181) );
  NOR2_X1 U15937 ( .A1(n12779), .A2(n19181), .ZN(n12764) );
  AOI21_X1 U15938 ( .B1(n12809), .B2(P2_EAX_REG_21__SCAN_IN), .A(n12764), .ZN(
        n12727) );
  OAI21_X1 U15939 ( .B1(n12812), .B2(n12728), .A(n12727), .ZN(P2_U2957) );
  INV_X1 U15940 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12733) );
  INV_X1 U15941 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n12729) );
  OR2_X1 U15942 ( .A1(n14505), .A2(n12729), .ZN(n12731) );
  NAND2_X1 U15943 ( .A1(n14505), .A2(BUF2_REG_0__SCAN_IN), .ZN(n12730) );
  AND2_X1 U15944 ( .A1(n12731), .A2(n12730), .ZN(n19091) );
  NOR2_X1 U15945 ( .A1(n12779), .A2(n19091), .ZN(n12734) );
  AOI21_X1 U15946 ( .B1(n12809), .B2(P2_EAX_REG_0__SCAN_IN), .A(n12734), .ZN(
        n12732) );
  OAI21_X1 U15947 ( .B1(n12812), .B2(n12733), .A(n12732), .ZN(P2_U2967) );
  INV_X1 U15948 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12736) );
  AOI21_X1 U15949 ( .B1(n12809), .B2(P2_EAX_REG_16__SCAN_IN), .A(n12734), .ZN(
        n12735) );
  OAI21_X1 U15950 ( .B1(n12812), .B2(n12736), .A(n12735), .ZN(P2_U2952) );
  INV_X1 U15951 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n12740) );
  INV_X1 U15952 ( .A(n14505), .ZN(n14507) );
  INV_X1 U15953 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n12737) );
  NOR2_X1 U15954 ( .A1(n14507), .A2(n12737), .ZN(n12738) );
  AOI21_X1 U15955 ( .B1(n14507), .B2(BUF1_REG_12__SCAN_IN), .A(n12738), .ZN(
        n14677) );
  NOR2_X1 U15956 ( .A1(n12779), .A2(n14677), .ZN(n12773) );
  AOI21_X1 U15957 ( .B1(n12809), .B2(P2_EAX_REG_12__SCAN_IN), .A(n12773), .ZN(
        n12739) );
  OAI21_X1 U15958 ( .B1(n12812), .B2(n12740), .A(n12739), .ZN(P2_U2979) );
  INV_X1 U15959 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n12745) );
  INV_X1 U15960 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n12741) );
  OR2_X1 U15961 ( .A1(n14505), .A2(n12741), .ZN(n12743) );
  NAND2_X1 U15962 ( .A1(n14505), .A2(BUF2_REG_1__SCAN_IN), .ZN(n12742) );
  AND2_X1 U15963 ( .A1(n12743), .A2(n12742), .ZN(n15340) );
  NOR2_X1 U15964 ( .A1(n12779), .A2(n15340), .ZN(n12805) );
  AOI21_X1 U15965 ( .B1(n12809), .B2(P2_EAX_REG_17__SCAN_IN), .A(n12805), .ZN(
        n12744) );
  OAI21_X1 U15966 ( .B1(n12812), .B2(n12745), .A(n12744), .ZN(P2_U2953) );
  INV_X1 U15967 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n12750) );
  INV_X1 U15968 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n12746) );
  OR2_X1 U15969 ( .A1(n14505), .A2(n12746), .ZN(n12748) );
  NAND2_X1 U15970 ( .A1(n14505), .A2(BUF2_REG_4__SCAN_IN), .ZN(n12747) );
  AND2_X1 U15971 ( .A1(n12748), .A2(n12747), .ZN(n16081) );
  NOR2_X1 U15972 ( .A1(n12779), .A2(n16081), .ZN(n12770) );
  AOI21_X1 U15973 ( .B1(n12809), .B2(P2_EAX_REG_4__SCAN_IN), .A(n12770), .ZN(
        n12749) );
  OAI21_X1 U15974 ( .B1(n12812), .B2(n12750), .A(n12749), .ZN(P2_U2971) );
  INV_X1 U15975 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n12755) );
  INV_X1 U15976 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n12751) );
  OR2_X1 U15977 ( .A1(n14505), .A2(n12751), .ZN(n12753) );
  NAND2_X1 U15978 ( .A1(n14505), .A2(BUF2_REG_7__SCAN_IN), .ZN(n12752) );
  AND2_X1 U15979 ( .A1(n12753), .A2(n12752), .ZN(n15348) );
  NOR2_X1 U15980 ( .A1(n12779), .A2(n15348), .ZN(n12761) );
  AOI21_X1 U15981 ( .B1(n12809), .B2(P2_EAX_REG_23__SCAN_IN), .A(n12761), .ZN(
        n12754) );
  OAI21_X1 U15982 ( .B1(n12812), .B2(n12755), .A(n12754), .ZN(P2_U2959) );
  INV_X1 U15983 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n12760) );
  INV_X1 U15984 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n12756) );
  OR2_X1 U15985 ( .A1(n14505), .A2(n12756), .ZN(n12758) );
  NAND2_X1 U15986 ( .A1(n14505), .A2(BUF2_REG_3__SCAN_IN), .ZN(n12757) );
  AND2_X1 U15987 ( .A1(n12758), .A2(n12757), .ZN(n19173) );
  NOR2_X1 U15988 ( .A1(n12779), .A2(n19173), .ZN(n12767) );
  AOI21_X1 U15989 ( .B1(n12809), .B2(P2_EAX_REG_3__SCAN_IN), .A(n12767), .ZN(
        n12759) );
  OAI21_X1 U15990 ( .B1(n12812), .B2(n12760), .A(n12759), .ZN(P2_U2970) );
  INV_X1 U15991 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n12763) );
  AOI21_X1 U15992 ( .B1(n12809), .B2(P2_EAX_REG_7__SCAN_IN), .A(n12761), .ZN(
        n12762) );
  OAI21_X1 U15993 ( .B1(n12812), .B2(n12763), .A(n12762), .ZN(P2_U2974) );
  INV_X1 U15994 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n12766) );
  AOI21_X1 U15995 ( .B1(n12809), .B2(P2_EAX_REG_5__SCAN_IN), .A(n12764), .ZN(
        n12765) );
  OAI21_X1 U15996 ( .B1(n12812), .B2(n12766), .A(n12765), .ZN(P2_U2972) );
  INV_X1 U15997 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n12769) );
  AOI21_X1 U15998 ( .B1(n12809), .B2(P2_EAX_REG_19__SCAN_IN), .A(n12767), .ZN(
        n12768) );
  OAI21_X1 U15999 ( .B1(n12812), .B2(n12769), .A(n12768), .ZN(P2_U2955) );
  INV_X1 U16000 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n12772) );
  AOI21_X1 U16001 ( .B1(n12809), .B2(P2_EAX_REG_20__SCAN_IN), .A(n12770), .ZN(
        n12771) );
  OAI21_X1 U16002 ( .B1(n12812), .B2(n12772), .A(n12771), .ZN(P2_U2956) );
  INV_X1 U16003 ( .A(P2_UWORD_REG_12__SCAN_IN), .ZN(n12775) );
  AOI21_X1 U16004 ( .B1(n12809), .B2(P2_EAX_REG_28__SCAN_IN), .A(n12773), .ZN(
        n12774) );
  OAI21_X1 U16005 ( .B1(n12812), .B2(n12775), .A(n12774), .ZN(P2_U2964) );
  INV_X1 U16006 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n12781) );
  INV_X1 U16007 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n12776) );
  OR2_X1 U16008 ( .A1(n14505), .A2(n12776), .ZN(n12778) );
  NAND2_X1 U16009 ( .A1(n14505), .A2(BUF2_REG_2__SCAN_IN), .ZN(n12777) );
  AND2_X1 U16010 ( .A1(n12778), .A2(n12777), .ZN(n16089) );
  NOR2_X1 U16011 ( .A1(n12779), .A2(n16089), .ZN(n12808) );
  AOI21_X1 U16012 ( .B1(n12809), .B2(P2_EAX_REG_18__SCAN_IN), .A(n12808), .ZN(
        n12780) );
  OAI21_X1 U16013 ( .B1(n12812), .B2(n12781), .A(n12780), .ZN(P2_U2954) );
  INV_X1 U16014 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n12785) );
  INV_X1 U16015 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13631) );
  OR2_X1 U16016 ( .A1(n14505), .A2(n13631), .ZN(n12783) );
  NAND2_X1 U16017 ( .A1(n14505), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12782) );
  NAND2_X1 U16018 ( .A1(n12783), .A2(n12782), .ZN(n14512) );
  NAND2_X1 U16019 ( .A1(n12802), .A2(n14512), .ZN(n12816) );
  NAND2_X1 U16020 ( .A1(n12809), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n12784) );
  OAI211_X1 U16021 ( .C1(n12812), .C2(n12785), .A(n12816), .B(n12784), .ZN(
        P2_U2981) );
  INV_X1 U16022 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n12790) );
  INV_X1 U16023 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n12786) );
  OR2_X1 U16024 ( .A1(n14505), .A2(n12786), .ZN(n12788) );
  NAND2_X1 U16025 ( .A1(n14505), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12787) );
  NAND2_X1 U16026 ( .A1(n12788), .A2(n12787), .ZN(n13022) );
  NAND2_X1 U16027 ( .A1(n12802), .A2(n13022), .ZN(n12819) );
  NAND2_X1 U16028 ( .A1(n12809), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n12789) );
  OAI211_X1 U16029 ( .C1(n12812), .C2(n12790), .A(n12819), .B(n12789), .ZN(
        P2_U2976) );
  INV_X1 U16030 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n12792) );
  MUX2_X1 U16031 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n14505), .Z(n14697) );
  NAND2_X1 U16032 ( .A1(n12802), .A2(n14697), .ZN(n12821) );
  NAND2_X1 U16033 ( .A1(n12809), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n12791) );
  OAI211_X1 U16034 ( .C1(n12812), .C2(n12792), .A(n12821), .B(n12791), .ZN(
        P2_U2977) );
  INV_X1 U16035 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n12794) );
  MUX2_X1 U16036 ( .A(BUF1_REG_11__SCAN_IN), .B(BUF2_REG_11__SCAN_IN), .S(
        n14505), .Z(n14689) );
  NAND2_X1 U16037 ( .A1(n12802), .A2(n14689), .ZN(n12830) );
  NAND2_X1 U16038 ( .A1(n12809), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n12793) );
  OAI211_X1 U16039 ( .C1(n12812), .C2(n12794), .A(n12830), .B(n12793), .ZN(
        P2_U2978) );
  INV_X1 U16040 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n12796) );
  MUX2_X1 U16041 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n14505), .Z(n14715) );
  NAND2_X1 U16042 ( .A1(n12802), .A2(n14715), .ZN(n12824) );
  NAND2_X1 U16043 ( .A1(n12809), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n12795) );
  OAI211_X1 U16044 ( .C1(n12812), .C2(n12796), .A(n12824), .B(n12795), .ZN(
        P2_U2975) );
  INV_X1 U16045 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n12798) );
  MUX2_X1 U16046 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n14505), .Z(n14523) );
  NAND2_X1 U16047 ( .A1(n12802), .A2(n14523), .ZN(n12827) );
  NAND2_X1 U16048 ( .A1(n12809), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n12797) );
  OAI211_X1 U16049 ( .C1(n12812), .C2(n12798), .A(n12827), .B(n12797), .ZN(
        P2_U2980) );
  INV_X1 U16050 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n12804) );
  INV_X1 U16051 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n12799) );
  OR2_X1 U16052 ( .A1(n14505), .A2(n12799), .ZN(n12801) );
  NAND2_X1 U16053 ( .A1(n14505), .A2(BUF2_REG_6__SCAN_IN), .ZN(n12800) );
  AND2_X1 U16054 ( .A1(n12801), .A2(n12800), .ZN(n19191) );
  INV_X1 U16055 ( .A(n19191), .ZN(n14733) );
  NAND2_X1 U16056 ( .A1(n12802), .A2(n14733), .ZN(n12813) );
  NAND2_X1 U16057 ( .A1(n12809), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n12803) );
  OAI211_X1 U16058 ( .C1(n12812), .C2(n12804), .A(n12813), .B(n12803), .ZN(
        P2_U2973) );
  INV_X1 U16059 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n12807) );
  AOI21_X1 U16060 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n12809), .A(n12805), .ZN(
        n12806) );
  OAI21_X1 U16061 ( .B1(n12812), .B2(n12807), .A(n12806), .ZN(P2_U2968) );
  INV_X1 U16062 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n12811) );
  AOI21_X1 U16063 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n12809), .A(n12808), .ZN(
        n12810) );
  OAI21_X1 U16064 ( .B1(n12812), .B2(n12811), .A(n12810), .ZN(P2_U2969) );
  INV_X1 U16065 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12815) );
  NAND2_X1 U16066 ( .A1(n12829), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n12814) );
  OAI211_X1 U16067 ( .C1(n12833), .C2(n12815), .A(n12814), .B(n12813), .ZN(
        P2_U2958) );
  INV_X1 U16068 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12818) );
  NAND2_X1 U16069 ( .A1(n12829), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12817) );
  OAI211_X1 U16070 ( .C1(n12833), .C2(n12818), .A(n12817), .B(n12816), .ZN(
        P2_U2966) );
  INV_X1 U16071 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n12862) );
  NAND2_X1 U16072 ( .A1(n12829), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12820) );
  OAI211_X1 U16073 ( .C1(n12833), .C2(n12862), .A(n12820), .B(n12819), .ZN(
        P2_U2961) );
  INV_X1 U16074 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n12823) );
  NAND2_X1 U16075 ( .A1(n12829), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12822) );
  OAI211_X1 U16076 ( .C1(n12833), .C2(n12823), .A(n12822), .B(n12821), .ZN(
        P2_U2962) );
  INV_X1 U16077 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n12826) );
  NAND2_X1 U16078 ( .A1(n12829), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12825) );
  OAI211_X1 U16079 ( .C1(n12833), .C2(n12826), .A(n12825), .B(n12824), .ZN(
        P2_U2960) );
  INV_X1 U16080 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14521) );
  NAND2_X1 U16081 ( .A1(n12829), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n12828) );
  OAI211_X1 U16082 ( .C1(n12833), .C2(n14521), .A(n12828), .B(n12827), .ZN(
        P2_U2965) );
  INV_X1 U16083 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14686) );
  NAND2_X1 U16084 ( .A1(n12829), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12831) );
  OAI211_X1 U16085 ( .C1(n12833), .C2(n14686), .A(n12831), .B(n12830), .ZN(
        P2_U2963) );
  INV_X1 U16086 ( .A(n12832), .ZN(n12834) );
  OAI21_X1 U16087 ( .B1(n13312), .B2(n12834), .A(n12833), .ZN(n12836) );
  INV_X1 U16088 ( .A(n12835), .ZN(n19856) );
  OR2_X1 U16089 ( .A1(n19150), .A2(n12837), .ZN(n19113) );
  NAND2_X1 U16090 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n12876) );
  OR2_X1 U16091 ( .A1(n12876), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16210) );
  NAND2_X1 U16092 ( .A1(n16210), .A2(n19150), .ZN(n19117) );
  INV_X2 U16093 ( .A(n16210), .ZN(n19148) );
  AOI22_X1 U16094 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n19147), .B1(n19148), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12838) );
  OAI21_X1 U16095 ( .B1(n12823), .B2(n19113), .A(n12838), .ZN(P2_U2925) );
  INV_X1 U16096 ( .A(n12840), .ZN(n12845) );
  OR3_X1 U16097 ( .A1(n12843), .A2(n12842), .A3(n12841), .ZN(n12844) );
  NAND2_X1 U16098 ( .A1(n12845), .A2(n12844), .ZN(n12847) );
  NOR2_X1 U16099 ( .A1(n12979), .A2(n19870), .ZN(n12848) );
  NAND2_X1 U16100 ( .A1(n12839), .A2(n12848), .ZN(n12873) );
  INV_X1 U16101 ( .A(n12873), .ZN(n12851) );
  INV_X1 U16102 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20860) );
  AND2_X1 U16104 ( .A1(n20701), .A2(n20753), .ZN(n13511) );
  INV_X1 U16105 ( .A(n13511), .ZN(n12850) );
  OAI211_X1 U16106 ( .C1(n12851), .C2(n20860), .A(n13078), .B(n12850), .ZN(
        P1_U2801) );
  INV_X1 U16107 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14640) );
  AOI22_X1 U16108 ( .A1(P2_UWORD_REG_12__SCAN_IN), .A2(n19148), .B1(n19147), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12852) );
  OAI21_X1 U16109 ( .B1(n14640), .B2(n19113), .A(n12852), .ZN(P2_U2923) );
  INV_X1 U16110 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14564) );
  AOI22_X1 U16111 ( .A1(n19148), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12853) );
  OAI21_X1 U16112 ( .B1(n14564), .B2(n19113), .A(n12853), .ZN(P2_U2934) );
  INV_X1 U16113 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n12855) );
  AOI22_X1 U16114 ( .A1(n19148), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12854) );
  OAI21_X1 U16115 ( .B1(n12855), .B2(n19113), .A(n12854), .ZN(P2_U2933) );
  INV_X1 U16116 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n12857) );
  AOI22_X1 U16117 ( .A1(n19148), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12856) );
  OAI21_X1 U16118 ( .B1(n12857), .B2(n19113), .A(n12856), .ZN(P2_U2935) );
  INV_X1 U16119 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12859) );
  AOI22_X1 U16120 ( .A1(n19148), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12858) );
  OAI21_X1 U16121 ( .B1(n12859), .B2(n19113), .A(n12858), .ZN(P2_U2931) );
  AOI22_X1 U16122 ( .A1(n19148), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12860) );
  OAI21_X1 U16123 ( .B1(n12826), .B2(n19113), .A(n12860), .ZN(P2_U2927) );
  AOI22_X1 U16124 ( .A1(n19148), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12861) );
  OAI21_X1 U16125 ( .B1(n12862), .B2(n19113), .A(n12861), .ZN(P2_U2926) );
  INV_X1 U16126 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U16127 ( .A1(n19148), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12863) );
  OAI21_X1 U16128 ( .B1(n12864), .B2(n19113), .A(n12863), .ZN(P2_U2928) );
  AOI22_X1 U16129 ( .A1(n19148), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12865) );
  OAI21_X1 U16130 ( .B1(n14686), .B2(n19113), .A(n12865), .ZN(P2_U2924) );
  AOI22_X1 U16131 ( .A1(n19148), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12866) );
  OAI21_X1 U16132 ( .B1(n12815), .B2(n19113), .A(n12866), .ZN(P2_U2929) );
  INV_X1 U16133 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n12868) );
  AOI22_X1 U16134 ( .A1(n19148), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12867) );
  OAI21_X1 U16135 ( .B1(n12868), .B2(n19113), .A(n12867), .ZN(P2_U2932) );
  AOI22_X1 U16136 ( .A1(n19148), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12869) );
  OAI21_X1 U16137 ( .B1(n14521), .B2(n19113), .A(n12869), .ZN(P2_U2922) );
  AOI22_X1 U16138 ( .A1(n19148), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12870) );
  OAI21_X1 U16139 ( .B1(n12871), .B2(n19113), .A(n12870), .ZN(P2_U2930) );
  INV_X1 U16140 ( .A(n12872), .ZN(n12875) );
  OAI21_X1 U16141 ( .B1(n13511), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n20848), 
        .ZN(n12874) );
  OAI21_X1 U16142 ( .B1(n12875), .B2(n20848), .A(n12874), .ZN(P1_U3487) );
  OAI21_X1 U16143 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n19855), .ZN(n19859) );
  INV_X1 U16144 ( .A(n12876), .ZN(n13383) );
  NOR2_X1 U16145 ( .A1(n19859), .A2(n13383), .ZN(n12877) );
  NAND2_X1 U16146 ( .A1(n19838), .A2(n16220), .ZN(n12878) );
  NAND2_X1 U16147 ( .A1(n12879), .A2(n12878), .ZN(n12880) );
  NAND2_X1 U16148 ( .A1(n12880), .A2(n19700), .ZN(n18792) );
  OAI21_X1 U16149 ( .B1(n13582), .B2(n15009), .A(n12881), .ZN(n12882) );
  XNOR2_X1 U16150 ( .A(n12882), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n19154) );
  NAND2_X1 U16151 ( .A1(n19844), .A2(n19587), .ZN(n19799) );
  INV_X1 U16152 ( .A(n19799), .ZN(n19702) );
  OR2_X1 U16153 ( .A1(n19806), .A2(n19702), .ZN(n19848) );
  NAND2_X1 U16154 ( .A1(n19848), .A2(n19855), .ZN(n12883) );
  NAND2_X1 U16155 ( .A1(n19797), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12884) );
  NAND2_X1 U16156 ( .A1(n12885), .A2(n12884), .ZN(n15005) );
  INV_X1 U16157 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13586) );
  OAI21_X1 U16158 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12887), .A(
        n12886), .ZN(n12888) );
  INV_X1 U16159 ( .A(n12888), .ZN(n19161) );
  INV_X1 U16160 ( .A(n18966), .ZN(n18992) );
  NOR2_X1 U16161 ( .A1(n18974), .A2(n19731), .ZN(n19160) );
  NOR2_X1 U16162 ( .A1(n16161), .A2(n13586), .ZN(n12889) );
  AOI211_X1 U16163 ( .C1(n16146), .C2(n19161), .A(n19160), .B(n12889), .ZN(
        n12890) );
  OAI21_X1 U16164 ( .B1(n16150), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n12890), .ZN(n12891) );
  AOI21_X1 U16165 ( .B1(n16145), .B2(n19154), .A(n12891), .ZN(n12892) );
  OAI21_X1 U16166 ( .B1(n19158), .B2(n16138), .A(n12892), .ZN(P2_U3013) );
  AND2_X1 U16167 ( .A1(n12893), .A2(n19850), .ZN(n13372) );
  AOI22_X1 U16168 ( .A1(n13334), .A2(n13336), .B1(n13374), .B2(n13372), .ZN(
        n13317) );
  NAND2_X1 U16169 ( .A1(n13317), .A2(n12896), .ZN(n12897) );
  NOR2_X1 U16170 ( .A1(n15345), .A2(n19102), .ZN(n14509) );
  NAND2_X1 U16171 ( .A1(n14509), .A2(n10349), .ZN(n13398) );
  XNOR2_X1 U16172 ( .A(n12899), .B(n12898), .ZN(n18987) );
  OR2_X1 U16173 ( .A1(n12900), .A2(n19102), .ZN(n16085) );
  INV_X1 U16174 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19136) );
  OAI222_X1 U16175 ( .A1(n13398), .A2(n19191), .B1(n18987), .B2(n19111), .C1(
        n19136), .C2(n14687), .ZN(P2_U2913) );
  INV_X1 U16176 ( .A(n13149), .ZN(n13193) );
  NAND2_X1 U16177 ( .A1(n13193), .A2(n12901), .ZN(n12905) );
  AND2_X1 U16178 ( .A1(n20146), .A2(n9614), .ZN(n13274) );
  NAND2_X1 U16179 ( .A1(n13154), .A2(n20162), .ZN(n12903) );
  NAND2_X1 U16180 ( .A1(n12903), .A2(n12902), .ZN(n12904) );
  AOI21_X1 U16181 ( .B1(n12905), .B2(n13274), .A(n12904), .ZN(n12909) );
  INV_X1 U16182 ( .A(n12906), .ZN(n20169) );
  NAND2_X1 U16183 ( .A1(n12907), .A2(n13879), .ZN(n12908) );
  NAND2_X1 U16184 ( .A1(n12909), .A2(n12908), .ZN(n12995) );
  OR2_X1 U16185 ( .A1(n11152), .A2(n15548), .ZN(n13035) );
  NAND2_X1 U16186 ( .A1(n12974), .A2(n11171), .ZN(n13030) );
  NAND3_X1 U16187 ( .A1(n13030), .A2(n15541), .A3(n12910), .ZN(n12911) );
  NAND2_X1 U16188 ( .A1(n12911), .A2(n13006), .ZN(n12913) );
  NAND2_X1 U16189 ( .A1(n12839), .A2(n12979), .ZN(n12912) );
  OAI211_X1 U16190 ( .C1(n13006), .C2(n13045), .A(n12913), .B(n12912), .ZN(
        n12914) );
  NAND2_X1 U16191 ( .A1(n12914), .A2(n11154), .ZN(n15540) );
  OR2_X1 U16192 ( .A1(n12915), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15584) );
  INV_X1 U16193 ( .A(n15584), .ZN(n15547) );
  NOR3_X1 U16194 ( .A1(n11171), .A2(n13874), .A3(n15547), .ZN(n12916) );
  NAND2_X1 U16195 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20769) );
  INV_X1 U16196 ( .A(n20769), .ZN(n20851) );
  NOR2_X1 U16197 ( .A1(n12916), .A2(n20851), .ZN(n20852) );
  OAI21_X1 U16198 ( .B1(n9848), .B2(n12979), .A(n9782), .ZN(n12918) );
  OAI21_X1 U16199 ( .B1(n11171), .B2(n15553), .A(n12918), .ZN(n19869) );
  NOR2_X1 U16200 ( .A1(n20852), .A2(n19869), .ZN(n15538) );
  OR2_X1 U16201 ( .A1(n19870), .A2(n15538), .ZN(n19876) );
  INV_X1 U16202 ( .A(n19876), .ZN(n12920) );
  INV_X1 U16203 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12919) );
  OR2_X1 U16204 ( .A1(n12920), .A2(n12919), .ZN(n12921) );
  OAI21_X1 U16205 ( .B1(n15540), .B2(n19876), .A(n12921), .ZN(P1_U3484) );
  MUX2_X1 U16206 ( .A(n19158), .B(n10398), .S(n19084), .Z(n12925) );
  OAI21_X1 U16207 ( .B1(n19808), .B2(n19075), .A(n12925), .ZN(P2_U2886) );
  NAND2_X1 U16208 ( .A1(n12927), .A2(n12926), .ZN(n12929) );
  AND2_X1 U16209 ( .A1(n12929), .A2(n10048), .ZN(n14422) );
  INV_X1 U16210 ( .A(n12930), .ZN(n13478) );
  OAI21_X1 U16211 ( .B1(n13478), .B2(n12931), .A(n13479), .ZN(n12945) );
  INV_X1 U16212 ( .A(n13480), .ZN(n12943) );
  NOR2_X1 U16213 ( .A1(n12932), .A2(n19163), .ZN(n12942) );
  XNOR2_X1 U16214 ( .A(n12934), .B(n12933), .ZN(n12951) );
  NAND2_X1 U16215 ( .A1(n9617), .A2(n16203), .ZN(n12940) );
  INV_X1 U16216 ( .A(n12935), .ZN(n12936) );
  AOI21_X1 U16217 ( .B1(n12938), .B2(n12937), .A(n12936), .ZN(n12954) );
  AOI22_X1 U16218 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n18992), .B1(n16200), 
        .B2(n12954), .ZN(n12939) );
  OAI211_X1 U16219 ( .C1(n16189), .C2(n12951), .A(n12940), .B(n12939), .ZN(
        n12941) );
  AOI211_X1 U16220 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n12943), .A(
        n12942), .B(n12941), .ZN(n12944) );
  OAI211_X1 U16221 ( .C1(n14422), .C2(n16184), .A(n12945), .B(n12944), .ZN(
        P2_U3044) );
  OR2_X1 U16222 ( .A1(n12947), .A2(n12946), .ZN(n12949) );
  NAND2_X1 U16223 ( .A1(n12949), .A2(n12948), .ZN(n18969) );
  INV_X1 U16224 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19134) );
  OAI222_X1 U16225 ( .A1(n13398), .A2(n15348), .B1(n18969), .B2(n19111), .C1(
        n19134), .C2(n14687), .ZN(P2_U2912) );
  AOI22_X1 U16226 ( .A1(n16142), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n18992), .B2(P2_REIP_REG_2__SCAN_IN), .ZN(n12950) );
  OAI21_X1 U16227 ( .B1(n16150), .B2(n14417), .A(n12950), .ZN(n12953) );
  OAI22_X1 U16228 ( .A1(n12969), .A2(n16138), .B1(n12951), .B2(n16154), .ZN(
        n12952) );
  AOI211_X1 U16229 ( .C1(n16145), .C2(n12954), .A(n12953), .B(n12952), .ZN(
        n12955) );
  INV_X1 U16230 ( .A(n12955), .ZN(P2_U3012) );
  NAND2_X1 U16231 ( .A1(n15338), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12956) );
  NAND4_X1 U16232 ( .A1(n19188), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12956), 
        .A4(n19587), .ZN(n12957) );
  AOI21_X1 U16233 ( .B1(n19826), .B2(n19105), .A(n19096), .ZN(n12963) );
  XNOR2_X1 U16234 ( .A(n12959), .B(n12958), .ZN(n19031) );
  NOR2_X1 U16235 ( .A1(n13398), .A2(n19091), .ZN(n12961) );
  INV_X1 U16236 ( .A(n19031), .ZN(n16198) );
  NOR3_X1 U16237 ( .A1(n19826), .A2(n16198), .A3(n16083), .ZN(n12960) );
  AOI211_X1 U16238 ( .C1(P2_EAX_REG_0__SCAN_IN), .C2(n19102), .A(n12961), .B(
        n12960), .ZN(n12962) );
  OAI21_X1 U16239 ( .B1(n12963), .B2(n19031), .A(n12962), .ZN(P2_U2919) );
  NOR2_X1 U16240 ( .A1(n19084), .A2(n19023), .ZN(n12964) );
  AOI21_X1 U16241 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19084), .A(n12964), .ZN(
        n12965) );
  OAI21_X1 U16242 ( .B1(n19826), .B2(n19075), .A(n12965), .ZN(P2_U2887) );
  MUX2_X1 U16243 ( .A(n12969), .B(n10420), .S(n19084), .Z(n12970) );
  OAI21_X1 U16244 ( .B1(n19807), .B2(n19075), .A(n12970), .ZN(P2_U2885) );
  NAND2_X1 U16245 ( .A1(n12839), .A2(n9614), .ZN(n15583) );
  NAND2_X1 U16246 ( .A1(n12971), .A2(n11154), .ZN(n13159) );
  NAND2_X1 U16247 ( .A1(n15583), .A2(n13159), .ZN(n12972) );
  NAND4_X1 U16248 ( .A1(n12972), .A2(n20769), .A3(n15547), .A4(n15553), .ZN(
        n12977) );
  NAND3_X1 U16249 ( .A1(n12973), .A2(n19976), .A3(n13035), .ZN(n12993) );
  NAND2_X1 U16250 ( .A1(n12974), .A2(n12993), .ZN(n12975) );
  NAND2_X1 U16251 ( .A1(n9848), .A2(n12975), .ZN(n13038) );
  NAND2_X1 U16252 ( .A1(n13274), .A2(n11776), .ZN(n12976) );
  NAND4_X1 U16253 ( .A1(n12977), .A2(n13038), .A3(n13404), .A4(n12976), .ZN(
        n12983) );
  NOR2_X1 U16254 ( .A1(n20851), .A2(n12979), .ZN(n13032) );
  INV_X1 U16255 ( .A(n13032), .ZN(n12982) );
  NAND3_X1 U16256 ( .A1(n12849), .A2(n20769), .A3(n9614), .ZN(n12980) );
  NOR2_X1 U16257 ( .A1(n12983), .A2(n13151), .ZN(n15529) );
  OR2_X1 U16258 ( .A1(n15529), .A2(n19870), .ZN(n12985) );
  NAND2_X1 U16259 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15980) );
  NOR2_X1 U16260 ( .A1(n20754), .A2(n15980), .ZN(n13210) );
  AOI22_X1 U16261 ( .A1(n20754), .A2(P1_STATE2_REG_3__SCAN_IN), .B1(n13210), 
        .B2(P1_FLUSH_REG_SCAN_IN), .ZN(n12984) );
  NAND2_X1 U16262 ( .A1(n12985), .A2(n12984), .ZN(n20836) );
  INV_X1 U16263 ( .A(n20305), .ZN(n20568) );
  NOR2_X1 U16264 ( .A1(n12986), .A2(n20568), .ZN(n12987) );
  XNOR2_X1 U16265 ( .A(n12987), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13205) );
  INV_X1 U16266 ( .A(n13205), .ZN(n19938) );
  INV_X1 U16267 ( .A(n12978), .ZN(n12988) );
  NAND4_X1 U16268 ( .A1(n19938), .A2(n14410), .A3(n12988), .A4(n20836), .ZN(
        n12989) );
  OAI21_X1 U16269 ( .B1(n12990), .B2(n20836), .A(n12989), .ZN(P1_U3468) );
  INV_X1 U16270 ( .A(n11161), .ZN(n12992) );
  NAND2_X1 U16271 ( .A1(n12992), .A2(n11171), .ZN(n12997) );
  INV_X1 U16272 ( .A(n12993), .ZN(n12994) );
  NOR2_X1 U16273 ( .A1(n12995), .A2(n12994), .ZN(n12996) );
  AND2_X1 U16274 ( .A1(n12997), .A2(n12996), .ZN(n13047) );
  AND2_X1 U16275 ( .A1(n13048), .A2(n13159), .ZN(n12998) );
  NAND3_X1 U16276 ( .A1(n13047), .A2(n12978), .A3(n12998), .ZN(n14409) );
  INV_X1 U16277 ( .A(n14409), .ZN(n13199) );
  XNOR2_X1 U16278 ( .A(n12999), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13000) );
  INV_X1 U16279 ( .A(n13000), .ZN(n13007) );
  AND2_X1 U16280 ( .A1(n13149), .A2(n13007), .ZN(n13004) );
  XNOR2_X1 U16281 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13002) );
  NAND2_X1 U16282 ( .A1(n13045), .A2(n13030), .ZN(n13196) );
  NAND2_X1 U16283 ( .A1(n13196), .A2(n13000), .ZN(n13001) );
  OAI21_X1 U16284 ( .B1(n15583), .B2(n13002), .A(n13001), .ZN(n13003) );
  AOI21_X1 U16285 ( .B1(n13199), .B2(n13004), .A(n13003), .ZN(n13005) );
  OAI21_X1 U16286 ( .B1(n12991), .B2(n13199), .A(n13005), .ZN(n13200) );
  INV_X1 U16287 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20110) );
  NOR2_X1 U16288 ( .A1(n20753), .A2(n20110), .ZN(n14412) );
  INV_X1 U16289 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15566) );
  OAI22_X1 U16290 ( .A1(n20135), .A2(n15566), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14413) );
  INV_X1 U16291 ( .A(n14413), .ZN(n13008) );
  INV_X1 U16292 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20570) );
  AOI222_X1 U16293 ( .A1(n13200), .A2(n14410), .B1(n14412), .B2(n13008), .C1(
        n13007), .C2(n13016), .ZN(n13010) );
  INV_X1 U16294 ( .A(n20836), .ZN(n13020) );
  NAND2_X1 U16295 ( .A1(n13020), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13009) );
  OAI21_X1 U16296 ( .B1(n13010), .B2(n13020), .A(n13009), .ZN(P1_U3472) );
  INV_X1 U16297 ( .A(n14715), .ZN(n13015) );
  OR2_X1 U16298 ( .A1(n13011), .A2(n10044), .ZN(n13013) );
  INV_X1 U16299 ( .A(n13025), .ZN(n13012) );
  AND2_X1 U16300 ( .A1(n13013), .A2(n13012), .ZN(n18958) );
  INV_X1 U16301 ( .A(n18958), .ZN(n13014) );
  INV_X1 U16302 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19132) );
  OAI222_X1 U16303 ( .A1(n13398), .A2(n13015), .B1(n13014), .B2(n19111), .C1(
        n19132), .C2(n14687), .ZN(P2_U2911) );
  INV_X1 U16304 ( .A(n11289), .ZN(n13213) );
  OAI22_X1 U16305 ( .A1(n13213), .A2(n13199), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14406), .ZN(n15526) );
  OAI22_X1 U16306 ( .A1(n20753), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20832), .ZN(n13017) );
  AOI21_X1 U16307 ( .B1(n15526), .B2(n14410), .A(n13017), .ZN(n13021) );
  NOR2_X1 U16308 ( .A1(n15583), .A2(n13018), .ZN(n15527) );
  AOI22_X1 U16309 ( .A1(n13020), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n14410), .B2(n15527), .ZN(n13019) );
  OAI21_X1 U16310 ( .B1(n13021), .B2(n13020), .A(n13019), .ZN(P1_U3474) );
  INV_X1 U16311 ( .A(n13022), .ZN(n14706) );
  INV_X1 U16312 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19130) );
  OAI21_X1 U16313 ( .B1(n13025), .B2(n13024), .A(n13023), .ZN(n18951) );
  OAI222_X1 U16314 ( .A1(n13398), .A2(n14706), .B1(n14687), .B2(n19130), .C1(
        n19111), .C2(n18951), .ZN(P2_U2910) );
  INV_X1 U16315 ( .A(n14697), .ZN(n13027) );
  INV_X1 U16316 ( .A(n13026), .ZN(n13073) );
  XNOR2_X1 U16317 ( .A(n13023), .B(n13073), .ZN(n18936) );
  INV_X1 U16318 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19128) );
  OAI222_X1 U16319 ( .A1(n13398), .A2(n13027), .B1(n18936), .B2(n19111), .C1(
        n19128), .C2(n14687), .ZN(P2_U2909) );
  XNOR2_X1 U16320 ( .A(n13028), .B(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20090) );
  OAI211_X1 U16321 ( .C1(n13054), .C2(n13053), .A(n15541), .B(n13030), .ZN(
        n13031) );
  NOR2_X1 U16322 ( .A1(n13029), .A2(n13031), .ZN(n13044) );
  NAND2_X1 U16323 ( .A1(n9614), .A2(n15584), .ZN(n13033) );
  NAND3_X1 U16324 ( .A1(n13033), .A2(n13032), .A3(n20162), .ZN(n13034) );
  OAI21_X1 U16325 ( .B1(n15553), .B2(n13035), .A(n13034), .ZN(n13036) );
  INV_X1 U16326 ( .A(n13036), .ZN(n13037) );
  NAND2_X1 U16327 ( .A1(n13038), .A2(n13037), .ZN(n13043) );
  OR2_X1 U16328 ( .A1(n9614), .A2(n15547), .ZN(n13268) );
  NAND2_X1 U16329 ( .A1(n13268), .A2(n20769), .ZN(n13039) );
  OAI211_X1 U16330 ( .C1(n13159), .C2(n13039), .A(n19976), .B(n13154), .ZN(
        n13040) );
  NAND2_X1 U16331 ( .A1(n13040), .A2(n11776), .ZN(n13041) );
  NOR2_X1 U16332 ( .A1(n15585), .A2(n13041), .ZN(n13042) );
  INV_X1 U16333 ( .A(n20092), .ZN(n20109) );
  OAI211_X1 U16334 ( .C1(n13048), .C2(n19976), .A(n13047), .B(n13046), .ZN(
        n13049) );
  INV_X1 U16335 ( .A(n13049), .ZN(n13050) );
  OR2_X1 U16336 ( .A1(n13050), .A2(n13058), .ZN(n14345) );
  NAND2_X1 U16337 ( .A1(n20109), .A2(n14345), .ZN(n13051) );
  AND2_X1 U16338 ( .A1(n20114), .A2(n13058), .ZN(n14348) );
  AOI21_X1 U16339 ( .B1(n20110), .B2(n13051), .A(n14348), .ZN(n20134) );
  INV_X1 U16340 ( .A(n20134), .ZN(n13052) );
  OAI22_X1 U16341 ( .A1(n13052), .A2(n14344), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13051), .ZN(n13064) );
  NAND2_X1 U16342 ( .A1(n12849), .A2(n15548), .ZN(n15582) );
  INV_X1 U16343 ( .A(n13053), .ZN(n13055) );
  NAND2_X1 U16344 ( .A1(n13055), .A2(n13054), .ZN(n13056) );
  AND2_X1 U16345 ( .A1(n15582), .A2(n13056), .ZN(n13057) );
  OR2_X1 U16346 ( .A1(n13879), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13061) );
  NAND2_X1 U16347 ( .A1(n13415), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13060) );
  INV_X1 U16348 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13284) );
  NAND2_X1 U16349 ( .A1(n13894), .A2(n13284), .ZN(n13059) );
  NAND2_X1 U16350 ( .A1(n13060), .A2(n13059), .ZN(n13409) );
  NAND2_X1 U16351 ( .A1(n13061), .A2(n13409), .ZN(n13604) );
  INV_X1 U16352 ( .A(n13604), .ZN(n13062) );
  AOI22_X1 U16353 ( .A1(n20131), .A2(n13062), .B1(n20128), .B2(
        P1_REIP_REG_0__SCAN_IN), .ZN(n13063) );
  OAI211_X1 U16354 ( .C1(n20090), .C2(n20120), .A(n13064), .B(n13063), .ZN(
        P1_U3031) );
  NOR2_X1 U16355 ( .A1(n19826), .A2(n19031), .ZN(n13069) );
  XNOR2_X1 U16356 ( .A(n13066), .B(n13065), .ZN(n19819) );
  INV_X1 U16357 ( .A(n19819), .ZN(n13067) );
  NAND2_X1 U16358 ( .A1(n19808), .A2(n13067), .ZN(n13166) );
  OAI21_X1 U16359 ( .B1(n19808), .B2(n13067), .A(n13166), .ZN(n13068) );
  NOR2_X1 U16360 ( .A1(n13068), .A2(n13069), .ZN(n13168) );
  AOI21_X1 U16361 ( .B1(n13069), .B2(n13068), .A(n13168), .ZN(n13072) );
  AOI22_X1 U16362 ( .A1(n19096), .A2(n19819), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19102), .ZN(n13071) );
  INV_X1 U16363 ( .A(n13398), .ZN(n19104) );
  INV_X1 U16364 ( .A(n15340), .ZN(n14754) );
  NAND2_X1 U16365 ( .A1(n19104), .A2(n14754), .ZN(n13070) );
  OAI211_X1 U16366 ( .C1(n13072), .C2(n16083), .A(n13071), .B(n13070), .ZN(
        P2_U2918) );
  INV_X1 U16367 ( .A(n14689), .ZN(n13076) );
  NOR2_X1 U16368 ( .A1(n13023), .A2(n13073), .ZN(n13075) );
  OAI21_X1 U16369 ( .B1(n13075), .B2(n13074), .A(n9649), .ZN(n18920) );
  INV_X1 U16370 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19126) );
  OAI222_X1 U16371 ( .A1(n13398), .A2(n13076), .B1(n18920), .B2(n19111), .C1(
        n19126), .C2(n14687), .ZN(P2_U2908) );
  AND2_X1 U16372 ( .A1(n11172), .A2(n20851), .ZN(n13077) );
  AND2_X2 U16373 ( .A1(n13138), .A2(n15548), .ZN(n13133) );
  INV_X2 U16374 ( .A(n13138), .ZN(n20064) );
  AOI22_X1 U16375 ( .A1(n13133), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13081) );
  NAND2_X1 U16376 ( .A1(n13138), .A2(n9614), .ZN(n13139) );
  INV_X1 U16377 ( .A(DATAI_5_), .ZN(n13080) );
  NAND2_X1 U16378 ( .A1(n14158), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13079) );
  OAI21_X1 U16379 ( .B1(n14158), .B2(n13080), .A(n13079), .ZN(n20184) );
  NAND2_X1 U16380 ( .A1(n20052), .A2(n20184), .ZN(n13093) );
  NAND2_X1 U16381 ( .A1(n13081), .A2(n13093), .ZN(P1_U2942) );
  AOI22_X1 U16382 ( .A1(n13133), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13084) );
  INV_X1 U16383 ( .A(DATAI_6_), .ZN(n13083) );
  NAND2_X1 U16384 ( .A1(n14158), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13082) );
  OAI21_X1 U16385 ( .B1(n14158), .B2(n13083), .A(n13082), .ZN(n20190) );
  NAND2_X1 U16386 ( .A1(n20052), .A2(n20190), .ZN(n13101) );
  NAND2_X1 U16387 ( .A1(n13084), .A2(n13101), .ZN(P1_U2943) );
  AOI22_X1 U16388 ( .A1(n13133), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13087) );
  INV_X1 U16389 ( .A(DATAI_7_), .ZN(n13086) );
  NAND2_X1 U16390 ( .A1(n14158), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13085) );
  OAI21_X1 U16391 ( .B1(n14158), .B2(n13086), .A(n13085), .ZN(n20198) );
  NAND2_X1 U16392 ( .A1(n20052), .A2(n20198), .ZN(n13091) );
  NAND2_X1 U16393 ( .A1(n13087), .A2(n13091), .ZN(P1_U2944) );
  AOI22_X1 U16394 ( .A1(n13133), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13090) );
  INV_X1 U16395 ( .A(DATAI_1_), .ZN(n13089) );
  NAND2_X1 U16396 ( .A1(n14158), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13088) );
  OAI21_X1 U16397 ( .B1(n14158), .B2(n13089), .A(n13088), .ZN(n20159) );
  NAND2_X1 U16398 ( .A1(n20052), .A2(n20159), .ZN(n13431) );
  NAND2_X1 U16399 ( .A1(n13090), .A2(n13431), .ZN(P1_U2938) );
  AOI22_X1 U16400 ( .A1(n13133), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20064), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13092) );
  NAND2_X1 U16401 ( .A1(n13092), .A2(n13091), .ZN(P1_U2959) );
  AOI22_X1 U16402 ( .A1(n13133), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20064), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13094) );
  NAND2_X1 U16403 ( .A1(n13094), .A2(n13093), .ZN(P1_U2957) );
  AOI22_X1 U16404 ( .A1(n13133), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13097) );
  INV_X1 U16405 ( .A(DATAI_0_), .ZN(n13096) );
  NAND2_X1 U16406 ( .A1(n14158), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13095) );
  OAI21_X1 U16407 ( .B1(n14158), .B2(n13096), .A(n13095), .ZN(n20150) );
  NAND2_X1 U16408 ( .A1(n20052), .A2(n20150), .ZN(n13433) );
  NAND2_X1 U16409 ( .A1(n13097), .A2(n13433), .ZN(P1_U2937) );
  AOI22_X1 U16410 ( .A1(n13133), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13100) );
  INV_X1 U16411 ( .A(DATAI_3_), .ZN(n13099) );
  NAND2_X1 U16412 ( .A1(n14158), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13098) );
  OAI21_X1 U16413 ( .B1(n14158), .B2(n13099), .A(n13098), .ZN(n20172) );
  NAND2_X1 U16414 ( .A1(n20052), .A2(n20172), .ZN(n13112) );
  NAND2_X1 U16415 ( .A1(n13100), .A2(n13112), .ZN(P1_U2940) );
  AOI22_X1 U16416 ( .A1(n13133), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20064), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13102) );
  NAND2_X1 U16417 ( .A1(n13102), .A2(n13101), .ZN(P1_U2958) );
  AOI22_X1 U16418 ( .A1(n13133), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13105) );
  INV_X1 U16419 ( .A(DATAI_4_), .ZN(n13104) );
  NAND2_X1 U16420 ( .A1(n14158), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13103) );
  OAI21_X1 U16421 ( .B1(n14158), .B2(n13104), .A(n13103), .ZN(n20178) );
  NAND2_X1 U16422 ( .A1(n20052), .A2(n20178), .ZN(n13114) );
  NAND2_X1 U16423 ( .A1(n13105), .A2(n13114), .ZN(P1_U2941) );
  AOI22_X1 U16424 ( .A1(n13133), .A2(P1_EAX_REG_24__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13108) );
  INV_X1 U16425 ( .A(DATAI_8_), .ZN(n13107) );
  NAND2_X1 U16426 ( .A1(n14158), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13106) );
  OAI21_X1 U16427 ( .B1(n14158), .B2(n13107), .A(n13106), .ZN(n14121) );
  NAND2_X1 U16428 ( .A1(n20052), .A2(n14121), .ZN(n13134) );
  NAND2_X1 U16429 ( .A1(n13108), .A2(n13134), .ZN(P1_U2945) );
  AOI22_X1 U16430 ( .A1(n13133), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13111) );
  INV_X1 U16431 ( .A(DATAI_2_), .ZN(n13110) );
  NAND2_X1 U16432 ( .A1(n14158), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13109) );
  OAI21_X1 U16433 ( .B1(n14158), .B2(n13110), .A(n13109), .ZN(n20164) );
  NAND2_X1 U16434 ( .A1(n20052), .A2(n20164), .ZN(n13429) );
  NAND2_X1 U16435 ( .A1(n13111), .A2(n13429), .ZN(P1_U2939) );
  AOI22_X1 U16436 ( .A1(n13133), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20064), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13113) );
  NAND2_X1 U16437 ( .A1(n13113), .A2(n13112), .ZN(P1_U2955) );
  AOI22_X1 U16438 ( .A1(n13133), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20064), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13115) );
  NAND2_X1 U16439 ( .A1(n13115), .A2(n13114), .ZN(P1_U2956) );
  INV_X1 U16440 ( .A(n19073), .ZN(n13394) );
  XOR2_X1 U16441 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13394), .Z(n13120)
         );
  NAND2_X1 U16442 ( .A1(n19084), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n13119) );
  OR2_X1 U16443 ( .A1(n13482), .A2(n13116), .ZN(n13117) );
  AND2_X1 U16444 ( .A1(n13125), .A2(n13117), .ZN(n18997) );
  NAND2_X1 U16445 ( .A1(n18997), .A2(n19070), .ZN(n13118) );
  OAI211_X1 U16446 ( .C1(n13120), .C2(n19075), .A(n13119), .B(n13118), .ZN(
        P2_U2882) );
  NOR2_X1 U16447 ( .A1(n13394), .A2(n13121), .ZN(n13123) );
  OR2_X1 U16448 ( .A1(n13394), .A2(n13122), .ZN(n13140) );
  OAI211_X1 U16449 ( .C1(n13123), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n19081), .B(n13140), .ZN(n13128) );
  NAND2_X1 U16450 ( .A1(n13125), .A2(n13124), .ZN(n13126) );
  AND2_X1 U16451 ( .A1(n13142), .A2(n13126), .ZN(n18983) );
  NAND2_X1 U16452 ( .A1(n18983), .A2(n19070), .ZN(n13127) );
  OAI211_X1 U16453 ( .C1(n19070), .C2(n18976), .A(n13128), .B(n13127), .ZN(
        P2_U2881) );
  XOR2_X1 U16454 ( .A(n19060), .B(n19062), .Z(n13132) );
  INV_X1 U16455 ( .A(n16103), .ZN(n13129) );
  AOI21_X1 U16456 ( .B1(n9734), .B2(n16135), .A(n13129), .ZN(n18947) );
  NOR2_X1 U16457 ( .A1(n19070), .A2(n10988), .ZN(n13130) );
  AOI21_X1 U16458 ( .B1(n18947), .B2(n19070), .A(n13130), .ZN(n13131) );
  OAI21_X1 U16459 ( .B1(n13132), .B2(n19075), .A(n13131), .ZN(P2_U2878) );
  INV_X1 U16460 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20019) );
  NAND2_X1 U16461 ( .A1(n20064), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13135) );
  OAI211_X1 U16462 ( .C1(n13428), .C2(n20019), .A(n13135), .B(n13134), .ZN(
        P1_U2960) );
  INV_X1 U16463 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13644) );
  NOR2_X1 U16464 ( .A1(n20147), .A2(n13136), .ZN(n13137) );
  AOI21_X1 U16465 ( .B1(DATAI_15_), .B2(n20147), .A(n13137), .ZN(n13643) );
  INV_X1 U16466 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20007) );
  OAI222_X1 U16467 ( .A1(n13428), .A2(n13644), .B1(n13139), .B2(n13643), .C1(
        n13138), .C2(n20007), .ZN(P1_U2967) );
  XOR2_X1 U16468 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13140), .Z(n13145)
         );
  AND2_X1 U16469 ( .A1(n13142), .A2(n13141), .ZN(n13143) );
  OR2_X1 U16470 ( .A1(n16137), .A2(n13143), .ZN(n18968) );
  MUX2_X1 U16471 ( .A(n18968), .B(n10981), .S(n19084), .Z(n13144) );
  OAI21_X1 U16472 ( .B1(n13145), .B2(n19075), .A(n13144), .ZN(P2_U2880) );
  AOI21_X1 U16473 ( .B1(n10046), .B2(n9649), .A(n9725), .ZN(n18915) );
  INV_X1 U16474 ( .A(n18915), .ZN(n13147) );
  INV_X1 U16475 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19124) );
  OAI222_X1 U16476 ( .A1(n13398), .A2(n14677), .B1(n13147), .B2(n19111), .C1(
        n19124), .C2(n14687), .ZN(P2_U2907) );
  NOR2_X1 U16477 ( .A1(n20182), .A2(n20176), .ZN(n13148) );
  NAND4_X1 U16478 ( .A1(n13149), .A2(n13810), .A3(n13148), .A4(n20188), .ZN(
        n13402) );
  INV_X1 U16479 ( .A(n11171), .ZN(n13261) );
  NOR2_X1 U16480 ( .A1(n13402), .A2(n13261), .ZN(n13150) );
  AND2_X1 U16481 ( .A1(n13159), .A2(n13154), .ZN(n13155) );
  INV_X1 U16482 ( .A(n13156), .ZN(n13157) );
  AOI21_X1 U16483 ( .B1(n13158), .B2(n13399), .A(n13157), .ZN(n13179) );
  INV_X1 U16484 ( .A(n13179), .ZN(n14011) );
  INV_X1 U16485 ( .A(n20164), .ZN(n13163) );
  INV_X1 U16486 ( .A(n13159), .ZN(n13160) );
  NAND2_X1 U16487 ( .A1(n19972), .A2(n13161), .ZN(n13813) );
  INV_X1 U16488 ( .A(n13813), .ZN(n13162) );
  INV_X1 U16489 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20032) );
  OAI222_X1 U16490 ( .A1(n19975), .A2(n14011), .B1(n13163), .B2(n19974), .C1(
        n19972), .C2(n20032), .ZN(P1_U2902) );
  INV_X1 U16491 ( .A(n14523), .ZN(n13165) );
  OAI21_X1 U16492 ( .B1(n9725), .B2(n13164), .A(n13221), .ZN(n18909) );
  INV_X1 U16493 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19122) );
  OAI222_X1 U16494 ( .A1(n13398), .A2(n13165), .B1(n18909), .B2(n19111), .C1(
        n19122), .C2(n14687), .ZN(P2_U2906) );
  INV_X1 U16495 ( .A(n13166), .ZN(n13167) );
  NOR2_X1 U16496 ( .A1(n13168), .A2(n13167), .ZN(n13170) );
  NAND2_X1 U16497 ( .A1(n19807), .A2(n14422), .ZN(n13224) );
  OAI21_X1 U16498 ( .B1(n19807), .B2(n14422), .A(n13224), .ZN(n13169) );
  NOR2_X1 U16499 ( .A1(n13170), .A2(n13169), .ZN(n13226) );
  AOI21_X1 U16500 ( .B1(n13170), .B2(n13169), .A(n13226), .ZN(n13174) );
  INV_X1 U16501 ( .A(n16089), .ZN(n13171) );
  AOI22_X1 U16502 ( .A1(n19104), .A2(n13171), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19102), .ZN(n13173) );
  INV_X1 U16503 ( .A(n14422), .ZN(n19811) );
  NAND2_X1 U16504 ( .A1(n19811), .A2(n19096), .ZN(n13172) );
  OAI211_X1 U16505 ( .C1(n13174), .C2(n16083), .A(n13173), .B(n13172), .ZN(
        P2_U2917) );
  XNOR2_X1 U16506 ( .A(n13175), .B(n13176), .ZN(n20121) );
  AOI22_X1 U16507 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13177) );
  OAI21_X1 U16508 ( .B1(n20075), .B2(n14000), .A(n13177), .ZN(n13178) );
  AOI21_X1 U16509 ( .B1(n13179), .B2(n20070), .A(n13178), .ZN(n13180) );
  OAI21_X1 U16510 ( .B1(n20121), .B2(n20089), .A(n13180), .ZN(P1_U2997) );
  INV_X1 U16511 ( .A(n13249), .ZN(n13181) );
  OAI21_X1 U16512 ( .B1(n13183), .B2(n13182), .A(n13181), .ZN(n13999) );
  INV_X1 U16513 ( .A(n20172), .ZN(n13184) );
  INV_X1 U16514 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20030) );
  OAI222_X1 U16515 ( .A1(n19975), .A2(n13999), .B1(n13184), .B2(n19974), .C1(
        n19972), .C2(n20030), .ZN(P1_U2901) );
  INV_X1 U16516 ( .A(n20428), .ZN(n14401) );
  MUX2_X1 U16517 ( .A(n13185), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n12999), .Z(n13187) );
  NOR2_X1 U16518 ( .A1(n13187), .A2(n13186), .ZN(n13197) );
  NAND2_X1 U16519 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13189) );
  INV_X1 U16520 ( .A(n13189), .ZN(n13188) );
  MUX2_X1 U16521 ( .A(n13189), .B(n13188), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13190) );
  NOR2_X1 U16522 ( .A1(n15583), .A2(n13190), .ZN(n13195) );
  INV_X1 U16523 ( .A(n13185), .ZN(n13191) );
  OAI211_X1 U16524 ( .C1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n12999), .A(
        n13192), .B(n13191), .ZN(n20833) );
  NOR3_X1 U16525 ( .A1(n14409), .A2(n13193), .A3(n20833), .ZN(n13194) );
  AOI211_X1 U16526 ( .C1(n13197), .C2(n13196), .A(n13195), .B(n13194), .ZN(
        n13198) );
  OAI21_X1 U16527 ( .B1(n14401), .B2(n13199), .A(n13198), .ZN(n20831) );
  MUX2_X1 U16528 ( .A(n20831), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15529), .Z(n15534) );
  NOR2_X1 U16529 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20753), .ZN(n13206) );
  AOI22_X1 U16530 ( .A1(n15534), .A2(n20753), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13206), .ZN(n13202) );
  INV_X1 U16531 ( .A(n15529), .ZN(n13204) );
  MUX2_X1 U16532 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13200), .S(
        n13204), .Z(n15532) );
  AOI22_X1 U16533 ( .A1(n13206), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15532), .B2(n20753), .ZN(n13201) );
  NOR2_X1 U16534 ( .A1(n13202), .A2(n13201), .ZN(n15544) );
  INV_X1 U16535 ( .A(n15544), .ZN(n13209) );
  INV_X1 U16536 ( .A(n13203), .ZN(n14405) );
  OAI21_X1 U16537 ( .B1(n13205), .B2(n12978), .A(n13204), .ZN(n13208) );
  AOI21_X1 U16538 ( .B1(n15529), .B2(n12990), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13207) );
  AOI22_X1 U16539 ( .A1(n13208), .A2(n13207), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13206), .ZN(n15542) );
  OAI21_X1 U16540 ( .B1(n13209), .B2(n13203), .A(n15542), .ZN(n13212) );
  OAI21_X1 U16541 ( .B1(n13212), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13210), .ZN(
        n13211) );
  INV_X1 U16542 ( .A(n15980), .ZN(n15975) );
  NAND2_X1 U16543 ( .A1(n11268), .A2(n20753), .ZN(n15977) );
  NAND2_X1 U16544 ( .A1(n20754), .A2(n15977), .ZN(n20853) );
  INV_X1 U16545 ( .A(n20197), .ZN(n20310) );
  NAND2_X1 U16546 ( .A1(n13211), .A2(n20310), .ZN(n20137) );
  NOR2_X1 U16547 ( .A1(n13212), .A2(n15980), .ZN(n15556) );
  INV_X1 U16548 ( .A(n20617), .ZN(n20693) );
  AND2_X1 U16549 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20570), .ZN(n14400) );
  OAI22_X1 U16550 ( .A1(n11869), .A2(n20693), .B1(n13213), .B2(n14400), .ZN(
        n13214) );
  OAI21_X1 U16551 ( .B1(n15556), .B2(n13214), .A(n20137), .ZN(n13215) );
  OAI21_X1 U16552 ( .B1(n20137), .B2(n20611), .A(n13215), .ZN(P1_U3478) );
  AOI21_X1 U16553 ( .B1(n13249), .B2(n13250), .A(n13217), .ZN(n13218) );
  OR2_X1 U16554 ( .A1(n13216), .A2(n13218), .ZN(n15840) );
  INV_X1 U16555 ( .A(n20184), .ZN(n13219) );
  INV_X1 U16556 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20026) );
  OAI222_X1 U16557 ( .A1(n19975), .A2(n15840), .B1(n13219), .B2(n19974), .C1(
        n19972), .C2(n20026), .ZN(P1_U2899) );
  INV_X1 U16558 ( .A(n14512), .ZN(n13223) );
  AND2_X1 U16559 ( .A1(n13221), .A2(n13220), .ZN(n13222) );
  OR2_X1 U16560 ( .A1(n13222), .A2(n13239), .ZN(n15212) );
  INV_X1 U16561 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19120) );
  OAI222_X1 U16562 ( .A1(n13398), .A2(n13223), .B1(n15212), .B2(n19111), .C1(
        n19120), .C2(n14687), .ZN(P2_U2905) );
  INV_X1 U16563 ( .A(n13224), .ZN(n13225) );
  NOR2_X1 U16564 ( .A1(n13226), .A2(n13225), .ZN(n13234) );
  OR2_X1 U16565 ( .A1(n13231), .A2(n13230), .ZN(n13232) );
  NAND2_X1 U16566 ( .A1(n13232), .A2(n13384), .ZN(n16185) );
  XNOR2_X1 U16567 ( .A(n19791), .B(n16185), .ZN(n13233) );
  NOR2_X1 U16568 ( .A1(n13234), .A2(n13233), .ZN(n13390) );
  AOI21_X1 U16569 ( .B1(n13234), .B2(n13233), .A(n13390), .ZN(n13237) );
  INV_X1 U16570 ( .A(n19173), .ZN(n14746) );
  AOI22_X1 U16571 ( .A1(n19104), .A2(n14746), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19102), .ZN(n13236) );
  INV_X1 U16572 ( .A(n16185), .ZN(n19802) );
  NAND2_X1 U16573 ( .A1(n19802), .A2(n19096), .ZN(n13235) );
  OAI211_X1 U16574 ( .C1(n13237), .C2(n16083), .A(n13236), .B(n13235), .ZN(
        P2_U2916) );
  NOR2_X1 U16575 ( .A1(n13239), .A2(n13238), .ZN(n13240) );
  OR2_X1 U16576 ( .A1(n15187), .A2(n13240), .ZN(n18889) );
  OAI222_X1 U16577 ( .A1(n18889), .A2(n19111), .B1(n13398), .B2(n13241), .C1(
        n12722), .C2(n14687), .ZN(P2_U2904) );
  AND2_X1 U16578 ( .A1(n16105), .A2(n13242), .ZN(n13243) );
  OR2_X1 U16579 ( .A1(n13243), .A2(n14970), .ZN(n18929) );
  INV_X1 U16580 ( .A(n18929), .ZN(n15248) );
  NOR2_X1 U16581 ( .A1(n19070), .A2(n13244), .ZN(n13247) );
  AOI211_X1 U16582 ( .C1(n13245), .C2(n19063), .A(n19075), .B(n19054), .ZN(
        n13246) );
  AOI211_X1 U16583 ( .C1(n15248), .C2(n19070), .A(n13247), .B(n13246), .ZN(
        n13248) );
  INV_X1 U16584 ( .A(n13248), .ZN(P2_U2876) );
  XOR2_X1 U16585 ( .A(n13250), .B(n13249), .Z(n20069) );
  INV_X1 U16586 ( .A(n20069), .ZN(n13439) );
  INV_X1 U16587 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20028) );
  INV_X1 U16588 ( .A(n20178), .ZN(n13251) );
  OAI222_X1 U16589 ( .A1(n19975), .A2(n13439), .B1(n20028), .B2(n19972), .C1(
        n13251), .C2(n19974), .ZN(P1_U2900) );
  OAI21_X1 U16590 ( .B1(n13216), .B2(n13252), .A(n13446), .ZN(n19919) );
  INV_X1 U16591 ( .A(n20190), .ZN(n13253) );
  INV_X1 U16592 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20024) );
  OAI222_X1 U16593 ( .A1(n19975), .A2(n19919), .B1(n19974), .B2(n13253), .C1(
        n19972), .C2(n20024), .ZN(P1_U2898) );
  NAND2_X1 U16594 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20754), .ZN(n13255) );
  NOR2_X1 U16595 ( .A1(n20570), .A2(n15977), .ZN(n15555) );
  NAND2_X1 U16596 ( .A1(n15555), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13254) );
  OAI211_X1 U16597 ( .C1(n13255), .C2(n13797), .A(n13254), .B(n20114), .ZN(
        n13256) );
  INV_X1 U16598 ( .A(n13256), .ZN(n13257) );
  INV_X1 U16599 ( .A(n13803), .ZN(n13258) );
  NAND2_X1 U16600 ( .A1(n13258), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13259) );
  XNOR2_X1 U16601 ( .A(n13259), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13824) );
  AND2_X1 U16602 ( .A1(n13824), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13260) );
  OR2_X1 U16603 ( .A1(n13276), .A2(n13261), .ZN(n13262) );
  INV_X1 U16604 ( .A(n13263), .ZN(n13267) );
  INV_X1 U16605 ( .A(n13264), .ZN(n13266) );
  OAI21_X1 U16606 ( .B1(n13267), .B2(n13266), .A(n13265), .ZN(n20083) );
  OR2_X1 U16607 ( .A1(n13276), .A2(n20146), .ZN(n13281) );
  NAND2_X1 U16608 ( .A1(n20769), .A2(n14399), .ZN(n13271) );
  INV_X1 U16609 ( .A(n13271), .ZN(n15546) );
  NAND2_X1 U16610 ( .A1(n13268), .A2(n15546), .ZN(n13278) );
  INV_X1 U16611 ( .A(n13278), .ZN(n13269) );
  NAND2_X1 U16612 ( .A1(n19958), .A2(n19931), .ZN(n15681) );
  INV_X1 U16613 ( .A(n15681), .ZN(n13970) );
  INV_X1 U16614 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20844) );
  AND2_X1 U16615 ( .A1(n9614), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13277) );
  NAND2_X1 U16616 ( .A1(n13277), .A2(n13271), .ZN(n13272) );
  NOR2_X2 U16617 ( .A1(n13281), .A2(n13272), .ZN(n19926) );
  OAI22_X1 U16618 ( .A1(n13970), .A2(n20844), .B1(n19952), .B2(n13604), .ZN(
        n13273) );
  INV_X1 U16619 ( .A(n13273), .ZN(n13287) );
  INV_X1 U16620 ( .A(n13274), .ZN(n13275) );
  OR2_X1 U16621 ( .A1(n13276), .A2(n13275), .ZN(n14005) );
  INV_X1 U16622 ( .A(n14005), .ZN(n19953) );
  INV_X1 U16623 ( .A(n13277), .ZN(n13279) );
  NAND2_X1 U16624 ( .A1(n13279), .A2(n13278), .ZN(n13280) );
  NOR2_X2 U16625 ( .A1(n13281), .A2(n13280), .ZN(n19937) );
  NOR2_X1 U16626 ( .A1(n13824), .A2(n20753), .ZN(n13282) );
  OAI21_X1 U16627 ( .B1(n19955), .B2(n19961), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13283) );
  OAI21_X1 U16628 ( .B1(n19950), .B2(n13284), .A(n13283), .ZN(n13285) );
  AOI21_X1 U16629 ( .B1(n11289), .B2(n19953), .A(n13285), .ZN(n13286) );
  OAI211_X1 U16630 ( .C1(n19963), .C2(n20083), .A(n13287), .B(n13286), .ZN(
        P1_U2840) );
  AOI21_X1 U16631 ( .B1(n13288), .B2(n14972), .A(n9720), .ZN(n18905) );
  INV_X1 U16632 ( .A(n18905), .ZN(n14961) );
  INV_X1 U16633 ( .A(n9709), .ZN(n19048) );
  OAI211_X1 U16634 ( .C1(n13289), .C2(n13290), .A(n19048), .B(n19081), .ZN(
        n13292) );
  NAND2_X1 U16635 ( .A1(n19084), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13291) );
  OAI211_X1 U16636 ( .C1(n14961), .C2(n19084), .A(n13292), .B(n13291), .ZN(
        P2_U2874) );
  INV_X1 U16637 ( .A(n13356), .ZN(n13350) );
  NAND2_X1 U16638 ( .A1(n13293), .A2(n13350), .ZN(n13311) );
  NAND2_X1 U16639 ( .A1(n13294), .A2(n11023), .ZN(n13331) );
  INV_X1 U16640 ( .A(n13295), .ZN(n13296) );
  OAI21_X1 U16641 ( .B1(n13297), .B2(n10259), .A(n13296), .ZN(n13309) );
  INV_X1 U16642 ( .A(n13336), .ZN(n13298) );
  NAND2_X1 U16643 ( .A1(n13299), .A2(n13298), .ZN(n13323) );
  INV_X1 U16644 ( .A(n13300), .ZN(n13302) );
  NAND2_X1 U16645 ( .A1(n13302), .A2(n13301), .ZN(n13320) );
  XNOR2_X1 U16646 ( .A(n13320), .B(n10259), .ZN(n13303) );
  NAND2_X1 U16647 ( .A1(n13323), .A2(n13303), .ZN(n13307) );
  INV_X1 U16648 ( .A(n13304), .ZN(n13305) );
  OAI211_X1 U16649 ( .C1(n10315), .C2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11022), .B(n13305), .ZN(n13306) );
  NAND2_X1 U16650 ( .A1(n13307), .A2(n13306), .ZN(n13308) );
  AOI21_X1 U16651 ( .B1(n13331), .B2(n13309), .A(n13308), .ZN(n13310) );
  NAND2_X1 U16652 ( .A1(n13311), .A2(n13310), .ZN(n19788) );
  INV_X1 U16653 ( .A(n13312), .ZN(n13315) );
  NOR2_X1 U16654 ( .A1(n15492), .A2(n13313), .ZN(n13314) );
  NAND2_X1 U16655 ( .A1(n13315), .A2(n13314), .ZN(n13318) );
  AND4_X1 U16656 ( .A1(n13319), .A2(n13318), .A3(n13317), .A4(n13316), .ZN(
        n13563) );
  INV_X1 U16657 ( .A(n13563), .ZN(n13357) );
  MUX2_X1 U16658 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n19788), .S(
        n13357), .Z(n13380) );
  NAND2_X1 U16659 ( .A1(n14425), .A2(n13350), .ZN(n13333) );
  NAND2_X1 U16660 ( .A1(n13321), .A2(n13320), .ZN(n13322) );
  INV_X1 U16661 ( .A(n13322), .ZN(n13330) );
  NAND2_X1 U16662 ( .A1(n13323), .A2(n13322), .ZN(n13328) );
  INV_X1 U16663 ( .A(n13324), .ZN(n13326) );
  NAND3_X1 U16664 ( .A1(n11022), .A2(n13326), .A3(n13325), .ZN(n13327) );
  NAND2_X1 U16665 ( .A1(n13328), .A2(n13327), .ZN(n13329) );
  AOI21_X1 U16666 ( .B1(n13331), .B2(n13330), .A(n13329), .ZN(n13332) );
  NAND2_X1 U16667 ( .A1(n13333), .A2(n13332), .ZN(n15320) );
  MUX2_X1 U16668 ( .A(n15320), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n13563), .Z(n13379) );
  NAND2_X1 U16669 ( .A1(n13563), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13377) );
  NAND2_X1 U16670 ( .A1(n13335), .A2(n13334), .ZN(n13343) );
  NAND2_X1 U16671 ( .A1(n13337), .A2(n13336), .ZN(n13342) );
  INV_X1 U16672 ( .A(n13338), .ZN(n13339) );
  NAND2_X1 U16673 ( .A1(n13340), .A2(n13339), .ZN(n13341) );
  AND3_X1 U16674 ( .A1(n13343), .A2(n13342), .A3(n13341), .ZN(n19840) );
  INV_X1 U16675 ( .A(n10374), .ZN(n13370) );
  NAND2_X1 U16676 ( .A1(n19852), .A2(n15490), .ZN(n13367) );
  AND2_X1 U16677 ( .A1(n13379), .A2(n19805), .ZN(n13365) );
  INV_X1 U16678 ( .A(n13380), .ZN(n13363) );
  INV_X1 U16679 ( .A(n11022), .ZN(n13354) );
  NAND2_X1 U16680 ( .A1(n13345), .A2(n13344), .ZN(n13352) );
  OAI21_X1 U16681 ( .B1(n13347), .B2(n13346), .A(n13352), .ZN(n13348) );
  OAI21_X1 U16682 ( .B1(n13354), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13348), .ZN(n13349) );
  AOI21_X1 U16683 ( .B1(n13351), .B2(n13350), .A(n13349), .ZN(n13577) );
  INV_X1 U16684 ( .A(n13352), .ZN(n13353) );
  MUX2_X1 U16685 ( .A(n13354), .B(n13353), .S(n10170), .Z(n13355) );
  OAI21_X1 U16686 ( .B1(n19023), .B2(n13356), .A(n13355), .ZN(n13561) );
  OAI21_X1 U16687 ( .B1(n19830), .B2(n13561), .A(n19821), .ZN(n13360) );
  NOR2_X1 U16688 ( .A1(n13365), .A2(n19813), .ZN(n13359) );
  OAI21_X1 U16689 ( .B1(n13561), .B2(n19511), .A(n13357), .ZN(n13358) );
  AOI211_X1 U16690 ( .C1(n13577), .C2(n13360), .A(n13359), .B(n13358), .ZN(
        n13361) );
  OAI21_X1 U16691 ( .B1(n13380), .B2(n19805), .A(n13361), .ZN(n13362) );
  OAI21_X1 U16692 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13363), .A(
        n13362), .ZN(n13364) );
  AOI21_X1 U16693 ( .B1(n13365), .B2(n19813), .A(n13364), .ZN(n13366) );
  OAI22_X1 U16694 ( .A1(n15492), .A2(n13367), .B1(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n13366), .ZN(n13368) );
  AOI21_X1 U16695 ( .B1(n13370), .B2(n13369), .A(n13368), .ZN(n13376) );
  NOR2_X1 U16696 ( .A1(n13372), .A2(n13371), .ZN(n13373) );
  AND2_X1 U16697 ( .A1(n13374), .A2(n13373), .ZN(n18791) );
  OAI21_X1 U16698 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18791), .ZN(n13375) );
  NAND4_X1 U16699 ( .A1(n13377), .A2(n19840), .A3(n13376), .A4(n13375), .ZN(
        n13378) );
  AOI21_X1 U16700 ( .B1(n13380), .B2(n13379), .A(n13378), .ZN(n16217) );
  OAI211_X1 U16701 ( .C1(n13382), .C2(n13381), .A(n16217), .B(n19700), .ZN(
        n16211) );
  NAND2_X1 U16702 ( .A1(n19855), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13562) );
  NAND2_X1 U16703 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13383), .ZN(n15599) );
  OAI211_X1 U16704 ( .C1(n16211), .C2(n19587), .A(n13562), .B(n15599), .ZN(
        P2_U3593) );
  INV_X1 U16705 ( .A(n19791), .ZN(n19803) );
  NOR2_X1 U16706 ( .A1(n19803), .A2(n19802), .ZN(n13389) );
  INV_X1 U16707 ( .A(n13384), .ZN(n13385) );
  OR2_X1 U16708 ( .A1(n13386), .A2(n13385), .ZN(n13388) );
  INV_X1 U16709 ( .A(n15306), .ZN(n13387) );
  NAND2_X1 U16710 ( .A1(n13388), .A2(n13387), .ZN(n13486) );
  OAI21_X1 U16711 ( .B1(n13390), .B2(n13389), .A(n13486), .ZN(n19107) );
  OR2_X1 U16712 ( .A1(n13391), .A2(n13392), .ZN(n13393) );
  NAND2_X1 U16713 ( .A1(n13394), .A2(n13393), .ZN(n19080) );
  XNOR2_X1 U16714 ( .A(n19107), .B(n19080), .ZN(n13395) );
  NAND2_X1 U16715 ( .A1(n13395), .A2(n19105), .ZN(n13397) );
  INV_X1 U16716 ( .A(n13486), .ZN(n19009) );
  AOI22_X1 U16717 ( .A1(n19096), .A2(n19009), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19102), .ZN(n13396) );
  OAI211_X1 U16718 ( .C1(n16081), .C2(n13398), .A(n13397), .B(n13396), .ZN(
        P2_U2915) );
  OAI21_X1 U16719 ( .B1(n13401), .B2(n13400), .A(n13399), .ZN(n20082) );
  NAND2_X2 U16720 ( .A1(n19970), .A2(n11154), .ZN(n14078) );
  INV_X1 U16721 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n19949) );
  NAND2_X1 U16722 ( .A1(n13868), .A2(n19949), .ZN(n13408) );
  NAND2_X1 U16723 ( .A1(n13415), .A2(n20135), .ZN(n13406) );
  NAND2_X1 U16724 ( .A1(n13874), .A2(n19949), .ZN(n13405) );
  NAND3_X1 U16725 ( .A1(n13406), .A2(n13894), .A3(n13405), .ZN(n13407) );
  NAND2_X1 U16726 ( .A1(n13408), .A2(n13407), .ZN(n13413) );
  XNOR2_X1 U16727 ( .A(n13413), .B(n13409), .ZN(n13410) );
  NAND2_X1 U16728 ( .A1(n13410), .A2(n13874), .ZN(n13414) );
  OR2_X1 U16729 ( .A1(n13410), .A2(n13874), .ZN(n13411) );
  NAND2_X1 U16730 ( .A1(n13414), .A2(n13411), .ZN(n20132) );
  AOI22_X1 U16731 ( .A1(n19965), .A2(n20132), .B1(n14068), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13412) );
  OAI21_X1 U16732 ( .B1(n20082), .B2(n14078), .A(n13412), .ZN(P1_U2871) );
  NAND2_X1 U16733 ( .A1(n13414), .A2(n13413), .ZN(n13553) );
  INV_X1 U16734 ( .A(n13415), .ZN(n13416) );
  NAND2_X1 U16735 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n9777), .ZN(
        n13417) );
  MUX2_X1 U16736 ( .A(n13867), .B(n13894), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13419) );
  OAI21_X1 U16737 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13879), .A(
        n13419), .ZN(n13601) );
  MUX2_X1 U16738 ( .A(n13877), .B(n13415), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13422) );
  NAND2_X1 U16739 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n9777), .ZN(
        n13420) );
  AND2_X1 U16740 ( .A1(n13857), .A2(n13420), .ZN(n13421) );
  NAND2_X1 U16741 ( .A1(n13422), .A2(n13421), .ZN(n13438) );
  MUX2_X1 U16742 ( .A(n13867), .B(n13894), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n13423) );
  OAI21_X1 U16743 ( .B1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n13879), .A(
        n13423), .ZN(n13550) );
  MUX2_X1 U16744 ( .A(n13877), .B(n13415), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13426) );
  NAND2_X1 U16745 ( .A1(n9777), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13424) );
  AND2_X1 U16746 ( .A1(n13857), .A2(n13424), .ZN(n13425) );
  NAND2_X1 U16747 ( .A1(n13426), .A2(n13425), .ZN(n13591) );
  XNOR2_X1 U16748 ( .A(n13594), .B(n13591), .ZN(n19917) );
  AOI22_X1 U16749 ( .A1(n19917), .A2(n19965), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14068), .ZN(n13427) );
  OAI21_X1 U16750 ( .B1(n19919), .B2(n14078), .A(n13427), .ZN(P1_U2866) );
  AOI22_X1 U16751 ( .A1(n13133), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20064), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13430) );
  NAND2_X1 U16752 ( .A1(n13430), .A2(n13429), .ZN(P1_U2954) );
  AOI22_X1 U16753 ( .A1(n13133), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20064), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13432) );
  NAND2_X1 U16754 ( .A1(n13432), .A2(n13431), .ZN(P1_U2953) );
  AOI22_X1 U16755 ( .A1(n13133), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20064), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13434) );
  NAND2_X1 U16756 ( .A1(n13434), .A2(n13433), .ZN(P1_U2952) );
  AOI21_X1 U16757 ( .B1(n13436), .B2(n10078), .A(n10164), .ZN(n14260) );
  INV_X1 U16758 ( .A(n14260), .ZN(n13988) );
  AOI22_X1 U16759 ( .A1(n15759), .A2(n14121), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15760), .ZN(n13437) );
  OAI21_X1 U16760 ( .B1(n13988), .B2(n19975), .A(n13437), .ZN(P1_U2896) );
  OAI21_X1 U16761 ( .B1(n13600), .B2(n13438), .A(n13549), .ZN(n20094) );
  INV_X1 U16762 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13440) );
  OAI222_X1 U16763 ( .A1(n14098), .A2(n20094), .B1(n13440), .B2(n19970), .C1(
        n14078), .C2(n13439), .ZN(P1_U2868) );
  OAI21_X1 U16764 ( .B1(n10164), .B2(n13442), .A(n13497), .ZN(n15828) );
  INV_X1 U16765 ( .A(DATAI_9_), .ZN(n13444) );
  NAND2_X1 U16766 ( .A1(n14158), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13443) );
  OAI21_X1 U16767 ( .B1(n14158), .B2(n13444), .A(n13443), .ZN(n20040) );
  AOI22_X1 U16768 ( .A1(n15759), .A2(n20040), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15760), .ZN(n13445) );
  OAI21_X1 U16769 ( .B1(n15828), .B2(n19975), .A(n13445), .ZN(P1_U2895) );
  AOI21_X1 U16770 ( .B1(n13447), .B2(n13446), .A(n13435), .ZN(n19906) );
  INV_X1 U16771 ( .A(n19906), .ZN(n13598) );
  INV_X1 U16772 ( .A(n20198), .ZN(n13448) );
  INV_X1 U16773 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20021) );
  OAI222_X1 U16774 ( .A1(n19975), .A2(n13598), .B1(n13448), .B2(n19974), .C1(
        n19972), .C2(n20021), .ZN(P1_U2897) );
  XNOR2_X1 U16775 ( .A(n13449), .B(n13450), .ZN(n16190) );
  XNOR2_X1 U16776 ( .A(n13451), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13452) );
  XNOR2_X1 U16777 ( .A(n13453), .B(n13452), .ZN(n16192) );
  NAND2_X1 U16778 ( .A1(n16192), .A2(n16145), .ZN(n13459) );
  INV_X1 U16779 ( .A(n16138), .ZN(n16157) );
  NAND2_X1 U16780 ( .A1(n16151), .A2(n13522), .ZN(n13456) );
  NOR2_X1 U16781 ( .A1(n18974), .A2(n13454), .ZN(n16187) );
  INV_X1 U16782 ( .A(n16187), .ZN(n13455) );
  OAI211_X1 U16783 ( .C1(n13524), .C2(n16161), .A(n13456), .B(n13455), .ZN(
        n13457) );
  AOI21_X1 U16784 ( .B1(n13293), .B2(n16157), .A(n13457), .ZN(n13458) );
  OAI211_X1 U16785 ( .C1(n16190), .C2(n16154), .A(n13459), .B(n13458), .ZN(
        P2_U3011) );
  NOR2_X1 U16786 ( .A1(n19048), .A2(n19049), .ZN(n13463) );
  INV_X1 U16787 ( .A(n13460), .ZN(n13462) );
  OR2_X1 U16788 ( .A1(n19048), .A2(n13461), .ZN(n19044) );
  OAI211_X1 U16789 ( .C1(n13463), .C2(n13462), .A(n19081), .B(n19044), .ZN(
        n13466) );
  AOI21_X1 U16790 ( .B1(n13464), .B2(n14944), .A(n14923), .ZN(n18886) );
  NAND2_X1 U16791 ( .A1(n18886), .A2(n19070), .ZN(n13465) );
  OAI211_X1 U16792 ( .C1(n19070), .C2(n11010), .A(n13466), .B(n13465), .ZN(
        P2_U2872) );
  AOI21_X1 U16793 ( .B1(n13469), .B2(n13468), .A(n13467), .ZN(n20104) );
  NAND2_X1 U16794 ( .A1(n20104), .A2(n20071), .ZN(n13472) );
  AND2_X1 U16795 ( .A1(n20128), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20101) );
  NOR2_X1 U16796 ( .A1(n20075), .A2(n13990), .ZN(n13470) );
  AOI211_X1 U16797 ( .C1(n20086), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20101), .B(n13470), .ZN(n13471) );
  OAI211_X1 U16798 ( .C1(n20149), .C2(n13999), .A(n13472), .B(n13471), .ZN(
        P1_U2996) );
  XNOR2_X1 U16799 ( .A(n13474), .B(n13473), .ZN(n13495) );
  OR2_X1 U16800 ( .A1(n16195), .A2(n16196), .ZN(n15305) );
  AOI21_X1 U16801 ( .B1(n13479), .B2(n13478), .A(n13477), .ZN(n16194) );
  INV_X1 U16802 ( .A(n16194), .ZN(n15272) );
  NAND2_X1 U16803 ( .A1(n16209), .A2(n13480), .ZN(n15058) );
  OAI21_X1 U16804 ( .B1(n16195), .B2(n15272), .A(n15058), .ZN(n15309) );
  NAND2_X1 U16805 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n18992), .ZN(n13481) );
  OAI221_X1 U16806 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15305), .C1(
        n13475), .C2(n15309), .A(n13481), .ZN(n13488) );
  INV_X1 U16807 ( .A(n13482), .ZN(n13483) );
  OAI21_X1 U16808 ( .B1(n13485), .B2(n13484), .A(n13483), .ZN(n19083) );
  OAI22_X1 U16809 ( .A1(n19083), .A2(n19157), .B1(n16184), .B2(n13486), .ZN(
        n13487) );
  AOI211_X1 U16810 ( .C1(n13493), .C2(n19162), .A(n13488), .B(n13487), .ZN(
        n13489) );
  OAI21_X1 U16811 ( .B1(n13495), .B2(n19155), .A(n13489), .ZN(P2_U3042) );
  OAI22_X1 U16812 ( .A1(n10972), .A2(n18974), .B1(n16150), .B2(n19014), .ZN(
        n13492) );
  INV_X1 U16813 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13490) );
  OAI22_X1 U16814 ( .A1(n19083), .A2(n16138), .B1(n16161), .B2(n13490), .ZN(
        n13491) );
  AOI211_X1 U16815 ( .C1(n13493), .C2(n16146), .A(n13492), .B(n13491), .ZN(
        n13494) );
  OAI21_X1 U16816 ( .B1(n13495), .B2(n16152), .A(n13494), .ZN(P2_U3010) );
  INV_X1 U16817 ( .A(n13964), .ZN(n13496) );
  AOI21_X1 U16818 ( .B1(n13498), .B2(n13497), .A(n13496), .ZN(n14251) );
  INV_X1 U16819 ( .A(n14251), .ZN(n13556) );
  INV_X1 U16820 ( .A(n14249), .ZN(n13515) );
  MUX2_X1 U16821 ( .A(n13867), .B(n13894), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n13499) );
  OAI21_X1 U16822 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n13879), .A(
        n13499), .ZN(n13592) );
  INV_X1 U16823 ( .A(n13592), .ZN(n13500) );
  MUX2_X1 U16824 ( .A(n13877), .B(n13415), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13503) );
  NAND2_X1 U16825 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n9777), .ZN(
        n13501) );
  AND2_X1 U16826 ( .A1(n13857), .A2(n13501), .ZN(n13502) );
  NAND2_X1 U16827 ( .A1(n13503), .A2(n13502), .ZN(n13558) );
  INV_X1 U16828 ( .A(n13867), .ZN(n13859) );
  INV_X1 U16829 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n19969) );
  NAND2_X1 U16830 ( .A1(n13859), .A2(n19969), .ZN(n13506) );
  NAND2_X1 U16831 ( .A1(n13894), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13504) );
  OAI211_X1 U16832 ( .C1(n9777), .C2(P1_EBX_REG_9__SCAN_IN), .A(n13415), .B(
        n13504), .ZN(n13505) );
  MUX2_X1 U16833 ( .A(n13877), .B(n13415), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13508) );
  NAND2_X1 U16834 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n9777), .ZN(
        n13507) );
  INV_X1 U16835 ( .A(n13509), .ZN(n13510) );
  OAI21_X1 U16836 ( .B1(n9721), .B2(n13510), .A(n15731), .ZN(n15932) );
  AOI22_X1 U16837 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n19937), .B1(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19955), .ZN(n13512) );
  NAND2_X1 U16838 ( .A1(n19931), .A2(n13511), .ZN(n19910) );
  OAI211_X1 U16839 ( .C1(n15932), .C2(n19952), .A(n13512), .B(n19910), .ZN(
        n13514) );
  INV_X1 U16840 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15931) );
  INV_X1 U16841 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20787) );
  INV_X1 U16842 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20784) );
  INV_X1 U16843 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20781) );
  NAND3_X1 U16844 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19942) );
  NOR2_X1 U16845 ( .A1(n20781), .A2(n19942), .ZN(n19932) );
  NAND2_X1 U16846 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19932), .ZN(n19914) );
  NOR2_X1 U16847 ( .A1(n20784), .A2(n19914), .ZN(n19904) );
  NAND2_X1 U16848 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19904), .ZN(n13984) );
  NOR2_X1 U16849 ( .A1(n20787), .A2(n13984), .ZN(n19893) );
  OAI211_X1 U16850 ( .C1(n19893), .C2(n19958), .A(P1_REIP_REG_9__SCAN_IN), .B(
        n19931), .ZN(n19894) );
  INV_X1 U16851 ( .A(n19931), .ZN(n19954) );
  NAND3_X1 U16852 ( .A1(n19893), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_9__SCAN_IN), .ZN(n13827) );
  NOR2_X1 U16853 ( .A1(n19954), .A2(n13827), .ZN(n13971) );
  OR2_X1 U16854 ( .A1(n13970), .A2(n13971), .ZN(n15728) );
  AOI21_X1 U16855 ( .B1(n15931), .B2(n19894), .A(n15728), .ZN(n13513) );
  AOI211_X1 U16856 ( .C1(n19961), .C2(n13515), .A(n13514), .B(n13513), .ZN(
        n13516) );
  OAI21_X1 U16857 ( .B1(n13556), .B2(n19920), .A(n13516), .ZN(P1_U2830) );
  INV_X1 U16858 ( .A(DATAI_10_), .ZN(n13518) );
  NAND2_X1 U16859 ( .A1(n14158), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13517) );
  OAI21_X1 U16860 ( .B1(n14158), .B2(n13518), .A(n13517), .ZN(n20042) );
  AOI22_X1 U16861 ( .A1(n15759), .A2(n20042), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15760), .ZN(n13519) );
  OAI21_X1 U16862 ( .B1(n13556), .B2(n19975), .A(n13519), .ZN(P1_U2894) );
  NAND2_X1 U16863 ( .A1(n18994), .A2(n13520), .ZN(n13521) );
  XNOR2_X1 U16864 ( .A(n13522), .B(n13521), .ZN(n13530) );
  OAI22_X1 U16865 ( .A1(n13454), .A2(n19004), .B1(n13523), .B2(n18989), .ZN(
        n13526) );
  OAI22_X1 U16866 ( .A1(n13524), .A2(n18850), .B1(n19032), .B2(n16185), .ZN(
        n13525) );
  AOI211_X1 U16867 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19028), .A(n13526), .B(
        n13525), .ZN(n13528) );
  NAND2_X1 U16868 ( .A1(n13293), .A2(n18998), .ZN(n13527) );
  OAI211_X1 U16869 ( .C1(n19012), .C2(n19791), .A(n13528), .B(n13527), .ZN(
        n13529) );
  AOI21_X1 U16870 ( .B1(n13530), .B2(n14419), .A(n13529), .ZN(n13531) );
  INV_X1 U16871 ( .A(n13531), .ZN(P2_U2852) );
  NOR2_X1 U16872 ( .A1(n19791), .A2(n19797), .ZN(n19516) );
  INV_X1 U16873 ( .A(n19808), .ZN(n19817) );
  INV_X1 U16874 ( .A(n19796), .ZN(n13532) );
  NAND2_X1 U16875 ( .A1(n19516), .A2(n13532), .ZN(n13536) );
  OR2_X1 U16876 ( .A1(n19805), .A2(n15367), .ZN(n15378) );
  INV_X1 U16877 ( .A(n19660), .ZN(n19689) );
  AND2_X1 U16878 ( .A1(n19660), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13533) );
  NAND2_X1 U16879 ( .A1(n13534), .A2(n13533), .ZN(n13538) );
  OAI211_X1 U16880 ( .C1(n19689), .C2(n19587), .A(n19593), .B(n13538), .ZN(
        n13535) );
  INV_X1 U16881 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19843) );
  OAI21_X1 U16882 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n15378), .A(n19843), 
        .ZN(n13537) );
  NAND2_X1 U16883 ( .A1(n13538), .A2(n13537), .ZN(n19669) );
  INV_X1 U16884 ( .A(n13539), .ZN(n13544) );
  AOI22_X1 U16885 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19193), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19192), .ZN(n19524) );
  INV_X1 U16886 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16299) );
  INV_X1 U16887 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18120) );
  AOI22_X1 U16888 ( .A1(n19693), .A2(n19595), .B1(n19695), .B2(n19521), .ZN(
        n13543) );
  NAND2_X1 U16889 ( .A1(n19586), .A2(n19689), .ZN(n13542) );
  OAI211_X1 U16890 ( .C1(n19669), .C2(n13544), .A(n13543), .B(n13542), .ZN(
        n13545) );
  INV_X1 U16891 ( .A(n13545), .ZN(n13546) );
  OAI21_X1 U16892 ( .B1(n19699), .B2(n13547), .A(n13546), .ZN(P2_U3168) );
  INV_X1 U16893 ( .A(n13594), .ZN(n13548) );
  AOI21_X1 U16894 ( .B1(n13550), .B2(n13549), .A(n13548), .ZN(n19927) );
  AOI22_X1 U16895 ( .A1(n19927), .A2(n19965), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14068), .ZN(n13551) );
  OAI21_X1 U16896 ( .B1(n15840), .B2(n14078), .A(n13551), .ZN(P1_U2867) );
  NAND2_X1 U16897 ( .A1(n13553), .A2(n13552), .ZN(n13554) );
  NAND2_X1 U16898 ( .A1(n13602), .A2(n13554), .ZN(n20115) );
  OAI222_X1 U16899 ( .A1(n14011), .A2(n14078), .B1(n14091), .B2(n9967), .C1(
        n20115), .C2(n14098), .ZN(P1_U2870) );
  INV_X1 U16900 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13555) );
  OAI222_X1 U16901 ( .A1(n13556), .A2(n14078), .B1(n19970), .B2(n13555), .C1(
        n15932), .C2(n14098), .ZN(P1_U2862) );
  INV_X1 U16902 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13559) );
  INV_X1 U16903 ( .A(n13557), .ZN(n15940) );
  OAI21_X1 U16904 ( .B1(n13596), .B2(n13558), .A(n15940), .ZN(n15950) );
  OAI222_X1 U16905 ( .A1(n13988), .A2(n14078), .B1(n14091), .B2(n13559), .C1(
        n15950), .C2(n14098), .ZN(P1_U2864) );
  OAI22_X1 U16906 ( .A1(n18994), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n13575), .B2(n19016), .ZN(n13576) );
  AOI222_X1 U16907 ( .A1(n13561), .A2(n19702), .B1(n13560), .B2(n15321), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n13576), .ZN(n13566) );
  INV_X1 U16908 ( .A(n15599), .ZN(n16221) );
  OAI21_X1 U16909 ( .B1(n13563), .B2(n19849), .A(n13562), .ZN(n13564) );
  AOI21_X1 U16910 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16221), .A(n13564), .ZN(
        n19792) );
  NAND2_X1 U16911 ( .A1(n19792), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13565) );
  OAI21_X1 U16912 ( .B1(n13566), .B2(n19792), .A(n13565), .ZN(P2_U3601) );
  INV_X1 U16913 ( .A(n13567), .ZN(n13570) );
  AOI22_X1 U16914 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19193), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19192), .ZN(n19530) );
  INV_X1 U16915 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16295) );
  INV_X1 U16916 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18133) );
  OAI22_X1 U16917 ( .A1(n16295), .A2(n19186), .B1(n18133), .B2(n19184), .ZN(
        n19629) );
  AOI22_X1 U16918 ( .A1(n19693), .A2(n19630), .B1(n19695), .B2(n19629), .ZN(
        n13569) );
  NOR2_X2 U16919 ( .A1(n19189), .A2(n10372), .ZN(n19628) );
  NAND2_X1 U16920 ( .A1(n19628), .A2(n19689), .ZN(n13568) );
  OAI211_X1 U16921 ( .C1(n19669), .C2(n13570), .A(n13569), .B(n13568), .ZN(
        n13571) );
  INV_X1 U16922 ( .A(n13571), .ZN(n13572) );
  OAI21_X1 U16923 ( .B1(n19699), .B2(n13573), .A(n13572), .ZN(P2_U3170) );
  AOI211_X1 U16924 ( .C1(n13575), .C2(n13574), .A(n19016), .B(n14416), .ZN(
        n13581) );
  AOI21_X1 U16925 ( .B1(n19016), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13581), .ZN(n15324) );
  NOR2_X1 U16926 ( .A1(n19844), .A2(n13576), .ZN(n15319) );
  INV_X1 U16927 ( .A(n15321), .ZN(n19790) );
  OAI22_X1 U16928 ( .A1(n19808), .A2(n19790), .B1(n19799), .B2(n13577), .ZN(
        n13578) );
  AOI21_X1 U16929 ( .B1(n15324), .B2(n15319), .A(n13578), .ZN(n13580) );
  NAND2_X1 U16930 ( .A1(n19792), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13579) );
  OAI21_X1 U16931 ( .B1(n13580), .B2(n19792), .A(n13579), .ZN(P2_U3600) );
  NOR2_X1 U16932 ( .A1(n19705), .A2(n18994), .ZN(n19037) );
  AOI22_X1 U16933 ( .A1(n13581), .A2(n19000), .B1(n19037), .B2(n13586), .ZN(
        n13590) );
  INV_X1 U16934 ( .A(n13582), .ZN(n13584) );
  OAI22_X1 U16935 ( .A1(n19006), .A2(n10398), .B1(n19731), .B2(n19004), .ZN(
        n13583) );
  AOI21_X1 U16936 ( .B1(n19026), .B2(n13584), .A(n13583), .ZN(n13585) );
  OAI21_X1 U16937 ( .B1(n19158), .B2(n19022), .A(n13585), .ZN(n13588) );
  NOR2_X1 U16938 ( .A1(n18850), .A2(n13586), .ZN(n13587) );
  AOI211_X1 U16939 ( .C1(n19819), .C2(n19008), .A(n13588), .B(n13587), .ZN(
        n13589) );
  OAI211_X1 U16940 ( .C1(n19808), .C2(n19012), .A(n13590), .B(n13589), .ZN(
        P2_U2854) );
  INV_X1 U16941 ( .A(n13591), .ZN(n13593) );
  OAI21_X1 U16942 ( .B1(n13594), .B2(n13593), .A(n13592), .ZN(n13595) );
  INV_X1 U16943 ( .A(n13595), .ZN(n13597) );
  OR2_X1 U16944 ( .A1(n13597), .A2(n13596), .ZN(n15958) );
  INV_X1 U16945 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13599) );
  OAI222_X1 U16946 ( .A1(n15958), .A2(n14098), .B1(n13599), .B2(n19970), .C1(
        n13598), .C2(n14078), .ZN(P1_U2865) );
  AOI21_X1 U16947 ( .B1(n13602), .B2(n13601), .A(n13600), .ZN(n20102) );
  INV_X1 U16948 ( .A(n20102), .ZN(n13603) );
  INV_X1 U16949 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13991) );
  OAI222_X1 U16950 ( .A1(n13603), .A2(n14098), .B1(n14091), .B2(n13991), .C1(
        n13999), .C2(n14078), .ZN(P1_U2869) );
  OAI222_X1 U16951 ( .A1(n13604), .A2(n14098), .B1(n13284), .B2(n19970), .C1(
        n20083), .C2(n14078), .ZN(P1_U2872) );
  OAI21_X1 U16952 ( .B1(n13606), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13605), .ZN(n13608) );
  XNOR2_X1 U16953 ( .A(n13608), .B(n13607), .ZN(n14263) );
  INV_X1 U16954 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15954) );
  NAND2_X1 U16955 ( .A1(n20110), .A2(n14329), .ZN(n20126) );
  NAND3_X1 U16956 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20113), .A3(
        n20126), .ZN(n20125) );
  NAND2_X1 U16957 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20097) );
  NOR2_X1 U16958 ( .A1(n20097), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15966) );
  NAND2_X1 U16959 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20093) );
  AOI21_X1 U16960 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20091) );
  NOR2_X1 U16961 ( .A1(n15970), .A2(n20097), .ZN(n13610) );
  INV_X1 U16962 ( .A(n13610), .ZN(n14271) );
  NOR2_X1 U16963 ( .A1(n20091), .A2(n14271), .ZN(n14342) );
  AOI21_X1 U16964 ( .B1(n14328), .B2(n20110), .A(n14348), .ZN(n14270) );
  OAI21_X1 U16965 ( .B1(n14342), .B2(n20109), .A(n14270), .ZN(n14371) );
  AOI221_X1 U16966 ( .B1(n20097), .B2(n20113), .C1(n20093), .C2(n20113), .A(
        n14371), .ZN(n15971) );
  INV_X1 U16967 ( .A(n15971), .ZN(n13609) );
  AOI21_X1 U16968 ( .B1(n14378), .B2(n15966), .A(n13609), .ZN(n15947) );
  OAI22_X1 U16969 ( .A1(n15954), .A2(n15947), .B1(n15953), .B2(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13611) );
  INV_X1 U16970 ( .A(n13611), .ZN(n13613) );
  NOR2_X1 U16971 ( .A1(n20114), .A2(n20784), .ZN(n14265) );
  AOI21_X1 U16972 ( .B1(n19917), .B2(n20131), .A(n14265), .ZN(n13612) );
  OAI211_X1 U16973 ( .C1(n14263), .C2(n20120), .A(n13613), .B(n13612), .ZN(
        P1_U3025) );
  NOR2_X1 U16974 ( .A1(n13967), .A2(n13614), .ZN(n13615) );
  OR2_X1 U16975 ( .A1(n13635), .A2(n13615), .ZN(n15808) );
  INV_X1 U16976 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14370) );
  INV_X1 U16977 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15743) );
  NAND2_X1 U16978 ( .A1(n13874), .A2(n15743), .ZN(n13616) );
  OAI211_X1 U16979 ( .C1(n11170), .C2(n14370), .A(n13616), .B(n13415), .ZN(
        n13617) );
  OAI21_X1 U16980 ( .B1(n13867), .B2(P1_EBX_REG_11__SCAN_IN), .A(n13617), .ZN(
        n15730) );
  MUX2_X1 U16981 ( .A(n13877), .B(n13415), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n13619) );
  NAND2_X1 U16982 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n9777), .ZN(
        n13618) );
  MUX2_X1 U16983 ( .A(n13867), .B(n13894), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13622) );
  INV_X1 U16984 ( .A(n13879), .ZN(n13620) );
  NAND2_X1 U16985 ( .A1(n15916), .A2(n13620), .ZN(n13621) );
  NAND2_X1 U16986 ( .A1(n14096), .A2(n13974), .ZN(n13975) );
  INV_X1 U16987 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15708) );
  NAND2_X1 U16988 ( .A1(n13868), .A2(n15708), .ZN(n13626) );
  NAND2_X1 U16989 ( .A1(n13415), .A2(n15895), .ZN(n13624) );
  NAND2_X1 U16990 ( .A1(n13874), .A2(n15708), .ZN(n13623) );
  NAND3_X1 U16991 ( .A1(n13624), .A2(n13894), .A3(n13623), .ZN(n13625) );
  NAND2_X1 U16992 ( .A1(n13975), .A2(n13627), .ZN(n13628) );
  NAND2_X1 U16993 ( .A1(n13639), .A2(n13628), .ZN(n15709) );
  OAI22_X1 U16994 ( .A1(n15709), .A2(n14098), .B1(n15708), .B2(n19970), .ZN(
        n13629) );
  INV_X1 U16995 ( .A(n13629), .ZN(n13630) );
  OAI21_X1 U16996 ( .B1(n15808), .B2(n14078), .A(n13630), .ZN(P1_U2858) );
  INV_X1 U16997 ( .A(DATAI_14_), .ZN(n13632) );
  MUX2_X1 U16998 ( .A(n13632), .B(n13631), .S(n14158), .Z(n20050) );
  INV_X1 U16999 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n13633) );
  OAI222_X1 U17000 ( .A1(n15808), .A2(n19975), .B1(n20050), .B2(n19974), .C1(
        n13633), .C2(n19972), .ZN(P1_U2890) );
  OR2_X1 U17001 ( .A1(n13635), .A2(n13634), .ZN(n13636) );
  NAND2_X1 U17002 ( .A1(n9656), .A2(n13636), .ZN(n15694) );
  INV_X1 U17003 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n13642) );
  MUX2_X1 U17004 ( .A(n13867), .B(n13894), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13637) );
  OAI21_X1 U17005 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n13879), .A(
        n13637), .ZN(n13638) );
  INV_X1 U17006 ( .A(n14083), .ZN(n13641) );
  NAND2_X1 U17007 ( .A1(n13639), .A2(n13638), .ZN(n13640) );
  NAND2_X1 U17008 ( .A1(n13641), .A2(n13640), .ZN(n15905) );
  OAI222_X1 U17009 ( .A1(n15694), .A2(n14078), .B1(n19970), .B2(n13642), .C1(
        n15905), .C2(n14098), .ZN(P1_U2857) );
  OAI222_X1 U17010 ( .A1(n15694), .A2(n19975), .B1(n19972), .B2(n13644), .C1(
        n19974), .C2(n13643), .ZN(P1_U2889) );
  NAND2_X1 U17011 ( .A1(n15483), .A2(n18607), .ZN(n13645) );
  NAND2_X1 U17012 ( .A1(n18571), .A2(n13645), .ZN(n18557) );
  NOR2_X1 U17013 ( .A1(n18729), .A2(n18557), .ZN(n13662) );
  INV_X1 U17014 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18628) );
  INV_X2 U17015 ( .A(n18777), .ZN(n18758) );
  NOR2_X1 U17016 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16379) );
  INV_X1 U17017 ( .A(n16379), .ZN(n18627) );
  NAND3_X1 U17018 ( .A1(n18628), .A2(n18705), .A3(n18627), .ZN(n18635) );
  INV_X1 U17019 ( .A(n18635), .ZN(n18762) );
  NAND2_X1 U17020 ( .A1(n17348), .A2(n17347), .ZN(n18611) );
  NAND2_X1 U17021 ( .A1(n13646), .A2(n18611), .ZN(n13647) );
  INV_X1 U17022 ( .A(n16381), .ZN(n18551) );
  NAND2_X1 U17023 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18773) );
  NAND2_X1 U17024 ( .A1(n18551), .A2(n18773), .ZN(n13660) );
  AOI21_X1 U17025 ( .B1(n13652), .B2(n13651), .A(n13650), .ZN(n13653) );
  NOR2_X1 U17026 ( .A1(n13654), .A2(n13653), .ZN(n15506) );
  INV_X1 U17027 ( .A(n18773), .ZN(n18764) );
  AOI22_X1 U17028 ( .A1(n13656), .A2(n13655), .B1(n17347), .B2(n18128), .ZN(
        n13657) );
  NOR2_X1 U17029 ( .A1(n15603), .A2(n15397), .ZN(n13659) );
  OAI211_X1 U17030 ( .C1(n17309), .C2(n13660), .A(n15506), .B(n13659), .ZN(
        n18582) );
  NOR3_X1 U17031 ( .A1(n18726), .A2(n18767), .A3(n18779), .ZN(n18623) );
  INV_X1 U17032 ( .A(n18623), .ZN(n18716) );
  INV_X1 U17033 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18114) );
  OAI22_X1 U17034 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18743), .B1(n18716), 
        .B2(n18114), .ZN(n13661) );
  MUX2_X1 U17035 ( .A(n13662), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18748), .Z(P3_U3284) );
  NOR2_X1 U17036 ( .A1(n19070), .A2(n13663), .ZN(n13664) );
  AOI21_X1 U17037 ( .B1(n13293), .B2(n19070), .A(n13664), .ZN(n13665) );
  OAI21_X1 U17038 ( .B1(n19791), .B2(n19075), .A(n13665), .ZN(P2_U2884) );
  NOR2_X1 U17039 ( .A1(n13666), .A2(n13709), .ZN(n13667) );
  INV_X1 U17040 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15048) );
  NOR2_X1 U17041 ( .A1(n13706), .A2(n14466), .ZN(n13668) );
  NAND2_X1 U17042 ( .A1(n19180), .A2(n13668), .ZN(n13669) );
  AND2_X1 U17043 ( .A1(n13712), .A2(n13669), .ZN(n13670) );
  NAND2_X1 U17044 ( .A1(n13708), .A2(n13670), .ZN(n16035) );
  INV_X1 U17045 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15073) );
  NAND2_X1 U17046 ( .A1(n19180), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13673) );
  MUX2_X1 U17047 ( .A(n19180), .B(n13673), .S(n13672), .Z(n13674) );
  NAND2_X1 U17048 ( .A1(n13674), .A2(n13682), .ZN(n18826) );
  OR2_X1 U17049 ( .A1(n18826), .A2(n10733), .ZN(n13675) );
  INV_X1 U17050 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14866) );
  NAND2_X1 U17051 ( .A1(n13675), .A2(n14866), .ZN(n14870) );
  XNOR2_X1 U17052 ( .A(n13676), .B(n9724), .ZN(n18836) );
  NAND2_X1 U17053 ( .A1(n18836), .A2(n13728), .ZN(n13688) );
  INV_X1 U17054 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14882) );
  NAND2_X1 U17055 ( .A1(n13688), .A2(n14882), .ZN(n14884) );
  INV_X1 U17056 ( .A(n13677), .ZN(n13678) );
  XNOR2_X1 U17057 ( .A(n13679), .B(n13678), .ZN(n18847) );
  NAND2_X1 U17058 ( .A1(n18847), .A2(n13728), .ZN(n13680) );
  INV_X1 U17059 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15176) );
  NAND2_X1 U17060 ( .A1(n13680), .A2(n15176), .ZN(n14897) );
  AND2_X1 U17061 ( .A1(n14884), .A2(n14897), .ZN(n14871) );
  AND2_X1 U17062 ( .A1(n14870), .A2(n14871), .ZN(n14855) );
  AND4_X1 U17063 ( .A1(n14850), .A2(n14918), .A3(n14931), .A4(n14940), .ZN(
        n13686) );
  INV_X1 U17064 ( .A(n13681), .ZN(n13684) );
  NAND3_X1 U17065 ( .A1(n13682), .A2(n19180), .A3(P2_EBX_REG_21__SCAN_IN), 
        .ZN(n13683) );
  NAND2_X1 U17066 ( .A1(n13684), .A2(n13683), .ZN(n18814) );
  OR2_X1 U17067 ( .A1(n18814), .A2(n10733), .ZN(n13685) );
  NAND2_X1 U17068 ( .A1(n13685), .A2(n14860), .ZN(n14857) );
  NAND2_X1 U17069 ( .A1(n13728), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13687) );
  OR2_X1 U17070 ( .A1(n18814), .A2(n13687), .ZN(n14856) );
  OR2_X1 U17071 ( .A1(n13688), .A2(n14882), .ZN(n14885) );
  AND2_X1 U17072 ( .A1(n13728), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13689) );
  NAND2_X1 U17073 ( .A1(n18847), .A2(n13689), .ZN(n14896) );
  AND2_X1 U17074 ( .A1(n14885), .A2(n14896), .ZN(n14853) );
  AND4_X1 U17075 ( .A1(n13692), .A2(n13691), .A3(n13690), .A4(n14952), .ZN(
        n13693) );
  AND4_X1 U17076 ( .A1(n14856), .A2(n14853), .A3(n13693), .A4(n14869), .ZN(
        n13694) );
  NAND3_X1 U17077 ( .A1(n13695), .A2(n19180), .A3(P2_EBX_REG_22__SCAN_IN), 
        .ZN(n13696) );
  AND2_X1 U17078 ( .A1(n13700), .A2(n13696), .ZN(n15518) );
  NAND2_X1 U17079 ( .A1(n15518), .A2(n13728), .ZN(n13697) );
  INV_X1 U17080 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15099) );
  NAND2_X1 U17081 ( .A1(n13697), .A2(n15099), .ZN(n15122) );
  OR2_X1 U17082 ( .A1(n13697), .A2(n15099), .ZN(n15123) );
  INV_X1 U17083 ( .A(n13698), .ZN(n13699) );
  XNOR2_X1 U17084 ( .A(n13700), .B(n13699), .ZN(n16057) );
  NAND2_X1 U17085 ( .A1(n16057), .A2(n13728), .ZN(n13701) );
  XNOR2_X1 U17086 ( .A(n13701), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14844) );
  INV_X1 U17087 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15098) );
  OR2_X1 U17088 ( .A1(n13701), .A2(n15098), .ZN(n13702) );
  NAND2_X1 U17089 ( .A1(n19180), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n13703) );
  OAI21_X1 U17090 ( .B1(n13704), .B2(n13703), .A(n13712), .ZN(n13705) );
  OR2_X1 U17091 ( .A1(n13706), .A2(n13705), .ZN(n16046) );
  INV_X1 U17092 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14831) );
  NOR2_X1 U17093 ( .A1(n13707), .A2(n14831), .ZN(n14827) );
  NAND2_X1 U17094 ( .A1(n13707), .A2(n14831), .ZN(n14826) );
  AND2_X1 U17095 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n13708), .ZN(n13710) );
  AOI21_X1 U17096 ( .B1(n19180), .B2(n13710), .A(n13709), .ZN(n13711) );
  AND2_X1 U17097 ( .A1(n13712), .A2(n13711), .ZN(n16025) );
  NAND2_X1 U17098 ( .A1(n13713), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13719) );
  INV_X1 U17099 ( .A(n13713), .ZN(n13714) );
  INV_X1 U17100 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15059) );
  NAND2_X1 U17101 ( .A1(n13714), .A2(n15059), .ZN(n13715) );
  NAND2_X1 U17102 ( .A1(n13719), .A2(n13715), .ZN(n14807) );
  NOR2_X2 U17103 ( .A1(n13716), .A2(n14786), .ZN(n13721) );
  INV_X1 U17104 ( .A(n13717), .ZN(n13718) );
  NAND2_X1 U17105 ( .A1(n13718), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14814) );
  NAND2_X1 U17106 ( .A1(n14814), .A2(n13719), .ZN(n14785) );
  XOR2_X1 U17107 ( .A(n13723), .B(n13722), .Z(n16003) );
  NAND2_X1 U17108 ( .A1(n16003), .A2(n13728), .ZN(n14790) );
  AOI21_X1 U17109 ( .B1(n15992), .B2(n13728), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14774) );
  INV_X1 U17110 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15015) );
  OAI21_X1 U17111 ( .B1(n13727), .B2(n10733), .A(n15015), .ZN(n14763) );
  NAND2_X1 U17112 ( .A1(n13728), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13726) );
  INV_X1 U17113 ( .A(n13731), .ZN(n13734) );
  NOR2_X1 U17114 ( .A1(n13732), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13733) );
  MUX2_X1 U17115 ( .A(n13734), .B(n13733), .S(n10302), .Z(n15985) );
  NAND2_X1 U17116 ( .A1(n15985), .A2(n13728), .ZN(n13735) );
  XOR2_X1 U17117 ( .A(n13735), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(
        n13736) );
  XNOR2_X1 U17118 ( .A(n13737), .B(n13736), .ZN(n13770) );
  NOR2_X1 U17119 ( .A1(n14431), .A2(n13738), .ZN(n13745) );
  INV_X1 U17120 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19779) );
  AOI22_X1 U17121 ( .A1(n13739), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13740) );
  OAI21_X1 U17122 ( .B1(n13741), .B2(n19779), .A(n13740), .ZN(n13742) );
  AOI21_X1 U17123 ( .B1(n13743), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n13742), .ZN(n13744) );
  XNOR2_X1 U17124 ( .A(n13745), .B(n13744), .ZN(n16068) );
  NOR2_X1 U17125 ( .A1(n18974), .A2(n19779), .ZN(n13762) );
  AOI21_X1 U17126 ( .B1(n16142), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13762), .ZN(n13746) );
  OAI21_X1 U17127 ( .B1(n16150), .B2(n13747), .A(n13746), .ZN(n13751) );
  NOR2_X1 U17128 ( .A1(n13748), .A2(n11033), .ZN(n15177) );
  AND2_X1 U17129 ( .A1(n15177), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15145) );
  NAND2_X1 U17130 ( .A1(n15145), .A2(n13749), .ZN(n15130) );
  NAND2_X1 U17131 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15149) );
  OR2_X1 U17132 ( .A1(n15130), .A2(n15149), .ZN(n14838) );
  NOR2_X1 U17133 ( .A1(n14838), .A2(n14860), .ZN(n15096) );
  AND2_X1 U17134 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13750) );
  AND2_X1 U17135 ( .A1(n15096), .A2(n13750), .ZN(n13754) );
  NAND2_X1 U17136 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15026) );
  OAI21_X1 U17137 ( .B1(n13770), .B2(n16152), .A(n13752), .ZN(P2_U2983) );
  INV_X1 U17138 ( .A(n13754), .ZN(n13753) );
  NOR2_X1 U17139 ( .A1(n13753), .A2(n15261), .ZN(n15084) );
  NAND2_X1 U17140 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15084), .ZN(
        n15078) );
  NAND2_X1 U17141 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13755) );
  NOR2_X1 U17142 ( .A1(n15078), .A2(n13755), .ZN(n13760) );
  NAND2_X1 U17143 ( .A1(n13760), .A2(n15048), .ZN(n15052) );
  OAI211_X1 U17144 ( .C1(n13754), .C2(n16209), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15257), .ZN(n15083) );
  OAI21_X1 U17145 ( .B1(n13755), .B2(n15083), .A(n15058), .ZN(n15049) );
  NAND2_X1 U17146 ( .A1(n15052), .A2(n15049), .ZN(n15044) );
  AOI21_X1 U17147 ( .B1(n15026), .B2(n19164), .A(n15044), .ZN(n15016) );
  OAI21_X1 U17148 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16209), .A(
        n15016), .ZN(n13768) );
  INV_X1 U17149 ( .A(n16068), .ZN(n13764) );
  AOI222_X1 U17150 ( .A1(n11999), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n13756), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n10823), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13757) );
  NAND2_X1 U17151 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n13760), .ZN(
        n15037) );
  NOR4_X1 U17152 ( .A1(n15026), .A2(n15015), .A3(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A4(n15037), .ZN(n13761) );
  AOI211_X1 U17153 ( .C1(n19086), .C2(n19152), .A(n13762), .B(n13761), .ZN(
        n13763) );
  OAI21_X1 U17154 ( .B1(n13764), .B2(n19157), .A(n13763), .ZN(n13767) );
  NOR2_X1 U17155 ( .A1(n13765), .A2(n16189), .ZN(n13766) );
  OAI21_X1 U17156 ( .B1(n13770), .B2(n19155), .A(n13769), .ZN(P2_U3015) );
  INV_X1 U17157 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n13816) );
  AOI22_X1 U17158 ( .A1(n13772), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13771), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13780) );
  AOI22_X1 U17159 ( .A1(n13773), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11693), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13779) );
  AOI22_X1 U17160 ( .A1(n13775), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13774), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13778) );
  AOI22_X1 U17161 ( .A1(n9603), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13776), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13777) );
  NAND4_X1 U17162 ( .A1(n13780), .A2(n13779), .A3(n13778), .A4(n13777), .ZN(
        n13791) );
  AOI22_X1 U17163 ( .A1(n13782), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13781), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13789) );
  AOI22_X1 U17164 ( .A1(n11708), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9605), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U17165 ( .A1(n13784), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11694), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13787) );
  AOI22_X1 U17166 ( .A1(n13785), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13786) );
  NAND4_X1 U17167 ( .A1(n13789), .A2(n13788), .A3(n13787), .A4(n13786), .ZN(
        n13790) );
  NOR2_X1 U17168 ( .A1(n13791), .A2(n13790), .ZN(n13795) );
  NOR2_X1 U17169 ( .A1(n13793), .A2(n13792), .ZN(n13794) );
  XOR2_X1 U17170 ( .A(n13795), .B(n13794), .Z(n13802) );
  NAND2_X1 U17171 ( .A1(n11268), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13796) );
  NAND2_X1 U17172 ( .A1(n13797), .A2(n13796), .ZN(n13798) );
  AOI21_X1 U17173 ( .B1(n13799), .B2(P1_EAX_REG_30__SCAN_IN), .A(n13798), .ZN(
        n13800) );
  OAI21_X1 U17174 ( .B1(n13802), .B2(n13801), .A(n13800), .ZN(n13806) );
  XNOR2_X1 U17175 ( .A(n13803), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14168) );
  NAND2_X1 U17176 ( .A1(n14168), .A2(n13804), .ZN(n13805) );
  AOI22_X1 U17177 ( .A1(n13799), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13808), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13809) );
  INV_X1 U17178 ( .A(n13817), .ZN(n13812) );
  AND2_X1 U17179 ( .A1(n19972), .A2(n13810), .ZN(n13811) );
  NAND2_X1 U17180 ( .A1(n13812), .A2(n13811), .ZN(n13815) );
  AOI22_X1 U17181 ( .A1(n15752), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15760), .ZN(n13814) );
  OAI211_X1 U17182 ( .C1(n15756), .C2(n13816), .A(n13815), .B(n13814), .ZN(
        P1_U2873) );
  AND2_X1 U17183 ( .A1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15568) );
  INV_X1 U17184 ( .A(n13818), .ZN(n13819) );
  NOR2_X1 U17185 ( .A1(n15819), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14162) );
  INV_X1 U17186 ( .A(n14162), .ZN(n13820) );
  OAI21_X1 U17187 ( .B1(n14163), .B2(n15568), .A(n13821), .ZN(n13822) );
  XNOR2_X1 U17188 ( .A(n13822), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15563) );
  NAND2_X1 U17189 ( .A1(n15563), .A2(n20071), .ZN(n13826) );
  INV_X1 U17190 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13834) );
  INV_X1 U17191 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n13831) );
  OAI22_X1 U17192 ( .A1(n15800), .A2(n13834), .B1(n20114), .B2(n13831), .ZN(
        n13823) );
  AOI21_X1 U17193 ( .B1(n20079), .B2(n13824), .A(n13823), .ZN(n13825) );
  OAI211_X1 U17194 ( .C1(n13817), .C2(n20149), .A(n13826), .B(n13825), .ZN(
        P1_U2968) );
  INV_X1 U17195 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20809) );
  INV_X1 U17196 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20804) );
  INV_X1 U17197 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20802) );
  INV_X1 U17198 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20799) );
  INV_X1 U17199 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20792) );
  INV_X1 U17200 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15729) );
  NOR3_X1 U17201 ( .A1(n20792), .A2(n13827), .A3(n15729), .ZN(n13973) );
  NAND3_X1 U17202 ( .A1(n13973), .A2(P1_REIP_REG_14__SCAN_IN), .A3(
        P1_REIP_REG_13__SCAN_IN), .ZN(n13954) );
  NAND2_X1 U17203 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15683) );
  NOR3_X1 U17204 ( .A1(n20799), .A2(n13954), .A3(n15683), .ZN(n13941) );
  NAND2_X1 U17205 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n13941), .ZN(n13946) );
  NOR2_X1 U17206 ( .A1(n20802), .A2(n13946), .ZN(n15666) );
  NAND2_X1 U17207 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n15666), .ZN(n15656) );
  NOR2_X1 U17208 ( .A1(n20804), .A2(n15656), .ZN(n15650) );
  NAND2_X1 U17209 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15650), .ZN(n13928) );
  NOR2_X1 U17210 ( .A1(n14192), .A2(n13928), .ZN(n15640) );
  NAND2_X1 U17211 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15640), .ZN(n13919) );
  NOR2_X1 U17212 ( .A1(n20809), .A2(n13919), .ZN(n13830) );
  NAND3_X1 U17213 ( .A1(n13830), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n19931), 
        .ZN(n15634) );
  NAND2_X1 U17214 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n13828) );
  OAI21_X1 U17215 ( .B1(n15634), .B2(n13828), .A(n15681), .ZN(n15627) );
  INV_X1 U17216 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20815) );
  INV_X1 U17217 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20817) );
  OAI21_X1 U17218 ( .B1(n20815), .B2(n20817), .A(n15681), .ZN(n13829) );
  NAND2_X1 U17219 ( .A1(n15627), .A2(n13829), .ZN(n13897) );
  NAND2_X1 U17220 ( .A1(n19937), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13833) );
  INV_X1 U17221 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n15626) );
  INV_X1 U17222 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15633) );
  NAND2_X1 U17223 ( .A1(n19925), .A2(n13830), .ZN(n15632) );
  NOR2_X1 U17224 ( .A1(n15633), .A2(n15632), .ZN(n13911) );
  NAND2_X1 U17225 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n13911), .ZN(n15625) );
  NOR3_X1 U17226 ( .A1(n15626), .A2(n20815), .A3(n15625), .ZN(n13898) );
  NAND3_X1 U17227 ( .A1(n13898), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n13831), 
        .ZN(n13832) );
  OAI211_X1 U17228 ( .C1(n13834), .C2(n19913), .A(n13833), .B(n13832), .ZN(
        n13835) );
  AOI21_X1 U17229 ( .B1(n13897), .B2(P1_REIP_REG_31__SCAN_IN), .A(n13835), 
        .ZN(n13884) );
  AOI22_X1 U17230 ( .A1(n13879), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n9777), .ZN(n13882) );
  INV_X1 U17231 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14086) );
  NAND2_X1 U17232 ( .A1(n13868), .A2(n14086), .ZN(n13839) );
  NAND2_X1 U17233 ( .A1(n13415), .A2(n15896), .ZN(n13837) );
  NAND2_X1 U17234 ( .A1(n13874), .A2(n14086), .ZN(n13836) );
  NAND3_X1 U17235 ( .A1(n13837), .A2(n13894), .A3(n13836), .ZN(n13838) );
  NAND2_X1 U17236 ( .A1(n13839), .A2(n13838), .ZN(n14082) );
  MUX2_X1 U17237 ( .A(n13867), .B(n13894), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n13840) );
  OAI21_X1 U17238 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n13879), .A(
        n13840), .ZN(n13841) );
  INV_X1 U17239 ( .A(n13841), .ZN(n13955) );
  INV_X1 U17240 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15673) );
  NAND2_X1 U17241 ( .A1(n13868), .A2(n15673), .ZN(n13845) );
  NAND2_X1 U17242 ( .A1(n13415), .A2(n15894), .ZN(n13843) );
  NAND2_X1 U17243 ( .A1(n13874), .A2(n15673), .ZN(n13842) );
  NAND3_X1 U17244 ( .A1(n13843), .A2(n13894), .A3(n13842), .ZN(n13844) );
  NAND2_X1 U17245 ( .A1(n13894), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13846) );
  OAI211_X1 U17246 ( .C1(n9777), .C2(P1_EBX_REG_19__SCAN_IN), .A(n13415), .B(
        n13846), .ZN(n13847) );
  OAI21_X1 U17247 ( .B1(n13867), .B2(P1_EBX_REG_19__SCAN_IN), .A(n13847), .ZN(
        n13942) );
  MUX2_X1 U17248 ( .A(n13877), .B(n13415), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n13850) );
  NAND2_X1 U17249 ( .A1(n9777), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13848) );
  AND2_X1 U17250 ( .A1(n13857), .A2(n13848), .ZN(n13849) );
  NAND2_X1 U17251 ( .A1(n13850), .A2(n13849), .ZN(n14062) );
  MUX2_X1 U17252 ( .A(n13867), .B(n13894), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n13851) );
  OAI21_X1 U17253 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13879), .A(
        n13851), .ZN(n13852) );
  INV_X1 U17254 ( .A(n13852), .ZN(n14056) );
  MUX2_X1 U17255 ( .A(n13877), .B(n13415), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n13854) );
  NAND2_X1 U17256 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n9777), .ZN(
        n13853) );
  AND3_X1 U17257 ( .A1(n13854), .A2(n13857), .A3(n13853), .ZN(n14049) );
  MUX2_X1 U17258 ( .A(n13867), .B(n13894), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13855) );
  OAI21_X1 U17259 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n13879), .A(
        n13855), .ZN(n13929) );
  MUX2_X1 U17260 ( .A(n13877), .B(n13415), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n13858) );
  NAND2_X1 U17261 ( .A1(n9777), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13856) );
  AND3_X1 U17262 ( .A1(n13858), .A2(n13857), .A3(n13856), .ZN(n14039) );
  INV_X1 U17263 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14036) );
  NAND2_X1 U17264 ( .A1(n13859), .A2(n14036), .ZN(n13862) );
  NAND2_X1 U17265 ( .A1(n13874), .A2(n14036), .ZN(n13860) );
  OAI211_X1 U17266 ( .C1(n11170), .C2(n15853), .A(n13860), .B(n13415), .ZN(
        n13861) );
  AND2_X1 U17267 ( .A1(n13862), .A2(n13861), .ZN(n13917) );
  NAND2_X1 U17268 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n9777), .ZN(
        n13864) );
  MUX2_X1 U17269 ( .A(n13877), .B(n13415), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n13863) );
  AND2_X1 U17270 ( .A1(n13864), .A2(n13863), .ZN(n14028) );
  INV_X1 U17271 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n13908) );
  NAND2_X1 U17272 ( .A1(n13874), .A2(n13908), .ZN(n13865) );
  OAI211_X1 U17273 ( .C1(n11170), .C2(n14289), .A(n13865), .B(n13415), .ZN(
        n13866) );
  OAI21_X1 U17274 ( .B1(n13867), .B2(P1_EBX_REG_27__SCAN_IN), .A(n13866), .ZN(
        n13912) );
  INV_X1 U17275 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n13869) );
  NAND2_X1 U17276 ( .A1(n13868), .A2(n13869), .ZN(n13873) );
  NAND2_X1 U17277 ( .A1(n13415), .A2(n14290), .ZN(n13871) );
  NAND2_X1 U17278 ( .A1(n13874), .A2(n13869), .ZN(n13870) );
  NAND3_X1 U17279 ( .A1(n13871), .A2(n13894), .A3(n13870), .ZN(n13872) );
  NAND2_X1 U17280 ( .A1(n13873), .A2(n13872), .ZN(n14020) );
  OR2_X1 U17281 ( .A1(n13879), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13876) );
  INV_X1 U17282 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14019) );
  NAND2_X1 U17283 ( .A1(n13874), .A2(n14019), .ZN(n13875) );
  NAND2_X1 U17284 ( .A1(n13876), .A2(n13875), .ZN(n13892) );
  OAI22_X1 U17285 ( .A1(n13892), .A2(n11170), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n13877), .ZN(n14017) );
  AND2_X1 U17286 ( .A1(n9777), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13878) );
  AOI21_X1 U17287 ( .B1(n13879), .B2(P1_EBX_REG_30__SCAN_IN), .A(n13878), .ZN(
        n13895) );
  NAND2_X1 U17288 ( .A1(n15562), .A2(n19926), .ZN(n13883) );
  OAI211_X1 U17289 ( .C1(n13817), .C2(n19920), .A(n13884), .B(n13883), .ZN(
        P1_U2809) );
  INV_X1 U17290 ( .A(n13885), .ZN(n13889) );
  INV_X1 U17291 ( .A(n13886), .ZN(n13887) );
  OAI21_X1 U17292 ( .B1(n13889), .B2(n13888), .A(n13887), .ZN(n13890) );
  INV_X1 U17293 ( .A(n14023), .ZN(n13893) );
  OAI22_X1 U17294 ( .A1(n14015), .A2(n13894), .B1(n13893), .B2(n13892), .ZN(
        n13896) );
  XNOR2_X1 U17295 ( .A(n13896), .B(n13895), .ZN(n14276) );
  INV_X1 U17296 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n13901) );
  OAI21_X1 U17297 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n13898), .A(n13897), 
        .ZN(n13900) );
  AOI22_X1 U17298 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19955), .B1(
        n19961), .B2(n14168), .ZN(n13899) );
  OAI211_X1 U17299 ( .C1(n19950), .C2(n13901), .A(n13900), .B(n13899), .ZN(
        n13902) );
  AOI21_X1 U17300 ( .B1(n14276), .B2(n19926), .A(n13902), .ZN(n13903) );
  OAI21_X1 U17301 ( .B1(n14171), .B2(n19920), .A(n13903), .ZN(P1_U2810) );
  AOI21_X1 U17302 ( .B1(n13904), .B2(n9660), .A(n11772), .ZN(n13905) );
  INV_X1 U17303 ( .A(n13905), .ZN(n14179) );
  INV_X1 U17304 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n13910) );
  NAND3_X1 U17305 ( .A1(n15634), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n15681), 
        .ZN(n13907) );
  AOI22_X1 U17306 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19955), .B1(
        n19961), .B2(n14176), .ZN(n13906) );
  OAI211_X1 U17307 ( .C1(n13908), .C2(n19950), .A(n13907), .B(n13906), .ZN(
        n13909) );
  AOI21_X1 U17308 ( .B1(n13911), .B2(n13910), .A(n13909), .ZN(n13914) );
  AOI21_X1 U17309 ( .B1(n13912), .B2(n9662), .A(n14021), .ZN(n15844) );
  NAND2_X1 U17310 ( .A1(n15844), .A2(n19926), .ZN(n13913) );
  OAI211_X1 U17311 ( .C1(n14179), .C2(n19920), .A(n13914), .B(n13913), .ZN(
        P1_U2813) );
  OAI21_X1 U17312 ( .B1(n13915), .B2(n13916), .A(n14032), .ZN(n14189) );
  OR2_X1 U17313 ( .A1(n14042), .A2(n13917), .ZN(n13918) );
  AND2_X1 U17314 ( .A1(n13918), .A2(n14029), .ZN(n15848) );
  NOR3_X1 U17315 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n19958), .A3(n13919), 
        .ZN(n13925) );
  INV_X1 U17316 ( .A(n14186), .ZN(n13921) );
  NOR2_X1 U17317 ( .A1(n19958), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15641) );
  OAI21_X1 U17318 ( .B1(n15640), .B2(n19958), .A(n19931), .ZN(n15646) );
  OAI21_X1 U17319 ( .B1(n15641), .B2(n15646), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n13920) );
  OAI21_X1 U17320 ( .B1(n19948), .B2(n13921), .A(n13920), .ZN(n13922) );
  AOI21_X1 U17321 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19955), .A(
        n13922), .ZN(n13923) );
  OAI21_X1 U17322 ( .B1(n14036), .B2(n19950), .A(n13923), .ZN(n13924) );
  AOI211_X1 U17323 ( .C1(n15848), .C2(n19926), .A(n13925), .B(n13924), .ZN(
        n13926) );
  OAI21_X1 U17324 ( .B1(n14189), .B2(n19920), .A(n13926), .ZN(P1_U2815) );
  OAI21_X1 U17325 ( .B1(n13927), .B2(n9661), .A(n9625), .ZN(n14198) );
  OAI21_X1 U17326 ( .B1(n19958), .B2(n13928), .A(n14192), .ZN(n13934) );
  INV_X1 U17327 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14046) );
  NAND2_X1 U17328 ( .A1(n14051), .A2(n13929), .ZN(n13930) );
  NAND2_X1 U17329 ( .A1(n14040), .A2(n13930), .ZN(n14045) );
  INV_X1 U17330 ( .A(n14045), .ZN(n15857) );
  NAND2_X1 U17331 ( .A1(n15857), .A2(n19926), .ZN(n13932) );
  AOI22_X1 U17332 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19955), .B1(
        n19961), .B2(n14195), .ZN(n13931) );
  OAI211_X1 U17333 ( .C1(n14046), .C2(n19950), .A(n13932), .B(n13931), .ZN(
        n13933) );
  AOI21_X1 U17334 ( .B1(n13934), .B2(n15646), .A(n13933), .ZN(n13935) );
  OAI21_X1 U17335 ( .B1(n14198), .B2(n19920), .A(n13935), .ZN(P1_U2817) );
  INV_X1 U17336 ( .A(n13937), .ZN(n13938) );
  OAI21_X1 U17337 ( .B1(n13939), .B2(n13936), .A(n13938), .ZN(n14207) );
  INV_X1 U17338 ( .A(n14207), .ZN(n14137) );
  NAND2_X1 U17339 ( .A1(n14137), .A2(n19905), .ZN(n13950) );
  INV_X1 U17340 ( .A(n13941), .ZN(n13940) );
  NOR3_X1 U17341 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n19958), .A3(n13940), 
        .ZN(n15677) );
  OAI21_X1 U17342 ( .B1(n13941), .B2(n19958), .A(n19931), .ZN(n15678) );
  OAI21_X1 U17343 ( .B1(n15677), .B2(n15678), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n13949) );
  AND2_X1 U17344 ( .A1(n9657), .A2(n13942), .ZN(n13943) );
  NOR2_X1 U17345 ( .A1(n14063), .A2(n13943), .ZN(n15880) );
  AOI22_X1 U17346 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(n19937), .B1(n19961), 
        .B2(n14204), .ZN(n13944) );
  OAI211_X1 U17347 ( .C1(n19913), .C2(n14202), .A(n13944), .B(n19910), .ZN(
        n13945) );
  AOI21_X1 U17348 ( .B1(n15880), .B2(n19926), .A(n13945), .ZN(n13948) );
  OR3_X1 U17349 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n19958), .A3(n13946), .ZN(
        n13947) );
  NAND4_X1 U17350 ( .A1(n13950), .A2(n13949), .A3(n13948), .A4(n13947), .ZN(
        P1_U2821) );
  NAND2_X1 U17351 ( .A1(n14081), .A2(n13952), .ZN(n13953) );
  NAND2_X1 U17352 ( .A1(n14070), .A2(n13953), .ZN(n14220) );
  OR2_X1 U17353 ( .A1(n19958), .A2(n13954), .ZN(n15702) );
  OAI21_X1 U17354 ( .B1(n15683), .B2(n15702), .A(n20799), .ZN(n13961) );
  OR2_X1 U17355 ( .A1(n14085), .A2(n13955), .ZN(n13956) );
  AND2_X1 U17356 ( .A1(n9692), .A2(n13956), .ZN(n15899) );
  INV_X1 U17357 ( .A(n15899), .ZN(n14076) );
  OAI21_X1 U17358 ( .B1(n19948), .B2(n14215), .A(n19910), .ZN(n13958) );
  INV_X1 U17359 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14077) );
  NOR2_X1 U17360 ( .A1(n19950), .A2(n14077), .ZN(n13957) );
  AOI211_X1 U17361 ( .C1(n19955), .C2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n13958), .B(n13957), .ZN(n13959) );
  OAI21_X1 U17362 ( .B1(n14076), .B2(n19952), .A(n13959), .ZN(n13960) );
  AOI21_X1 U17363 ( .B1(n13961), .B2(n15678), .A(n13960), .ZN(n13962) );
  OAI21_X1 U17364 ( .B1(n14220), .B2(n19920), .A(n13962), .ZN(P1_U2823) );
  NAND2_X1 U17365 ( .A1(n13964), .A2(n13963), .ZN(n13965) );
  NAND2_X1 U17366 ( .A1(n9694), .A2(n13965), .ZN(n15727) );
  OR2_X1 U17367 ( .A1(n15727), .A2(n15725), .ZN(n13966) );
  NAND2_X1 U17368 ( .A1(n13966), .A2(n9694), .ZN(n14093) );
  INV_X1 U17369 ( .A(n13967), .ZN(n13968) );
  NOR2_X1 U17370 ( .A1(n20792), .A2(n15729), .ZN(n13972) );
  AOI21_X1 U17371 ( .B1(n13972), .B2(n13971), .A(n13970), .ZN(n15722) );
  NAND2_X1 U17372 ( .A1(n19925), .A2(n13973), .ZN(n15706) );
  INV_X1 U17373 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14090) );
  OAI22_X1 U17374 ( .A1(n15706), .A2(P1_REIP_REG_13__SCAN_IN), .B1(n14090), 
        .B2(n19950), .ZN(n13979) );
  OR2_X1 U17375 ( .A1(n14096), .A2(n13974), .ZN(n13976) );
  AND2_X1 U17376 ( .A1(n13976), .A2(n13975), .ZN(n15914) );
  AOI22_X1 U17377 ( .A1(n14244), .A2(n19961), .B1(n19926), .B2(n15914), .ZN(
        n13977) );
  OAI211_X1 U17378 ( .C1(n19913), .C2(n14242), .A(n13977), .B(n19910), .ZN(
        n13978) );
  AOI211_X1 U17379 ( .C1(n15722), .C2(P1_REIP_REG_13__SCAN_IN), .A(n13979), 
        .B(n13978), .ZN(n13980) );
  OAI21_X1 U17380 ( .B1(n14246), .B2(n19920), .A(n13980), .ZN(P1_U2827) );
  NOR2_X1 U17381 ( .A1(n19952), .A2(n15950), .ZN(n13981) );
  AOI211_X1 U17382 ( .C1(n19954), .C2(P1_REIP_REG_8__SCAN_IN), .A(n13981), .B(
        n19941), .ZN(n13983) );
  NAND2_X1 U17383 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13982) );
  OAI211_X1 U17384 ( .C1(n14258), .C2(n19948), .A(n13983), .B(n13982), .ZN(
        n13986) );
  AOI211_X1 U17385 ( .C1(n20787), .C2(n13984), .A(n19893), .B(n19958), .ZN(
        n13985) );
  AOI211_X1 U17386 ( .C1(n19937), .C2(P1_EBX_REG_8__SCAN_IN), .A(n13986), .B(
        n13985), .ZN(n13987) );
  OAI21_X1 U17387 ( .B1(n13988), .B2(n19920), .A(n13987), .ZN(P1_U2832) );
  NAND2_X1 U17388 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13995) );
  NAND2_X1 U17389 ( .A1(n19925), .A2(n13995), .ZN(n14006) );
  NAND2_X1 U17390 ( .A1(n14006), .A2(n19931), .ZN(n14009) );
  OAI22_X1 U17391 ( .A1(n13990), .A2(n19948), .B1(n19913), .B2(n13989), .ZN(
        n13993) );
  NOR2_X1 U17392 ( .A1(n19950), .A2(n13991), .ZN(n13992) );
  AOI211_X1 U17393 ( .C1(n20102), .C2(n19926), .A(n13993), .B(n13992), .ZN(
        n13994) );
  OAI21_X1 U17394 ( .B1(n14401), .B2(n14005), .A(n13994), .ZN(n13997) );
  NOR3_X1 U17395 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n19958), .A3(n13995), .ZN(
        n13996) );
  AOI211_X1 U17396 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(n14009), .A(n13997), .B(
        n13996), .ZN(n13998) );
  OAI21_X1 U17397 ( .B1(n19963), .B2(n13999), .A(n13998), .ZN(P1_U2837) );
  OAI22_X1 U17398 ( .A1(n14001), .A2(n19913), .B1(n19948), .B2(n14000), .ZN(
        n14003) );
  NOR2_X1 U17399 ( .A1(n19952), .A2(n20115), .ZN(n14002) );
  AOI211_X1 U17400 ( .C1(n19937), .C2(P1_EBX_REG_2__SCAN_IN), .A(n14003), .B(
        n14002), .ZN(n14004) );
  OAI21_X1 U17401 ( .B1(n12991), .B2(n14005), .A(n14004), .ZN(n14008) );
  INV_X1 U17402 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20838) );
  NOR2_X1 U17403 ( .A1(n14006), .A2(n20838), .ZN(n14007) );
  AOI211_X1 U17404 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(n14009), .A(n14008), .B(
        n14007), .ZN(n14010) );
  OAI21_X1 U17405 ( .B1(n19963), .B2(n14011), .A(n14010), .ZN(P1_U2838) );
  INV_X1 U17406 ( .A(n15562), .ZN(n14013) );
  INV_X1 U17407 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14012) );
  OAI22_X1 U17408 ( .A1(n14013), .A2(n14098), .B1(n19970), .B2(n14012), .ZN(
        P1_U2841) );
  AOI22_X1 U17409 ( .A1(n14276), .A2(n19965), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n14068), .ZN(n14014) );
  OAI21_X1 U17410 ( .B1(n14171), .B2(n14078), .A(n14014), .ZN(P1_U2842) );
  INV_X1 U17411 ( .A(n14015), .ZN(n14016) );
  OAI21_X1 U17412 ( .B1(n14023), .B2(n14017), .A(n14016), .ZN(n15616) );
  INV_X1 U17413 ( .A(n15744), .ZN(n14018) );
  OAI222_X1 U17414 ( .A1(n14098), .A2(n15616), .B1(n14019), .B2(n19970), .C1(
        n14018), .C2(n14078), .ZN(P1_U2843) );
  NOR2_X1 U17415 ( .A1(n14021), .A2(n14020), .ZN(n14022) );
  OR2_X1 U17416 ( .A1(n14023), .A2(n14022), .ZN(n15621) );
  INV_X1 U17417 ( .A(n15621), .ZN(n14024) );
  AOI22_X1 U17418 ( .A1(n14024), .A2(n19965), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14068), .ZN(n14025) );
  OAI21_X1 U17419 ( .B1(n14026), .B2(n14078), .A(n14025), .ZN(P1_U2844) );
  AOI22_X1 U17420 ( .A1(n15844), .A2(n19965), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14068), .ZN(n14027) );
  OAI21_X1 U17421 ( .B1(n14179), .B2(n14078), .A(n14027), .ZN(P1_U2845) );
  NAND2_X1 U17422 ( .A1(n14029), .A2(n14028), .ZN(n14030) );
  NAND2_X1 U17423 ( .A1(n9662), .A2(n14030), .ZN(n15639) );
  INV_X1 U17424 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14035) );
  NAND2_X1 U17425 ( .A1(n14032), .A2(n14031), .ZN(n14033) );
  INV_X1 U17426 ( .A(n15763), .ZN(n14034) );
  OAI222_X1 U17427 ( .A1(n14098), .A2(n15639), .B1(n14035), .B2(n19970), .C1(
        n14034), .C2(n14078), .ZN(P1_U2846) );
  NOR2_X1 U17428 ( .A1(n19970), .A2(n14036), .ZN(n14037) );
  AOI21_X1 U17429 ( .B1(n15848), .B2(n19965), .A(n14037), .ZN(n14038) );
  OAI21_X1 U17430 ( .B1(n14189), .B2(n14078), .A(n14038), .ZN(P1_U2847) );
  AND2_X1 U17431 ( .A1(n14040), .A2(n14039), .ZN(n14041) );
  NOR2_X1 U17432 ( .A1(n14042), .A2(n14041), .ZN(n14315) );
  INV_X1 U17433 ( .A(n14315), .ZN(n15642) );
  INV_X1 U17434 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14044) );
  AOI21_X1 U17435 ( .B1(n10073), .B2(n9625), .A(n13915), .ZN(n15768) );
  INV_X1 U17436 ( .A(n15768), .ZN(n15643) );
  OAI222_X1 U17437 ( .A1(n14098), .A2(n15642), .B1(n14091), .B2(n14044), .C1(
        n15643), .C2(n14078), .ZN(P1_U2848) );
  OAI222_X1 U17438 ( .A1(n14078), .A2(n14198), .B1(n14091), .B2(n14046), .C1(
        n14045), .C2(n14098), .ZN(P1_U2849) );
  OR2_X1 U17439 ( .A1(n14047), .A2(n14055), .ZN(n14053) );
  AOI21_X1 U17440 ( .B1(n14048), .B2(n14053), .A(n9661), .ZN(n15776) );
  INV_X1 U17441 ( .A(n15776), .ZN(n14052) );
  INV_X1 U17442 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15654) );
  NAND2_X1 U17443 ( .A1(n14058), .A2(n14049), .ZN(n14050) );
  NAND2_X1 U17444 ( .A1(n14051), .A2(n14050), .ZN(n15869) );
  OAI222_X1 U17445 ( .A1(n14078), .A2(n14052), .B1(n15654), .B2(n19970), .C1(
        n15869), .C2(n14098), .ZN(P1_U2850) );
  INV_X1 U17446 ( .A(n14053), .ZN(n14054) );
  AOI21_X1 U17447 ( .B1(n14055), .B2(n14047), .A(n14054), .ZN(n15781) );
  INV_X1 U17448 ( .A(n15781), .ZN(n14136) );
  OR2_X1 U17449 ( .A1(n14065), .A2(n14056), .ZN(n14057) );
  AND2_X1 U17450 ( .A1(n14058), .A2(n14057), .ZN(n15660) );
  AOI22_X1 U17451 ( .A1(n15660), .A2(n19965), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14068), .ZN(n14059) );
  OAI21_X1 U17452 ( .B1(n14136), .B2(n14078), .A(n14059), .ZN(P1_U2851) );
  OR2_X1 U17453 ( .A1(n13937), .A2(n14060), .ZN(n14061) );
  INV_X1 U17454 ( .A(n15787), .ZN(n14067) );
  INV_X1 U17455 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14066) );
  NOR2_X1 U17456 ( .A1(n14063), .A2(n14062), .ZN(n14064) );
  OR2_X1 U17457 ( .A1(n14065), .A2(n14064), .ZN(n15667) );
  OAI222_X1 U17458 ( .A1(n14078), .A2(n14067), .B1(n14066), .B2(n19970), .C1(
        n15667), .C2(n14098), .ZN(P1_U2852) );
  AOI22_X1 U17459 ( .A1(n15880), .A2(n19965), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14068), .ZN(n14069) );
  OAI21_X1 U17460 ( .B1(n14207), .B2(n14078), .A(n14069), .ZN(P1_U2853) );
  AOI21_X1 U17461 ( .B1(n14071), .B2(n14070), .A(n13936), .ZN(n15796) );
  INV_X1 U17462 ( .A(n15796), .ZN(n15674) );
  NAND2_X1 U17463 ( .A1(n9692), .A2(n14072), .ZN(n14073) );
  NAND2_X1 U17464 ( .A1(n9657), .A2(n14073), .ZN(n15888) );
  OAI22_X1 U17465 ( .A1(n15888), .A2(n14098), .B1(n15673), .B2(n19970), .ZN(
        n14074) );
  INV_X1 U17466 ( .A(n14074), .ZN(n14075) );
  OAI21_X1 U17467 ( .B1(n15674), .B2(n14078), .A(n14075), .ZN(P1_U2854) );
  OAI222_X1 U17468 ( .A1(n14078), .A2(n14220), .B1(n14091), .B2(n14077), .C1(
        n14076), .C2(n14098), .ZN(P1_U2855) );
  NAND2_X1 U17469 ( .A1(n9656), .A2(n14079), .ZN(n14080) );
  AND2_X1 U17470 ( .A1(n14081), .A2(n14080), .ZN(n15802) );
  NOR2_X1 U17471 ( .A1(n14083), .A2(n14082), .ZN(n14084) );
  OR2_X1 U17472 ( .A1(n14085), .A2(n14084), .ZN(n15690) );
  OAI22_X1 U17473 ( .A1(n15690), .A2(n14098), .B1(n14086), .B2(n19970), .ZN(
        n14087) );
  AOI21_X1 U17474 ( .B1(n15802), .B2(n19966), .A(n14087), .ZN(n14088) );
  INV_X1 U17475 ( .A(n14088), .ZN(P1_U2856) );
  INV_X1 U17476 ( .A(n15914), .ZN(n14089) );
  OAI222_X1 U17477 ( .A1(n14246), .A2(n14078), .B1(n14091), .B2(n14090), .C1(
        n14089), .C2(n14098), .ZN(P1_U2859) );
  NOR2_X1 U17478 ( .A1(n14093), .A2(n14092), .ZN(n14094) );
  NOR2_X1 U17479 ( .A1(n14095), .A2(n14094), .ZN(n15813) );
  INV_X1 U17480 ( .A(n15813), .ZN(n15758) );
  INV_X1 U17481 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15718) );
  AOI21_X1 U17482 ( .B1(n14097), .B2(n15733), .A(n14096), .ZN(n15720) );
  INV_X1 U17483 ( .A(n15720), .ZN(n14099) );
  OAI222_X1 U17484 ( .A1(n15758), .A2(n14078), .B1(n19970), .B2(n15718), .C1(
        n14099), .C2(n14098), .ZN(P1_U2860) );
  INV_X1 U17485 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n19187) );
  NOR2_X1 U17486 ( .A1(n15756), .A2(n19187), .ZN(n14103) );
  INV_X1 U17487 ( .A(n15751), .ZN(n14101) );
  INV_X1 U17488 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14100) );
  OAI22_X1 U17489 ( .A1(n14101), .A2(n20050), .B1(n19972), .B2(n14100), .ZN(
        n14102) );
  AOI211_X1 U17490 ( .C1(n15752), .C2(DATAI_30_), .A(n14103), .B(n14102), .ZN(
        n14104) );
  OAI21_X1 U17491 ( .B1(n14171), .B2(n19975), .A(n14104), .ZN(P1_U2874) );
  NAND2_X1 U17492 ( .A1(n15623), .A2(n15753), .ZN(n14110) );
  INV_X1 U17493 ( .A(DATAI_12_), .ZN(n14106) );
  NAND2_X1 U17494 ( .A1(n14158), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14105) );
  OAI21_X1 U17495 ( .B1(n14158), .B2(n14106), .A(n14105), .ZN(n20046) );
  AOI22_X1 U17496 ( .A1(n15751), .A2(n20046), .B1(n15760), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n14109) );
  NAND2_X1 U17497 ( .A1(n14151), .A2(BUF1_REG_28__SCAN_IN), .ZN(n14108) );
  NAND2_X1 U17498 ( .A1(n15752), .A2(DATAI_28_), .ZN(n14107) );
  NAND4_X1 U17499 ( .A1(n14110), .A2(n14109), .A3(n14108), .A4(n14107), .ZN(
        P1_U2876) );
  INV_X1 U17500 ( .A(DATAI_27_), .ZN(n14114) );
  INV_X1 U17501 ( .A(DATAI_11_), .ZN(n14112) );
  NAND2_X1 U17502 ( .A1(n14158), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14111) );
  OAI21_X1 U17503 ( .B1(n14158), .B2(n14112), .A(n14111), .ZN(n20044) );
  AOI22_X1 U17504 ( .A1(n15751), .A2(n20044), .B1(n15760), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n14113) );
  OAI21_X1 U17505 ( .B1(n14133), .B2(n14114), .A(n14113), .ZN(n14115) );
  AOI21_X1 U17506 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14151), .A(n14115), .ZN(
        n14116) );
  OAI21_X1 U17507 ( .B1(n14179), .B2(n19975), .A(n14116), .ZN(P1_U2877) );
  INV_X1 U17508 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16297) );
  NAND2_X1 U17509 ( .A1(n15752), .A2(DATAI_25_), .ZN(n14118) );
  AOI22_X1 U17510 ( .A1(n15751), .A2(n20040), .B1(n15760), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n14117) );
  OAI211_X1 U17511 ( .C1(n16297), .C2(n15756), .A(n14118), .B(n14117), .ZN(
        n14119) );
  INV_X1 U17512 ( .A(n14119), .ZN(n14120) );
  OAI21_X1 U17513 ( .B1(n14189), .B2(n19975), .A(n14120), .ZN(P1_U2879) );
  NAND2_X1 U17514 ( .A1(n15768), .A2(n15753), .ZN(n14125) );
  AOI22_X1 U17515 ( .A1(n15751), .A2(n14121), .B1(n15760), .B2(
        P1_EAX_REG_24__SCAN_IN), .ZN(n14124) );
  NAND2_X1 U17516 ( .A1(n14151), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14123) );
  NAND2_X1 U17517 ( .A1(n15752), .A2(DATAI_24_), .ZN(n14122) );
  NAND4_X1 U17518 ( .A1(n14125), .A2(n14124), .A3(n14123), .A4(n14122), .ZN(
        P1_U2880) );
  INV_X1 U17519 ( .A(n14198), .ZN(n14126) );
  NAND2_X1 U17520 ( .A1(n14126), .A2(n15753), .ZN(n14130) );
  AOI22_X1 U17521 ( .A1(n15751), .A2(n20198), .B1(n15760), .B2(
        P1_EAX_REG_23__SCAN_IN), .ZN(n14129) );
  NAND2_X1 U17522 ( .A1(n14151), .A2(BUF1_REG_23__SCAN_IN), .ZN(n14128) );
  NAND2_X1 U17523 ( .A1(n15752), .A2(DATAI_23_), .ZN(n14127) );
  NAND4_X1 U17524 ( .A1(n14130), .A2(n14129), .A3(n14128), .A4(n14127), .ZN(
        P1_U2881) );
  INV_X1 U17525 ( .A(DATAI_21_), .ZN(n14132) );
  AOI22_X1 U17526 ( .A1(n15751), .A2(n20184), .B1(n15760), .B2(
        P1_EAX_REG_21__SCAN_IN), .ZN(n14131) );
  OAI21_X1 U17527 ( .B1(n14133), .B2(n14132), .A(n14131), .ZN(n14134) );
  AOI21_X1 U17528 ( .B1(n14151), .B2(BUF1_REG_21__SCAN_IN), .A(n14134), .ZN(
        n14135) );
  OAI21_X1 U17529 ( .B1(n14136), .B2(n19975), .A(n14135), .ZN(P1_U2883) );
  NAND2_X1 U17530 ( .A1(n14137), .A2(n15753), .ZN(n14141) );
  AOI22_X1 U17531 ( .A1(n15751), .A2(n20172), .B1(n15760), .B2(
        P1_EAX_REG_19__SCAN_IN), .ZN(n14140) );
  NAND2_X1 U17532 ( .A1(n14151), .A2(BUF1_REG_19__SCAN_IN), .ZN(n14139) );
  NAND2_X1 U17533 ( .A1(n15752), .A2(DATAI_19_), .ZN(n14138) );
  NAND4_X1 U17534 ( .A1(n14141), .A2(n14140), .A3(n14139), .A4(n14138), .ZN(
        P1_U2885) );
  NAND2_X1 U17535 ( .A1(n15796), .A2(n15753), .ZN(n14145) );
  AOI22_X1 U17536 ( .A1(n15751), .A2(n20164), .B1(n15760), .B2(
        P1_EAX_REG_18__SCAN_IN), .ZN(n14144) );
  NAND2_X1 U17537 ( .A1(n14151), .A2(BUF1_REG_18__SCAN_IN), .ZN(n14143) );
  NAND2_X1 U17538 ( .A1(n15752), .A2(DATAI_18_), .ZN(n14142) );
  NAND4_X1 U17539 ( .A1(n14145), .A2(n14144), .A3(n14143), .A4(n14142), .ZN(
        P1_U2886) );
  INV_X1 U17540 ( .A(n14220), .ZN(n14146) );
  NAND2_X1 U17541 ( .A1(n14146), .A2(n15753), .ZN(n14150) );
  AOI22_X1 U17542 ( .A1(n15751), .A2(n20159), .B1(n15760), .B2(
        P1_EAX_REG_17__SCAN_IN), .ZN(n14149) );
  NAND2_X1 U17543 ( .A1(n14151), .A2(BUF1_REG_17__SCAN_IN), .ZN(n14148) );
  NAND2_X1 U17544 ( .A1(n15752), .A2(DATAI_17_), .ZN(n14147) );
  NAND4_X1 U17545 ( .A1(n14150), .A2(n14149), .A3(n14148), .A4(n14147), .ZN(
        P1_U2887) );
  NAND2_X1 U17546 ( .A1(n15802), .A2(n15753), .ZN(n14155) );
  AOI22_X1 U17547 ( .A1(n15751), .A2(n20150), .B1(n15760), .B2(
        P1_EAX_REG_16__SCAN_IN), .ZN(n14154) );
  NAND2_X1 U17548 ( .A1(n14151), .A2(BUF1_REG_16__SCAN_IN), .ZN(n14153) );
  NAND2_X1 U17549 ( .A1(n15752), .A2(DATAI_16_), .ZN(n14152) );
  NAND4_X1 U17550 ( .A1(n14155), .A2(n14154), .A3(n14153), .A4(n14152), .ZN(
        P1_U2888) );
  INV_X1 U17551 ( .A(DATAI_13_), .ZN(n14157) );
  NAND2_X1 U17552 ( .A1(n14158), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14156) );
  OAI21_X1 U17553 ( .B1(n14158), .B2(n14157), .A(n14156), .ZN(n20048) );
  INV_X1 U17554 ( .A(n20048), .ZN(n14160) );
  OAI222_X1 U17555 ( .A1(n19975), .A2(n14246), .B1(n19974), .B2(n14160), .C1(
        n14159), .C2(n19972), .ZN(P1_U2891) );
  NOR2_X1 U17556 ( .A1(n9618), .A2(n14285), .ZN(n14161) );
  INV_X1 U17557 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14164) );
  NAND2_X1 U17558 ( .A1(n14267), .A2(n20071), .ZN(n14170) );
  INV_X1 U17559 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14166) );
  NAND2_X1 U17560 ( .A1(n20128), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14278) );
  OAI21_X1 U17561 ( .B1(n15800), .B2(n14166), .A(n14278), .ZN(n14167) );
  AOI21_X1 U17562 ( .B1(n14168), .B2(n20079), .A(n14167), .ZN(n14169) );
  OAI211_X1 U17563 ( .C1(n20149), .C2(n14171), .A(n14170), .B(n14169), .ZN(
        P1_U2969) );
  NAND2_X1 U17564 ( .A1(n15845), .A2(n20071), .ZN(n14178) );
  OAI22_X1 U17565 ( .A1(n15800), .A2(n14174), .B1(n20114), .B2(n13910), .ZN(
        n14175) );
  AOI21_X1 U17566 ( .B1(n20079), .B2(n14176), .A(n14175), .ZN(n14177) );
  OAI211_X1 U17567 ( .C1(n20149), .C2(n14179), .A(n14178), .B(n14177), .ZN(
        P1_U2972) );
  NAND2_X1 U17568 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n14180), .ZN(
        n14310) );
  INV_X1 U17569 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15862) );
  NAND2_X1 U17570 ( .A1(n9618), .A2(n14191), .ZN(n14181) );
  OAI221_X1 U17571 ( .B1(n9618), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C1(
        n15819), .C2(n15862), .A(n14181), .ZN(n14182) );
  AOI21_X1 U17572 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14310), .A(
        n14182), .ZN(n14183) );
  XOR2_X1 U17573 ( .A(n14183), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n15849) );
  NAND2_X1 U17574 ( .A1(n15849), .A2(n20071), .ZN(n14188) );
  OAI22_X1 U17575 ( .A1(n15800), .A2(n14184), .B1(n20114), .B2(n20809), .ZN(
        n14185) );
  AOI21_X1 U17576 ( .B1(n20079), .B2(n14186), .A(n14185), .ZN(n14187) );
  OAI211_X1 U17577 ( .C1(n20149), .C2(n14189), .A(n14188), .B(n14187), .ZN(
        P1_U2974) );
  AOI22_X1 U17578 ( .A1(n9618), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n15862), .B2(n15819), .ZN(n14190) );
  XOR2_X1 U17579 ( .A(n14191), .B(n14190), .Z(n15858) );
  NAND2_X1 U17580 ( .A1(n15858), .A2(n20071), .ZN(n14197) );
  INV_X1 U17581 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14192) );
  OAI22_X1 U17582 ( .A1(n15800), .A2(n14193), .B1(n20114), .B2(n14192), .ZN(
        n14194) );
  AOI21_X1 U17583 ( .B1(n20079), .B2(n14195), .A(n14194), .ZN(n14196) );
  OAI211_X1 U17584 ( .C1(n20149), .C2(n14198), .A(n14197), .B(n14196), .ZN(
        P1_U2976) );
  INV_X1 U17585 ( .A(n14199), .ZN(n14320) );
  NOR2_X1 U17586 ( .A1(n14320), .A2(n15819), .ZN(n14200) );
  AOI22_X1 U17587 ( .A1(n15894), .A2(n14200), .B1(n14320), .B2(n15819), .ZN(
        n14201) );
  XOR2_X1 U17588 ( .A(n14201), .B(n15884), .Z(n15881) );
  NAND2_X1 U17589 ( .A1(n15881), .A2(n20071), .ZN(n14206) );
  OAI22_X1 U17590 ( .A1(n15800), .A2(n14202), .B1(n20114), .B2(n20802), .ZN(
        n14203) );
  AOI21_X1 U17591 ( .B1(n20079), .B2(n14204), .A(n14203), .ZN(n14205) );
  OAI211_X1 U17592 ( .C1(n20149), .C2(n14207), .A(n14206), .B(n14205), .ZN(
        P1_U2980) );
  INV_X1 U17593 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14214) );
  INV_X1 U17594 ( .A(n14208), .ZN(n14358) );
  OAI21_X1 U17595 ( .B1(n14358), .B2(n14210), .A(n14209), .ZN(n14212) );
  OAI21_X1 U17596 ( .B1(n15819), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n14212), .ZN(n14211) );
  OAI21_X1 U17597 ( .B1(n15819), .B2(n14212), .A(n14211), .ZN(n14213) );
  XOR2_X1 U17598 ( .A(n14214), .B(n14213), .Z(n15900) );
  INV_X1 U17599 ( .A(n14215), .ZN(n14218) );
  OAI22_X1 U17600 ( .A1(n15800), .A2(n14216), .B1(n20114), .B2(n20799), .ZN(
        n14217) );
  AOI21_X1 U17601 ( .B1(n20079), .B2(n14218), .A(n14217), .ZN(n14219) );
  OAI21_X1 U17602 ( .B1(n14220), .B2(n20149), .A(n14219), .ZN(n14221) );
  AOI21_X1 U17603 ( .B1(n15900), .B2(n20071), .A(n14221), .ZN(n14222) );
  INV_X1 U17604 ( .A(n14222), .ZN(P1_U2982) );
  AOI21_X1 U17605 ( .B1(n14208), .B2(n14224), .A(n14223), .ZN(n14335) );
  NOR2_X1 U17606 ( .A1(n14335), .A2(n14225), .ZN(n14227) );
  AOI21_X1 U17607 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n9618), .A(
        n14336), .ZN(n14226) );
  XNOR2_X1 U17608 ( .A(n14227), .B(n14226), .ZN(n15907) );
  NAND2_X1 U17609 ( .A1(n15907), .A2(n20071), .ZN(n14233) );
  INV_X1 U17610 ( .A(n14228), .ZN(n15695) );
  INV_X1 U17611 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n14229) );
  OAI22_X1 U17612 ( .A1(n15800), .A2(n14230), .B1(n20114), .B2(n14229), .ZN(
        n14231) );
  AOI21_X1 U17613 ( .B1(n15695), .B2(n20079), .A(n14231), .ZN(n14232) );
  OAI211_X1 U17614 ( .C1(n20149), .C2(n15694), .A(n14233), .B(n14232), .ZN(
        P1_U2984) );
  NAND2_X1 U17615 ( .A1(n14235), .A2(n14234), .ZN(n14369) );
  OAI21_X1 U17616 ( .B1(n14237), .B2(n14208), .A(n14236), .ZN(n14368) );
  NOR2_X1 U17617 ( .A1(n14369), .A2(n14368), .ZN(n14367) );
  NOR2_X1 U17618 ( .A1(n14238), .A2(n14367), .ZN(n14240) );
  XNOR2_X1 U17619 ( .A(n14240), .B(n14239), .ZN(n15919) );
  AOI22_X1 U17620 ( .A1(n20071), .A2(n15919), .B1(n20128), .B2(
        P1_REIP_REG_13__SCAN_IN), .ZN(n14241) );
  OAI21_X1 U17621 ( .B1(n15800), .B2(n14242), .A(n14241), .ZN(n14243) );
  AOI21_X1 U17622 ( .B1(n14244), .B2(n20079), .A(n14243), .ZN(n14245) );
  OAI21_X1 U17623 ( .B1(n14246), .B2(n20149), .A(n14245), .ZN(P1_U2986) );
  AOI22_X1 U17624 ( .A1(n9618), .A2(n15818), .B1(n14208), .B2(n15819), .ZN(
        n14247) );
  XOR2_X1 U17625 ( .A(n14247), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(
        n15934) );
  INV_X1 U17626 ( .A(n15934), .ZN(n14253) );
  AOI22_X1 U17627 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14248) );
  OAI21_X1 U17628 ( .B1(n20075), .B2(n14249), .A(n14248), .ZN(n14250) );
  AOI21_X1 U17629 ( .B1(n14251), .B2(n20070), .A(n14250), .ZN(n14252) );
  OAI21_X1 U17630 ( .B1(n14253), .B2(n20089), .A(n14252), .ZN(P1_U2989) );
  AOI21_X1 U17631 ( .B1(n14255), .B2(n15957), .A(n14254), .ZN(n14256) );
  XOR2_X1 U17632 ( .A(n9677), .B(n14256), .Z(n15952) );
  INV_X1 U17633 ( .A(n15952), .ZN(n14262) );
  AOI22_X1 U17634 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14257) );
  OAI21_X1 U17635 ( .B1(n20075), .B2(n14258), .A(n14257), .ZN(n14259) );
  AOI21_X1 U17636 ( .B1(n14260), .B2(n20070), .A(n14259), .ZN(n14261) );
  OAI21_X1 U17637 ( .B1(n14262), .B2(n20089), .A(n14261), .ZN(P1_U2991) );
  OAI22_X1 U17638 ( .A1(n14263), .A2(n20089), .B1(n20075), .B2(n19924), .ZN(
        n14264) );
  AOI211_X1 U17639 ( .C1(n20086), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n14265), .B(n14264), .ZN(n14266) );
  OAI21_X1 U17640 ( .B1(n19919), .B2(n20149), .A(n14266), .ZN(P1_U2993) );
  NAND2_X1 U17641 ( .A1(n14267), .A2(n20130), .ZN(n14280) );
  INV_X1 U17642 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15867) );
  INV_X1 U17643 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15938) );
  NAND3_X1 U17644 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15935) );
  NOR3_X1 U17645 ( .A1(n15938), .A2(n15945), .A3(n15935), .ZN(n14374) );
  NAND2_X1 U17646 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14374), .ZN(
        n14372) );
  NOR2_X1 U17647 ( .A1(n14268), .A2(n14372), .ZN(n14341) );
  NAND4_X1 U17648 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15886) );
  NOR3_X1 U17649 ( .A1(n15894), .A2(n15916), .A3(n15886), .ZN(n14324) );
  NAND2_X1 U17650 ( .A1(n14341), .A2(n14324), .ZN(n14272) );
  NAND2_X1 U17651 ( .A1(n14313), .A2(n15863), .ZN(n15850) );
  NOR2_X1 U17652 ( .A1(n15853), .A2(n15850), .ZN(n14304) );
  NAND2_X1 U17653 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n14304), .ZN(
        n15847) );
  NOR2_X1 U17654 ( .A1(n14294), .A2(n15847), .ZN(n15567) );
  NOR2_X1 U17655 ( .A1(n20127), .A2(n20111), .ZN(n14275) );
  INV_X1 U17656 ( .A(n14275), .ZN(n15565) );
  NAND2_X1 U17657 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15872) );
  NOR2_X1 U17658 ( .A1(n15596), .A2(n15884), .ZN(n14323) );
  NOR2_X1 U17659 ( .A1(n14271), .A2(n20093), .ZN(n14375) );
  AOI21_X1 U17660 ( .B1(n14342), .B2(n14376), .A(n14375), .ZN(n15930) );
  OAI21_X1 U17661 ( .B1(n14323), .B2(n15948), .A(n9630), .ZN(n15866) );
  AOI21_X1 U17662 ( .B1(n20127), .B2(n15872), .A(n15866), .ZN(n15859) );
  OAI21_X1 U17663 ( .B1(n14273), .B2(n15948), .A(n15859), .ZN(n15852) );
  NOR2_X1 U17664 ( .A1(n14303), .A2(n15852), .ZN(n14274) );
  NOR2_X1 U17665 ( .A1(n14275), .A2(n14274), .ZN(n15843) );
  AOI21_X1 U17666 ( .B1(n14294), .B2(n15565), .A(n15843), .ZN(n14282) );
  OAI211_X1 U17667 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15948), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n14282), .ZN(n15564) );
  OAI221_X1 U17668 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n15567), .A(n15564), .ZN(
        n14279) );
  NAND2_X1 U17669 ( .A1(n14276), .A2(n20131), .ZN(n14277) );
  NAND4_X1 U17670 ( .A1(n14280), .A2(n14279), .A3(n14278), .A4(n14277), .ZN(
        P1_U3001) );
  INV_X1 U17671 ( .A(n14281), .ZN(n14287) );
  NOR2_X1 U17672 ( .A1(n14282), .A2(n14285), .ZN(n14284) );
  OAI22_X1 U17673 ( .A1(n15616), .A2(n20116), .B1(n20114), .B2(n20815), .ZN(
        n14283) );
  AOI211_X1 U17674 ( .C1(n15567), .C2(n14285), .A(n14284), .B(n14283), .ZN(
        n14286) );
  OAI21_X1 U17675 ( .B1(n14287), .B2(n20120), .A(n14286), .ZN(P1_U3002) );
  NAND2_X1 U17676 ( .A1(n14288), .A2(n20130), .ZN(n14297) );
  AOI21_X1 U17677 ( .B1(n14290), .B2(n14289), .A(n15847), .ZN(n14295) );
  NAND2_X1 U17678 ( .A1(n20128), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14292) );
  NAND2_X1 U17679 ( .A1(n15843), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14291) );
  OAI211_X1 U17680 ( .C1(n15621), .C2(n20116), .A(n14292), .B(n14291), .ZN(
        n14293) );
  AOI21_X1 U17681 ( .B1(n14295), .B2(n14294), .A(n14293), .ZN(n14296) );
  NAND2_X1 U17682 ( .A1(n14297), .A2(n14296), .ZN(P1_U3003) );
  NOR2_X1 U17683 ( .A1(n14298), .A2(n14299), .ZN(n14301) );
  OAI21_X1 U17684 ( .B1(n9618), .B2(n14301), .A(n14300), .ZN(n14302) );
  XOR2_X1 U17685 ( .A(n14302), .B(n14303), .Z(n15764) );
  AOI22_X1 U17686 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15852), .B1(
        n14304), .B2(n14303), .ZN(n14306) );
  NAND2_X1 U17687 ( .A1(n20128), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14305) );
  OAI211_X1 U17688 ( .C1(n20116), .C2(n15639), .A(n14306), .B(n14305), .ZN(
        n14307) );
  AOI21_X1 U17689 ( .B1(n15764), .B2(n20130), .A(n14307), .ZN(n14308) );
  INV_X1 U17690 ( .A(n14308), .ZN(P1_U3005) );
  NAND3_X1 U17691 ( .A1(n9618), .A2(n14310), .A3(n14298), .ZN(n14309) );
  OAI21_X1 U17692 ( .B1(n9618), .B2(n14310), .A(n14309), .ZN(n14311) );
  XOR2_X1 U17693 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14311), .Z(
        n15769) );
  AOI221_X1 U17694 ( .B1(n14313), .B2(n15859), .C1(n14343), .C2(n15859), .A(
        n14312), .ZN(n14314) );
  OAI21_X1 U17695 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15863), .A(
        n14314), .ZN(n14317) );
  AOI22_X1 U17696 ( .A1(n14315), .A2(n20131), .B1(n20128), .B2(
        P1_REIP_REG_24__SCAN_IN), .ZN(n14316) );
  NAND2_X1 U17697 ( .A1(n14317), .A2(n14316), .ZN(n14318) );
  AOI21_X1 U17698 ( .B1(n15769), .B2(n20130), .A(n14318), .ZN(n14319) );
  INV_X1 U17699 ( .A(n14319), .ZN(P1_U3007) );
  NAND3_X1 U17700 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n14320), .A3(
        n15819), .ZN(n15590) );
  NAND3_X1 U17701 ( .A1(n9618), .A2(n14321), .A3(n15884), .ZN(n15591) );
  AOI22_X1 U17702 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15590), .B1(
        n15591), .B2(n15596), .ZN(n14322) );
  XOR2_X1 U17703 ( .A(n11905), .B(n14322), .Z(n15784) );
  OR2_X1 U17704 ( .A1(n15784), .A2(n20120), .ZN(n14334) );
  AOI22_X1 U17705 ( .A1(n15660), .A2(n20131), .B1(n20128), .B2(
        P1_REIP_REG_21__SCAN_IN), .ZN(n14333) );
  NAND2_X1 U17706 ( .A1(n15866), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14332) );
  INV_X1 U17707 ( .A(n14323), .ZN(n14330) );
  NAND2_X1 U17708 ( .A1(n14375), .A2(n14341), .ZN(n15923) );
  NAND3_X1 U17709 ( .A1(n20092), .A2(n14342), .A3(n14341), .ZN(n14326) );
  INV_X1 U17710 ( .A(n14324), .ZN(n14325) );
  AOI21_X1 U17711 ( .B1(n15923), .B2(n14326), .A(n14325), .ZN(n15879) );
  NOR2_X1 U17712 ( .A1(n20110), .A2(n15923), .ZN(n14346) );
  INV_X1 U17713 ( .A(n14326), .ZN(n14327) );
  AOI21_X1 U17714 ( .B1(n14328), .B2(n14346), .A(n14327), .ZN(n15912) );
  NAND2_X1 U17715 ( .A1(n15912), .A2(n14329), .ZN(n15588) );
  NAND2_X1 U17716 ( .A1(n15879), .A2(n15588), .ZN(n15589) );
  NOR2_X1 U17717 ( .A1(n14330), .A2(n15589), .ZN(n15873) );
  NAND2_X1 U17718 ( .A1(n15873), .A2(n11905), .ZN(n14331) );
  NAND4_X1 U17719 ( .A1(n14334), .A2(n14333), .A3(n14332), .A4(n14331), .ZN(
        P1_U3010) );
  INV_X1 U17720 ( .A(n14335), .ZN(n14337) );
  AOI21_X1 U17721 ( .B1(n14338), .B2(n14337), .A(n14336), .ZN(n14339) );
  XNOR2_X1 U17722 ( .A(n14340), .B(n14339), .ZN(n15803) );
  INV_X1 U17723 ( .A(n15803), .ZN(n14355) );
  INV_X1 U17724 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15910) );
  NAND2_X1 U17725 ( .A1(n14342), .A2(n14341), .ZN(n14349) );
  NOR3_X1 U17726 ( .A1(n14343), .A2(n15916), .A3(n14349), .ZN(n15897) );
  INV_X1 U17727 ( .A(n15897), .ZN(n15887) );
  NOR4_X1 U17728 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15895), .A3(
        n15910), .A4(n15887), .ZN(n14353) );
  OAI21_X1 U17729 ( .B1(n15916), .B2(n15923), .A(n14344), .ZN(n15922) );
  OAI21_X1 U17730 ( .B1(n14346), .B2(n14345), .A(n15922), .ZN(n14347) );
  AOI211_X1 U17731 ( .C1(n20092), .C2(n14349), .A(n14348), .B(n14347), .ZN(
        n15917) );
  OAI21_X1 U17732 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15912), .A(
        n15917), .ZN(n15885) );
  AOI21_X1 U17733 ( .B1(n15895), .B2(n20127), .A(n15885), .ZN(n15911) );
  NAND3_X1 U17734 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15897), .A3(
        n15910), .ZN(n15908) );
  AOI21_X1 U17735 ( .B1(n15911), .B2(n15908), .A(n15896), .ZN(n14352) );
  INV_X1 U17736 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14350) );
  OAI22_X1 U17737 ( .A1(n15690), .A2(n20116), .B1(n20114), .B2(n14350), .ZN(
        n14351) );
  NOR3_X1 U17738 ( .A1(n14353), .A2(n14352), .A3(n14351), .ZN(n14354) );
  OAI21_X1 U17739 ( .B1(n14355), .B2(n20120), .A(n14354), .ZN(P1_U3015) );
  INV_X1 U17740 ( .A(n14356), .ZN(n14361) );
  NOR2_X1 U17741 ( .A1(n14358), .A2(n14357), .ZN(n14360) );
  OAI21_X1 U17742 ( .B1(n14361), .B2(n14360), .A(n14359), .ZN(n14363) );
  AOI22_X1 U17743 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n9618), .B1(
        n15819), .B2(n15895), .ZN(n14362) );
  XNOR2_X1 U17744 ( .A(n14363), .B(n14362), .ZN(n15812) );
  INV_X1 U17745 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20794) );
  OAI22_X1 U17746 ( .A1(n15709), .A2(n20116), .B1(n20794), .B2(n20114), .ZN(
        n14364) );
  AOI21_X1 U17747 ( .B1(n15885), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n14364), .ZN(n14366) );
  NAND2_X1 U17748 ( .A1(n15897), .A2(n15895), .ZN(n14365) );
  OAI211_X1 U17749 ( .C1(n15812), .C2(n20120), .A(n14366), .B(n14365), .ZN(
        P1_U3017) );
  AOI21_X1 U17750 ( .B1(n14369), .B2(n14368), .A(n14367), .ZN(n15817) );
  NOR2_X1 U17751 ( .A1(n20114), .A2(n20792), .ZN(n14383) );
  NOR2_X1 U17752 ( .A1(n14372), .A2(n15953), .ZN(n14381) );
  NAND2_X1 U17753 ( .A1(n14374), .A2(n14370), .ZN(n15929) );
  INV_X1 U17754 ( .A(n15929), .ZN(n14377) );
  AOI21_X1 U17755 ( .B1(n20092), .B2(n14372), .A(n14371), .ZN(n14373) );
  OAI221_X1 U17756 ( .B1(n14376), .B2(n14375), .C1(n14376), .C2(n14374), .A(
        n14373), .ZN(n15925) );
  AOI21_X1 U17757 ( .B1(n14378), .B2(n14377), .A(n15925), .ZN(n14379) );
  INV_X1 U17758 ( .A(n14379), .ZN(n14380) );
  MUX2_X1 U17759 ( .A(n14381), .B(n14380), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n14382) );
  AOI211_X1 U17760 ( .C1(n20131), .C2(n15720), .A(n14383), .B(n14382), .ZN(
        n14384) );
  OAI21_X1 U17761 ( .B1(n15817), .B2(n20120), .A(n14384), .ZN(P1_U3019) );
  NAND2_X1 U17762 ( .A1(n20617), .A2(n14399), .ZN(n20566) );
  NAND2_X1 U17763 ( .A1(n14387), .A2(n20566), .ZN(n20696) );
  OAI21_X1 U17764 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9620), .A(n20696), 
        .ZN(n14388) );
  OAI21_X1 U17765 ( .B1(n14400), .B2(n14385), .A(n14388), .ZN(n14389) );
  MUX2_X1 U17766 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14389), .S(
        n20137), .Z(P1_U3477) );
  NAND3_X1 U17767 ( .A1(n9620), .A2(n20701), .A3(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14391) );
  MUX2_X1 U17768 ( .A(n14391), .B(n20538), .S(n20139), .Z(n14392) );
  OAI21_X1 U17769 ( .B1(n14400), .B2(n12991), .A(n14392), .ZN(n14393) );
  MUX2_X1 U17770 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14393), .S(
        n20137), .Z(P1_U3476) );
  NAND2_X1 U17771 ( .A1(n20139), .A2(n14395), .ZN(n20403) );
  MUX2_X1 U17772 ( .A(n20642), .B(n20403), .S(n9620), .Z(n14397) );
  INV_X1 U17773 ( .A(n20139), .ZN(n14396) );
  AOI21_X1 U17774 ( .B1(n14397), .B2(n20541), .A(n14399), .ZN(n14398) );
  AOI21_X1 U17775 ( .B1(n14399), .B2(n20140), .A(n14398), .ZN(n14402) );
  OAI22_X1 U17776 ( .A1(n14402), .A2(n20693), .B1(n14401), .B2(n14400), .ZN(
        n14403) );
  MUX2_X1 U17777 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n14403), .S(
        n20137), .Z(P1_U3475) );
  INV_X1 U17778 ( .A(n14385), .ZN(n20638) );
  INV_X1 U17779 ( .A(n12999), .ZN(n14404) );
  NAND2_X1 U17780 ( .A1(n14405), .A2(n14404), .ZN(n14407) );
  OAI22_X1 U17781 ( .A1(n15583), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n14407), .B2(n14406), .ZN(n14408) );
  AOI21_X1 U17782 ( .B1(n20638), .B2(n14409), .A(n14408), .ZN(n15528) );
  INV_X1 U17783 ( .A(n14410), .ZN(n20834) );
  NOR3_X1 U17784 ( .A1(n13203), .A2(n12999), .A3(n20832), .ZN(n14411) );
  AOI21_X1 U17785 ( .B1(n14413), .B2(n14412), .A(n14411), .ZN(n14414) );
  OAI21_X1 U17786 ( .B1(n15528), .B2(n20834), .A(n14414), .ZN(n14415) );
  MUX2_X1 U17787 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14415), .S(
        n20836), .Z(P1_U3473) );
  NOR2_X1 U17788 ( .A1(n19016), .A2(n14416), .ZN(n14418) );
  XNOR2_X1 U17789 ( .A(n14418), .B(n14417), .ZN(n14420) );
  NAND2_X1 U17790 ( .A1(n14420), .A2(n14419), .ZN(n14428) );
  OAI22_X1 U17791 ( .A1(n19733), .A2(n19004), .B1(n14421), .B2(n18989), .ZN(
        n14424) );
  OAI22_X1 U17792 ( .A1(n19006), .A2(n10420), .B1(n14422), .B2(n19032), .ZN(
        n14423) );
  AOI211_X1 U17793 ( .C1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n19038), .A(
        n14424), .B(n14423), .ZN(n14427) );
  AOI22_X1 U17794 ( .A1(n15366), .A2(n19035), .B1(n18998), .B2(n14425), .ZN(
        n14426) );
  NAND3_X1 U17795 ( .A1(n14428), .A2(n14427), .A3(n14426), .ZN(P2_U2853) );
  OR2_X1 U17796 ( .A1(n14439), .A2(n14429), .ZN(n14430) );
  NAND2_X1 U17797 ( .A1(n14431), .A2(n14430), .ZN(n15994) );
  OR2_X1 U17798 ( .A1(n14433), .A2(n14432), .ZN(n14517) );
  NAND3_X1 U17799 ( .A1(n14517), .A2(n14434), .A3(n19081), .ZN(n14436) );
  NAND2_X1 U17800 ( .A1(n19084), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14435) );
  OAI211_X1 U17801 ( .C1(n19084), .C2(n15994), .A(n14436), .B(n14435), .ZN(
        P2_U2858) );
  AND2_X1 U17802 ( .A1(n14451), .A2(n14437), .ZN(n14438) );
  OR2_X1 U17803 ( .A1(n14439), .A2(n14438), .ZN(n14793) );
  NAND2_X1 U17804 ( .A1(n14441), .A2(n14440), .ZN(n14443) );
  XNOR2_X1 U17805 ( .A(n14443), .B(n14442), .ZN(n14679) );
  NAND2_X1 U17806 ( .A1(n14679), .A2(n19081), .ZN(n14445) );
  NAND2_X1 U17807 ( .A1(n19084), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14444) );
  OAI211_X1 U17808 ( .C1(n14793), .C2(n19084), .A(n14445), .B(n14444), .ZN(
        P2_U2859) );
  OAI21_X1 U17809 ( .B1(n14448), .B2(n14447), .A(n14446), .ZN(n14692) );
  NAND2_X1 U17810 ( .A1(n19084), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14453) );
  NAND2_X1 U17811 ( .A1(n14454), .A2(n14449), .ZN(n14450) );
  NAND2_X1 U17812 ( .A1(n16018), .A2(n19070), .ZN(n14452) );
  OAI211_X1 U17813 ( .C1(n14692), .C2(n19075), .A(n14453), .B(n14452), .ZN(
        P2_U2860) );
  OAI21_X1 U17814 ( .B1(n9690), .B2(n14455), .A(n14454), .ZN(n15063) );
  AOI21_X1 U17815 ( .B1(n14458), .B2(n14457), .A(n14456), .ZN(n14693) );
  NAND2_X1 U17816 ( .A1(n14693), .A2(n19081), .ZN(n14460) );
  NAND2_X1 U17817 ( .A1(n19084), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14459) );
  OAI211_X1 U17818 ( .C1(n15063), .C2(n19084), .A(n14460), .B(n14459), .ZN(
        P2_U2861) );
  OAI21_X1 U17819 ( .B1(n14463), .B2(n14462), .A(n14461), .ZN(n14709) );
  AND2_X1 U17820 ( .A1(n14471), .A2(n14464), .ZN(n14465) );
  OR2_X1 U17821 ( .A1(n14465), .A2(n9690), .ZN(n14818) );
  MUX2_X1 U17822 ( .A(n14818), .B(n14466), .S(n19084), .Z(n14467) );
  OAI21_X1 U17823 ( .B1(n14709), .B2(n19075), .A(n14467), .ZN(P2_U2862) );
  NAND2_X1 U17824 ( .A1(n9705), .A2(n14468), .ZN(n14710) );
  NAND3_X1 U17825 ( .A1(n14711), .A2(n19081), .A3(n14710), .ZN(n14473) );
  NAND2_X1 U17826 ( .A1(n14476), .A2(n14469), .ZN(n14470) );
  NAND2_X1 U17827 ( .A1(n14471), .A2(n14470), .ZN(n16056) );
  INV_X1 U17828 ( .A(n16056), .ZN(n15086) );
  NAND2_X1 U17829 ( .A1(n15086), .A2(n19070), .ZN(n14472) );
  OAI211_X1 U17830 ( .C1(n19070), .C2(n12054), .A(n14473), .B(n14472), .ZN(
        P2_U2863) );
  OR2_X1 U17831 ( .A1(n14474), .A2(n15112), .ZN(n14475) );
  AND2_X1 U17832 ( .A1(n14476), .A2(n14475), .ZN(n16060) );
  INV_X1 U17833 ( .A(n16060), .ZN(n14482) );
  AOI21_X1 U17834 ( .B1(n14479), .B2(n14478), .A(n14477), .ZN(n14727) );
  NAND2_X1 U17835 ( .A1(n14727), .A2(n19081), .ZN(n14481) );
  NAND2_X1 U17836 ( .A1(n19084), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14480) );
  OAI211_X1 U17837 ( .C1(n14482), .C2(n19084), .A(n14481), .B(n14480), .ZN(
        P2_U2864) );
  OR2_X1 U17838 ( .A1(n14484), .A2(n14485), .ZN(n14486) );
  NAND2_X1 U17839 ( .A1(n14483), .A2(n14486), .ZN(n14744) );
  AND2_X1 U17840 ( .A1(n9695), .A2(n14487), .ZN(n14488) );
  OR2_X1 U17841 ( .A1(n15111), .A2(n14488), .ZN(n15134) );
  NOR2_X1 U17842 ( .A1(n15134), .A2(n19084), .ZN(n14489) );
  AOI21_X1 U17843 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n19084), .A(n14489), .ZN(
        n14490) );
  OAI21_X1 U17844 ( .B1(n14744), .B2(n19075), .A(n14490), .ZN(P2_U2866) );
  NOR2_X1 U17845 ( .A1(n14902), .A2(n14491), .ZN(n14492) );
  OR2_X1 U17846 ( .A1(n14873), .A2(n14492), .ZN(n15158) );
  AOI21_X1 U17847 ( .B1(n14495), .B2(n16077), .A(n14494), .ZN(n14751) );
  NAND2_X1 U17848 ( .A1(n14751), .A2(n19081), .ZN(n14497) );
  NAND2_X1 U17849 ( .A1(n19084), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14496) );
  OAI211_X1 U17850 ( .C1(n15158), .C2(n19084), .A(n14497), .B(n14496), .ZN(
        P2_U2868) );
  AND2_X1 U17851 ( .A1(n9709), .A2(n14499), .ZN(n19043) );
  OR2_X1 U17852 ( .A1(n19043), .A2(n14500), .ZN(n14501) );
  NAND2_X1 U17853 ( .A1(n14498), .A2(n14501), .ZN(n14761) );
  NAND2_X1 U17854 ( .A1(n19084), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14503) );
  NAND2_X1 U17855 ( .A1(n18863), .A2(n19070), .ZN(n14502) );
  OAI211_X1 U17856 ( .C1(n14761), .C2(n19075), .A(n14503), .B(n14502), .ZN(
        P2_U2870) );
  NAND2_X1 U17857 ( .A1(n14504), .A2(n19105), .ZN(n14516) );
  AOI22_X1 U17858 ( .A1(n9658), .A2(n19096), .B1(P2_EAX_REG_30__SCAN_IN), .B2(
        n19102), .ZN(n14515) );
  AND2_X1 U17859 ( .A1(n10362), .A2(n14505), .ZN(n14506) );
  NAND2_X1 U17860 ( .A1(n14509), .A2(n14506), .ZN(n19101) );
  AND2_X1 U17861 ( .A1(n10362), .A2(n14507), .ZN(n14508) );
  AOI22_X1 U17862 ( .A1(n19085), .A2(BUF2_REG_30__SCAN_IN), .B1(n19087), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n14514) );
  INV_X1 U17863 ( .A(n14510), .ZN(n14511) );
  NAND2_X1 U17864 ( .A1(n14755), .A2(n14512), .ZN(n14513) );
  NAND4_X1 U17865 ( .A1(n14516), .A2(n14515), .A3(n14514), .A4(n14513), .ZN(
        P2_U2889) );
  NAND3_X1 U17866 ( .A1(n14517), .A2(n14434), .A3(n19105), .ZN(n14526) );
  AND2_X1 U17867 ( .A1(n14674), .A2(n14518), .ZN(n14519) );
  OAI22_X1 U17868 ( .A1(n15993), .A2(n16085), .B1(n14687), .B2(n14521), .ZN(
        n14522) );
  AOI21_X1 U17869 ( .B1(n14755), .B2(n14523), .A(n14522), .ZN(n14525) );
  AOI22_X1 U17870 ( .A1(n19085), .A2(BUF2_REG_29__SCAN_IN), .B1(n19087), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14524) );
  NAND3_X1 U17871 ( .A1(n14526), .A2(n14525), .A3(n14524), .ZN(P2_U2890) );
  NAND2_X1 U17872 ( .A1(keyinput59), .A2(keyinput3), .ZN(n14530) );
  NOR3_X1 U17873 ( .A1(keyinput57), .A2(keyinput16), .A3(keyinput12), .ZN(
        n14528) );
  NOR3_X1 U17874 ( .A1(keyinput21), .A2(keyinput13), .A3(keyinput35), .ZN(
        n14527) );
  NAND4_X1 U17875 ( .A1(keyinput22), .A2(n14528), .A3(keyinput25), .A4(n14527), 
        .ZN(n14529) );
  NOR4_X1 U17876 ( .A1(keyinput26), .A2(keyinput39), .A3(n14530), .A4(n14529), 
        .ZN(n14532) );
  INV_X1 U17877 ( .A(keyinput60), .ZN(n14531) );
  NAND4_X1 U17878 ( .A1(keyinput19), .A2(keyinput27), .A3(n14532), .A4(n14531), 
        .ZN(n14547) );
  NOR2_X1 U17879 ( .A1(keyinput1), .A2(keyinput55), .ZN(n14538) );
  NAND2_X1 U17880 ( .A1(keyinput29), .A2(keyinput18), .ZN(n14536) );
  NOR3_X1 U17881 ( .A1(keyinput36), .A2(keyinput14), .A3(keyinput15), .ZN(
        n14534) );
  INV_X1 U17882 ( .A(keyinput30), .ZN(n14654) );
  INV_X1 U17883 ( .A(keyinput56), .ZN(n14663) );
  AND3_X1 U17884 ( .A1(n14654), .A2(n14663), .A3(keyinput47), .ZN(n14533) );
  NAND4_X1 U17885 ( .A1(keyinput8), .A2(n14534), .A3(keyinput11), .A4(n14533), 
        .ZN(n14535) );
  NOR4_X1 U17886 ( .A1(keyinput54), .A2(keyinput40), .A3(n14536), .A4(n14535), 
        .ZN(n14537) );
  NAND4_X1 U17887 ( .A1(keyinput17), .A2(keyinput38), .A3(n14538), .A4(n14537), 
        .ZN(n14546) );
  INV_X1 U17888 ( .A(keyinput37), .ZN(n14539) );
  NAND4_X1 U17889 ( .A1(keyinput2), .A2(keyinput52), .A3(keyinput9), .A4(
        n14539), .ZN(n14545) );
  NOR4_X1 U17890 ( .A1(keyinput61), .A2(keyinput46), .A3(keyinput48), .A4(
        keyinput23), .ZN(n14543) );
  NAND3_X1 U17891 ( .A1(keyinput28), .A2(keyinput33), .A3(keyinput63), .ZN(
        n14541) );
  NAND3_X1 U17892 ( .A1(keyinput34), .A2(keyinput45), .A3(keyinput44), .ZN(
        n14540) );
  NOR4_X1 U17893 ( .A1(keyinput42), .A2(keyinput5), .A3(n14541), .A4(n14540), 
        .ZN(n14542) );
  NAND2_X1 U17894 ( .A1(n14543), .A2(n14542), .ZN(n14544) );
  NOR4_X1 U17895 ( .A1(n14547), .A2(n14546), .A3(n14545), .A4(n14544), .ZN(
        n14555) );
  NAND3_X1 U17896 ( .A1(keyinput41), .A2(keyinput7), .A3(keyinput20), .ZN(
        n14553) );
  INV_X1 U17897 ( .A(keyinput62), .ZN(n14548) );
  NAND4_X1 U17898 ( .A1(keyinput43), .A2(keyinput0), .A3(keyinput32), .A4(
        n14548), .ZN(n14552) );
  NOR3_X1 U17899 ( .A1(keyinput10), .A2(keyinput53), .A3(keyinput51), .ZN(
        n14550) );
  NOR3_X1 U17900 ( .A1(keyinput4), .A2(keyinput31), .A3(keyinput50), .ZN(
        n14549) );
  NAND4_X1 U17901 ( .A1(keyinput49), .A2(n14550), .A3(keyinput58), .A4(n14549), 
        .ZN(n14551) );
  NOR4_X1 U17902 ( .A1(keyinput24), .A2(n14553), .A3(n14552), .A4(n14551), 
        .ZN(n14554) );
  AOI21_X1 U17903 ( .B1(n14555), .B2(n14554), .A(keyinput6), .ZN(n14671) );
  INV_X1 U17904 ( .A(keyinput49), .ZN(n14557) );
  OAI22_X1 U17905 ( .A1(keyinput51), .A2(n14558), .B1(n14557), .B2(
        P1_REIP_REG_8__SCAN_IN), .ZN(n14556) );
  AOI221_X1 U17906 ( .B1(n14558), .B2(keyinput51), .C1(n14557), .C2(
        P1_REIP_REG_8__SCAN_IN), .A(n14556), .ZN(n14570) );
  INV_X1 U17907 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14561) );
  INV_X1 U17908 ( .A(keyinput53), .ZN(n14560) );
  OAI22_X1 U17909 ( .A1(n14561), .A2(keyinput24), .B1(n14560), .B2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n14559) );
  AOI221_X1 U17910 ( .B1(n14561), .B2(keyinput24), .C1(
        P3_DATAWIDTH_REG_11__SCAN_IN), .C2(n14560), .A(n14559), .ZN(n14569) );
  INV_X1 U17911 ( .A(keyinput20), .ZN(n14563) );
  OAI22_X1 U17912 ( .A1(n14564), .A2(keyinput0), .B1(n14563), .B2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n14562) );
  AOI221_X1 U17913 ( .B1(n14564), .B2(keyinput0), .C1(
        P3_DATAWIDTH_REG_2__SCAN_IN), .C2(n14563), .A(n14562), .ZN(n14568) );
  INV_X1 U17914 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18129) );
  INV_X1 U17915 ( .A(keyinput7), .ZN(n14566) );
  OAI22_X1 U17916 ( .A1(keyinput41), .A2(n18129), .B1(n14566), .B2(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n14565) );
  AOI221_X1 U17917 ( .B1(n18129), .B2(keyinput41), .C1(n14566), .C2(
        P1_ADDRESS_REG_8__SCAN_IN), .A(n14565), .ZN(n14567) );
  NAND4_X1 U17918 ( .A1(n14570), .A2(n14569), .A3(n14568), .A4(n14567), .ZN(
        n14585) );
  INV_X1 U17919 ( .A(DATAI_17_), .ZN(n14573) );
  INV_X1 U17920 ( .A(keyinput35), .ZN(n14572) );
  OAI22_X1 U17921 ( .A1(keyinput13), .A2(n14573), .B1(n14572), .B2(
        P3_ADDRESS_REG_22__SCAN_IN), .ZN(n14571) );
  AOI221_X1 U17922 ( .B1(n14573), .B2(keyinput13), .C1(n14572), .C2(
        P3_ADDRESS_REG_22__SCAN_IN), .A(n14571), .ZN(n14583) );
  INV_X1 U17923 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19747) );
  INV_X1 U17924 ( .A(keyinput25), .ZN(n14575) );
  OAI22_X1 U17925 ( .A1(n19747), .A2(keyinput26), .B1(n14575), .B2(
        P3_EAX_REG_7__SCAN_IN), .ZN(n14574) );
  AOI221_X1 U17926 ( .B1(n19747), .B2(keyinput26), .C1(P3_EAX_REG_7__SCAN_IN), 
        .C2(n14575), .A(n14574), .ZN(n14582) );
  INV_X1 U17927 ( .A(P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n19709) );
  INV_X1 U17928 ( .A(keyinput39), .ZN(n14577) );
  OAI22_X1 U17929 ( .A1(keyinput59), .A2(n19709), .B1(n14577), .B2(
        P1_M_IO_N_REG_SCAN_IN), .ZN(n14576) );
  AOI221_X1 U17930 ( .B1(n19709), .B2(keyinput59), .C1(n14577), .C2(
        P1_M_IO_N_REG_SCAN_IN), .A(n14576), .ZN(n14581) );
  INV_X1 U17931 ( .A(keyinput17), .ZN(n14579) );
  OAI22_X1 U17932 ( .A1(keyinput3), .A2(n20689), .B1(n14579), .B2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .ZN(n14578) );
  AOI221_X1 U17933 ( .B1(n20689), .B2(keyinput3), .C1(n14579), .C2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A(n14578), .ZN(n14580) );
  NAND4_X1 U17934 ( .A1(n14583), .A2(n14582), .A3(n14581), .A4(n14580), .ZN(
        n14584) );
  NOR2_X1 U17935 ( .A1(n14585), .A2(n14584), .ZN(n14589) );
  INV_X1 U17936 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14587) );
  OAI22_X1 U17937 ( .A1(n14587), .A2(keyinput32), .B1(n14821), .B2(keyinput62), 
        .ZN(n14586) );
  AOI221_X1 U17938 ( .B1(n14587), .B2(keyinput32), .C1(keyinput62), .C2(n14821), .A(n14586), .ZN(n14588) );
  NAND2_X1 U17939 ( .A1(n14589), .A2(n14588), .ZN(n14623) );
  INV_X1 U17940 ( .A(keyinput28), .ZN(n14591) );
  OAI22_X1 U17941 ( .A1(keyinput9), .A2(n17685), .B1(n14591), .B2(
        P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14590) );
  AOI221_X1 U17942 ( .B1(n17685), .B2(keyinput9), .C1(n14591), .C2(
        P1_INSTQUEUE_REG_6__4__SCAN_IN), .A(n14590), .ZN(n14600) );
  INV_X1 U17943 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20816) );
  INV_X1 U17944 ( .A(keyinput52), .ZN(n14593) );
  OAI22_X1 U17945 ( .A1(keyinput37), .A2(n20816), .B1(n14593), .B2(
        P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14592) );
  AOI221_X1 U17946 ( .B1(n20816), .B2(keyinput37), .C1(n14593), .C2(
        P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(n14592), .ZN(n14599) );
  INV_X1 U17947 ( .A(keyinput61), .ZN(n14595) );
  OAI22_X1 U17948 ( .A1(n19737), .A2(keyinput33), .B1(n14595), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n14594) );
  AOI221_X1 U17949 ( .B1(n19737), .B2(keyinput33), .C1(
        P1_DATAO_REG_12__SCAN_IN), .C2(n14595), .A(n14594), .ZN(n14598) );
  INV_X1 U17950 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19764) );
  INV_X1 U17951 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19761) );
  OAI22_X1 U17952 ( .A1(n19764), .A2(keyinput42), .B1(n19761), .B2(keyinput63), 
        .ZN(n14596) );
  AOI221_X1 U17953 ( .B1(n19764), .B2(keyinput42), .C1(keyinput63), .C2(n19761), .A(n14596), .ZN(n14597) );
  NAND4_X1 U17954 ( .A1(n14600), .A2(n14599), .A3(n14598), .A4(n14597), .ZN(
        n14622) );
  INV_X1 U17955 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17385) );
  INV_X1 U17956 ( .A(keyinput23), .ZN(n14602) );
  OAI22_X1 U17957 ( .A1(keyinput48), .A2(n17385), .B1(n14602), .B2(
        P3_EAX_REG_19__SCAN_IN), .ZN(n14601) );
  AOI221_X1 U17958 ( .B1(n17385), .B2(keyinput48), .C1(n14602), .C2(
        P3_EAX_REG_19__SCAN_IN), .A(n14601), .ZN(n14613) );
  OAI22_X1 U17959 ( .A1(n19587), .A2(keyinput46), .B1(n19760), .B2(keyinput34), 
        .ZN(n14603) );
  AOI221_X1 U17960 ( .B1(n19587), .B2(keyinput46), .C1(keyinput34), .C2(n19760), .A(n14603), .ZN(n14612) );
  INV_X1 U17961 ( .A(keyinput10), .ZN(n14605) );
  OAI22_X1 U17962 ( .A1(keyinput44), .A2(n14606), .B1(n14605), .B2(
        P2_DATAO_REG_26__SCAN_IN), .ZN(n14604) );
  AOI221_X1 U17963 ( .B1(n14606), .B2(keyinput44), .C1(n14605), .C2(
        P2_DATAO_REG_26__SCAN_IN), .A(n14604), .ZN(n14611) );
  INV_X1 U17964 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n14609) );
  INV_X1 U17965 ( .A(keyinput45), .ZN(n14608) );
  OAI22_X1 U17966 ( .A1(keyinput5), .A2(n14609), .B1(n14608), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n14607) );
  AOI221_X1 U17967 ( .B1(n14609), .B2(keyinput5), .C1(n14608), .C2(
        P1_EBX_REG_12__SCAN_IN), .A(n14607), .ZN(n14610) );
  NAND4_X1 U17968 ( .A1(n14613), .A2(n14612), .A3(n14611), .A4(n14610), .ZN(
        n14621) );
  INV_X1 U17969 ( .A(keyinput31), .ZN(n14614) );
  XOR2_X1 U17970 ( .A(P1_DATAWIDTH_REG_17__SCAN_IN), .B(n14614), .Z(n14619) );
  INV_X1 U17971 ( .A(keyinput36), .ZN(n14615) );
  XOR2_X1 U17972 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B(n14615), .Z(n14618) );
  XNOR2_X1 U17973 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B(keyinput14), .ZN(
        n14617) );
  XNOR2_X1 U17974 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B(keyinput50), .ZN(
        n14616) );
  NAND4_X1 U17975 ( .A1(n14619), .A2(n14618), .A3(n14617), .A4(n14616), .ZN(
        n14620) );
  NOR4_X1 U17976 ( .A1(n14623), .A2(n14622), .A3(n14621), .A4(n14620), .ZN(
        n14669) );
  INV_X1 U17977 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16598) );
  INV_X1 U17978 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20824) );
  OAI22_X1 U17979 ( .A1(n20824), .A2(keyinput6), .B1(n16598), .B2(keyinput60), 
        .ZN(n14624) );
  AOI21_X1 U17980 ( .B1(n16598), .B2(keyinput60), .A(n14624), .ZN(n14634) );
  INV_X1 U17981 ( .A(keyinput57), .ZN(n14626) );
  OAI22_X1 U17982 ( .A1(keyinput19), .A2(n16986), .B1(n14626), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n14625) );
  AOI221_X1 U17983 ( .B1(n16986), .B2(keyinput19), .C1(n14626), .C2(
        BUF1_REG_17__SCAN_IN), .A(n14625), .ZN(n14633) );
  INV_X1 U17984 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17401) );
  INV_X1 U17985 ( .A(keyinput12), .ZN(n14628) );
  OAI22_X1 U17986 ( .A1(keyinput16), .A2(n17401), .B1(n14628), .B2(
        P3_UWORD_REG_8__SCAN_IN), .ZN(n14627) );
  AOI221_X1 U17987 ( .B1(n17401), .B2(keyinput16), .C1(n14628), .C2(
        P3_UWORD_REG_8__SCAN_IN), .A(n14627), .ZN(n14632) );
  INV_X1 U17988 ( .A(keyinput21), .ZN(n14630) );
  OAI22_X1 U17989 ( .A1(keyinput22), .A2(n15896), .B1(n14630), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n14629) );
  AOI221_X1 U17990 ( .B1(n15896), .B2(keyinput22), .C1(n14630), .C2(
        BUF1_REG_18__SCAN_IN), .A(n14629), .ZN(n14631) );
  NAND4_X1 U17991 ( .A1(n14634), .A2(n14633), .A3(n14632), .A4(n14631), .ZN(
        n14650) );
  INV_X1 U17992 ( .A(keyinput55), .ZN(n14636) );
  OAI22_X1 U17993 ( .A1(keyinput1), .A2(n14637), .B1(n14636), .B2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14635) );
  AOI221_X1 U17994 ( .B1(n14637), .B2(keyinput1), .C1(n14636), .C2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n14635), .ZN(n14648) );
  INV_X1 U17995 ( .A(keyinput54), .ZN(n14639) );
  OAI22_X1 U17996 ( .A1(n14640), .A2(keyinput38), .B1(n14639), .B2(
        P1_DATAO_REG_2__SCAN_IN), .ZN(n14638) );
  AOI221_X1 U17997 ( .B1(n14640), .B2(keyinput38), .C1(P1_DATAO_REG_2__SCAN_IN), .C2(n14639), .A(n14638), .ZN(n14647) );
  INV_X1 U17998 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16307) );
  INV_X1 U17999 ( .A(keyinput29), .ZN(n14642) );
  OAI22_X1 U18000 ( .A1(keyinput40), .A2(n16307), .B1(n14642), .B2(
        P2_UWORD_REG_12__SCAN_IN), .ZN(n14641) );
  AOI221_X1 U18001 ( .B1(n16307), .B2(keyinput40), .C1(n14642), .C2(
        P2_UWORD_REG_12__SCAN_IN), .A(n14641), .ZN(n14646) );
  INV_X1 U18002 ( .A(P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20758) );
  INV_X1 U18003 ( .A(keyinput8), .ZN(n14644) );
  OAI22_X1 U18004 ( .A1(keyinput18), .A2(n20758), .B1(n14644), .B2(
        P3_EBX_REG_6__SCAN_IN), .ZN(n14643) );
  AOI221_X1 U18005 ( .B1(n20758), .B2(keyinput18), .C1(n14644), .C2(
        P3_EBX_REG_6__SCAN_IN), .A(n14643), .ZN(n14645) );
  NAND4_X1 U18006 ( .A1(n14648), .A2(n14647), .A3(n14646), .A4(n14645), .ZN(
        n14649) );
  NOR2_X1 U18007 ( .A1(n14650), .A2(n14649), .ZN(n14661) );
  INV_X1 U18008 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19865) );
  INV_X1 U18009 ( .A(keyinput2), .ZN(n14652) );
  OAI22_X1 U18010 ( .A1(keyinput47), .A2(n19865), .B1(n14652), .B2(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14651) );
  AOI221_X1 U18011 ( .B1(n19865), .B2(keyinput47), .C1(n14652), .C2(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .A(n14651), .ZN(n14660) );
  INV_X1 U18012 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n19832) );
  OAI22_X1 U18013 ( .A1(keyinput15), .A2(n19832), .B1(n14654), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n14653) );
  AOI221_X1 U18014 ( .B1(n19832), .B2(keyinput15), .C1(n14654), .C2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(n14653), .ZN(n14659) );
  INV_X1 U18015 ( .A(keyinput4), .ZN(n14656) );
  OAI22_X1 U18016 ( .A1(keyinput43), .A2(n14657), .B1(n14656), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n14655) );
  AOI221_X1 U18017 ( .B1(n14657), .B2(keyinput43), .C1(n14656), .C2(
        P1_EBX_REG_3__SCAN_IN), .A(n14655), .ZN(n14658) );
  AND4_X1 U18018 ( .A1(n14661), .A2(n14660), .A3(n14659), .A4(n14658), .ZN(
        n14668) );
  INV_X1 U18019 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19144) );
  OAI22_X1 U18020 ( .A1(n19144), .A2(keyinput11), .B1(n14663), .B2(
        P3_REIP_REG_21__SCAN_IN), .ZN(n14662) );
  AOI221_X1 U18021 ( .B1(n19144), .B2(keyinput11), .C1(P3_REIP_REG_21__SCAN_IN), .C2(n14663), .A(n14662), .ZN(n14667) );
  INV_X1 U18022 ( .A(DATAI_31_), .ZN(n14665) );
  OAI22_X1 U18023 ( .A1(keyinput27), .A2(n14665), .B1(n20792), .B2(keyinput58), 
        .ZN(n14664) );
  AOI221_X1 U18024 ( .B1(n14665), .B2(keyinput27), .C1(n20792), .C2(keyinput58), .A(n14664), .ZN(n14666) );
  AND4_X1 U18025 ( .A1(n14669), .A2(n14668), .A3(n14667), .A4(n14666), .ZN(
        n14670) );
  OAI21_X1 U18026 ( .B1(n14671), .B2(P1_BE_N_REG_1__SCAN_IN), .A(n14670), .ZN(
        n14681) );
  AOI22_X1 U18027 ( .A1(n19085), .A2(BUF2_REG_28__SCAN_IN), .B1(n19087), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14676) );
  NAND2_X1 U18028 ( .A1(n14685), .A2(n14672), .ZN(n14673) );
  AOI22_X1 U18029 ( .A1(n19096), .A2(n16004), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n19102), .ZN(n14675) );
  OAI211_X1 U18030 ( .C1(n14677), .C2(n19090), .A(n14676), .B(n14675), .ZN(
        n14678) );
  AOI21_X1 U18031 ( .B1(n14679), .B2(n19105), .A(n14678), .ZN(n14680) );
  XOR2_X1 U18032 ( .A(n14681), .B(n14680), .Z(P2_U2891) );
  NAND2_X1 U18033 ( .A1(n14682), .A2(n14683), .ZN(n14684) );
  NAND2_X1 U18034 ( .A1(n14685), .A2(n14684), .ZN(n16024) );
  OAI22_X1 U18035 ( .A1(n16024), .A2(n16085), .B1(n14687), .B2(n14686), .ZN(
        n14688) );
  AOI21_X1 U18036 ( .B1(n14755), .B2(n14689), .A(n14688), .ZN(n14691) );
  AOI22_X1 U18037 ( .A1(n19085), .A2(BUF2_REG_27__SCAN_IN), .B1(n19087), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14690) );
  OAI211_X1 U18038 ( .C1(n14692), .C2(n16083), .A(n14691), .B(n14690), .ZN(
        P2_U2892) );
  NAND2_X1 U18039 ( .A1(n14693), .A2(n19105), .ZN(n14701) );
  OR2_X1 U18040 ( .A1(n14695), .A2(n14694), .ZN(n14696) );
  AND2_X1 U18041 ( .A1(n14682), .A2(n14696), .ZN(n16026) );
  AOI22_X1 U18042 ( .A1(n19096), .A2(n16026), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19102), .ZN(n14700) );
  AOI22_X1 U18043 ( .A1(n19085), .A2(BUF2_REG_26__SCAN_IN), .B1(n19087), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14699) );
  NAND2_X1 U18044 ( .A1(n14755), .A2(n14697), .ZN(n14698) );
  NAND4_X1 U18045 ( .A1(n14701), .A2(n14700), .A3(n14699), .A4(n14698), .ZN(
        P2_U2893) );
  AOI22_X1 U18046 ( .A1(n19085), .A2(BUF2_REG_25__SCAN_IN), .B1(n19087), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14705) );
  INV_X1 U18047 ( .A(n14702), .ZN(n14703) );
  XNOR2_X1 U18048 ( .A(n14713), .B(n14703), .ZN(n16037) );
  AOI22_X1 U18049 ( .A1(n19096), .A2(n16037), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n19102), .ZN(n14704) );
  OAI211_X1 U18050 ( .C1(n14706), .C2(n19090), .A(n14705), .B(n14704), .ZN(
        n14707) );
  INV_X1 U18051 ( .A(n14707), .ZN(n14708) );
  OAI21_X1 U18052 ( .B1(n14709), .B2(n16083), .A(n14708), .ZN(P2_U2894) );
  NAND3_X1 U18053 ( .A1(n14711), .A2(n19105), .A3(n14710), .ZN(n14719) );
  OAI21_X1 U18054 ( .B1(n14712), .B2(n14714), .A(n14713), .ZN(n15089) );
  INV_X1 U18055 ( .A(n15089), .ZN(n16050) );
  AOI22_X1 U18056 ( .A1(n19096), .A2(n16050), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19102), .ZN(n14718) );
  AOI22_X1 U18057 ( .A1(n19085), .A2(BUF2_REG_24__SCAN_IN), .B1(n19087), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14717) );
  NAND2_X1 U18058 ( .A1(n14755), .A2(n14715), .ZN(n14716) );
  NAND4_X1 U18059 ( .A1(n14719), .A2(n14718), .A3(n14717), .A4(n14716), .ZN(
        P2_U2895) );
  NOR2_X1 U18060 ( .A1(n14721), .A2(n14720), .ZN(n14722) );
  OR2_X1 U18061 ( .A1(n14712), .A2(n14722), .ZN(n16058) );
  AOI22_X1 U18062 ( .A1(n19085), .A2(BUF2_REG_23__SCAN_IN), .B1(n19087), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14725) );
  INV_X1 U18063 ( .A(n15348), .ZN(n14723) );
  AOI22_X1 U18064 ( .A1(n14755), .A2(n14723), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n19102), .ZN(n14724) );
  OAI211_X1 U18065 ( .C1(n16085), .C2(n16058), .A(n14725), .B(n14724), .ZN(
        n14726) );
  AOI21_X1 U18066 ( .B1(n14727), .B2(n19105), .A(n14726), .ZN(n14728) );
  INV_X1 U18067 ( .A(n14728), .ZN(P2_U2896) );
  AOI21_X1 U18068 ( .B1(n14730), .B2(n14483), .A(n14729), .ZN(n16070) );
  XNOR2_X1 U18069 ( .A(n14732), .B(n14731), .ZN(n15118) );
  AOI22_X1 U18070 ( .A1(n19085), .A2(BUF2_REG_22__SCAN_IN), .B1(n19087), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n14735) );
  AOI22_X1 U18071 ( .A1(n14755), .A2(n14733), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19102), .ZN(n14734) );
  OAI211_X1 U18072 ( .C1(n16085), .C2(n15118), .A(n14735), .B(n14734), .ZN(
        n14736) );
  AOI21_X1 U18073 ( .B1(n16070), .B2(n19105), .A(n14736), .ZN(n14737) );
  INV_X1 U18074 ( .A(n14737), .ZN(P2_U2897) );
  INV_X1 U18075 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n14739) );
  INV_X1 U18076 ( .A(n19181), .ZN(n19103) );
  AOI22_X1 U18077 ( .A1(n14755), .A2(n19103), .B1(P2_EAX_REG_21__SCAN_IN), 
        .B2(n19102), .ZN(n14738) );
  OAI21_X1 U18078 ( .B1(n19101), .B2(n14739), .A(n14738), .ZN(n14742) );
  OAI21_X1 U18079 ( .B1(n15144), .B2(n14740), .A(n14731), .ZN(n18823) );
  NOR2_X1 U18080 ( .A1(n18823), .A2(n16085), .ZN(n14741) );
  AOI211_X1 U18081 ( .C1(BUF1_REG_21__SCAN_IN), .C2(n19087), .A(n14742), .B(
        n14741), .ZN(n14743) );
  OAI21_X1 U18082 ( .B1(n16083), .B2(n14744), .A(n14743), .ZN(P2_U2898) );
  XNOR2_X1 U18083 ( .A(n15169), .B(n14745), .ZN(n18839) );
  INV_X1 U18084 ( .A(n18839), .ZN(n14753) );
  INV_X1 U18085 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n14749) );
  NAND2_X1 U18086 ( .A1(n19087), .A2(BUF1_REG_19__SCAN_IN), .ZN(n14748) );
  AOI22_X1 U18087 ( .A1(n14755), .A2(n14746), .B1(n19102), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n14747) );
  OAI211_X1 U18088 ( .C1(n19101), .C2(n14749), .A(n14748), .B(n14747), .ZN(
        n14750) );
  AOI21_X1 U18089 ( .B1(n14751), .B2(n19105), .A(n14750), .ZN(n14752) );
  OAI21_X1 U18090 ( .B1(n14753), .B2(n16085), .A(n14752), .ZN(P2_U2900) );
  INV_X1 U18091 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14757) );
  AOI22_X1 U18092 ( .A1(n14755), .A2(n14754), .B1(P2_EAX_REG_17__SCAN_IN), 
        .B2(n19102), .ZN(n14756) );
  OAI21_X1 U18093 ( .B1(n19101), .B2(n14757), .A(n14756), .ZN(n14759) );
  NOR2_X1 U18094 ( .A1(n18869), .A2(n16085), .ZN(n14758) );
  AOI211_X1 U18095 ( .C1(BUF1_REG_17__SCAN_IN), .C2(n19087), .A(n14759), .B(
        n14758), .ZN(n14760) );
  OAI21_X1 U18096 ( .B1(n16083), .B2(n14761), .A(n14760), .ZN(P2_U2902) );
  NOR2_X1 U18097 ( .A1(n14762), .A2(n14773), .ZN(n14765) );
  NAND2_X1 U18098 ( .A1(n10160), .A2(n14763), .ZN(n14764) );
  XNOR2_X1 U18099 ( .A(n14765), .B(n14764), .ZN(n15025) );
  INV_X1 U18100 ( .A(n14777), .ZN(n14768) );
  INV_X1 U18101 ( .A(n14766), .ZN(n14767) );
  AOI21_X1 U18102 ( .B1(n15015), .B2(n14768), .A(n14767), .ZN(n15023) );
  NOR2_X1 U18103 ( .A1(n18974), .A2(n19777), .ZN(n15018) );
  NOR2_X1 U18104 ( .A1(n16150), .A2(n15983), .ZN(n14769) );
  AOI211_X1 U18105 ( .C1(n16142), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15018), .B(n14769), .ZN(n14770) );
  OAI21_X1 U18106 ( .B1(n15020), .B2(n16138), .A(n14770), .ZN(n14771) );
  AOI21_X1 U18107 ( .B1(n15023), .B2(n16146), .A(n14771), .ZN(n14772) );
  OAI21_X1 U18108 ( .B1(n15025), .B2(n16152), .A(n14772), .ZN(P2_U2984) );
  NOR2_X1 U18109 ( .A1(n14774), .A2(n14773), .ZN(n14776) );
  XOR2_X1 U18110 ( .A(n14776), .B(n14775), .Z(n15035) );
  INV_X1 U18111 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14778) );
  NOR2_X1 U18112 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15027) );
  AOI211_X1 U18113 ( .C1(n14778), .C2(n14802), .A(n15027), .B(n14777), .ZN(
        n15032) );
  NAND2_X1 U18114 ( .A1(n18992), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15029) );
  OAI21_X1 U18115 ( .B1(n16161), .B2(n14779), .A(n15029), .ZN(n14780) );
  AOI21_X1 U18116 ( .B1(n16151), .B2(n14781), .A(n14780), .ZN(n14782) );
  OAI21_X1 U18117 ( .B1(n15994), .B2(n16138), .A(n14782), .ZN(n14783) );
  AOI21_X1 U18118 ( .B1(n15032), .B2(n16146), .A(n14783), .ZN(n14784) );
  OAI21_X1 U18119 ( .B1(n15035), .B2(n16152), .A(n14784), .ZN(P2_U2985) );
  OAI21_X2 U18120 ( .B1(n14786), .B2(n14813), .A(n13720), .ZN(n14787) );
  XOR2_X1 U18121 ( .A(n14788), .B(n14787), .Z(n14798) );
  INV_X1 U18122 ( .A(n14787), .ZN(n14789) );
  OAI22_X1 U18123 ( .A1(n14798), .A2(n15048), .B1(n14789), .B2(n14788), .ZN(
        n14792) );
  XNOR2_X1 U18124 ( .A(n14790), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14791) );
  XNOR2_X1 U18125 ( .A(n14792), .B(n14791), .ZN(n15046) );
  NAND2_X1 U18126 ( .A1(n18992), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15036) );
  NAND2_X1 U18127 ( .A1(n16142), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14794) );
  OAI211_X1 U18128 ( .C1(n16150), .C2(n16008), .A(n15036), .B(n14794), .ZN(
        n14796) );
  XOR2_X1 U18129 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14802), .Z(
        n15041) );
  NOR2_X1 U18130 ( .A1(n15041), .A2(n16154), .ZN(n14795) );
  AOI211_X1 U18131 ( .C1(n16157), .C2(n16005), .A(n14796), .B(n14795), .ZN(
        n14797) );
  OAI21_X1 U18132 ( .B1(n15046), .B2(n16152), .A(n14797), .ZN(P2_U2986) );
  XNOR2_X1 U18133 ( .A(n14798), .B(n15048), .ZN(n15057) );
  NAND2_X1 U18134 ( .A1(n16151), .A2(n14799), .ZN(n14800) );
  NAND2_X1 U18135 ( .A1(n18992), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15047) );
  OAI211_X1 U18136 ( .C1(n16161), .C2(n16014), .A(n14800), .B(n15047), .ZN(
        n14804) );
  NAND2_X1 U18137 ( .A1(n14809), .A2(n15048), .ZN(n14801) );
  NAND2_X1 U18138 ( .A1(n14802), .A2(n14801), .ZN(n15054) );
  NOR2_X1 U18139 ( .A1(n15054), .A2(n16154), .ZN(n14803) );
  AOI211_X1 U18140 ( .C1(n16157), .C2(n16018), .A(n14804), .B(n14803), .ZN(
        n14805) );
  OAI21_X1 U18141 ( .B1(n15057), .B2(n16152), .A(n14805), .ZN(P2_U2987) );
  OAI21_X1 U18142 ( .B1(n14816), .B2(n14813), .A(n14814), .ZN(n14806) );
  XOR2_X1 U18143 ( .A(n14807), .B(n14806), .Z(n15070) );
  INV_X1 U18144 ( .A(n15063), .ZN(n16027) );
  NOR2_X1 U18145 ( .A1(n18974), .A2(n19768), .ZN(n15061) );
  AOI21_X1 U18146 ( .B1(n16142), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15061), .ZN(n14808) );
  OAI21_X1 U18147 ( .B1(n16150), .B2(n16030), .A(n14808), .ZN(n14811) );
  OAI21_X1 U18148 ( .B1(n9659), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14809), .ZN(n15064) );
  NOR2_X1 U18149 ( .A1(n15064), .A2(n16154), .ZN(n14810) );
  AOI211_X1 U18150 ( .C1(n16157), .C2(n16027), .A(n14811), .B(n14810), .ZN(
        n14812) );
  OAI21_X1 U18151 ( .B1(n15070), .B2(n16152), .A(n14812), .ZN(P2_U2988) );
  INV_X1 U18152 ( .A(n14813), .ZN(n14815) );
  NAND2_X1 U18153 ( .A1(n14815), .A2(n14814), .ZN(n14817) );
  XOR2_X1 U18154 ( .A(n14817), .B(n14816), .Z(n15081) );
  INV_X1 U18155 ( .A(n15081), .ZN(n14825) );
  INV_X1 U18156 ( .A(n14818), .ZN(n16038) );
  NAND2_X1 U18157 ( .A1(n16151), .A2(n14819), .ZN(n14820) );
  INV_X1 U18158 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19766) );
  OR2_X1 U18159 ( .A1(n18974), .A2(n19766), .ZN(n15072) );
  OAI211_X1 U18160 ( .C1(n16161), .C2(n14821), .A(n14820), .B(n15072), .ZN(
        n14823) );
  NOR2_X1 U18161 ( .A1(n14830), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15071) );
  NOR3_X1 U18162 ( .A1(n15071), .A2(n9659), .A3(n16154), .ZN(n14822) );
  AOI211_X1 U18163 ( .C1(n16038), .C2(n16157), .A(n14823), .B(n14822), .ZN(
        n14824) );
  OAI21_X1 U18164 ( .B1(n14825), .B2(n16152), .A(n14824), .ZN(P2_U2989) );
  NOR2_X1 U18165 ( .A1(n14827), .A2(n9901), .ZN(n14828) );
  XNOR2_X1 U18166 ( .A(n14829), .B(n14828), .ZN(n15093) );
  AOI21_X1 U18167 ( .B1(n14831), .B2(n14839), .A(n14830), .ZN(n15091) );
  NOR2_X1 U18168 ( .A1(n18974), .A2(n14832), .ZN(n15085) );
  NOR2_X1 U18169 ( .A1(n16150), .A2(n16053), .ZN(n14833) );
  AOI211_X1 U18170 ( .C1(n16142), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15085), .B(n14833), .ZN(n14834) );
  OAI21_X1 U18171 ( .B1(n16138), .B2(n16056), .A(n14834), .ZN(n14835) );
  AOI21_X1 U18172 ( .B1(n15091), .B2(n16146), .A(n14835), .ZN(n14836) );
  OAI21_X1 U18173 ( .B1(n15093), .B2(n16152), .A(n14836), .ZN(P2_U2990) );
  INV_X1 U18174 ( .A(n14838), .ZN(n15129) );
  INV_X1 U18175 ( .A(n14839), .ZN(n14840) );
  AOI21_X1 U18176 ( .B1(n15108), .B2(n15098), .A(n14840), .ZN(n15106) );
  NAND2_X1 U18177 ( .A1(n15106), .A2(n16146), .ZN(n14849) );
  OAI22_X1 U18178 ( .A1(n16161), .A2(n14841), .B1(n19763), .B2(n18974), .ZN(
        n14842) );
  AOI21_X1 U18179 ( .B1(n16151), .B2(n14843), .A(n14842), .ZN(n14848) );
  OR2_X1 U18180 ( .A1(n14845), .A2(n14844), .ZN(n15095) );
  NAND3_X1 U18181 ( .A1(n15095), .A2(n15094), .A3(n16145), .ZN(n14847) );
  NAND2_X1 U18182 ( .A1(n16157), .A2(n16060), .ZN(n14846) );
  NAND4_X1 U18183 ( .A1(n14849), .A2(n14848), .A3(n14847), .A4(n14846), .ZN(
        P2_U2991) );
  INV_X1 U18184 ( .A(n14869), .ZN(n14854) );
  AOI21_X1 U18185 ( .B1(n14872), .B2(n14855), .A(n14854), .ZN(n14859) );
  NAND2_X1 U18186 ( .A1(n14857), .A2(n14856), .ZN(n14858) );
  XNOR2_X1 U18187 ( .A(n14859), .B(n14858), .ZN(n15140) );
  AOI21_X1 U18188 ( .B1(n14860), .B2(n14867), .A(n15109), .ZN(n15138) );
  NOR2_X1 U18189 ( .A1(n18974), .A2(n19760), .ZN(n15132) );
  NOR2_X1 U18190 ( .A1(n16161), .A2(n18813), .ZN(n14861) );
  AOI211_X1 U18191 ( .C1(n14862), .C2(n16151), .A(n15132), .B(n14861), .ZN(
        n14863) );
  OAI21_X1 U18192 ( .B1(n15134), .B2(n16138), .A(n14863), .ZN(n14864) );
  AOI21_X1 U18193 ( .B1(n15138), .B2(n16146), .A(n14864), .ZN(n14865) );
  OAI21_X1 U18194 ( .B1(n15140), .B2(n16152), .A(n14865), .ZN(P2_U2993) );
  NAND3_X1 U18195 ( .A1(n14909), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14894) );
  OAI21_X1 U18196 ( .B1(n14894), .B2(n14882), .A(n14866), .ZN(n14868) );
  NAND2_X1 U18197 ( .A1(n14868), .A2(n14867), .ZN(n15157) );
  INV_X1 U18198 ( .A(n14873), .ZN(n14876) );
  INV_X1 U18199 ( .A(n14874), .ZN(n14875) );
  NAND2_X1 U18200 ( .A1(n14876), .A2(n14875), .ZN(n14877) );
  NAND2_X1 U18201 ( .A1(n9695), .A2(n14877), .ZN(n18835) );
  NOR2_X1 U18202 ( .A1(n18966), .A2(n19758), .ZN(n15152) );
  NOR2_X1 U18203 ( .A1(n16150), .A2(n18832), .ZN(n14878) );
  AOI211_X1 U18204 ( .C1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n16142), .A(
        n15152), .B(n14878), .ZN(n14879) );
  OAI21_X1 U18205 ( .B1(n18835), .B2(n16138), .A(n14879), .ZN(n14880) );
  AOI21_X1 U18206 ( .B1(n15155), .B2(n16145), .A(n14880), .ZN(n14881) );
  OAI21_X1 U18207 ( .B1(n16154), .B2(n15157), .A(n14881), .ZN(P2_U2994) );
  XNOR2_X1 U18208 ( .A(n14894), .B(n14882), .ZN(n15168) );
  INV_X1 U18209 ( .A(n14897), .ZN(n14883) );
  NAND2_X1 U18210 ( .A1(n14885), .A2(n14884), .ZN(n14886) );
  XNOR2_X1 U18211 ( .A(n14887), .B(n14886), .ZN(n15165) );
  NOR2_X1 U18212 ( .A1(n18966), .A2(n19756), .ZN(n15159) );
  NOR2_X1 U18213 ( .A1(n16161), .A2(n14888), .ZN(n14889) );
  AOI211_X1 U18214 ( .C1(n14890), .C2(n16151), .A(n15159), .B(n14889), .ZN(
        n14891) );
  OAI21_X1 U18215 ( .B1(n15158), .B2(n16138), .A(n14891), .ZN(n14892) );
  AOI21_X1 U18216 ( .B1(n15165), .B2(n16145), .A(n14892), .ZN(n14893) );
  OAI21_X1 U18217 ( .B1(n15168), .B2(n16154), .A(n14893), .ZN(P2_U2995) );
  OAI21_X1 U18218 ( .B1(n14921), .B2(n11033), .A(n15176), .ZN(n14895) );
  NAND2_X1 U18219 ( .A1(n14895), .A2(n14894), .ZN(n15184) );
  NAND2_X1 U18220 ( .A1(n14897), .A2(n14896), .ZN(n14899) );
  XOR2_X1 U18221 ( .A(n14899), .B(n14898), .Z(n15182) );
  AND2_X1 U18222 ( .A1(n14901), .A2(n14900), .ZN(n14903) );
  OR2_X1 U18223 ( .A1(n14903), .A2(n14902), .ZN(n18858) );
  NOR2_X1 U18224 ( .A1(n18966), .A2(n14904), .ZN(n15174) );
  NOR2_X1 U18225 ( .A1(n18855), .A2(n16150), .ZN(n14905) );
  AOI211_X1 U18226 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n16142), .A(
        n15174), .B(n14905), .ZN(n14906) );
  OAI21_X1 U18227 ( .B1(n18858), .B2(n16138), .A(n14906), .ZN(n14907) );
  AOI21_X1 U18228 ( .B1(n15182), .B2(n16145), .A(n14907), .ZN(n14908) );
  OAI21_X1 U18229 ( .B1(n15184), .B2(n16154), .A(n14908), .ZN(P2_U2996) );
  XNOR2_X1 U18230 ( .A(n14909), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14916) );
  NAND2_X1 U18231 ( .A1(n18863), .A2(n16157), .ZN(n14912) );
  AOI21_X1 U18232 ( .B1(n16142), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n14910), .ZN(n14911) );
  OAI211_X1 U18233 ( .C1(n16150), .C2(n18866), .A(n14912), .B(n14911), .ZN(
        n14913) );
  AOI21_X1 U18234 ( .B1(n14914), .B2(n16145), .A(n14913), .ZN(n14915) );
  OAI21_X1 U18235 ( .B1(n14916), .B2(n16154), .A(n14915), .ZN(P2_U2997) );
  OAI21_X1 U18236 ( .B1(n14919), .B2(n14918), .A(n14917), .ZN(n15190) );
  INV_X1 U18237 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15197) );
  OAI21_X1 U18238 ( .B1(n15193), .B2(n15203), .A(n15197), .ZN(n14920) );
  NAND3_X1 U18239 ( .A1(n14921), .A2(n16146), .A3(n14920), .ZN(n14928) );
  OAI21_X1 U18240 ( .B1(n14923), .B2(n14922), .A(n11019), .ZN(n19047) );
  INV_X1 U18241 ( .A(n19047), .ZN(n14926) );
  NAND2_X1 U18242 ( .A1(n18992), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15189) );
  NAND2_X1 U18243 ( .A1(n16142), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14924) );
  OAI211_X1 U18244 ( .C1(n18876), .C2(n16150), .A(n15189), .B(n14924), .ZN(
        n14925) );
  AOI21_X1 U18245 ( .B1(n14926), .B2(n16157), .A(n14925), .ZN(n14927) );
  OAI211_X1 U18246 ( .C1(n15190), .C2(n16152), .A(n14928), .B(n14927), .ZN(
        P2_U2998) );
  XNOR2_X1 U18247 ( .A(n15193), .B(n15203), .ZN(n15209) );
  NAND2_X1 U18248 ( .A1(n14929), .A2(n14939), .ZN(n14933) );
  NAND2_X1 U18249 ( .A1(n14931), .A2(n14930), .ZN(n14932) );
  XNOR2_X1 U18250 ( .A(n14933), .B(n14932), .ZN(n15207) );
  NAND2_X1 U18251 ( .A1(n18886), .A2(n16157), .ZN(n14935) );
  NOR2_X1 U18252 ( .A1(n18966), .A2(n19750), .ZN(n15199) );
  AOI21_X1 U18253 ( .B1(n16142), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15199), .ZN(n14934) );
  OAI211_X1 U18254 ( .C1(n16150), .C2(n14936), .A(n14935), .B(n14934), .ZN(
        n14937) );
  AOI21_X1 U18255 ( .B1(n15207), .B2(n16145), .A(n14937), .ZN(n14938) );
  OAI21_X1 U18256 ( .B1(n15209), .B2(n16154), .A(n14938), .ZN(P2_U2999) );
  OAI21_X1 U18257 ( .B1(n14950), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15193), .ZN(n15223) );
  NAND2_X1 U18258 ( .A1(n14940), .A2(n14939), .ZN(n14941) );
  XNOR2_X1 U18259 ( .A(n14942), .B(n14941), .ZN(n15221) );
  OAI21_X1 U18260 ( .B1(n9720), .B2(n10124), .A(n14944), .ZN(n19052) );
  NOR2_X1 U18261 ( .A1(n18966), .A2(n14945), .ZN(n15215) );
  NOR2_X1 U18262 ( .A1(n16150), .A2(n18893), .ZN(n14946) );
  AOI211_X1 U18263 ( .C1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n16142), .A(
        n15215), .B(n14946), .ZN(n14947) );
  OAI21_X1 U18264 ( .B1(n19052), .B2(n16138), .A(n14947), .ZN(n14948) );
  AOI21_X1 U18265 ( .B1(n15221), .B2(n16145), .A(n14948), .ZN(n14949) );
  OAI21_X1 U18266 ( .B1(n15223), .B2(n16154), .A(n14949), .ZN(P2_U3000) );
  INV_X1 U18267 ( .A(n15234), .ZN(n14951) );
  OAI21_X1 U18268 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14951), .A(
        n9948), .ZN(n15233) );
  INV_X1 U18269 ( .A(n14952), .ZN(n14953) );
  NOR2_X1 U18270 ( .A1(n14954), .A2(n14953), .ZN(n14955) );
  XNOR2_X1 U18271 ( .A(n14956), .B(n14955), .ZN(n15231) );
  NOR2_X1 U18272 ( .A1(n18966), .A2(n14957), .ZN(n15228) );
  NOR2_X1 U18273 ( .A1(n16161), .A2(n14958), .ZN(n14959) );
  AOI211_X1 U18274 ( .C1(n16151), .C2(n18906), .A(n15228), .B(n14959), .ZN(
        n14960) );
  OAI21_X1 U18275 ( .B1(n14961), .B2(n16138), .A(n14960), .ZN(n14962) );
  AOI21_X1 U18276 ( .B1(n15231), .B2(n16145), .A(n14962), .ZN(n14963) );
  OAI21_X1 U18277 ( .B1(n15233), .B2(n16154), .A(n14963), .ZN(P2_U3001) );
  XNOR2_X1 U18278 ( .A(n14964), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14965) );
  XNOR2_X1 U18279 ( .A(n14966), .B(n14965), .ZN(n15244) );
  INV_X1 U18280 ( .A(n14967), .ZN(n14978) );
  NAND2_X1 U18281 ( .A1(n14978), .A2(n14968), .ZN(n15235) );
  NAND3_X1 U18282 ( .A1(n15235), .A2(n16146), .A3(n15234), .ZN(n14977) );
  OR2_X1 U18283 ( .A1(n14970), .A2(n14969), .ZN(n14971) );
  AND2_X1 U18284 ( .A1(n14972), .A2(n14971), .ZN(n19055) );
  NOR2_X1 U18285 ( .A1(n18966), .A2(n14973), .ZN(n15236) );
  AOI21_X1 U18286 ( .B1(n16142), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15236), .ZN(n14974) );
  OAI21_X1 U18287 ( .B1(n16150), .B2(n18911), .A(n14974), .ZN(n14975) );
  AOI21_X1 U18288 ( .B1(n19055), .B2(n16157), .A(n14975), .ZN(n14976) );
  OAI211_X1 U18289 ( .C1(n15244), .C2(n16152), .A(n14977), .B(n14976), .ZN(
        P2_U3002) );
  INV_X1 U18290 ( .A(n16112), .ZN(n14979) );
  OAI21_X1 U18291 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n14979), .A(
        n14978), .ZN(n15255) );
  NAND2_X1 U18292 ( .A1(n14981), .A2(n14980), .ZN(n15264) );
  INV_X1 U18293 ( .A(n15262), .ZN(n14982) );
  INV_X1 U18294 ( .A(n16107), .ZN(n14983) );
  OAI211_X1 U18295 ( .C1(n16109), .C2(n14983), .A(n16106), .B(n16108), .ZN(
        n14987) );
  NAND2_X1 U18296 ( .A1(n14985), .A2(n14984), .ZN(n14986) );
  XNOR2_X1 U18297 ( .A(n14987), .B(n14986), .ZN(n15253) );
  NOR2_X1 U18298 ( .A1(n18966), .A2(n19745), .ZN(n15247) );
  NOR2_X1 U18299 ( .A1(n16161), .A2(n14988), .ZN(n14989) );
  AOI211_X1 U18300 ( .C1(n10153), .C2(n16151), .A(n15247), .B(n14989), .ZN(
        n14990) );
  OAI21_X1 U18301 ( .B1(n16138), .B2(n18929), .A(n14990), .ZN(n14991) );
  AOI21_X1 U18302 ( .B1(n15253), .B2(n16145), .A(n14991), .ZN(n14992) );
  OAI21_X1 U18303 ( .B1(n15255), .B2(n16154), .A(n14992), .ZN(P2_U3003) );
  XNOR2_X1 U18304 ( .A(n14993), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14994) );
  XNOR2_X1 U18305 ( .A(n14995), .B(n14994), .ZN(n15281) );
  NAND2_X1 U18306 ( .A1(n16129), .A2(n16127), .ZN(n14996) );
  XNOR2_X1 U18307 ( .A(n16130), .B(n14996), .ZN(n15279) );
  OAI22_X1 U18308 ( .A1(n16161), .A2(n14997), .B1(n19739), .B2(n18974), .ZN(
        n14998) );
  AOI21_X1 U18309 ( .B1(n16151), .B2(n18963), .A(n14998), .ZN(n14999) );
  OAI21_X1 U18310 ( .B1(n18968), .B2(n16138), .A(n14999), .ZN(n15000) );
  AOI21_X1 U18311 ( .B1(n15279), .B2(n16145), .A(n15000), .ZN(n15001) );
  OAI21_X1 U18312 ( .B1(n15281), .B2(n16154), .A(n15001), .ZN(P2_U3007) );
  NAND2_X1 U18313 ( .A1(n16204), .A2(n16157), .ZN(n15014) );
  AOI21_X1 U18314 ( .B1(n15004), .B2(n15003), .A(n15002), .ZN(n16201) );
  NOR2_X1 U18315 ( .A1(n18974), .A2(n19024), .ZN(n16202) );
  AOI21_X1 U18316 ( .B1(n16146), .B2(n16201), .A(n16202), .ZN(n15013) );
  INV_X1 U18317 ( .A(n15005), .ZN(n15006) );
  NAND2_X1 U18318 ( .A1(n16161), .A2(n15006), .ZN(n15007) );
  NAND2_X1 U18319 ( .A1(n15007), .A2(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15012) );
  INV_X1 U18320 ( .A(n19025), .ZN(n15008) );
  NAND2_X1 U18321 ( .A1(n15008), .A2(n15003), .ZN(n15010) );
  AND2_X1 U18322 ( .A1(n15010), .A2(n15009), .ZN(n16199) );
  NAND2_X1 U18323 ( .A1(n16145), .A2(n16199), .ZN(n15011) );
  NAND4_X1 U18324 ( .A1(n15014), .A2(n15013), .A3(n15012), .A4(n15011), .ZN(
        P2_U3014) );
  NOR2_X1 U18325 ( .A1(n15016), .A2(n15015), .ZN(n15022) );
  NOR3_X1 U18326 ( .A1(n15026), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15037), .ZN(n15017) );
  OAI21_X1 U18327 ( .B1(n15020), .B2(n19157), .A(n15019), .ZN(n15021) );
  AOI211_X1 U18328 ( .C1(n15023), .C2(n19162), .A(n15022), .B(n15021), .ZN(
        n15024) );
  OAI21_X1 U18329 ( .B1(n15025), .B2(n19155), .A(n15024), .ZN(P2_U3016) );
  NOR2_X1 U18330 ( .A1(n15994), .A2(n19157), .ZN(n15031) );
  OR3_X1 U18331 ( .A1(n15027), .A2(n15037), .A3(n9754), .ZN(n15028) );
  OAI211_X1 U18332 ( .C1(n16184), .C2(n15993), .A(n15029), .B(n15028), .ZN(
        n15030) );
  AOI211_X1 U18333 ( .C1(n15044), .C2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15031), .B(n15030), .ZN(n15034) );
  NAND2_X1 U18334 ( .A1(n15032), .A2(n19162), .ZN(n15033) );
  OAI211_X1 U18335 ( .C1(n15035), .C2(n19155), .A(n15034), .B(n15033), .ZN(
        P2_U3017) );
  INV_X1 U18336 ( .A(n16004), .ZN(n15040) );
  OAI21_X1 U18337 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n15037), .A(
        n15036), .ZN(n15038) );
  AOI21_X1 U18338 ( .B1(n16005), .B2(n16203), .A(n15038), .ZN(n15039) );
  OAI21_X1 U18339 ( .B1(n15040), .B2(n16184), .A(n15039), .ZN(n15043) );
  NOR2_X1 U18340 ( .A1(n15041), .A2(n16189), .ZN(n15042) );
  AOI211_X1 U18341 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15044), .A(
        n15043), .B(n15042), .ZN(n15045) );
  OAI21_X1 U18342 ( .B1(n15046), .B2(n19155), .A(n15045), .ZN(P2_U3018) );
  OAI21_X1 U18343 ( .B1(n15049), .B2(n15048), .A(n15047), .ZN(n15051) );
  NOR2_X1 U18344 ( .A1(n16184), .A2(n16024), .ZN(n15050) );
  AOI211_X1 U18345 ( .C1(n16018), .C2(n16203), .A(n15051), .B(n15050), .ZN(
        n15053) );
  OAI211_X1 U18346 ( .C1(n15054), .C2(n16189), .A(n15053), .B(n15052), .ZN(
        n15055) );
  INV_X1 U18347 ( .A(n15055), .ZN(n15056) );
  OAI21_X1 U18348 ( .B1(n15057), .B2(n19155), .A(n15056), .ZN(P2_U3019) );
  XNOR2_X1 U18349 ( .A(n15059), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15068) );
  INV_X1 U18350 ( .A(n15078), .ZN(n15067) );
  NAND2_X1 U18351 ( .A1(n15058), .A2(n15083), .ZN(n15074) );
  NOR2_X1 U18352 ( .A1(n15059), .A2(n15074), .ZN(n15060) );
  AOI211_X1 U18353 ( .C1(n19152), .C2(n16026), .A(n15061), .B(n15060), .ZN(
        n15062) );
  OAI21_X1 U18354 ( .B1(n15063), .B2(n19157), .A(n15062), .ZN(n15066) );
  NOR2_X1 U18355 ( .A1(n15064), .A2(n16189), .ZN(n15065) );
  AOI211_X1 U18356 ( .C1(n15068), .C2(n15067), .A(n15066), .B(n15065), .ZN(
        n15069) );
  OAI21_X1 U18357 ( .B1(n15070), .B2(n19155), .A(n15069), .ZN(P2_U3020) );
  NOR3_X1 U18358 ( .A1(n15071), .A2(n9659), .A3(n16189), .ZN(n15080) );
  OAI21_X1 U18359 ( .B1(n15074), .B2(n15073), .A(n15072), .ZN(n15075) );
  AOI21_X1 U18360 ( .B1(n16038), .B2(n16203), .A(n15075), .ZN(n15077) );
  NAND2_X1 U18361 ( .A1(n19152), .A2(n16037), .ZN(n15076) );
  OAI211_X1 U18362 ( .C1(n15078), .C2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15077), .B(n15076), .ZN(n15079) );
  AOI211_X1 U18363 ( .C1(n15081), .C2(n16200), .A(n15080), .B(n15079), .ZN(
        n15082) );
  INV_X1 U18364 ( .A(n15082), .ZN(P2_U3021) );
  OAI21_X1 U18365 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15084), .A(
        n15083), .ZN(n15088) );
  AOI21_X1 U18366 ( .B1(n16203), .B2(n15086), .A(n15085), .ZN(n15087) );
  OAI211_X1 U18367 ( .C1(n16184), .C2(n15089), .A(n15088), .B(n15087), .ZN(
        n15090) );
  AOI21_X1 U18368 ( .B1(n15091), .B2(n19162), .A(n15090), .ZN(n15092) );
  OAI21_X1 U18369 ( .B1(n15093), .B2(n19155), .A(n15092), .ZN(P2_U3022) );
  NAND3_X1 U18370 ( .A1(n15095), .A2(n15094), .A3(n16200), .ZN(n15104) );
  OAI21_X1 U18371 ( .B1(n15096), .B2(n16209), .A(n15257), .ZN(n15115) );
  INV_X1 U18372 ( .A(n15261), .ZN(n15097) );
  NAND2_X1 U18373 ( .A1(n15097), .A2(n15096), .ZN(n15121) );
  AOI221_X1 U18374 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C1(n15099), .C2(n15098), .A(
        n15121), .ZN(n15100) );
  AOI21_X1 U18375 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15115), .A(
        n15100), .ZN(n15101) );
  OAI21_X1 U18376 ( .B1(n18974), .B2(n19763), .A(n15101), .ZN(n15102) );
  AOI21_X1 U18377 ( .B1(n16203), .B2(n16060), .A(n15102), .ZN(n15103) );
  OAI211_X1 U18378 ( .C1(n16184), .C2(n16058), .A(n15104), .B(n15103), .ZN(
        n15105) );
  AOI21_X1 U18379 ( .B1(n19162), .B2(n15106), .A(n15105), .ZN(n15107) );
  INV_X1 U18380 ( .A(n15107), .ZN(P2_U3023) );
  OR2_X1 U18381 ( .A1(n15111), .A2(n15110), .ZN(n15114) );
  AND2_X1 U18382 ( .A1(n15114), .A2(n15113), .ZN(n16097) );
  NOR2_X1 U18383 ( .A1(n12045), .A2(n18974), .ZN(n15117) );
  AND2_X1 U18384 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15115), .ZN(
        n15116) );
  NOR2_X1 U18385 ( .A1(n15117), .A2(n15116), .ZN(n15120) );
  INV_X1 U18386 ( .A(n15118), .ZN(n15519) );
  NAND2_X1 U18387 ( .A1(n19152), .A2(n15519), .ZN(n15119) );
  OAI211_X1 U18388 ( .C1(n15121), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15120), .B(n15119), .ZN(n15127) );
  NAND2_X1 U18389 ( .A1(n15123), .A2(n15122), .ZN(n15125) );
  XOR2_X1 U18390 ( .A(n15125), .B(n15124), .Z(n16094) );
  NOR2_X1 U18391 ( .A1(n16094), .A2(n19155), .ZN(n15126) );
  AOI211_X1 U18392 ( .C1(n16097), .C2(n16203), .A(n15127), .B(n15126), .ZN(
        n15128) );
  OAI21_X1 U18393 ( .B1(n16189), .B2(n16095), .A(n15128), .ZN(P2_U3024) );
  OAI21_X1 U18394 ( .B1(n15129), .B2(n16209), .A(n15257), .ZN(n15133) );
  OR2_X1 U18395 ( .A1(n15261), .A2(n15130), .ZN(n15163) );
  NOR3_X1 U18396 ( .A1(n15163), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15149), .ZN(n15131) );
  AOI211_X1 U18397 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15133), .A(
        n15132), .B(n15131), .ZN(n15136) );
  INV_X1 U18398 ( .A(n15134), .ZN(n18817) );
  NAND2_X1 U18399 ( .A1(n18817), .A2(n16203), .ZN(n15135) );
  OAI211_X1 U18400 ( .C1(n18823), .C2(n16184), .A(n15136), .B(n15135), .ZN(
        n15137) );
  AOI21_X1 U18401 ( .B1(n15138), .B2(n19162), .A(n15137), .ZN(n15139) );
  OAI21_X1 U18402 ( .B1(n15140), .B2(n19155), .A(n15139), .ZN(P2_U3025) );
  NOR2_X1 U18403 ( .A1(n15142), .A2(n15141), .ZN(n15143) );
  OR2_X1 U18404 ( .A1(n15144), .A2(n15143), .ZN(n18824) );
  INV_X1 U18405 ( .A(n15145), .ZN(n15146) );
  AND2_X1 U18406 ( .A1(n19164), .A2(n15146), .ZN(n15147) );
  OR2_X1 U18407 ( .A1(n15148), .A2(n15147), .ZN(n15160) );
  OAI21_X1 U18408 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n15149), .ZN(n15150) );
  OAI22_X1 U18409 ( .A1(n18835), .A2(n19157), .B1(n15150), .B2(n15163), .ZN(
        n15151) );
  AOI211_X1 U18410 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15160), .A(
        n15152), .B(n15151), .ZN(n15153) );
  OAI21_X1 U18411 ( .B1(n18824), .B2(n16184), .A(n15153), .ZN(n15154) );
  AOI21_X1 U18412 ( .B1(n15155), .B2(n16200), .A(n15154), .ZN(n15156) );
  OAI21_X1 U18413 ( .B1(n16189), .B2(n15157), .A(n15156), .ZN(P2_U3026) );
  INV_X1 U18414 ( .A(n15158), .ZN(n18840) );
  AOI21_X1 U18415 ( .B1(n18840), .B2(n16203), .A(n15159), .ZN(n15162) );
  NAND2_X1 U18416 ( .A1(n15160), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15161) );
  OAI211_X1 U18417 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15163), .A(
        n15162), .B(n15161), .ZN(n15164) );
  AOI21_X1 U18418 ( .B1(n18839), .B2(n19152), .A(n15164), .ZN(n15167) );
  NAND2_X1 U18419 ( .A1(n15165), .A2(n16200), .ZN(n15166) );
  OAI211_X1 U18420 ( .C1(n15168), .C2(n16189), .A(n15167), .B(n15166), .ZN(
        P2_U3027) );
  INV_X1 U18421 ( .A(n15169), .ZN(n15170) );
  AOI21_X1 U18422 ( .B1(n15172), .B2(n15171), .A(n15170), .ZN(n18852) );
  INV_X1 U18423 ( .A(n18852), .ZN(n15180) );
  OAI21_X1 U18424 ( .B1(n15177), .B2(n16209), .A(n15201), .ZN(n15175) );
  NOR2_X1 U18425 ( .A1(n18858), .A2(n19157), .ZN(n15173) );
  AOI211_X1 U18426 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15175), .A(
        n15174), .B(n15173), .ZN(n15179) );
  NAND3_X1 U18427 ( .A1(n15204), .A2(n15177), .A3(n15176), .ZN(n15178) );
  OAI211_X1 U18428 ( .C1(n15180), .C2(n16184), .A(n15179), .B(n15178), .ZN(
        n15181) );
  AOI21_X1 U18429 ( .B1(n15182), .B2(n16200), .A(n15181), .ZN(n15183) );
  OAI21_X1 U18430 ( .B1(n15184), .B2(n16189), .A(n15183), .ZN(P2_U3028) );
  INV_X1 U18431 ( .A(n15185), .ZN(n15198) );
  INV_X1 U18432 ( .A(n15187), .ZN(n15188) );
  AOI21_X1 U18433 ( .B1(n10061), .B2(n15188), .A(n9686), .ZN(n19097) );
  OAI21_X1 U18434 ( .B1(n19047), .B2(n19157), .A(n15189), .ZN(n15192) );
  NOR2_X1 U18435 ( .A1(n15190), .A2(n19155), .ZN(n15191) );
  AOI211_X1 U18436 ( .C1(n19152), .C2(n19097), .A(n15192), .B(n15191), .ZN(
        n15196) );
  NOR2_X1 U18437 ( .A1(n15193), .A2(n16189), .ZN(n15194) );
  OAI211_X1 U18438 ( .C1(n15194), .C2(n15204), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n15197), .ZN(n15195) );
  OAI211_X1 U18439 ( .C1(n15198), .C2(n15197), .A(n15196), .B(n15195), .ZN(
        P2_U3030) );
  AOI21_X1 U18440 ( .B1(n18886), .B2(n16203), .A(n15199), .ZN(n15200) );
  OAI21_X1 U18441 ( .B1(n15201), .B2(n15203), .A(n15200), .ZN(n15202) );
  AOI21_X1 U18442 ( .B1(n15204), .B2(n15203), .A(n15202), .ZN(n15205) );
  OAI21_X1 U18443 ( .B1(n18889), .B2(n16184), .A(n15205), .ZN(n15206) );
  AOI21_X1 U18444 ( .B1(n15207), .B2(n16200), .A(n15206), .ZN(n15208) );
  OAI21_X1 U18445 ( .B1(n15209), .B2(n16189), .A(n15208), .ZN(P2_U3031) );
  OR2_X1 U18446 ( .A1(n15261), .A2(n15210), .ZN(n15240) );
  INV_X1 U18447 ( .A(n15240), .ZN(n15224) );
  OAI21_X1 U18448 ( .B1(n16209), .B2(n15211), .A(n15257), .ZN(n15237) );
  AOI21_X1 U18449 ( .B1(n15224), .B2(n15213), .A(n15237), .ZN(n15226) );
  INV_X1 U18450 ( .A(n15212), .ZN(n18895) );
  NAND2_X1 U18451 ( .A1(n18895), .A2(n19152), .ZN(n15218) );
  INV_X1 U18452 ( .A(n19052), .ZN(n15216) );
  NOR3_X1 U18453 ( .A1(n15240), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n15213), .ZN(n15214) );
  AOI211_X1 U18454 ( .C1(n15216), .C2(n16203), .A(n15215), .B(n15214), .ZN(
        n15217) );
  OAI211_X1 U18455 ( .C1(n15226), .C2(n15219), .A(n15218), .B(n15217), .ZN(
        n15220) );
  AOI21_X1 U18456 ( .B1(n15221), .B2(n16200), .A(n15220), .ZN(n15222) );
  OAI21_X1 U18457 ( .B1(n15223), .B2(n16189), .A(n15222), .ZN(P2_U3032) );
  AOI21_X1 U18458 ( .B1(n15224), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15225) );
  NOR2_X1 U18459 ( .A1(n15226), .A2(n15225), .ZN(n15227) );
  AOI211_X1 U18460 ( .C1(n16203), .C2(n18905), .A(n15228), .B(n15227), .ZN(
        n15229) );
  OAI21_X1 U18461 ( .B1(n18909), .B2(n16184), .A(n15229), .ZN(n15230) );
  AOI21_X1 U18462 ( .B1(n15231), .B2(n16200), .A(n15230), .ZN(n15232) );
  OAI21_X1 U18463 ( .B1(n15233), .B2(n16189), .A(n15232), .ZN(P2_U3033) );
  NAND3_X1 U18464 ( .A1(n15235), .A2(n19162), .A3(n15234), .ZN(n15243) );
  AOI21_X1 U18465 ( .B1(n19055), .B2(n16203), .A(n15236), .ZN(n15239) );
  NAND2_X1 U18466 ( .A1(n15237), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15238) );
  OAI211_X1 U18467 ( .C1(n15240), .C2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15239), .B(n15238), .ZN(n15241) );
  AOI21_X1 U18468 ( .B1(n18915), .B2(n19152), .A(n15241), .ZN(n15242) );
  OAI211_X1 U18469 ( .C1(n15244), .C2(n19155), .A(n15243), .B(n15242), .ZN(
        P2_U3034) );
  NOR4_X1 U18470 ( .A1(n15261), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n14587), .A4(n15245), .ZN(n15246) );
  AOI211_X1 U18471 ( .C1(n15248), .C2(n16203), .A(n15247), .B(n15246), .ZN(
        n15251) );
  NOR3_X1 U18472 ( .A1(n15261), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n14587), .ZN(n16162) );
  NAND2_X1 U18473 ( .A1(n19164), .A2(n14587), .ZN(n15249) );
  NAND2_X1 U18474 ( .A1(n15257), .A2(n15249), .ZN(n16166) );
  OAI21_X1 U18475 ( .B1(n16162), .B2(n16166), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15250) );
  OAI211_X1 U18476 ( .C1(n18920), .C2(n16184), .A(n15251), .B(n15250), .ZN(
        n15252) );
  AOI21_X1 U18477 ( .B1(n15253), .B2(n16200), .A(n15252), .ZN(n15254) );
  OAI21_X1 U18478 ( .B1(n15255), .B2(n16189), .A(n15254), .ZN(P2_U3035) );
  INV_X1 U18479 ( .A(n16113), .ZN(n15256) );
  OAI21_X1 U18480 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n14837), .A(
        n15256), .ZN(n16118) );
  INV_X1 U18481 ( .A(n18951), .ZN(n15269) );
  INV_X1 U18482 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19742) );
  NOR2_X1 U18483 ( .A1(n19742), .A2(n18974), .ZN(n15259) );
  NOR2_X1 U18484 ( .A1(n15257), .A2(n14587), .ZN(n15258) );
  AOI211_X1 U18485 ( .C1(n16203), .C2(n18947), .A(n15259), .B(n15258), .ZN(
        n15260) );
  OAI21_X1 U18486 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15261), .A(
        n15260), .ZN(n15268) );
  INV_X1 U18487 ( .A(n16108), .ZN(n15266) );
  NAND2_X1 U18488 ( .A1(n16108), .A2(n15262), .ZN(n15263) );
  NAND2_X1 U18489 ( .A1(n15264), .A2(n15263), .ZN(n15265) );
  OAI21_X1 U18490 ( .B1(n16109), .B2(n15266), .A(n15265), .ZN(n16117) );
  NOR2_X1 U18491 ( .A1(n16117), .A2(n19155), .ZN(n15267) );
  AOI211_X1 U18492 ( .C1(n19152), .C2(n15269), .A(n15268), .B(n15267), .ZN(
        n15270) );
  OAI21_X1 U18493 ( .B1(n16118), .B2(n16189), .A(n15270), .ZN(P2_U3037) );
  NAND2_X1 U18494 ( .A1(n16172), .A2(n10669), .ZN(n16174) );
  INV_X1 U18495 ( .A(n16174), .ZN(n15278) );
  INV_X1 U18496 ( .A(n18968), .ZN(n15271) );
  NAND2_X1 U18497 ( .A1(n15271), .A2(n16203), .ZN(n15276) );
  NOR2_X1 U18498 ( .A1(n15273), .A2(n15272), .ZN(n16175) );
  INV_X1 U18499 ( .A(n16175), .ZN(n15274) );
  AOI22_X1 U18500 ( .A1(n18992), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15274), .ZN(n15275) );
  OAI211_X1 U18501 ( .C1(n16184), .C2(n18969), .A(n15276), .B(n15275), .ZN(
        n15277) );
  AOI211_X1 U18502 ( .C1(n15279), .C2(n16200), .A(n15278), .B(n15277), .ZN(
        n15280) );
  OAI21_X1 U18503 ( .B1(n15281), .B2(n16189), .A(n15280), .ZN(P2_U3039) );
  OAI21_X1 U18504 ( .B1(n15283), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15282), .ZN(n16143) );
  OAI21_X1 U18505 ( .B1(n15285), .B2(n16209), .A(n16194), .ZN(n15292) );
  NAND2_X1 U18506 ( .A1(n15285), .A2(n15284), .ZN(n15290) );
  NAND2_X1 U18507 ( .A1(n18983), .A2(n16203), .ZN(n15289) );
  INV_X1 U18508 ( .A(n18987), .ZN(n15287) );
  NOR2_X1 U18509 ( .A1(n19737), .A2(n18974), .ZN(n15286) );
  AOI21_X1 U18510 ( .B1(n19152), .B2(n15287), .A(n15286), .ZN(n15288) );
  OAI211_X1 U18511 ( .C1(n16196), .C2(n15290), .A(n15289), .B(n15288), .ZN(
        n15291) );
  AOI21_X1 U18512 ( .B1(n15292), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15291), .ZN(n15297) );
  INV_X1 U18513 ( .A(n15293), .ZN(n15295) );
  XNOR2_X1 U18514 ( .A(n15295), .B(n15294), .ZN(n16144) );
  NAND2_X1 U18515 ( .A1(n16144), .A2(n16200), .ZN(n15296) );
  OAI211_X1 U18516 ( .C1(n16143), .C2(n16189), .A(n15297), .B(n15296), .ZN(
        P2_U3040) );
  XNOR2_X1 U18517 ( .A(n15299), .B(n15298), .ZN(n16153) );
  AND2_X1 U18518 ( .A1(n15301), .A2(n15300), .ZN(n15302) );
  OAI22_X1 U18519 ( .A1(n15304), .A2(n15303), .B1(n9713), .B2(n15302), .ZN(
        n16155) );
  INV_X1 U18520 ( .A(n16155), .ZN(n15317) );
  AOI221_X1 U18521 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n13475), .C2(n15308), .A(
        n15305), .ZN(n15316) );
  NAND2_X1 U18522 ( .A1(n18997), .A2(n16203), .ZN(n15314) );
  XNOR2_X1 U18523 ( .A(n15307), .B(n15306), .ZN(n19110) );
  INV_X1 U18524 ( .A(n19110), .ZN(n15312) );
  OAI22_X1 U18525 ( .A1(n18974), .A2(n15310), .B1(n15309), .B2(n15308), .ZN(
        n15311) );
  AOI21_X1 U18526 ( .B1(n19152), .B2(n15312), .A(n15311), .ZN(n15313) );
  NAND2_X1 U18527 ( .A1(n15314), .A2(n15313), .ZN(n15315) );
  AOI211_X1 U18528 ( .C1(n15317), .C2(n19162), .A(n15316), .B(n15315), .ZN(
        n15318) );
  OAI21_X1 U18529 ( .B1(n19155), .B2(n16153), .A(n15318), .ZN(P2_U3041) );
  INV_X1 U18530 ( .A(n15319), .ZN(n15323) );
  AOI22_X1 U18531 ( .A1(n15366), .A2(n15321), .B1(n19702), .B2(n15320), .ZN(
        n15322) );
  OAI21_X1 U18532 ( .B1(n15324), .B2(n15323), .A(n15322), .ZN(n15325) );
  MUX2_X1 U18533 ( .A(n15325), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n19792), .Z(P2_U3599) );
  OAI21_X1 U18534 ( .B1(n19693), .B2(n19194), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n15326) );
  NAND2_X1 U18535 ( .A1(n15326), .A2(n19806), .ZN(n15328) );
  NAND2_X1 U18536 ( .A1(n19805), .A2(n19813), .ZN(n19245) );
  NOR2_X1 U18537 ( .A1(n19405), .A2(n19245), .ZN(n19190) );
  INV_X1 U18538 ( .A(n19190), .ZN(n15346) );
  AND2_X1 U18539 ( .A1(n19660), .A2(n15346), .ZN(n15331) );
  OAI21_X1 U18540 ( .B1(n15329), .B2(n19190), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15327) );
  INV_X1 U18541 ( .A(n15328), .ZN(n15332) );
  AOI211_X1 U18542 ( .C1(n15329), .C2(n19587), .A(n19190), .B(n19806), .ZN(
        n15330) );
  INV_X1 U18543 ( .A(n19199), .ZN(n15333) );
  NAND2_X1 U18544 ( .A1(n15333), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n15335) );
  AOI22_X1 U18545 ( .A1(n19521), .A2(n19693), .B1(n19586), .B2(n19190), .ZN(
        n15334) );
  OAI211_X1 U18546 ( .C1(n19524), .C2(n19225), .A(n15335), .B(n15334), .ZN(
        n15336) );
  AOI21_X1 U18547 ( .B1(n13539), .B2(n19195), .A(n15336), .ZN(n15337) );
  INV_X1 U18548 ( .A(n15337), .ZN(P2_U3048) );
  INV_X1 U18549 ( .A(n19189), .ZN(n19172) );
  NAND2_X1 U18550 ( .A1(n19172), .A2(n15338), .ZN(n19651) );
  AOI22_X1 U18551 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19193), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19192), .ZN(n19527) );
  OAI22_X1 U18552 ( .A1(n19651), .A2(n15346), .B1(n19527), .B2(n19225), .ZN(
        n15339) );
  AOI21_X1 U18553 ( .B1(n19654), .B2(n19693), .A(n15339), .ZN(n15343) );
  NAND2_X1 U18554 ( .A1(n19195), .A2(n15341), .ZN(n15342) );
  OAI211_X1 U18555 ( .C1(n19199), .C2(n15344), .A(n15343), .B(n15342), .ZN(
        P2_U3049) );
  AOI22_X1 U18556 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19193), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19192), .ZN(n19623) );
  INV_X1 U18557 ( .A(n19623), .ZN(n19694) );
  NOR2_X1 U18558 ( .A1(n19189), .A2(n15345), .ZN(n19688) );
  INV_X1 U18559 ( .A(n19688), .ZN(n19472) );
  AOI22_X1 U18560 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19193), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19192), .ZN(n19549) );
  OAI22_X1 U18561 ( .A1(n19472), .A2(n15346), .B1(n19549), .B2(n19225), .ZN(
        n15347) );
  AOI21_X1 U18562 ( .B1(n19693), .B2(n19694), .A(n15347), .ZN(n15350) );
  NOR2_X2 U18563 ( .A1(n15348), .A2(n19285), .ZN(n19690) );
  NAND2_X1 U18564 ( .A1(n19195), .A2(n19690), .ZN(n15349) );
  OAI211_X1 U18565 ( .C1(n19199), .C2(n15351), .A(n15350), .B(n15349), .ZN(
        P2_U3055) );
  INV_X1 U18566 ( .A(n15352), .ZN(n15357) );
  NOR3_X2 U18567 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19821), .A3(
        n19245), .ZN(n19238) );
  AOI21_X1 U18568 ( .B1(n15357), .B2(n19587), .A(n19238), .ZN(n15355) );
  NAND2_X1 U18569 ( .A1(n19791), .A2(n19036), .ZN(n19375) );
  NOR2_X2 U18570 ( .A1(n19442), .A2(n19375), .ZN(n19240) );
  NOR2_X1 U18571 ( .A1(n19481), .A2(n19245), .ZN(n15353) );
  AOI221_X1 U18572 ( .B1(n19255), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19240), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n15353), .ZN(n15354) );
  MUX2_X1 U18573 ( .A(n15355), .B(n15354), .S(n19806), .Z(n15356) );
  INV_X1 U18574 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15362) );
  AOI22_X1 U18575 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19193), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19192), .ZN(n19536) );
  AOI22_X1 U18576 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19192), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19193), .ZN(n19610) );
  INV_X1 U18577 ( .A(n19610), .ZN(n19672) );
  AOI22_X1 U18578 ( .A1(n19255), .A2(n19673), .B1(n19240), .B2(n19672), .ZN(
        n15361) );
  OAI21_X1 U18579 ( .B1(n15357), .B2(n19238), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15358) );
  OAI21_X1 U18580 ( .B1(n19245), .B2(n19481), .A(n15358), .ZN(n19239) );
  NOR2_X2 U18581 ( .A1(n16081), .A2(n19285), .ZN(n19671) );
  NOR2_X2 U18582 ( .A1(n19189), .A2(n15359), .ZN(n19670) );
  AOI22_X1 U18583 ( .A1(n19239), .A2(n19671), .B1(n19670), .B2(n19238), .ZN(
        n15360) );
  OAI211_X1 U18584 ( .C1(n19243), .C2(n15362), .A(n15361), .B(n15360), .ZN(
        P2_U3068) );
  INV_X1 U18585 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15365) );
  INV_X1 U18586 ( .A(n19549), .ZN(n19692) );
  AOI22_X1 U18587 ( .A1(n19240), .A2(n19694), .B1(n19255), .B2(n19692), .ZN(
        n15364) );
  AOI22_X1 U18588 ( .A1(n19239), .A2(n19690), .B1(n19238), .B2(n19688), .ZN(
        n15363) );
  OAI211_X1 U18589 ( .C1(n19243), .C2(n15365), .A(n15364), .B(n15363), .ZN(
        P2_U3071) );
  NOR3_X1 U18590 ( .A1(n19813), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19321) );
  INV_X1 U18591 ( .A(n19321), .ZN(n19326) );
  NOR2_X1 U18592 ( .A1(n19830), .A2(n19326), .ZN(n19346) );
  AOI21_X1 U18593 ( .B1(n19368), .B2(n19397), .A(n19797), .ZN(n15368) );
  NOR2_X1 U18594 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15367), .ZN(
        n19383) );
  INV_X1 U18595 ( .A(n19383), .ZN(n19379) );
  NOR2_X1 U18596 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19379), .ZN(
        n19369) );
  AOI221_X1 U18597 ( .B1(n19346), .B2(n19587), .C1(n15368), .C2(n19587), .A(
        n19369), .ZN(n15369) );
  NOR3_X1 U18598 ( .A1(n10509), .A2(n19369), .A3(n19843), .ZN(n15371) );
  INV_X1 U18599 ( .A(n19372), .ZN(n15376) );
  INV_X1 U18600 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15375) );
  INV_X1 U18601 ( .A(n19368), .ZN(n19371) );
  AOI22_X1 U18602 ( .A1(n19401), .A2(n19595), .B1(n19371), .B2(n19521), .ZN(
        n15374) );
  NOR2_X1 U18603 ( .A1(n19346), .A2(n19369), .ZN(n15370) );
  OR2_X1 U18604 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n15370), .ZN(n15372) );
  AOI21_X1 U18605 ( .B1(n19843), .B2(n15372), .A(n15371), .ZN(n19370) );
  AOI22_X1 U18606 ( .A1(n19370), .A2(n13539), .B1(n19586), .B2(n19369), .ZN(
        n15373) );
  OAI211_X1 U18607 ( .C1(n15376), .C2(n15375), .A(n15374), .B(n15373), .ZN(
        P2_U3096) );
  OAI21_X1 U18608 ( .B1(n19695), .B2(n19645), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n15377) );
  NAND2_X1 U18609 ( .A1(n15377), .A2(n19806), .ZN(n15380) );
  NOR2_X1 U18610 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15378), .ZN(
        n19644) );
  NAND3_X1 U18611 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19821), .ZN(n19589) );
  NOR2_X1 U18612 ( .A1(n19830), .A2(n19589), .ZN(n19617) );
  NOR2_X1 U18613 ( .A1(n19644), .A2(n19617), .ZN(n15383) );
  OAI21_X1 U18614 ( .B1(n15381), .B2(n19644), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15379) );
  INV_X1 U18615 ( .A(n19695), .ZN(n15390) );
  INV_X1 U18616 ( .A(n15380), .ZN(n15384) );
  AOI211_X1 U18617 ( .C1(n15381), .C2(n19587), .A(n19644), .B(n19806), .ZN(
        n15382) );
  AOI211_X2 U18618 ( .C1(n15384), .C2(n15383), .A(n15382), .B(n19285), .ZN(
        n19650) );
  INV_X1 U18619 ( .A(n19650), .ZN(n15392) );
  NAND2_X1 U18620 ( .A1(n15392), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n15386) );
  AOI22_X1 U18621 ( .A1(n19521), .A2(n19645), .B1(n19586), .B2(n19644), .ZN(
        n15385) );
  OAI211_X1 U18622 ( .C1(n19524), .C2(n15390), .A(n15386), .B(n15385), .ZN(
        n15387) );
  AOI21_X1 U18623 ( .B1(n13539), .B2(n19646), .A(n15387), .ZN(n15388) );
  INV_X1 U18624 ( .A(n15388), .ZN(P2_U3160) );
  INV_X1 U18625 ( .A(n19646), .ZN(n15395) );
  INV_X1 U18626 ( .A(n19690), .ZN(n15394) );
  AOI22_X1 U18627 ( .A1(n19645), .A2(n19694), .B1(n19688), .B2(n19644), .ZN(
        n15389) );
  OAI21_X1 U18628 ( .B1(n15390), .B2(n19549), .A(n15389), .ZN(n15391) );
  AOI21_X1 U18629 ( .B1(n15392), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n15391), .ZN(n15393) );
  OAI21_X1 U18630 ( .B1(n15395), .B2(n15394), .A(n15393), .ZN(P2_U3167) );
  NOR3_X1 U18631 ( .A1(n18158), .A2(n18143), .A3(n15396), .ZN(n15398) );
  AOI22_X1 U18632 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15400) );
  OAI21_X1 U18633 ( .B1(n10169), .B2(n17019), .A(n15400), .ZN(n15411) );
  INV_X1 U18634 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15409) );
  AOI22_X1 U18635 ( .A1(n17096), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15408) );
  INV_X1 U18636 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15402) );
  AOI22_X1 U18637 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15401) );
  OAI21_X1 U18638 ( .B1(n17005), .B2(n15402), .A(n15401), .ZN(n15406) );
  AOI22_X1 U18639 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16972), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15404) );
  AOI22_X1 U18640 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15403) );
  OAI211_X1 U18641 ( .C1(n17100), .C2(n16889), .A(n15404), .B(n15403), .ZN(
        n15405) );
  OAI211_X1 U18642 ( .C1(n12454), .C2(n15409), .A(n15408), .B(n15407), .ZN(
        n15410) );
  AOI211_X1 U18643 ( .C1(n17101), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n15411), .B(n15410), .ZN(n16837) );
  AOI22_X1 U18644 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15412) );
  OAI21_X1 U18645 ( .B1(n12420), .B2(n16919), .A(n15412), .ZN(n15421) );
  AOI22_X1 U18646 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15419) );
  OAI22_X1 U18647 ( .A1(n16918), .A2(n17038), .B1(n12454), .B2(n17063), .ZN(
        n15417) );
  AOI22_X1 U18648 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17115), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15415) );
  AOI22_X1 U18649 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15414) );
  AOI22_X1 U18650 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15413) );
  NAND3_X1 U18651 ( .A1(n15415), .A2(n15414), .A3(n15413), .ZN(n15416) );
  AOI211_X1 U18652 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n15417), .B(n15416), .ZN(n15418) );
  OAI211_X1 U18653 ( .C1(n10169), .C2(n17054), .A(n15419), .B(n15418), .ZN(
        n15420) );
  AOI211_X1 U18654 ( .C1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .C2(n17102), .A(
        n15421), .B(n15420), .ZN(n16845) );
  AOI22_X1 U18655 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15422) );
  OAI21_X1 U18656 ( .B1(n12445), .B2(n17105), .A(n15422), .ZN(n15433) );
  INV_X1 U18657 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15431) );
  AOI22_X1 U18658 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16906), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15430) );
  OAI22_X1 U18659 ( .A1(n17100), .A2(n15423), .B1(n17005), .B2(n17094), .ZN(
        n15428) );
  AOI22_X1 U18660 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15426) );
  AOI22_X1 U18661 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17101), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15425) );
  AOI22_X1 U18662 ( .A1(n16949), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15424) );
  NAND3_X1 U18663 ( .A1(n15426), .A2(n15425), .A3(n15424), .ZN(n15427) );
  AOI211_X1 U18664 ( .C1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .C2(n17074), .A(
        n15428), .B(n15427), .ZN(n15429) );
  OAI211_X1 U18665 ( .C1(n9596), .C2(n15431), .A(n15430), .B(n15429), .ZN(
        n15432) );
  AOI211_X1 U18666 ( .C1(n12442), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n15433), .B(n15432), .ZN(n16853) );
  AOI22_X1 U18667 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n17078), .ZN(n15434) );
  OAI21_X1 U18668 ( .B1(n10165), .B2(n15435), .A(n15434), .ZN(n15444) );
  AOI22_X1 U18669 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17096), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15442) );
  AOI22_X1 U18670 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17074), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15436) );
  OAI21_X1 U18671 ( .B1(n16968), .B2(n17106), .A(n15436), .ZN(n15440) );
  INV_X1 U18672 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U18673 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17070), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17095), .ZN(n15438) );
  AOI22_X1 U18674 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15437) );
  OAI211_X1 U18675 ( .C1(n16971), .C2(n17038), .A(n15438), .B(n15437), .ZN(
        n15439) );
  AOI211_X1 U18676 ( .C1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .C2(n12486), .A(
        n15440), .B(n15439), .ZN(n15441) );
  OAI211_X1 U18677 ( .C1(n17119), .C2(n17077), .A(n15442), .B(n15441), .ZN(
        n15443) );
  AOI211_X1 U18678 ( .C1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .C2(n17115), .A(
        n15444), .B(n15443), .ZN(n16854) );
  NOR2_X1 U18679 ( .A1(n16853), .A2(n16854), .ZN(n16852) );
  AOI22_X1 U18680 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n16972), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15455) );
  AOI22_X1 U18681 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15454) );
  AOI22_X1 U18682 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15453) );
  OAI22_X1 U18683 ( .A1(n9596), .A2(n17072), .B1(n12454), .B2(n15445), .ZN(
        n15451) );
  AOI22_X1 U18684 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15449) );
  AOI22_X1 U18685 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15448) );
  AOI22_X1 U18686 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15447) );
  NAND2_X1 U18687 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n15446) );
  NAND4_X1 U18688 ( .A1(n15449), .A2(n15448), .A3(n15447), .A4(n15446), .ZN(
        n15450) );
  AOI211_X1 U18689 ( .C1(n17096), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n15451), .B(n15450), .ZN(n15452) );
  NAND4_X1 U18690 ( .A1(n15455), .A2(n15454), .A3(n15453), .A4(n15452), .ZN(
        n16849) );
  NAND2_X1 U18691 ( .A1(n16852), .A2(n16849), .ZN(n16848) );
  NOR2_X1 U18692 ( .A1(n16845), .A2(n16848), .ZN(n17177) );
  AOI22_X1 U18693 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17101), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15467) );
  AOI22_X1 U18694 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17096), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15466) );
  OAI22_X1 U18695 ( .A1(n12445), .A2(n17134), .B1(n12454), .B2(n15456), .ZN(
        n15464) );
  AOI22_X1 U18696 ( .A1(n16949), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15462) );
  AOI22_X1 U18697 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17115), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15458) );
  AOI22_X1 U18698 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15457) );
  OAI211_X1 U18699 ( .C1(n17005), .C2(n15459), .A(n15458), .B(n15457), .ZN(
        n15460) );
  AOI21_X1 U18700 ( .B1(n17060), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n15460), .ZN(n15461) );
  OAI211_X1 U18701 ( .C1(n17077), .C2(n17037), .A(n15462), .B(n15461), .ZN(
        n15463) );
  AOI211_X1 U18702 ( .C1(n16812), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n15464), .B(n15463), .ZN(n15465) );
  NAND3_X1 U18703 ( .A1(n15467), .A2(n15466), .A3(n15465), .ZN(n17176) );
  NAND2_X1 U18704 ( .A1(n17177), .A2(n17176), .ZN(n17175) );
  NOR2_X1 U18705 ( .A1(n16837), .A2(n17175), .ZN(n16836) );
  INV_X1 U18706 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17004) );
  AOI22_X1 U18707 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15478) );
  INV_X1 U18708 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15470) );
  AOI22_X1 U18709 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15469) );
  AOI22_X1 U18710 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15468) );
  OAI211_X1 U18711 ( .C1(n17005), .C2(n15470), .A(n15469), .B(n15468), .ZN(
        n15476) );
  AOI22_X1 U18712 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16906), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15474) );
  AOI22_X1 U18713 ( .A1(n12405), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15473) );
  AOI22_X1 U18714 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15472) );
  NAND2_X1 U18715 ( .A1(n9600), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n15471) );
  NAND4_X1 U18716 ( .A1(n15474), .A2(n15473), .A3(n15472), .A4(n15471), .ZN(
        n15475) );
  AOI211_X1 U18717 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n15476), .B(n15475), .ZN(n15477) );
  OAI211_X1 U18718 ( .C1(n10165), .C2(n17004), .A(n15478), .B(n15477), .ZN(
        n15479) );
  NAND2_X1 U18719 ( .A1(n16836), .A2(n15479), .ZN(n16828) );
  OAI21_X1 U18720 ( .B1(n16836), .B2(n15479), .A(n16828), .ZN(n17169) );
  AND2_X1 U18721 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16832) );
  NAND2_X1 U18722 ( .A1(n17199), .A2(n17143), .ZN(n17149) );
  INV_X1 U18723 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16902) );
  INV_X1 U18724 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16930) );
  INV_X1 U18725 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16999) );
  INV_X1 U18726 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17067) );
  INV_X1 U18727 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n16707) );
  INV_X1 U18728 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16728) );
  INV_X1 U18729 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17132) );
  NAND2_X1 U18730 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16780) );
  INV_X1 U18731 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16855) );
  INV_X1 U18732 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16519) );
  INV_X1 U18733 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16887) );
  NOR3_X1 U18734 ( .A1(n16855), .A2(n16519), .A3(n16887), .ZN(n16841) );
  AND4_X1 U18735 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(n16841), .ZN(n16833) );
  NAND2_X1 U18736 ( .A1(n16885), .A2(n16833), .ZN(n15480) );
  NAND2_X1 U18737 ( .A1(n17139), .A2(n15480), .ZN(n16843) );
  OAI21_X1 U18738 ( .B1(n16832), .B2(n17149), .A(n16843), .ZN(n16830) );
  INV_X1 U18739 ( .A(n15480), .ZN(n16838) );
  INV_X1 U18740 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16840) );
  NOR2_X1 U18741 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16840), .ZN(n15481) );
  AOI22_X1 U18742 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16830), .B1(n16838), 
        .B2(n15481), .ZN(n15482) );
  OAI21_X1 U18743 ( .B1(n17139), .B2(n17169), .A(n15482), .ZN(P3_U2675) );
  NOR2_X1 U18744 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18743), .ZN(
        n18386) );
  NAND3_X1 U18745 ( .A1(n17077), .A2(n15483), .A3(n18607), .ZN(n18113) );
  AOI221_X1 U18746 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n18623), .C1(n18113), .C2(
        n18623), .A(n18410), .ZN(n15484) );
  NOR2_X1 U18747 ( .A1(n18386), .A2(n15484), .ZN(n15486) );
  INV_X1 U18748 ( .A(n15484), .ZN(n18119) );
  INV_X1 U18749 ( .A(n17728), .ZN(n17600) );
  OAI22_X1 U18750 ( .A1(n17600), .A2(n18770), .B1(n18589), .B2(n18743), .ZN(
        n15489) );
  NAND3_X1 U18751 ( .A1(n18591), .A2(n18119), .A3(n15489), .ZN(n15485) );
  OAI221_X1 U18752 ( .B1(n18591), .B2(n15486), .C1(n18591), .C2(n18408), .A(
        n15485), .ZN(P3_U2864) );
  NAND2_X1 U18753 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18272) );
  NOR2_X1 U18754 ( .A1(n17600), .A2(n18770), .ZN(n15488) );
  INV_X1 U18755 ( .A(n15486), .ZN(n15487) );
  AOI221_X1 U18756 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18272), .C1(n15488), 
        .C2(n18272), .A(n15487), .ZN(n18118) );
  INV_X1 U18757 ( .A(n18408), .ZN(n18123) );
  OAI221_X1 U18758 ( .B1(n18123), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18123), .C2(n15489), .A(n18119), .ZN(n18116) );
  AOI22_X1 U18759 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18118), .B1(
        n18116), .B2(n18596), .ZN(P3_U2865) );
  INV_X1 U18760 ( .A(n19792), .ZN(n19794) );
  NAND3_X1 U18761 ( .A1(n19852), .A2(n19702), .A3(n15490), .ZN(n15491) );
  OR3_X1 U18762 ( .A1(n19792), .A2(n15492), .A3(n15491), .ZN(n15493) );
  OAI21_X1 U18763 ( .B1(n19794), .B2(n15494), .A(n15493), .ZN(P2_U3595) );
  NAND2_X1 U18764 ( .A1(n9932), .A2(n18585), .ZN(n17959) );
  INV_X1 U18765 ( .A(n17959), .ZN(n17993) );
  INV_X1 U18766 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18045) );
  NOR3_X1 U18767 ( .A1(n18065), .A2(n18045), .A3(n17715), .ZN(n17893) );
  NAND3_X1 U18768 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n17893), .ZN(n18013) );
  NAND3_X1 U18769 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17951) );
  NOR2_X1 U18770 ( .A1(n18013), .A2(n17951), .ZN(n17991) );
  NAND2_X1 U18771 ( .A1(n17894), .A2(n17991), .ZN(n17934) );
  NOR2_X1 U18772 ( .A1(n17895), .A2(n17934), .ZN(n17884) );
  NAND2_X1 U18773 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17884), .ZN(
        n17909) );
  NOR2_X1 U18774 ( .A1(n15495), .A2(n17909), .ZN(n17777) );
  NAND3_X1 U18775 ( .A1(n16268), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17777), .ZN(n15498) );
  AOI21_X1 U18776 ( .B1(n16257), .B2(n17884), .A(n18585), .ZN(n15497) );
  AOI21_X1 U18777 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17892) );
  INV_X1 U18778 ( .A(n17892), .ZN(n18072) );
  NAND2_X1 U18779 ( .A1(n17893), .A2(n18072), .ZN(n18014) );
  NOR2_X1 U18780 ( .A1(n17951), .A2(n18014), .ZN(n17956) );
  NAND2_X1 U18781 ( .A1(n17606), .A2(n17956), .ZN(n17935) );
  NOR2_X1 U18782 ( .A1(n15496), .A2(n17935), .ZN(n17840) );
  AOI21_X1 U18783 ( .B1(n16257), .B2(n17840), .A(n9932), .ZN(n17786) );
  AOI211_X1 U18784 ( .C1(n18583), .C2(n15498), .A(n15497), .B(n17786), .ZN(
        n15576) );
  OAI21_X1 U18785 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17993), .A(
        n15576), .ZN(n16273) );
  AOI21_X1 U18786 ( .B1(n15500), .B2(n15499), .A(n18548), .ZN(n15509) );
  INV_X1 U18787 ( .A(n15501), .ZN(n15507) );
  AOI21_X1 U18788 ( .B1(n17348), .B2(n18132), .A(n18762), .ZN(n15503) );
  AOI21_X1 U18789 ( .B1(n15503), .B2(n15502), .A(n18764), .ZN(n16380) );
  NAND3_X1 U18790 ( .A1(n16380), .A2(n15504), .A3(n18551), .ZN(n15505) );
  OAI21_X1 U18791 ( .B1(n9622), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18101), .ZN(n15510) );
  NOR2_X1 U18792 ( .A1(n16239), .A2(n16254), .ZN(n16240) );
  NAND2_X1 U18793 ( .A1(n17276), .A2(n18050), .ZN(n18027) );
  OAI22_X1 U18794 ( .A1(n16236), .A2(n18110), .B1(n16240), .B2(n18027), .ZN(
        n15577) );
  AOI221_X1 U18795 ( .B1(n16273), .B2(n17988), .C1(n15510), .C2(n17988), .A(
        n15577), .ZN(n15517) );
  NOR3_X4 U18796 ( .A1(n17276), .A2(n18555), .A3(n18016), .ZN(n18009) );
  NOR2_X1 U18797 ( .A1(n15512), .A2(n15511), .ZN(n15513) );
  XOR2_X1 U18798 ( .A(n15513), .B(n16242), .Z(n16245) );
  AOI21_X1 U18799 ( .B1(n18583), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18559), .ZN(n18073) );
  INV_X1 U18800 ( .A(n18073), .ZN(n15514) );
  AOI22_X1 U18801 ( .A1(n18581), .A2(n17840), .B1(n15514), .B2(n17884), .ZN(
        n17808) );
  INV_X1 U18802 ( .A(n18555), .ZN(n15515) );
  NAND2_X1 U18803 ( .A1(n17276), .A2(n15515), .ZN(n17846) );
  INV_X1 U18804 ( .A(n17846), .ZN(n17976) );
  AOI22_X1 U18805 ( .A1(n18549), .A2(n17845), .B1(n17847), .B2(n17976), .ZN(
        n17896) );
  NAND2_X1 U18806 ( .A1(n17808), .A2(n17896), .ZN(n17850) );
  NAND3_X1 U18807 ( .A1(n16268), .A2(n17833), .A3(n17850), .ZN(n17776) );
  NOR3_X1 U18808 ( .A1(n16238), .A2(n18016), .A3(n17776), .ZN(n15574) );
  AOI22_X1 U18809 ( .A1(n18009), .A2(n16245), .B1(n15574), .B2(n16242), .ZN(
        n15516) );
  NAND2_X1 U18810 ( .A1(n9611), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16252) );
  OAI211_X1 U18811 ( .C1(n15517), .C2(n16242), .A(n15516), .B(n16252), .ZN(
        P3_U2833) );
  AOI22_X1 U18812 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19027), .B1(n15518), 
        .B2(n19026), .ZN(n15525) );
  AOI22_X1 U18813 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19038), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n19028), .ZN(n15524) );
  AOI22_X1 U18814 ( .A1(n19008), .A2(n15519), .B1(n18998), .B2(n16097), .ZN(
        n15523) );
  OAI211_X1 U18815 ( .C1(n16101), .C2(n15521), .A(n19000), .B(n15520), .ZN(
        n15522) );
  NAND4_X1 U18816 ( .A1(n15525), .A2(n15524), .A3(n15523), .A4(n15522), .ZN(
        P2_U2833) );
  INV_X1 U18817 ( .A(n15534), .ZN(n15537) );
  NOR3_X1 U18818 ( .A1(n15527), .A2(n15526), .A3(n20611), .ZN(n15531) );
  OR2_X1 U18819 ( .A1(n15529), .A2(n15528), .ZN(n15530) );
  AOI222_X1 U18820 ( .A1(n15531), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .B1(n15531), .B2(n15530), .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C2(n15530), .ZN(n15535) );
  AND2_X1 U18821 ( .A1(n20429), .A2(n15535), .ZN(n15533) );
  OAI222_X1 U18822 ( .A1(n20429), .A2(n15535), .B1(n20234), .B2(n15534), .C1(
        n15533), .C2(n15532), .ZN(n15536) );
  OAI21_X1 U18823 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15537), .A(
        n15536), .ZN(n15545) );
  OAI21_X1 U18824 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15538), .ZN(n15539) );
  NAND4_X1 U18825 ( .A1(n15542), .A2(n15541), .A3(n15540), .A4(n15539), .ZN(
        n15543) );
  AOI211_X1 U18826 ( .C1(n15545), .C2(n20138), .A(n15544), .B(n15543), .ZN(
        n15561) );
  INV_X1 U18827 ( .A(n15561), .ZN(n15552) );
  NOR3_X1 U18828 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11268), .A3(n20769), 
        .ZN(n15550) );
  NAND4_X1 U18829 ( .A1(n12849), .A2(n15548), .A3(n15547), .A4(n15546), .ZN(
        n15549) );
  OAI21_X1 U18830 ( .B1(n15551), .B2(n15550), .A(n15549), .ZN(n15974) );
  AOI221_X1 U18831 ( .B1(n20754), .B2(n20753), .C1(n15552), .C2(n20753), .A(
        n15974), .ZN(n15979) );
  AND2_X1 U18832 ( .A1(n15553), .A2(n15555), .ZN(n15554) );
  NOR2_X1 U18833 ( .A1(n15979), .A2(n15554), .ZN(n15559) );
  AOI211_X1 U18834 ( .C1(n20851), .C2(n11268), .A(n15556), .B(n15555), .ZN(
        n15557) );
  NAND2_X1 U18835 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15557), .ZN(n15558) );
  OAI22_X1 U18836 ( .A1(n15559), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n15979), 
        .B2(n15558), .ZN(n15560) );
  OAI21_X1 U18837 ( .B1(n15561), .B2(n19870), .A(n15560), .ZN(P1_U3161) );
  NAND2_X1 U18838 ( .A1(n20128), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n15570) );
  NAND3_X1 U18839 ( .A1(n15568), .A2(n15567), .A3(n15566), .ZN(n15569) );
  NAND2_X1 U18840 ( .A1(n15572), .A2(n15571), .ZN(n15573) );
  XOR2_X1 U18841 ( .A(n15573), .B(n16255), .Z(n16234) );
  NOR2_X1 U18842 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16254), .ZN(
        n16230) );
  AOI22_X1 U18843 ( .A1(n9611), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n16230), 
        .B2(n15574), .ZN(n15579) );
  NOR2_X1 U18844 ( .A1(n18581), .A2(n18583), .ZN(n17938) );
  AOI21_X1 U18845 ( .B1(n18585), .B2(n17938), .A(n18016), .ZN(n16258) );
  AOI21_X1 U18846 ( .B1(n16254), .B2(n16258), .A(n18092), .ZN(n15575) );
  OAI21_X1 U18847 ( .B1(n15576), .B2(n18016), .A(n15575), .ZN(n16263) );
  OAI21_X1 U18848 ( .B1(n16263), .B2(n15577), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15578) );
  OAI211_X1 U18849 ( .C1(n16234), .C2(n18021), .A(n15579), .B(n15578), .ZN(
        P3_U2832) );
  INV_X1 U18850 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20775) );
  INV_X1 U18851 ( .A(HOLD), .ZN(n20761) );
  NOR2_X1 U18852 ( .A1(n20775), .A2(n20761), .ZN(n15581) );
  AOI22_X1 U18853 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15580) );
  NAND2_X1 U18854 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20851), .ZN(n20760) );
  OAI211_X1 U18855 ( .C1(n15581), .C2(n15580), .A(n15584), .B(n20760), .ZN(
        P1_U3195) );
  NAND2_X1 U18856 ( .A1(n15583), .A2(n15582), .ZN(n15587) );
  NOR2_X1 U18857 ( .A1(n15585), .A2(n15584), .ZN(n15586) );
  NAND2_X1 U18858 ( .A1(n20754), .A2(n15975), .ZN(n20850) );
  INV_X2 U18859 ( .A(n20850), .ZN(n20036) );
  AND2_X1 U18860 ( .A1(n20022), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NAND2_X1 U18861 ( .A1(n15884), .A2(n15588), .ZN(n15877) );
  NOR3_X1 U18862 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15884), .A3(
        n15589), .ZN(n15594) );
  NAND2_X1 U18863 ( .A1(n15591), .A2(n15590), .ZN(n15592) );
  XOR2_X1 U18864 ( .A(n15592), .B(n15596), .Z(n15785) );
  OAI22_X1 U18865 ( .A1(n15785), .A2(n20120), .B1(n20116), .B2(n15667), .ZN(
        n15593) );
  AOI211_X1 U18866 ( .C1(P1_REIP_REG_20__SCAN_IN), .C2(n20128), .A(n15594), 
        .B(n15593), .ZN(n15595) );
  OAI221_X1 U18867 ( .B1(n15596), .B2(n9630), .C1(n15596), .C2(n15877), .A(
        n15595), .ZN(P1_U3011) );
  NOR2_X1 U18868 ( .A1(n19845), .A2(n19855), .ZN(n19701) );
  NAND2_X1 U18869 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATEBS16_REG_SCAN_IN), .ZN(n19814) );
  OAI21_X1 U18870 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n19814), .A(n19843), 
        .ZN(n15597) );
  AOI21_X1 U18871 ( .B1(n19701), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n15597), 
        .ZN(n15598) );
  NOR2_X1 U18872 ( .A1(n16221), .A2(n15598), .ZN(P2_U3178) );
  OAI221_X1 U18873 ( .B1(n10339), .B2(n15599), .C1(n16220), .C2(n15599), .A(
        n19285), .ZN(n19831) );
  NOR2_X1 U18874 ( .A1(n15600), .A2(n19831), .ZN(P2_U3047) );
  NAND2_X1 U18875 ( .A1(n15605), .A2(n17150), .ZN(n17300) );
  AOI22_X1 U18876 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17306), .B1(
        P3_EAX_REG_0__SCAN_IN), .B2(n17152), .ZN(n15606) );
  NOR2_X1 U18877 ( .A1(n18158), .A2(n17152), .ZN(n17301) );
  INV_X1 U18878 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17381) );
  NAND2_X1 U18879 ( .A1(n17301), .A2(n17381), .ZN(n17303) );
  OAI211_X1 U18880 ( .C1(n17769), .C2(n17308), .A(n15606), .B(n17303), .ZN(
        P3_U2735) );
  INV_X1 U18881 ( .A(n15607), .ZN(n15611) );
  NOR3_X1 U18882 ( .A1(n15626), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n15625), 
        .ZN(n15610) );
  INV_X1 U18883 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15608) );
  NOR2_X1 U18884 ( .A1(n19913), .A2(n15608), .ZN(n15609) );
  AOI211_X1 U18885 ( .C1(n19961), .C2(n15611), .A(n15610), .B(n15609), .ZN(
        n15613) );
  NAND2_X1 U18886 ( .A1(n19937), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n15612) );
  OAI211_X1 U18887 ( .C1(n15627), .C2(n20815), .A(n15613), .B(n15612), .ZN(
        n15614) );
  AOI21_X1 U18888 ( .B1(n15744), .B2(n19905), .A(n15614), .ZN(n15615) );
  OAI21_X1 U18889 ( .B1(n15616), .B2(n19952), .A(n15615), .ZN(P1_U2811) );
  INV_X1 U18890 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15618) );
  OAI22_X1 U18891 ( .A1(n15618), .A2(n19913), .B1(n19948), .B2(n15617), .ZN(
        n15619) );
  AOI21_X1 U18892 ( .B1(n19937), .B2(P1_EBX_REG_28__SCAN_IN), .A(n15619), .ZN(
        n15620) );
  OAI21_X1 U18893 ( .B1(n15621), .B2(n19952), .A(n15620), .ZN(n15622) );
  AOI21_X1 U18894 ( .B1(n15623), .B2(n19905), .A(n15622), .ZN(n15624) );
  OAI221_X1 U18895 ( .B1(n15627), .B2(n15626), .C1(n15627), .C2(n15625), .A(
        n15624), .ZN(P1_U2812) );
  NAND2_X1 U18896 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15630) );
  INV_X1 U18897 ( .A(n15767), .ZN(n15628) );
  NAND2_X1 U18898 ( .A1(n19961), .A2(n15628), .ZN(n15629) );
  NAND2_X1 U18899 ( .A1(n15630), .A2(n15629), .ZN(n15631) );
  AOI21_X1 U18900 ( .B1(n19937), .B2(P1_EBX_REG_26__SCAN_IN), .A(n15631), .ZN(
        n15638) );
  NAND2_X1 U18901 ( .A1(n15633), .A2(n15632), .ZN(n15635) );
  AND3_X1 U18902 ( .A1(n15635), .A2(n15681), .A3(n15634), .ZN(n15636) );
  AOI21_X1 U18903 ( .B1(n15763), .B2(n19905), .A(n15636), .ZN(n15637) );
  OAI211_X1 U18904 ( .C1(n19952), .C2(n15639), .A(n15638), .B(n15637), .ZN(
        P1_U2814) );
  AOI22_X1 U18905 ( .A1(n15641), .A2(n15640), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n19937), .ZN(n15648) );
  NOR2_X1 U18906 ( .A1(n15772), .A2(n19948), .ZN(n15645) );
  OAI22_X1 U18907 ( .A1(n15643), .A2(n19920), .B1(n15642), .B2(n19952), .ZN(
        n15644) );
  AOI211_X1 U18908 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(n15646), .A(n15645), 
        .B(n15644), .ZN(n15647) );
  OAI211_X1 U18909 ( .C1(n15649), .C2(n19913), .A(n15648), .B(n15647), .ZN(
        P1_U2816) );
  INV_X1 U18910 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n15876) );
  NAND3_X1 U18911 ( .A1(n19925), .A2(n15650), .A3(n15876), .ZN(n15653) );
  INV_X1 U18912 ( .A(n15779), .ZN(n15651) );
  AOI22_X1 U18913 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19955), .B1(
        n19961), .B2(n15651), .ZN(n15652) );
  OAI211_X1 U18914 ( .C1(n19950), .C2(n15654), .A(n15653), .B(n15652), .ZN(
        n15655) );
  AOI21_X1 U18915 ( .B1(n15776), .B2(n19905), .A(n15655), .ZN(n15658) );
  NOR3_X1 U18916 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n19958), .A3(n15656), 
        .ZN(n15661) );
  AOI21_X1 U18917 ( .B1(n15656), .B2(n19925), .A(n19954), .ZN(n15669) );
  INV_X1 U18918 ( .A(n15669), .ZN(n15659) );
  OAI21_X1 U18919 ( .B1(n15661), .B2(n15659), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15657) );
  OAI211_X1 U18920 ( .C1(n15869), .C2(n19952), .A(n15658), .B(n15657), .ZN(
        P1_U2818) );
  AOI22_X1 U18921 ( .A1(n15780), .A2(n19961), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n15659), .ZN(n15665) );
  AOI22_X1 U18922 ( .A1(n19937), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19955), .ZN(n15664) );
  AOI22_X1 U18923 ( .A1(n15781), .A2(n19905), .B1(n15660), .B2(n19926), .ZN(
        n15663) );
  INV_X1 U18924 ( .A(n15661), .ZN(n15662) );
  NAND4_X1 U18925 ( .A1(n15665), .A2(n15664), .A3(n15663), .A4(n15662), .ZN(
        P1_U2819) );
  AOI22_X1 U18926 ( .A1(n19937), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19955), .ZN(n15672) );
  AOI21_X1 U18927 ( .B1(n19925), .B2(n15666), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15668) );
  OAI22_X1 U18928 ( .A1(n15669), .A2(n15668), .B1(n15667), .B2(n19952), .ZN(
        n15670) );
  AOI21_X1 U18929 ( .B1(n15787), .B2(n19905), .A(n15670), .ZN(n15671) );
  OAI211_X1 U18930 ( .C1(n15786), .C2(n19948), .A(n15672), .B(n15671), .ZN(
        P1_U2820) );
  INV_X1 U18931 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15801) );
  OAI22_X1 U18932 ( .A1(n19950), .A2(n15673), .B1(n15801), .B2(n19913), .ZN(
        n15676) );
  OAI22_X1 U18933 ( .A1(n15674), .A2(n19920), .B1(n19952), .B2(n15888), .ZN(
        n15675) );
  NOR4_X1 U18934 ( .A1(n15677), .A2(n19941), .A3(n15676), .A4(n15675), .ZN(
        n15680) );
  NAND2_X1 U18935 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15678), .ZN(n15679) );
  OAI211_X1 U18936 ( .C1(n19948), .C2(n15795), .A(n15680), .B(n15679), .ZN(
        P1_U2822) );
  NAND2_X1 U18937 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n15682) );
  AOI21_X1 U18938 ( .B1(n15682), .B2(n15681), .A(n15722), .ZN(n15716) );
  OAI21_X1 U18939 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n15683), .ZN(n15684) );
  NOR2_X1 U18940 ( .A1(n15702), .A2(n15684), .ZN(n15692) );
  INV_X1 U18941 ( .A(n15806), .ZN(n15685) );
  NAND2_X1 U18942 ( .A1(n19961), .A2(n15685), .ZN(n15687) );
  NAND2_X1 U18943 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15686) );
  NAND3_X1 U18944 ( .A1(n15687), .A2(n15686), .A3(n19910), .ZN(n15688) );
  AOI21_X1 U18945 ( .B1(n19937), .B2(P1_EBX_REG_16__SCAN_IN), .A(n15688), .ZN(
        n15689) );
  OAI21_X1 U18946 ( .B1(n15690), .B2(n19952), .A(n15689), .ZN(n15691) );
  AOI211_X1 U18947 ( .C1(n15802), .C2(n19905), .A(n15692), .B(n15691), .ZN(
        n15693) );
  OAI21_X1 U18948 ( .B1(n15716), .B2(n14350), .A(n15693), .ZN(P1_U2824) );
  INV_X1 U18949 ( .A(n15694), .ZN(n15704) );
  INV_X1 U18950 ( .A(n15905), .ZN(n15700) );
  NAND2_X1 U18951 ( .A1(n19937), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n15698) );
  NAND2_X1 U18952 ( .A1(n15695), .A2(n19961), .ZN(n15697) );
  NAND2_X1 U18953 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15696) );
  NAND4_X1 U18954 ( .A1(n15698), .A2(n19910), .A3(n15697), .A4(n15696), .ZN(
        n15699) );
  AOI21_X1 U18955 ( .B1(n15700), .B2(n19926), .A(n15699), .ZN(n15701) );
  OAI21_X1 U18956 ( .B1(n15702), .B2(P1_REIP_REG_15__SCAN_IN), .A(n15701), 
        .ZN(n15703) );
  AOI21_X1 U18957 ( .B1(n15704), .B2(n19905), .A(n15703), .ZN(n15705) );
  OAI21_X1 U18958 ( .B1(n15716), .B2(n14229), .A(n15705), .ZN(P1_U2825) );
  INV_X1 U18959 ( .A(n15706), .ZN(n15707) );
  AOI21_X1 U18960 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15707), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15715) );
  OAI22_X1 U18961 ( .A1(n15709), .A2(n19952), .B1(n15708), .B2(n19950), .ZN(
        n15710) );
  AOI211_X1 U18962 ( .C1(n19955), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n19941), .B(n15710), .ZN(n15714) );
  INV_X1 U18963 ( .A(n15711), .ZN(n15807) );
  OAI22_X1 U18964 ( .A1(n15808), .A2(n19920), .B1(n19948), .B2(n15807), .ZN(
        n15712) );
  INV_X1 U18965 ( .A(n15712), .ZN(n15713) );
  OAI211_X1 U18966 ( .C1(n15716), .C2(n15715), .A(n15714), .B(n15713), .ZN(
        P1_U2826) );
  OAI22_X1 U18967 ( .A1(n19950), .A2(n15718), .B1(n15717), .B2(n19913), .ZN(
        n15719) );
  AOI211_X1 U18968 ( .C1(n15720), .C2(n19926), .A(n19941), .B(n15719), .ZN(
        n15724) );
  NAND4_X1 U18969 ( .A1(n19925), .A2(n19893), .A3(P1_REIP_REG_10__SCAN_IN), 
        .A4(P1_REIP_REG_9__SCAN_IN), .ZN(n15741) );
  OAI21_X1 U18970 ( .B1(n15729), .B2(n15741), .A(n20792), .ZN(n15721) );
  AOI22_X1 U18971 ( .A1(n15814), .A2(n19961), .B1(n15722), .B2(n15721), .ZN(
        n15723) );
  OAI211_X1 U18972 ( .C1(n19920), .C2(n15758), .A(n15724), .B(n15723), .ZN(
        P1_U2828) );
  INV_X1 U18973 ( .A(n15725), .ZN(n15726) );
  XNOR2_X1 U18974 ( .A(n15727), .B(n15726), .ZN(n15821) );
  OAI22_X1 U18975 ( .A1(n15824), .A2(n19948), .B1(n15729), .B2(n15728), .ZN(
        n15739) );
  NAND2_X1 U18976 ( .A1(n15731), .A2(n15730), .ZN(n15732) );
  AND2_X1 U18977 ( .A1(n15733), .A2(n15732), .ZN(n15924) );
  NAND2_X1 U18978 ( .A1(n19937), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n15734) );
  OAI211_X1 U18979 ( .C1(n19913), .C2(n15735), .A(n15734), .B(n19910), .ZN(
        n15736) );
  AOI21_X1 U18980 ( .B1(n15924), .B2(n19926), .A(n15736), .ZN(n15737) );
  INV_X1 U18981 ( .A(n15737), .ZN(n15738) );
  AOI211_X1 U18982 ( .C1(n19905), .C2(n15821), .A(n15739), .B(n15738), .ZN(
        n15740) );
  OAI21_X1 U18983 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15741), .A(n15740), 
        .ZN(P1_U2829) );
  AOI22_X1 U18984 ( .A1(n15821), .A2(n19966), .B1(n19965), .B2(n15924), .ZN(
        n15742) );
  OAI21_X1 U18985 ( .B1(n19970), .B2(n15743), .A(n15742), .ZN(P1_U2861) );
  INV_X1 U18986 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16289) );
  AOI22_X1 U18987 ( .A1(P1_EAX_REG_29__SCAN_IN), .A2(n15760), .B1(n15751), 
        .B2(n20048), .ZN(n15746) );
  AOI22_X1 U18988 ( .A1(n15744), .A2(n15753), .B1(n15752), .B2(DATAI_29_), 
        .ZN(n15745) );
  OAI211_X1 U18989 ( .C1(n16289), .C2(n15756), .A(n15746), .B(n15745), .ZN(
        P1_U2875) );
  AOI22_X1 U18990 ( .A1(P1_EAX_REG_26__SCAN_IN), .A2(n15760), .B1(n15751), 
        .B2(n20042), .ZN(n15748) );
  AOI22_X1 U18991 ( .A1(n15763), .A2(n15753), .B1(n15752), .B2(DATAI_26_), 
        .ZN(n15747) );
  OAI211_X1 U18992 ( .C1(n16295), .C2(n15756), .A(n15748), .B(n15747), .ZN(
        P1_U2878) );
  INV_X1 U18993 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16303) );
  AOI22_X1 U18994 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(n15760), .B1(n15751), 
        .B2(n20190), .ZN(n15750) );
  AOI22_X1 U18995 ( .A1(n15776), .A2(n15753), .B1(n15752), .B2(DATAI_22_), 
        .ZN(n15749) );
  OAI211_X1 U18996 ( .C1(n15756), .C2(n16303), .A(n15750), .B(n15749), .ZN(
        P1_U2882) );
  AOI22_X1 U18997 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(n15760), .B1(n15751), 
        .B2(n20178), .ZN(n15755) );
  AOI22_X1 U18998 ( .A1(n15787), .A2(n15753), .B1(n15752), .B2(DATAI_20_), 
        .ZN(n15754) );
  OAI211_X1 U18999 ( .C1(n16307), .C2(n15756), .A(n15755), .B(n15754), .ZN(
        P1_U2884) );
  AOI22_X1 U19000 ( .A1(P1_EAX_REG_12__SCAN_IN), .A2(n15760), .B1(n20046), 
        .B2(n15759), .ZN(n15757) );
  OAI21_X1 U19001 ( .B1(n19975), .B2(n15758), .A(n15757), .ZN(P1_U2892) );
  INV_X1 U19002 ( .A(n15821), .ZN(n15762) );
  AOI22_X1 U19003 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(n15760), .B1(n20044), 
        .B2(n15759), .ZN(n15761) );
  OAI21_X1 U19004 ( .B1(n19975), .B2(n15762), .A(n15761), .ZN(P1_U2893) );
  AOI22_X1 U19005 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n15766) );
  AOI22_X1 U19006 ( .A1(n15764), .A2(n20071), .B1(n20070), .B2(n15763), .ZN(
        n15765) );
  OAI211_X1 U19007 ( .C1(n20075), .C2(n15767), .A(n15766), .B(n15765), .ZN(
        P1_U2973) );
  AOI22_X1 U19008 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n15771) );
  AOI22_X1 U19009 ( .A1(n15769), .A2(n20071), .B1(n20070), .B2(n15768), .ZN(
        n15770) );
  OAI211_X1 U19010 ( .C1(n20075), .C2(n15772), .A(n15771), .B(n15770), .ZN(
        P1_U2975) );
  AOI22_X1 U19011 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15778) );
  NAND2_X1 U19012 ( .A1(n15774), .A2(n15773), .ZN(n15775) );
  XOR2_X1 U19013 ( .A(n15775), .B(n15867), .Z(n15871) );
  AOI22_X1 U19014 ( .A1(n15871), .A2(n20071), .B1(n20070), .B2(n15776), .ZN(
        n15777) );
  OAI211_X1 U19015 ( .C1(n20075), .C2(n15779), .A(n15778), .B(n15777), .ZN(
        P1_U2977) );
  AOI22_X1 U19016 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15783) );
  AOI22_X1 U19017 ( .A1(n15781), .A2(n20070), .B1(n20079), .B2(n15780), .ZN(
        n15782) );
  OAI211_X1 U19018 ( .C1(n15784), .C2(n20089), .A(n15783), .B(n15782), .ZN(
        P1_U2978) );
  INV_X1 U19019 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15792) );
  INV_X1 U19020 ( .A(n15785), .ZN(n15789) );
  INV_X1 U19021 ( .A(n15786), .ZN(n15788) );
  AOI222_X1 U19022 ( .A1(n15789), .A2(n20071), .B1(n15788), .B2(n20079), .C1(
        n20070), .C2(n15787), .ZN(n15791) );
  NAND2_X1 U19023 ( .A1(n20128), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15790) );
  OAI211_X1 U19024 ( .C1(n15792), .C2(n15800), .A(n15791), .B(n15790), .ZN(
        P1_U2979) );
  OAI21_X1 U19025 ( .B1(n15794), .B2(n15793), .A(n14199), .ZN(n15889) );
  INV_X1 U19026 ( .A(n15889), .ZN(n15798) );
  INV_X1 U19027 ( .A(n15795), .ZN(n15797) );
  AOI222_X1 U19028 ( .A1(n15798), .A2(n20071), .B1(n15797), .B2(n20079), .C1(
        n20070), .C2(n15796), .ZN(n15799) );
  NAND2_X1 U19029 ( .A1(n20128), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15892) );
  OAI211_X1 U19030 ( .C1(n15801), .C2(n15800), .A(n15799), .B(n15892), .ZN(
        P1_U2981) );
  AOI22_X1 U19031 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15805) );
  AOI22_X1 U19032 ( .A1(n15803), .A2(n20071), .B1(n20070), .B2(n15802), .ZN(
        n15804) );
  OAI211_X1 U19033 ( .C1(n20075), .C2(n15806), .A(n15805), .B(n15804), .ZN(
        P1_U2983) );
  AOI22_X1 U19034 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15811) );
  OAI22_X1 U19035 ( .A1(n15808), .A2(n20149), .B1(n20075), .B2(n15807), .ZN(
        n15809) );
  INV_X1 U19036 ( .A(n15809), .ZN(n15810) );
  OAI211_X1 U19037 ( .C1(n15812), .C2(n20089), .A(n15811), .B(n15810), .ZN(
        P1_U2985) );
  AOI22_X1 U19038 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n20128), .B1(n20086), 
        .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15816) );
  AOI22_X1 U19039 ( .A1(n20079), .A2(n15814), .B1(n20070), .B2(n15813), .ZN(
        n15815) );
  OAI211_X1 U19040 ( .C1(n15817), .C2(n20089), .A(n15816), .B(n15815), .ZN(
        P1_U2987) );
  AOI22_X1 U19041 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15823) );
  OAI33_X1 U19042 ( .A1(n9618), .A2(n15938), .A3(n14208), .B1(n15819), .B2(
        n15818), .B3(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15820) );
  XOR2_X1 U19043 ( .A(n15820), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n15926) );
  AOI22_X1 U19044 ( .A1(n20071), .A2(n15926), .B1(n20070), .B2(n15821), .ZN(
        n15822) );
  OAI211_X1 U19045 ( .C1(n20075), .C2(n15824), .A(n15823), .B(n15822), .ZN(
        P1_U2988) );
  AOI22_X1 U19046 ( .A1(n9618), .A2(n15945), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15819), .ZN(n15826) );
  XOR2_X1 U19047 ( .A(n15827), .B(n15826), .Z(n15942) );
  INV_X1 U19048 ( .A(n15942), .ZN(n15831) );
  AOI22_X1 U19049 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n15830) );
  INV_X1 U19050 ( .A(n15828), .ZN(n19967) );
  AOI22_X1 U19051 ( .A1(n19967), .A2(n20070), .B1(n20079), .B2(n19892), .ZN(
        n15829) );
  OAI211_X1 U19052 ( .C1(n15831), .C2(n20089), .A(n15830), .B(n15829), .ZN(
        P1_U2990) );
  AOI21_X1 U19053 ( .B1(n15834), .B2(n15833), .A(n15832), .ZN(n15959) );
  AOI22_X1 U19054 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15837) );
  INV_X1 U19055 ( .A(n19909), .ZN(n15835) );
  AOI22_X1 U19056 ( .A1(n19906), .A2(n20070), .B1(n20079), .B2(n15835), .ZN(
        n15836) );
  OAI211_X1 U19057 ( .C1(n15959), .C2(n20089), .A(n15837), .B(n15836), .ZN(
        P1_U2992) );
  AOI22_X1 U19058 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15842) );
  AOI21_X1 U19059 ( .B1(n15839), .B2(n15838), .A(n9647), .ZN(n15967) );
  INV_X1 U19060 ( .A(n15840), .ZN(n19933) );
  AOI22_X1 U19061 ( .A1(n15967), .A2(n20071), .B1(n20070), .B2(n19933), .ZN(
        n15841) );
  OAI211_X1 U19062 ( .C1(n20075), .C2(n19936), .A(n15842), .B(n15841), .ZN(
        P1_U2994) );
  AOI22_X1 U19063 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15843), .B1(
        n20128), .B2(P1_REIP_REG_27__SCAN_IN), .ZN(n15846) );
  AOI22_X1 U19064 ( .A1(n15849), .A2(n20130), .B1(n20131), .B2(n15848), .ZN(
        n15856) );
  INV_X1 U19065 ( .A(n15850), .ZN(n15854) );
  NOR2_X1 U19066 ( .A1(n20114), .A2(n20809), .ZN(n15851) );
  AOI221_X1 U19067 ( .B1(n15854), .B2(n15853), .C1(n15852), .C2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15851), .ZN(n15855) );
  NAND2_X1 U19068 ( .A1(n15856), .A2(n15855), .ZN(P1_U3006) );
  AOI22_X1 U19069 ( .A1(n15858), .A2(n20130), .B1(n20131), .B2(n15857), .ZN(
        n15865) );
  INV_X1 U19070 ( .A(n15859), .ZN(n15861) );
  NOR2_X1 U19071 ( .A1(n20114), .A2(n14192), .ZN(n15860) );
  AOI221_X1 U19072 ( .B1(n15863), .B2(n15862), .C1(n15861), .C2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n15860), .ZN(n15864) );
  NAND2_X1 U19073 ( .A1(n15865), .A2(n15864), .ZN(P1_U3008) );
  INV_X1 U19074 ( .A(n15866), .ZN(n15868) );
  OAI22_X1 U19075 ( .A1(n15869), .A2(n20116), .B1(n15868), .B2(n15867), .ZN(
        n15870) );
  AOI21_X1 U19076 ( .B1(n15871), .B2(n20130), .A(n15870), .ZN(n15875) );
  OAI211_X1 U19077 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15873), .B(n15872), .ZN(
        n15874) );
  OAI211_X1 U19078 ( .C1(n15876), .C2(n20114), .A(n15875), .B(n15874), .ZN(
        P1_U3009) );
  INV_X1 U19079 ( .A(n15877), .ZN(n15878) );
  AOI22_X1 U19080 ( .A1(n20128), .A2(P1_REIP_REG_19__SCAN_IN), .B1(n15879), 
        .B2(n15878), .ZN(n15883) );
  AOI22_X1 U19081 ( .A1(n15881), .A2(n20130), .B1(n20131), .B2(n15880), .ZN(
        n15882) );
  OAI211_X1 U19082 ( .C1(n9630), .C2(n15884), .A(n15883), .B(n15882), .ZN(
        P1_U3012) );
  AOI21_X1 U19083 ( .B1(n20127), .B2(n15886), .A(n15885), .ZN(n15904) );
  NOR3_X1 U19084 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15887), .A3(
        n15886), .ZN(n15891) );
  OAI22_X1 U19085 ( .A1(n15889), .A2(n20120), .B1(n20116), .B2(n15888), .ZN(
        n15890) );
  NOR2_X1 U19086 ( .A1(n15891), .A2(n15890), .ZN(n15893) );
  OAI211_X1 U19087 ( .C1(n15904), .C2(n15894), .A(n15893), .B(n15892), .ZN(
        P1_U3013) );
  NOR3_X1 U19088 ( .A1(n15896), .A2(n15895), .A3(n15910), .ZN(n15898) );
  AOI21_X1 U19089 ( .B1(n15898), .B2(n15897), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15903) );
  AOI22_X1 U19090 ( .A1(n15900), .A2(n20130), .B1(n20131), .B2(n15899), .ZN(
        n15902) );
  NAND2_X1 U19091 ( .A1(n20128), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15901) );
  OAI211_X1 U19092 ( .C1(n15904), .C2(n15903), .A(n15902), .B(n15901), .ZN(
        P1_U3014) );
  OAI22_X1 U19093 ( .A1(n15905), .A2(n20116), .B1(n14229), .B2(n20114), .ZN(
        n15906) );
  AOI21_X1 U19094 ( .B1(n15907), .B2(n20130), .A(n15906), .ZN(n15909) );
  OAI211_X1 U19095 ( .C1(n15911), .C2(n15910), .A(n15909), .B(n15908), .ZN(
        P1_U3016) );
  NOR2_X1 U19096 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15912), .ZN(
        n15913) );
  AOI21_X1 U19097 ( .B1(n20131), .B2(n15914), .A(n15913), .ZN(n15915) );
  OAI21_X1 U19098 ( .B1(n15917), .B2(n15916), .A(n15915), .ZN(n15918) );
  AOI21_X1 U19099 ( .B1(n15919), .B2(n20130), .A(n15918), .ZN(n15921) );
  NAND2_X1 U19100 ( .A1(n20128), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15920) );
  OAI211_X1 U19101 ( .C1(n15923), .C2(n15922), .A(n15921), .B(n15920), .ZN(
        P1_U3018) );
  AOI22_X1 U19102 ( .A1(n15924), .A2(n20131), .B1(n20128), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15928) );
  AOI22_X1 U19103 ( .A1(n15926), .A2(n20130), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15925), .ZN(n15927) );
  OAI211_X1 U19104 ( .C1(n15953), .C2(n15929), .A(n15928), .B(n15927), .ZN(
        P1_U3020) );
  AOI221_X1 U19105 ( .B1(n15930), .B2(n20127), .C1(n15935), .C2(n20127), .A(
        n20111), .ZN(n15946) );
  OAI22_X1 U19106 ( .A1(n15932), .A2(n20116), .B1(n15931), .B2(n20114), .ZN(
        n15933) );
  AOI21_X1 U19107 ( .B1(n15934), .B2(n20130), .A(n15933), .ZN(n15937) );
  NOR2_X1 U19108 ( .A1(n15935), .A2(n15953), .ZN(n15941) );
  OAI221_X1 U19109 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n15938), .C2(n15945), .A(
        n15941), .ZN(n15936) );
  OAI211_X1 U19110 ( .C1(n15946), .C2(n15938), .A(n15937), .B(n15936), .ZN(
        P1_U3021) );
  AOI21_X1 U19111 ( .B1(n9976), .B2(n15940), .A(n9721), .ZN(n19964) );
  AOI22_X1 U19112 ( .A1(n19964), .A2(n20131), .B1(n20128), .B2(
        P1_REIP_REG_9__SCAN_IN), .ZN(n15944) );
  AOI22_X1 U19113 ( .A1(n15942), .A2(n20130), .B1(n15945), .B2(n15941), .ZN(
        n15943) );
  OAI211_X1 U19114 ( .C1(n15946), .C2(n15945), .A(n15944), .B(n15943), .ZN(
        P1_U3022) );
  OAI21_X1 U19115 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15948), .A(
        n15947), .ZN(n15949) );
  INV_X1 U19116 ( .A(n15949), .ZN(n15965) );
  INV_X1 U19117 ( .A(n15950), .ZN(n15951) );
  AOI222_X1 U19118 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20128), .B1(n20130), 
        .B2(n15952), .C1(n20131), .C2(n15951), .ZN(n15956) );
  INV_X1 U19119 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15964) );
  NOR2_X1 U19120 ( .A1(n15954), .A2(n15953), .ZN(n15960) );
  OAI221_X1 U19121 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n15957), .C2(n15964), .A(
        n15960), .ZN(n15955) );
  OAI211_X1 U19122 ( .C1(n15965), .C2(n15957), .A(n15956), .B(n15955), .ZN(
        P1_U3023) );
  INV_X1 U19123 ( .A(n15958), .ZN(n19900) );
  AOI22_X1 U19124 ( .A1(n19900), .A2(n20131), .B1(n20128), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n15963) );
  INV_X1 U19125 ( .A(n15959), .ZN(n15961) );
  AOI22_X1 U19126 ( .A1(n15961), .A2(n20130), .B1(n15964), .B2(n15960), .ZN(
        n15962) );
  OAI211_X1 U19127 ( .C1(n15965), .C2(n15964), .A(n15963), .B(n15962), .ZN(
        P1_U3024) );
  AOI22_X1 U19128 ( .A1(n19927), .A2(n20131), .B1(n20128), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n15969) );
  AOI22_X1 U19129 ( .A1(n15967), .A2(n20130), .B1(n20103), .B2(n15966), .ZN(
        n15968) );
  OAI211_X1 U19130 ( .C1(n15971), .C2(n15970), .A(n15969), .B(n15968), .ZN(
        P1_U3026) );
  NAND4_X1 U19131 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n11268), .A4(n20769), .ZN(n15972) );
  NAND2_X1 U19132 ( .A1(n15973), .A2(n15972), .ZN(n20755) );
  OAI21_X1 U19133 ( .B1(n15975), .B2(n20755), .A(n15974), .ZN(n15976) );
  OAI221_X1 U19134 ( .B1(n15977), .B2(n20570), .C1(n15977), .C2(n20769), .A(
        n15976), .ZN(n15978) );
  AOI221_X1 U19135 ( .B1(n15979), .B2(n20753), .C1(n20754), .C2(n20753), .A(
        n15978), .ZN(P1_U3162) );
  NOR2_X1 U19136 ( .A1(n15979), .A2(n20754), .ZN(n15981) );
  OAI22_X1 U19137 ( .A1(n20570), .A2(n15981), .B1(n15980), .B2(n20754), .ZN(
        P1_U3466) );
  AOI22_X1 U19138 ( .A1(P2_REIP_REG_31__SCAN_IN), .A2(n19027), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n18979), .ZN(n15991) );
  AOI22_X1 U19139 ( .A1(n19008), .A2(n19086), .B1(n18998), .B2(n16068), .ZN(
        n15990) );
  NAND4_X1 U19140 ( .A1(n19000), .A2(n15983), .A3(n18994), .A4(n15982), .ZN(
        n15989) );
  AND2_X1 U19141 ( .A1(n15985), .A2(n15984), .ZN(n15987) );
  OAI21_X1 U19142 ( .B1(n15987), .B2(n15986), .A(P2_EBX_REG_31__SCAN_IN), .ZN(
        n15988) );
  NAND4_X1 U19143 ( .A1(n15991), .A2(n15990), .A3(n15989), .A4(n15988), .ZN(
        P2_U2824) );
  AOI22_X1 U19144 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18979), .B1(
        n15992), .B2(n19026), .ZN(n16002) );
  AOI22_X1 U19145 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19027), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19028), .ZN(n16001) );
  OAI22_X1 U19146 ( .A1(n15994), .A2(n19022), .B1(n15993), .B2(n19032), .ZN(
        n15995) );
  INV_X1 U19147 ( .A(n15995), .ZN(n16000) );
  OAI211_X1 U19148 ( .C1(n15998), .C2(n15997), .A(n19000), .B(n15996), .ZN(
        n15999) );
  NAND4_X1 U19149 ( .A1(n16002), .A2(n16001), .A3(n16000), .A4(n15999), .ZN(
        P2_U2826) );
  AOI22_X1 U19150 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n19027), .B1(n16003), 
        .B2(n19026), .ZN(n16012) );
  AOI22_X1 U19151 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18979), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n19028), .ZN(n16011) );
  AOI22_X1 U19152 ( .A1(n16005), .A2(n18998), .B1(n16004), .B2(n19008), .ZN(
        n16010) );
  OAI211_X1 U19153 ( .C1(n16008), .C2(n16007), .A(n19000), .B(n16006), .ZN(
        n16009) );
  NAND4_X1 U19154 ( .A1(n16012), .A2(n16011), .A3(n16010), .A4(n16009), .ZN(
        P2_U2827) );
  OAI22_X1 U19155 ( .A1(n16014), .A2(n18850), .B1(n16013), .B2(n18989), .ZN(
        n16017) );
  AOI22_X1 U19156 ( .A1(n19028), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19027), .ZN(n16015) );
  INV_X1 U19157 ( .A(n16015), .ZN(n16016) );
  AOI211_X1 U19158 ( .C1(n16018), .C2(n18998), .A(n16017), .B(n16016), .ZN(
        n16023) );
  OAI211_X1 U19159 ( .C1(n16021), .C2(n16020), .A(n19000), .B(n16019), .ZN(
        n16022) );
  OAI211_X1 U19160 ( .C1(n19032), .C2(n16024), .A(n16023), .B(n16022), .ZN(
        P2_U2828) );
  AOI22_X1 U19161 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19027), .B1(n16025), 
        .B2(n19026), .ZN(n16034) );
  AOI22_X1 U19162 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18979), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19028), .ZN(n16033) );
  AOI22_X1 U19163 ( .A1(n16027), .A2(n18998), .B1(n16026), .B2(n19008), .ZN(
        n16032) );
  OAI211_X1 U19164 ( .C1(n16030), .C2(n16029), .A(n19000), .B(n16028), .ZN(
        n16031) );
  NAND4_X1 U19165 ( .A1(n16034), .A2(n16033), .A3(n16032), .A4(n16031), .ZN(
        P2_U2829) );
  OAI22_X1 U19166 ( .A1(n16035), .A2(n18989), .B1(n19766), .B2(n19004), .ZN(
        n16036) );
  INV_X1 U19167 ( .A(n16036), .ZN(n16045) );
  AOI22_X1 U19168 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18979), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19028), .ZN(n16044) );
  AOI22_X1 U19169 ( .A1(n16038), .A2(n18998), .B1(n16037), .B2(n19008), .ZN(
        n16043) );
  OAI211_X1 U19170 ( .C1(n16041), .C2(n16040), .A(n19000), .B(n16039), .ZN(
        n16042) );
  NAND4_X1 U19171 ( .A1(n16045), .A2(n16044), .A3(n16043), .A4(n16042), .ZN(
        P2_U2830) );
  OAI22_X1 U19172 ( .A1(n14832), .A2(n19004), .B1(n16046), .B2(n18989), .ZN(
        n16049) );
  AOI22_X1 U19173 ( .A1(n19028), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19038), .ZN(n16047) );
  INV_X1 U19174 ( .A(n16047), .ZN(n16048) );
  AOI211_X1 U19175 ( .C1(n16050), .C2(n19008), .A(n16049), .B(n16048), .ZN(
        n16055) );
  OAI211_X1 U19176 ( .C1(n16053), .C2(n16052), .A(n19000), .B(n16051), .ZN(
        n16054) );
  OAI211_X1 U19177 ( .C1(n19022), .C2(n16056), .A(n16055), .B(n16054), .ZN(
        P2_U2831) );
  AOI22_X1 U19178 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19038), .B1(
        n16057), .B2(n19026), .ZN(n16067) );
  AOI22_X1 U19179 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19027), .B1(
        P2_EBX_REG_23__SCAN_IN), .B2(n19028), .ZN(n16066) );
  INV_X1 U19180 ( .A(n16058), .ZN(n16059) );
  AOI22_X1 U19181 ( .A1(n16060), .A2(n18998), .B1(n16059), .B2(n19008), .ZN(
        n16065) );
  OAI211_X1 U19182 ( .C1(n16063), .C2(n16062), .A(n19000), .B(n16061), .ZN(
        n16064) );
  NAND4_X1 U19183 ( .A1(n16067), .A2(n16066), .A3(n16065), .A4(n16064), .ZN(
        P2_U2832) );
  OAI22_X1 U19184 ( .A1(n19084), .A2(n16068), .B1(P2_EBX_REG_31__SCAN_IN), 
        .B2(n19070), .ZN(n16069) );
  INV_X1 U19185 ( .A(n16069), .ZN(P2_U2856) );
  INV_X1 U19186 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16072) );
  AOI22_X1 U19187 ( .A1(n16070), .A2(n19081), .B1(n19070), .B2(n16097), .ZN(
        n16071) );
  OAI21_X1 U19188 ( .B1(n19070), .B2(n16072), .A(n16071), .ZN(P2_U2865) );
  NOR2_X1 U19189 ( .A1(n14494), .A2(n16073), .ZN(n16074) );
  OR2_X1 U19190 ( .A1(n14484), .A2(n16074), .ZN(n16084) );
  OAI22_X1 U19191 ( .A1(n16084), .A2(n19075), .B1(n19070), .B2(n9997), .ZN(
        n16075) );
  INV_X1 U19192 ( .A(n16075), .ZN(n16076) );
  OAI21_X1 U19193 ( .B1(n19084), .B2(n18835), .A(n16076), .ZN(P2_U2867) );
  INV_X1 U19194 ( .A(n16077), .ZN(n16078) );
  AOI21_X1 U19195 ( .B1(n16079), .B2(n14498), .A(n16078), .ZN(n16091) );
  AOI22_X1 U19196 ( .A1(n16091), .A2(n19081), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19084), .ZN(n16080) );
  OAI21_X1 U19197 ( .B1(n19084), .B2(n18858), .A(n16080), .ZN(P2_U2869) );
  INV_X1 U19198 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18145) );
  INV_X1 U19199 ( .A(n19087), .ZN(n19093) );
  OAI22_X1 U19200 ( .A1(n19093), .A2(n16307), .B1(n16081), .B2(n19090), .ZN(
        n16082) );
  AOI21_X1 U19201 ( .B1(P2_EAX_REG_20__SCAN_IN), .B2(n19102), .A(n16082), .ZN(
        n16088) );
  OAI22_X1 U19202 ( .A1(n18824), .A2(n16085), .B1(n16084), .B2(n16083), .ZN(
        n16086) );
  INV_X1 U19203 ( .A(n16086), .ZN(n16087) );
  OAI211_X1 U19204 ( .C1(n19101), .C2(n18145), .A(n16088), .B(n16087), .ZN(
        P2_U2899) );
  INV_X1 U19205 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18135) );
  INV_X1 U19206 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16311) );
  OAI22_X1 U19207 ( .A1(n19093), .A2(n16311), .B1(n16089), .B2(n19090), .ZN(
        n16090) );
  AOI21_X1 U19208 ( .B1(P2_EAX_REG_18__SCAN_IN), .B2(n19102), .A(n16090), .ZN(
        n16093) );
  AOI22_X1 U19209 ( .A1(n18852), .A2(n19096), .B1(n16091), .B2(n19105), .ZN(
        n16092) );
  OAI211_X1 U19210 ( .C1(n19101), .C2(n18135), .A(n16093), .B(n16092), .ZN(
        P2_U2901) );
  AOI22_X1 U19211 ( .A1(n16142), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18992), .ZN(n16100) );
  INV_X1 U19212 ( .A(n16094), .ZN(n16098) );
  AOI222_X1 U19213 ( .A1(n16098), .A2(n16145), .B1(n16157), .B2(n16097), .C1(
        n16146), .C2(n16096), .ZN(n16099) );
  OAI211_X1 U19214 ( .C1(n16150), .C2(n16101), .A(n16100), .B(n16099), .ZN(
        P2_U2992) );
  AOI22_X1 U19215 ( .A1(n16142), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n18992), .ZN(n16116) );
  NAND2_X1 U19216 ( .A1(n16103), .A2(n16102), .ZN(n16104) );
  NAND2_X1 U19217 ( .A1(n16105), .A2(n16104), .ZN(n19059) );
  NAND2_X1 U19218 ( .A1(n16107), .A2(n16106), .ZN(n16111) );
  NAND2_X1 U19219 ( .A1(n16109), .A2(n16108), .ZN(n16110) );
  XOR2_X1 U19220 ( .A(n16111), .B(n16110), .Z(n16171) );
  OAI21_X1 U19221 ( .B1(n16113), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16112), .ZN(n16167) );
  OAI222_X1 U19222 ( .A1(n19059), .A2(n16138), .B1(n16152), .B2(n16171), .C1(
        n16154), .C2(n16167), .ZN(n16114) );
  INV_X1 U19223 ( .A(n16114), .ZN(n16115) );
  OAI211_X1 U19224 ( .C1(n16150), .C2(n18932), .A(n16116), .B(n16115), .ZN(
        P2_U3004) );
  AOI22_X1 U19225 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18992), .B1(n16151), 
        .B2(n18946), .ZN(n16121) );
  OAI22_X1 U19226 ( .A1(n16118), .A2(n16154), .B1(n16152), .B2(n16117), .ZN(
        n16119) );
  AOI21_X1 U19227 ( .B1(n16157), .B2(n18947), .A(n16119), .ZN(n16120) );
  OAI211_X1 U19228 ( .C1(n16161), .C2(n16122), .A(n16121), .B(n16120), .ZN(
        P2_U3005) );
  AOI22_X1 U19229 ( .A1(n16142), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18992), .ZN(n16141) );
  INV_X1 U19230 ( .A(n16123), .ZN(n16124) );
  AOI21_X1 U19231 ( .B1(n16126), .B2(n16125), .A(n16124), .ZN(n16180) );
  INV_X1 U19232 ( .A(n16127), .ZN(n16128) );
  AOI21_X1 U19233 ( .B1(n16130), .B2(n16129), .A(n16128), .ZN(n16134) );
  NAND2_X1 U19234 ( .A1(n16132), .A2(n16131), .ZN(n16133) );
  XNOR2_X1 U19235 ( .A(n16134), .B(n16133), .ZN(n16183) );
  OAI21_X1 U19236 ( .B1(n16137), .B2(n16136), .A(n16135), .ZN(n19079) );
  OAI22_X1 U19237 ( .A1(n16183), .A2(n16152), .B1(n16138), .B2(n19079), .ZN(
        n16139) );
  AOI21_X1 U19238 ( .B1(n16180), .B2(n16146), .A(n16139), .ZN(n16140) );
  OAI211_X1 U19239 ( .C1(n16150), .C2(n18956), .A(n16141), .B(n16140), .ZN(
        P2_U3006) );
  AOI22_X1 U19240 ( .A1(n16142), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n18992), .ZN(n16149) );
  INV_X1 U19241 ( .A(n16143), .ZN(n16147) );
  AOI222_X1 U19242 ( .A1(n16147), .A2(n16146), .B1(n16145), .B2(n16144), .C1(
        n16157), .C2(n18983), .ZN(n16148) );
  OAI211_X1 U19243 ( .C1(n16150), .C2(n18981), .A(n16149), .B(n16148), .ZN(
        P2_U3008) );
  AOI22_X1 U19244 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n18992), .B1(n16151), 
        .B2(n18996), .ZN(n16159) );
  OAI22_X1 U19245 ( .A1(n16155), .A2(n16154), .B1(n16153), .B2(n16152), .ZN(
        n16156) );
  AOI21_X1 U19246 ( .B1(n16157), .B2(n18997), .A(n16156), .ZN(n16158) );
  OAI211_X1 U19247 ( .C1(n16161), .C2(n16160), .A(n16159), .B(n16158), .ZN(
        P2_U3009) );
  NOR2_X1 U19248 ( .A1(n10895), .A2(n18974), .ZN(n16165) );
  INV_X1 U19249 ( .A(n16162), .ZN(n16163) );
  OAI21_X1 U19250 ( .B1(n18936), .B2(n16184), .A(n16163), .ZN(n16164) );
  AOI211_X1 U19251 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16166), .A(
        n16165), .B(n16164), .ZN(n16170) );
  OAI22_X1 U19252 ( .A1(n16167), .A2(n16189), .B1(n19157), .B2(n19059), .ZN(
        n16168) );
  INV_X1 U19253 ( .A(n16168), .ZN(n16169) );
  OAI211_X1 U19254 ( .C1(n16171), .C2(n19155), .A(n16170), .B(n16169), .ZN(
        P2_U3036) );
  NOR2_X1 U19255 ( .A1(n18974), .A2(n10868), .ZN(n16178) );
  NAND3_X1 U19256 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n16172), .A3(
        n16176), .ZN(n16173) );
  OAI221_X1 U19257 ( .B1(n16176), .B2(n16175), .C1(n16176), .C2(n16174), .A(
        n16173), .ZN(n16177) );
  AOI211_X1 U19258 ( .C1(n19152), .C2(n18958), .A(n16178), .B(n16177), .ZN(
        n16182) );
  INV_X1 U19259 ( .A(n19079), .ZN(n16179) );
  AOI22_X1 U19260 ( .A1(n16180), .A2(n19162), .B1(n16203), .B2(n16179), .ZN(
        n16181) );
  OAI211_X1 U19261 ( .C1(n16183), .C2(n19155), .A(n16182), .B(n16181), .ZN(
        P2_U3038) );
  NOR2_X1 U19262 ( .A1(n16185), .A2(n16184), .ZN(n16186) );
  AOI211_X1 U19263 ( .C1(n16203), .C2(n13293), .A(n16187), .B(n16186), .ZN(
        n16188) );
  OAI21_X1 U19264 ( .B1(n16190), .B2(n16189), .A(n16188), .ZN(n16191) );
  AOI21_X1 U19265 ( .B1(n16200), .B2(n16192), .A(n16191), .ZN(n16193) );
  OAI221_X1 U19266 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16196), .C1(
        n16195), .C2(n16194), .A(n16193), .ZN(P2_U3043) );
  INV_X1 U19267 ( .A(n16197), .ZN(n19153) );
  AOI22_X1 U19268 ( .A1(n19153), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19152), .B2(n16198), .ZN(n16208) );
  AOI22_X1 U19269 ( .A1(n19162), .A2(n16201), .B1(n16200), .B2(n16199), .ZN(
        n16206) );
  AOI21_X1 U19270 ( .B1(n16204), .B2(n16203), .A(n16202), .ZN(n16205) );
  AND2_X1 U19271 ( .A1(n16206), .A2(n16205), .ZN(n16207) );
  OAI211_X1 U19272 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16209), .A(
        n16208), .B(n16207), .ZN(P2_U3046) );
  NOR2_X1 U19273 ( .A1(n19855), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19703) );
  INV_X1 U19274 ( .A(n19703), .ZN(n16224) );
  NAND2_X1 U19275 ( .A1(n16211), .A2(n16210), .ZN(n19706) );
  NAND2_X1 U19276 ( .A1(n19855), .A2(n19790), .ZN(n16212) );
  AOI22_X1 U19277 ( .A1(n19845), .A2(n19706), .B1(n19859), .B2(n16212), .ZN(
        n16219) );
  NAND2_X1 U19278 ( .A1(n19852), .A2(n16213), .ZN(n16214) );
  NOR2_X1 U19279 ( .A1(n16215), .A2(n16214), .ZN(n16216) );
  AOI21_X1 U19280 ( .B1(n16217), .B2(n16216), .A(n19849), .ZN(n16218) );
  AOI211_X1 U19281 ( .C1(n16221), .C2(n16220), .A(n16219), .B(n16218), .ZN(
        n16223) );
  OAI211_X1 U19282 ( .C1(n19850), .C2(n16224), .A(n16223), .B(n16222), .ZN(
        P2_U3176) );
  INV_X1 U19283 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16432) );
  XNOR2_X1 U19284 ( .A(n16432), .B(n16246), .ZN(n16431) );
  NAND2_X1 U19285 ( .A1(n9611), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16225) );
  OAI221_X1 U19286 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16227), .C1(
        n16432), .C2(n16226), .A(n16225), .ZN(n16228) );
  AOI21_X1 U19287 ( .B1(n17605), .B2(n16431), .A(n16228), .ZN(n16233) );
  OAI22_X1 U19288 ( .A1(n16240), .A2(n17678), .B1(n16236), .B2(n17775), .ZN(
        n16231) );
  NOR2_X1 U19289 ( .A1(n9613), .A2(n16229), .ZN(n17440) );
  AOI22_X1 U19290 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16231), .B1(
        n16230), .B2(n17440), .ZN(n16232) );
  OAI211_X1 U19291 ( .C1(n16234), .C2(n17682), .A(n16233), .B(n16232), .ZN(
        P3_U2800) );
  NOR2_X1 U19292 ( .A1(n16238), .A2(n16235), .ZN(n16270) );
  INV_X1 U19293 ( .A(n16270), .ZN(n16237) );
  AOI211_X1 U19294 ( .C1(n16242), .C2(n16237), .A(n16236), .B(n17775), .ZN(
        n16244) );
  NOR2_X1 U19295 ( .A1(n16239), .A2(n16238), .ZN(n16271) );
  INV_X1 U19296 ( .A(n16271), .ZN(n16241) );
  AOI211_X1 U19297 ( .C1(n16242), .C2(n16241), .A(n16240), .B(n17678), .ZN(
        n16243) );
  AOI211_X1 U19298 ( .C1(n17664), .C2(n16245), .A(n16244), .B(n16243), .ZN(
        n16253) );
  INV_X1 U19299 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16442) );
  AOI21_X1 U19300 ( .B1(n16442), .B2(n16408), .A(n16246), .ZN(n16441) );
  OAI21_X1 U19301 ( .B1(n16247), .B2(n17605), .A(n16441), .ZN(n16251) );
  OAI221_X1 U19302 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18493), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16249), .A(n16248), .ZN(
        n16250) );
  NAND4_X1 U19303 ( .A1(n16253), .A2(n16252), .A3(n16251), .A4(n16250), .ZN(
        P3_U2801) );
  NOR3_X1 U19304 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16255), .A3(
        n16254), .ZN(n16256) );
  NAND3_X1 U19305 ( .A1(n16257), .A2(n16256), .A3(n18101), .ZN(n16260) );
  INV_X1 U19306 ( .A(n16258), .ZN(n18090) );
  OAI22_X1 U19307 ( .A1(n17808), .A2(n16260), .B1(n18090), .B2(n16259), .ZN(
        n16261) );
  AOI211_X1 U19308 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16263), .A(
        n16262), .B(n16261), .ZN(n16266) );
  NAND3_X1 U19309 ( .A1(n18101), .A2(n17898), .A3(n17850), .ZN(n17876) );
  INV_X1 U19310 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17418) );
  NAND4_X1 U19311 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16268), .A3(
        n17803), .A4(n17418), .ZN(n17432) );
  NOR4_X1 U19312 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17792), .A3(
        n17670), .A4(n16269), .ZN(n16281) );
  OAI22_X1 U19313 ( .A1(n16271), .A2(n17846), .B1(n16270), .B2(n17844), .ZN(
        n16272) );
  NOR3_X1 U19314 ( .A1(n18092), .A2(n16273), .A3(n16272), .ZN(n16278) );
  NOR2_X1 U19315 ( .A1(n17276), .A2(n18555), .ZN(n16275) );
  AOI22_X1 U19316 ( .A1(n17662), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n17418), .B2(n17670), .ZN(n17429) );
  NAND2_X1 U19317 ( .A1(n17429), .A2(n17428), .ZN(n17427) );
  OAI211_X1 U19318 ( .C1(n17435), .C2(n16276), .A(n16275), .B(n17427), .ZN(
        n16277) );
  AOI211_X1 U19319 ( .C1(n16278), .C2(n16277), .A(n9611), .B(n17418), .ZN(
        n16280) );
  NOR3_X1 U19320 ( .A1(n17429), .A2(n18021), .A3(n17436), .ZN(n16279) );
  NAND2_X1 U19321 ( .A1(n9611), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17423) );
  OAI211_X1 U19322 ( .C1(n17876), .C2(n17432), .A(n16282), .B(n17423), .ZN(
        P3_U2834) );
  NOR3_X1 U19323 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16284) );
  NOR4_X1 U19324 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16283) );
  NAND4_X1 U19325 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16284), .A3(n16283), .A4(
        U215), .ZN(U213) );
  INV_X2 U19326 ( .A(U212), .ZN(n16335) );
  INV_X2 U19327 ( .A(U214), .ZN(n16336) );
  NOR2_X1 U19328 ( .A1(n16336), .A2(n16285), .ZN(n16287) );
  AOI222_X1 U19329 ( .A1(n16335), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(n16287), 
        .B2(BUF1_REG_31__SCAN_IN), .C1(n16336), .C2(P1_DATAO_REG_31__SCAN_IN), 
        .ZN(n16286) );
  INV_X1 U19330 ( .A(n16286), .ZN(U216) );
  INV_X1 U19331 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19116) );
  INV_X1 U19332 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16372) );
  OAI222_X1 U19333 ( .A1(U212), .A2(n19116), .B1(n16338), .B2(n19187), .C1(
        U214), .C2(n16372), .ZN(U217) );
  AOI22_X1 U19334 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16335), .ZN(n16288) );
  OAI21_X1 U19335 ( .B1(n16289), .B2(n16338), .A(n16288), .ZN(U218) );
  INV_X1 U19336 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16291) );
  AOI22_X1 U19337 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16335), .ZN(n16290) );
  OAI21_X1 U19338 ( .B1(n16291), .B2(n16338), .A(n16290), .ZN(U219) );
  INV_X1 U19339 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16293) );
  AOI22_X1 U19340 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16335), .ZN(n16292) );
  OAI21_X1 U19341 ( .B1(n16293), .B2(n16338), .A(n16292), .ZN(U220) );
  AOI22_X1 U19342 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16335), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16336), .ZN(n16294) );
  OAI21_X1 U19343 ( .B1(n16295), .B2(n16338), .A(n16294), .ZN(U221) );
  AOI22_X1 U19344 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16335), .ZN(n16296) );
  OAI21_X1 U19345 ( .B1(n16297), .B2(n16338), .A(n16296), .ZN(U222) );
  AOI22_X1 U19346 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16335), .ZN(n16298) );
  OAI21_X1 U19347 ( .B1(n16299), .B2(n16338), .A(n16298), .ZN(U223) );
  INV_X1 U19348 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16301) );
  AOI22_X1 U19349 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16335), .ZN(n16300) );
  OAI21_X1 U19350 ( .B1(n16301), .B2(n16338), .A(n16300), .ZN(U224) );
  AOI22_X1 U19351 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16335), .ZN(n16302) );
  OAI21_X1 U19352 ( .B1(n16303), .B2(n16338), .A(n16302), .ZN(U225) );
  INV_X1 U19353 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16305) );
  AOI22_X1 U19354 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16335), .ZN(n16304) );
  OAI21_X1 U19355 ( .B1(n16305), .B2(n16338), .A(n16304), .ZN(U226) );
  AOI22_X1 U19356 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16335), .ZN(n16306) );
  OAI21_X1 U19357 ( .B1(n16307), .B2(n16338), .A(n16306), .ZN(U227) );
  INV_X1 U19358 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16309) );
  AOI22_X1 U19359 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16335), .ZN(n16308) );
  OAI21_X1 U19360 ( .B1(n16309), .B2(n16338), .A(n16308), .ZN(U228) );
  AOI22_X1 U19361 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16335), .ZN(n16310) );
  OAI21_X1 U19362 ( .B1(n16311), .B2(n16338), .A(n16310), .ZN(U229) );
  INV_X1 U19363 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16313) );
  AOI22_X1 U19364 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16335), .ZN(n16312) );
  OAI21_X1 U19365 ( .B1(n16313), .B2(n16338), .A(n16312), .ZN(U230) );
  INV_X1 U19366 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n19092) );
  AOI22_X1 U19367 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16335), .ZN(n16314) );
  OAI21_X1 U19368 ( .B1(n19092), .B2(n16338), .A(n16314), .ZN(U231) );
  AOI22_X1 U19369 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16335), .ZN(n16315) );
  OAI21_X1 U19370 ( .B1(n13136), .B2(n16338), .A(n16315), .ZN(U232) );
  AOI22_X1 U19371 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16335), .ZN(n16316) );
  OAI21_X1 U19372 ( .B1(n13631), .B2(n16338), .A(n16316), .ZN(U233) );
  INV_X1 U19373 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16318) );
  AOI22_X1 U19374 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16335), .ZN(n16317) );
  OAI21_X1 U19375 ( .B1(n16318), .B2(n16338), .A(n16317), .ZN(U234) );
  INV_X1 U19376 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16320) );
  AOI22_X1 U19377 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16335), .ZN(n16319) );
  OAI21_X1 U19378 ( .B1(n16320), .B2(n16338), .A(n16319), .ZN(U235) );
  INV_X1 U19379 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16322) );
  AOI22_X1 U19380 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16335), .ZN(n16321) );
  OAI21_X1 U19381 ( .B1(n16322), .B2(n16338), .A(n16321), .ZN(U236) );
  INV_X1 U19382 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16324) );
  AOI22_X1 U19383 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16335), .ZN(n16323) );
  OAI21_X1 U19384 ( .B1(n16324), .B2(n16338), .A(n16323), .ZN(U237) );
  AOI22_X1 U19385 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16335), .ZN(n16325) );
  OAI21_X1 U19386 ( .B1(n12786), .B2(n16338), .A(n16325), .ZN(U238) );
  INV_X1 U19387 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16327) );
  AOI22_X1 U19388 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16335), .ZN(n16326) );
  OAI21_X1 U19389 ( .B1(n16327), .B2(n16338), .A(n16326), .ZN(U239) );
  AOI22_X1 U19390 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16335), .ZN(n16328) );
  OAI21_X1 U19391 ( .B1(n12751), .B2(n16338), .A(n16328), .ZN(U240) );
  AOI22_X1 U19392 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16335), .ZN(n16329) );
  OAI21_X1 U19393 ( .B1(n12799), .B2(n16338), .A(n16329), .ZN(U241) );
  AOI22_X1 U19394 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16335), .ZN(n16330) );
  OAI21_X1 U19395 ( .B1(n12724), .B2(n16338), .A(n16330), .ZN(U242) );
  AOI22_X1 U19396 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16335), .ZN(n16331) );
  OAI21_X1 U19397 ( .B1(n12746), .B2(n16338), .A(n16331), .ZN(U243) );
  AOI22_X1 U19398 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16335), .ZN(n16332) );
  OAI21_X1 U19399 ( .B1(n12756), .B2(n16338), .A(n16332), .ZN(U244) );
  AOI22_X1 U19400 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16335), .ZN(n16333) );
  OAI21_X1 U19401 ( .B1(n12776), .B2(n16338), .A(n16333), .ZN(U245) );
  AOI22_X1 U19402 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16335), .ZN(n16334) );
  OAI21_X1 U19403 ( .B1(n12741), .B2(n16338), .A(n16334), .ZN(U246) );
  AOI22_X1 U19404 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16336), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16335), .ZN(n16337) );
  OAI21_X1 U19405 ( .B1(n12729), .B2(n16338), .A(n16337), .ZN(U247) );
  OAI22_X1 U19406 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16370), .ZN(n16339) );
  INV_X1 U19407 ( .A(n16339), .ZN(U251) );
  OAI22_X1 U19408 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16370), .ZN(n16340) );
  INV_X1 U19409 ( .A(n16340), .ZN(U252) );
  OAI22_X1 U19410 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16370), .ZN(n16341) );
  INV_X1 U19411 ( .A(n16341), .ZN(U253) );
  OAI22_X1 U19412 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16370), .ZN(n16342) );
  INV_X1 U19413 ( .A(n16342), .ZN(U254) );
  OAI22_X1 U19414 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16370), .ZN(n16343) );
  INV_X1 U19415 ( .A(n16343), .ZN(U255) );
  OAI22_X1 U19416 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16370), .ZN(n16344) );
  INV_X1 U19417 ( .A(n16344), .ZN(U256) );
  OAI22_X1 U19418 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16370), .ZN(n16345) );
  INV_X1 U19419 ( .A(n16345), .ZN(U257) );
  OAI22_X1 U19420 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16370), .ZN(n16346) );
  INV_X1 U19421 ( .A(n16346), .ZN(U258) );
  OAI22_X1 U19422 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16370), .ZN(n16347) );
  INV_X1 U19423 ( .A(n16347), .ZN(U259) );
  OAI22_X1 U19424 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16362), .ZN(n16348) );
  INV_X1 U19425 ( .A(n16348), .ZN(U260) );
  OAI22_X1 U19426 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16362), .ZN(n16349) );
  INV_X1 U19427 ( .A(n16349), .ZN(U261) );
  OAI22_X1 U19428 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16370), .ZN(n16350) );
  INV_X1 U19429 ( .A(n16350), .ZN(U262) );
  OAI22_X1 U19430 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16362), .ZN(n16351) );
  INV_X1 U19431 ( .A(n16351), .ZN(U263) );
  OAI22_X1 U19432 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16370), .ZN(n16352) );
  INV_X1 U19433 ( .A(n16352), .ZN(U264) );
  OAI22_X1 U19434 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16370), .ZN(n16353) );
  INV_X1 U19435 ( .A(n16353), .ZN(U265) );
  OAI22_X1 U19436 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16362), .ZN(n16354) );
  INV_X1 U19437 ( .A(n16354), .ZN(U266) );
  OAI22_X1 U19438 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16362), .ZN(n16355) );
  INV_X1 U19439 ( .A(n16355), .ZN(U267) );
  OAI22_X1 U19440 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16362), .ZN(n16356) );
  INV_X1 U19441 ( .A(n16356), .ZN(U268) );
  OAI22_X1 U19442 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16362), .ZN(n16357) );
  INV_X1 U19443 ( .A(n16357), .ZN(U269) );
  OAI22_X1 U19444 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16362), .ZN(n16358) );
  INV_X1 U19445 ( .A(n16358), .ZN(U270) );
  OAI22_X1 U19446 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16362), .ZN(n16359) );
  INV_X1 U19447 ( .A(n16359), .ZN(U271) );
  OAI22_X1 U19448 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16370), .ZN(n16360) );
  INV_X1 U19449 ( .A(n16360), .ZN(U272) );
  OAI22_X1 U19450 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16370), .ZN(n16361) );
  INV_X1 U19451 ( .A(n16361), .ZN(U273) );
  OAI22_X1 U19452 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16362), .ZN(n16363) );
  INV_X1 U19453 ( .A(n16363), .ZN(U274) );
  OAI22_X1 U19454 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16370), .ZN(n16364) );
  INV_X1 U19455 ( .A(n16364), .ZN(U275) );
  OAI22_X1 U19456 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16370), .ZN(n16365) );
  INV_X1 U19457 ( .A(n16365), .ZN(U276) );
  OAI22_X1 U19458 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16370), .ZN(n16366) );
  INV_X1 U19459 ( .A(n16366), .ZN(U277) );
  OAI22_X1 U19460 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16370), .ZN(n16367) );
  INV_X1 U19461 ( .A(n16367), .ZN(U278) );
  OAI22_X1 U19462 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16370), .ZN(n16368) );
  INV_X1 U19463 ( .A(n16368), .ZN(U279) );
  OAI22_X1 U19464 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16370), .ZN(n16369) );
  INV_X1 U19465 ( .A(n16369), .ZN(U280) );
  INV_X1 U19466 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19185) );
  AOI22_X1 U19467 ( .A1(n16370), .A2(n19116), .B1(n19185), .B2(U215), .ZN(U281) );
  INV_X1 U19468 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19112) );
  INV_X1 U19469 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18162) );
  AOI22_X1 U19470 ( .A1(n16370), .A2(n19112), .B1(n18162), .B2(U215), .ZN(U282) );
  INV_X1 U19471 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n16371) );
  OAI222_X1 U19472 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n16372), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(n19116), .C1(P3_DATAO_REG_31__SCAN_IN), 
        .C2(n16371), .ZN(n16373) );
  INV_X1 U19473 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18662) );
  INV_X1 U19474 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19744) );
  AOI22_X1 U19475 ( .A1(n9612), .A2(n18662), .B1(n19744), .B2(n16374), .ZN(
        U347) );
  INV_X1 U19476 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18660) );
  INV_X1 U19477 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19743) );
  AOI22_X1 U19478 ( .A1(n9612), .A2(n18660), .B1(n19743), .B2(n16374), .ZN(
        U348) );
  INV_X1 U19479 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18658) );
  INV_X1 U19480 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19741) );
  AOI22_X1 U19481 ( .A1(n9612), .A2(n18658), .B1(n19741), .B2(n16374), .ZN(
        U349) );
  INV_X1 U19482 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18656) );
  INV_X1 U19483 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19740) );
  AOI22_X1 U19484 ( .A1(n9612), .A2(n18656), .B1(n19740), .B2(n16374), .ZN(
        U350) );
  INV_X1 U19485 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18654) );
  INV_X1 U19486 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19738) );
  AOI22_X1 U19487 ( .A1(n9612), .A2(n18654), .B1(n19738), .B2(n16374), .ZN(
        U351) );
  INV_X1 U19488 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18652) );
  INV_X1 U19489 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19736) );
  AOI22_X1 U19490 ( .A1(n9612), .A2(n18652), .B1(n19736), .B2(n16374), .ZN(
        U352) );
  INV_X1 U19491 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18650) );
  INV_X1 U19492 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19735) );
  AOI22_X1 U19493 ( .A1(n9612), .A2(n18650), .B1(n19735), .B2(n16374), .ZN(
        U353) );
  INV_X1 U19494 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18647) );
  INV_X1 U19495 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19734) );
  AOI22_X1 U19496 ( .A1(n9612), .A2(n18647), .B1(n19734), .B2(n16374), .ZN(
        U354) );
  INV_X1 U19497 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18703) );
  INV_X1 U19498 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19778) );
  AOI22_X1 U19499 ( .A1(n9612), .A2(n18703), .B1(n19778), .B2(n16373), .ZN(
        U355) );
  INV_X1 U19500 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18700) );
  INV_X1 U19501 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19775) );
  AOI22_X1 U19502 ( .A1(n9612), .A2(n18700), .B1(n19775), .B2(n16374), .ZN(
        U356) );
  INV_X1 U19503 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18697) );
  INV_X1 U19504 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19773) );
  AOI22_X1 U19505 ( .A1(n9612), .A2(n18697), .B1(n19773), .B2(n16374), .ZN(
        U357) );
  INV_X1 U19506 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18696) );
  INV_X1 U19507 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19770) );
  AOI22_X1 U19508 ( .A1(n9612), .A2(n18696), .B1(n19770), .B2(n16373), .ZN(
        U358) );
  INV_X1 U19509 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18694) );
  INV_X1 U19510 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19769) );
  AOI22_X1 U19511 ( .A1(n9612), .A2(n18694), .B1(n19769), .B2(n16373), .ZN(
        U359) );
  INV_X1 U19512 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18692) );
  INV_X1 U19513 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19767) );
  AOI22_X1 U19514 ( .A1(n9612), .A2(n18692), .B1(n19767), .B2(n16373), .ZN(
        U360) );
  INV_X1 U19515 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18690) );
  INV_X1 U19516 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19765) );
  AOI22_X1 U19517 ( .A1(n9612), .A2(n18690), .B1(n19765), .B2(n16373), .ZN(
        U361) );
  INV_X1 U19518 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18688) );
  AOI22_X1 U19519 ( .A1(n9612), .A2(n18688), .B1(n19764), .B2(n16374), .ZN(
        U362) );
  INV_X1 U19520 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18686) );
  INV_X1 U19521 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19762) );
  AOI22_X1 U19522 ( .A1(n9612), .A2(n18686), .B1(n19762), .B2(n16374), .ZN(
        U363) );
  INV_X1 U19523 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18684) );
  AOI22_X1 U19524 ( .A1(n9612), .A2(n18684), .B1(n19761), .B2(n16374), .ZN(
        U364) );
  INV_X1 U19525 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18646) );
  INV_X1 U19526 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19732) );
  AOI22_X1 U19527 ( .A1(n9612), .A2(n18646), .B1(n19732), .B2(n16374), .ZN(
        U365) );
  INV_X1 U19528 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18681) );
  INV_X1 U19529 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19759) );
  AOI22_X1 U19530 ( .A1(n9612), .A2(n18681), .B1(n19759), .B2(n16374), .ZN(
        U366) );
  INV_X1 U19531 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18679) );
  INV_X1 U19532 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19757) );
  AOI22_X1 U19533 ( .A1(n9612), .A2(n18679), .B1(n19757), .B2(n16374), .ZN(
        U367) );
  INV_X1 U19534 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18678) );
  INV_X1 U19535 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19755) );
  AOI22_X1 U19536 ( .A1(n9612), .A2(n18678), .B1(n19755), .B2(n16374), .ZN(
        U368) );
  INV_X1 U19537 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18675) );
  INV_X1 U19538 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19754) );
  AOI22_X1 U19539 ( .A1(n9612), .A2(n18675), .B1(n19754), .B2(n16374), .ZN(
        U369) );
  INV_X1 U19540 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18674) );
  INV_X1 U19541 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19752) );
  AOI22_X1 U19542 ( .A1(n9612), .A2(n18674), .B1(n19752), .B2(n16374), .ZN(
        U370) );
  INV_X1 U19543 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18672) );
  INV_X1 U19544 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19751) );
  AOI22_X1 U19545 ( .A1(n9612), .A2(n18672), .B1(n19751), .B2(n16374), .ZN(
        U371) );
  INV_X1 U19546 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18669) );
  INV_X1 U19547 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19749) );
  AOI22_X1 U19548 ( .A1(n9612), .A2(n18669), .B1(n19749), .B2(n16373), .ZN(
        U372) );
  INV_X1 U19549 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18668) );
  INV_X1 U19550 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19748) );
  AOI22_X1 U19551 ( .A1(n9612), .A2(n18668), .B1(n19748), .B2(n16374), .ZN(
        U373) );
  INV_X1 U19552 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18666) );
  AOI22_X1 U19553 ( .A1(n9612), .A2(n18666), .B1(n19747), .B2(n16373), .ZN(
        U374) );
  INV_X1 U19554 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18664) );
  INV_X1 U19555 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19746) );
  AOI22_X1 U19556 ( .A1(n9612), .A2(n18664), .B1(n19746), .B2(n16373), .ZN(
        U375) );
  INV_X1 U19557 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18644) );
  AOI22_X1 U19558 ( .A1(n9612), .A2(n18644), .B1(n19730), .B2(n16374), .ZN(
        U376) );
  INV_X1 U19559 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18643) );
  NAND2_X1 U19560 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18643), .ZN(n18632) );
  AOI22_X1 U19561 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18632), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18629), .ZN(n18715) );
  AOI21_X1 U19562 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18715), .ZN(n16375) );
  INV_X1 U19563 ( .A(n16375), .ZN(P3_U2633) );
  INV_X1 U19564 ( .A(n18729), .ZN(n18780) );
  NAND2_X1 U19565 ( .A1(n18780), .A2(n18779), .ZN(n16377) );
  OAI21_X1 U19566 ( .B1(n16382), .B2(n17345), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16376) );
  OAI21_X1 U19567 ( .B1(n16377), .B2(n18767), .A(n16376), .ZN(P3_U2634) );
  AOI21_X1 U19568 ( .B1(n18628), .B2(n18643), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16378) );
  AOI22_X1 U19569 ( .A1(n18758), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16378), 
        .B2(n18777), .ZN(P3_U2635) );
  INV_X1 U19570 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16406) );
  OAI21_X1 U19571 ( .B1(n16379), .B2(BS16), .A(n18715), .ZN(n18713) );
  OAI21_X1 U19572 ( .B1(n18715), .B2(n16406), .A(n18713), .ZN(P3_U2636) );
  NOR3_X1 U19573 ( .A1(n16382), .A2(n16381), .A3(n16380), .ZN(n18556) );
  NOR2_X1 U19574 ( .A1(n18556), .A2(n18617), .ZN(n18760) );
  OAI21_X1 U19575 ( .B1(n18760), .B2(n18114), .A(n16383), .ZN(P3_U2637) );
  NOR4_X1 U19576 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16387) );
  NOR4_X1 U19577 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16386) );
  NOR4_X1 U19578 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16385) );
  NOR4_X1 U19579 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16384) );
  NAND4_X1 U19580 ( .A1(n16387), .A2(n16386), .A3(n16385), .A4(n16384), .ZN(
        n16393) );
  NOR4_X1 U19581 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16391) );
  AOI211_X1 U19582 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_11__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16390) );
  NOR4_X1 U19583 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16389) );
  NOR4_X1 U19584 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16388) );
  NAND4_X1 U19585 ( .A1(n16391), .A2(n16390), .A3(n16389), .A4(n16388), .ZN(
        n16392) );
  NOR2_X1 U19586 ( .A1(n16393), .A2(n16392), .ZN(n18757) );
  INV_X1 U19587 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16395) );
  NOR3_X1 U19588 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16396) );
  OAI21_X1 U19589 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16396), .A(n18757), .ZN(
        n16394) );
  OAI21_X1 U19590 ( .B1(n18757), .B2(n16395), .A(n16394), .ZN(P3_U2638) );
  INV_X1 U19591 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18750) );
  INV_X1 U19592 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18714) );
  AOI21_X1 U19593 ( .B1(n18750), .B2(n18714), .A(n16396), .ZN(n16398) );
  INV_X1 U19594 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16397) );
  INV_X1 U19595 ( .A(n18757), .ZN(n18752) );
  AOI22_X1 U19596 ( .A1(n18757), .A2(n16398), .B1(n16397), .B2(n18752), .ZN(
        P3_U2639) );
  NAND2_X1 U19597 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18726), .ZN(n16400) );
  NOR2_X1 U19598 ( .A1(n18743), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18487) );
  INV_X1 U19599 ( .A(n18487), .ZN(n18613) );
  NOR3_X1 U19600 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18625) );
  NAND2_X1 U19601 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18625), .ZN(n16764) );
  NAND2_X1 U19602 ( .A1(n17988), .A2(n16764), .ZN(n16737) );
  INV_X1 U19603 ( .A(n16737), .ZN(n16638) );
  AOI211_X1 U19604 ( .C1(n18635), .C2(n17348), .A(n18764), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16402) );
  NAND2_X1 U19605 ( .A1(n18782), .A2(n18125), .ZN(n16405) );
  AOI211_X1 U19606 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18128), .A(n16402), .B(
        n16405), .ZN(n16401) );
  INV_X1 U19607 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18704) );
  INV_X1 U19608 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18695) );
  INV_X1 U19609 ( .A(n16402), .ZN(n18610) );
  INV_X1 U19610 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18693) );
  INV_X1 U19611 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18691) );
  INV_X1 U19612 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18683) );
  INV_X1 U19613 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18687) );
  INV_X1 U19614 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18685) );
  INV_X1 U19615 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18676) );
  INV_X1 U19616 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18667) );
  INV_X1 U19617 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18663) );
  INV_X1 U19618 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18659) );
  INV_X1 U19619 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18655) );
  NAND3_X1 U19620 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16696) );
  NAND3_X1 U19621 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(P3_REIP_REG_5__SCAN_IN), 
        .A3(P3_REIP_REG_4__SCAN_IN), .ZN(n16697) );
  NOR3_X1 U19622 ( .A1(n18655), .A2(n16696), .A3(n16697), .ZN(n16679) );
  NAND2_X1 U19623 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16679), .ZN(n16664) );
  NOR2_X1 U19624 ( .A1(n18659), .A2(n16664), .ZN(n16665) );
  NAND2_X1 U19625 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16665), .ZN(n16649) );
  NOR2_X1 U19626 ( .A1(n18663), .A2(n16649), .ZN(n16642) );
  NAND2_X1 U19627 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16642), .ZN(n16621) );
  NOR2_X1 U19628 ( .A1(n18667), .A2(n16621), .ZN(n16608) );
  NAND2_X1 U19629 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16608), .ZN(n16586) );
  NAND2_X1 U19630 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16587) );
  NOR3_X1 U19631 ( .A1(n18676), .A2(n16586), .A3(n16587), .ZN(n16571) );
  NAND4_X1 U19632 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16571), .A3(
        P3_REIP_REG_20__SCAN_IN), .A4(P3_REIP_REG_18__SCAN_IN), .ZN(n16515) );
  NOR4_X1 U19633 ( .A1(n18683), .A2(n18687), .A3(n18685), .A4(n16515), .ZN(
        n16495) );
  NAND2_X1 U19634 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16495), .ZN(n16471) );
  NOR3_X1 U19635 ( .A1(n18693), .A2(n18691), .A3(n16471), .ZN(n16419) );
  NAND2_X1 U19636 ( .A1(n16770), .A2(n16419), .ZN(n16465) );
  NOR2_X1 U19637 ( .A1(n18695), .A2(n16465), .ZN(n16451) );
  NAND3_X1 U19638 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(n16451), .ZN(n16421) );
  NOR3_X1 U19639 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18704), .A3(n16421), 
        .ZN(n16403) );
  AOI21_X1 U19640 ( .B1(n16758), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16403), .ZN(
        n16427) );
  NAND2_X1 U19641 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18128), .ZN(n16404) );
  AOI211_X4 U19642 ( .C1(n16406), .C2(n18773), .A(n16405), .B(n16404), .ZN(
        n16790) );
  NOR3_X1 U19643 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16762) );
  NAND2_X1 U19644 ( .A1(n16762), .A2(n17132), .ZN(n16752) );
  NOR2_X1 U19645 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16752), .ZN(n16731) );
  NAND2_X1 U19646 ( .A1(n16731), .A2(n16728), .ZN(n16727) );
  NOR2_X1 U19647 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16727), .ZN(n16706) );
  INV_X1 U19648 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16703) );
  NAND2_X1 U19649 ( .A1(n16706), .A2(n16703), .ZN(n16702) );
  NOR2_X1 U19650 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16702), .ZN(n16675) );
  INV_X1 U19651 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16407) );
  NAND2_X1 U19652 ( .A1(n16675), .A2(n16407), .ZN(n16658) );
  INV_X1 U19653 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16961) );
  NAND2_X1 U19654 ( .A1(n16657), .A2(n16961), .ZN(n16653) );
  INV_X1 U19655 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16627) );
  NAND2_X1 U19656 ( .A1(n16632), .A2(n16627), .ZN(n16626) );
  NAND2_X1 U19657 ( .A1(n16611), .A2(n16598), .ZN(n16596) );
  NAND2_X1 U19658 ( .A1(n16585), .A2(n16930), .ZN(n16578) );
  NAND2_X1 U19659 ( .A1(n16563), .A2(n16902), .ZN(n16553) );
  NOR2_X1 U19660 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16553), .ZN(n16540) );
  NAND2_X1 U19661 ( .A1(n16540), .A2(n16887), .ZN(n16534) );
  NOR2_X1 U19662 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16534), .ZN(n16518) );
  NAND2_X1 U19663 ( .A1(n16518), .A2(n16855), .ZN(n16511) );
  NOR2_X1 U19664 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16511), .ZN(n16498) );
  INV_X1 U19665 ( .A(n16498), .ZN(n16484) );
  NOR2_X1 U19666 ( .A1(n16484), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n16483) );
  INV_X1 U19667 ( .A(n16483), .ZN(n16473) );
  NOR2_X1 U19668 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16473), .ZN(n16472) );
  NAND2_X1 U19669 ( .A1(n16472), .A2(n16840), .ZN(n16468) );
  NOR2_X1 U19670 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16468), .ZN(n16453) );
  INV_X1 U19671 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16831) );
  NAND2_X1 U19672 ( .A1(n16453), .A2(n16831), .ZN(n16429) );
  NOR2_X1 U19673 ( .A1(n16782), .A2(n16429), .ZN(n16436) );
  INV_X1 U19674 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16425) );
  INV_X1 U19675 ( .A(n16411), .ZN(n16410) );
  INV_X1 U19676 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17438) );
  NOR2_X1 U19677 ( .A1(n16410), .A2(n17438), .ZN(n16409) );
  OAI21_X1 U19678 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16409), .A(
        n16408), .ZN(n17424) );
  INV_X1 U19679 ( .A(n17424), .ZN(n16456) );
  AOI21_X1 U19680 ( .B1(n16410), .B2(n17438), .A(n16409), .ZN(n17433) );
  INV_X1 U19681 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16476) );
  OR2_X1 U19682 ( .A1(n17763), .A2(n17458), .ZN(n16414) );
  NOR2_X1 U19683 ( .A1(n17459), .A2(n16414), .ZN(n17416) );
  INV_X1 U19684 ( .A(n17416), .ZN(n16412) );
  AOI21_X1 U19685 ( .B1(n16476), .B2(n16412), .A(n16411), .ZN(n17450) );
  INV_X1 U19686 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17471) );
  NOR2_X1 U19687 ( .A1(n17471), .A2(n16414), .ZN(n16413) );
  OAI21_X1 U19688 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16413), .A(
        n16412), .ZN(n17461) );
  INV_X1 U19689 ( .A(n17461), .ZN(n16487) );
  AOI21_X1 U19690 ( .B1(n17471), .B2(n16414), .A(n16413), .ZN(n17469) );
  NOR2_X1 U19691 ( .A1(n17763), .A2(n17497), .ZN(n16416) );
  INV_X1 U19692 ( .A(n16416), .ZN(n16417) );
  NOR2_X1 U19693 ( .A1(n17498), .A2(n16417), .ZN(n17456) );
  OAI21_X1 U19694 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17456), .A(
        n16414), .ZN(n17485) );
  INV_X1 U19695 ( .A(n17485), .ZN(n16507) );
  INV_X1 U19696 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16520) );
  NAND2_X1 U19697 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16416), .ZN(
        n16415) );
  AOI21_X1 U19698 ( .B1(n16520), .B2(n16415), .A(n17456), .ZN(n17496) );
  INV_X1 U19699 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17509) );
  AOI22_X1 U19700 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16417), .B1(
        n16416), .B2(n17509), .ZN(n17506) );
  INV_X1 U19701 ( .A(n17506), .ZN(n16531) );
  INV_X1 U19702 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16556) );
  NAND3_X1 U19703 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17589), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16606) );
  NOR2_X1 U19704 ( .A1(n17566), .A2(n16606), .ZN(n16582) );
  NAND2_X1 U19705 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16582), .ZN(
        n16569) );
  INV_X1 U19706 ( .A(n16569), .ZN(n17530) );
  NAND2_X1 U19707 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17530), .ZN(
        n16557) );
  NOR2_X1 U19708 ( .A1(n16556), .A2(n16557), .ZN(n17495) );
  OAI21_X1 U19709 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17495), .A(
        n16417), .ZN(n16418) );
  INV_X1 U19710 ( .A(n16418), .ZN(n17520) );
  INV_X1 U19711 ( .A(n16606), .ZN(n17563) );
  NAND2_X1 U19712 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17563), .ZN(
        n16595) );
  NOR2_X1 U19713 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16595), .ZN(
        n16591) );
  NOR2_X1 U19714 ( .A1(n17520), .A2(n16538), .ZN(n16537) );
  NOR2_X1 U19715 ( .A1(n16537), .A2(n16692), .ZN(n16530) );
  NOR2_X1 U19716 ( .A1(n16531), .A2(n16530), .ZN(n16529) );
  NOR2_X1 U19717 ( .A1(n16529), .A2(n16692), .ZN(n16517) );
  NOR2_X1 U19718 ( .A1(n17496), .A2(n16517), .ZN(n16516) );
  NOR2_X1 U19719 ( .A1(n16516), .A2(n16692), .ZN(n16506) );
  NOR2_X1 U19720 ( .A1(n16507), .A2(n16506), .ZN(n16505) );
  NOR2_X1 U19721 ( .A1(n16505), .A2(n16692), .ZN(n16497) );
  NOR2_X1 U19722 ( .A1(n17469), .A2(n16497), .ZN(n16496) );
  NOR2_X1 U19723 ( .A1(n16496), .A2(n16692), .ZN(n16486) );
  NOR2_X1 U19724 ( .A1(n16487), .A2(n16486), .ZN(n16485) );
  NOR2_X1 U19725 ( .A1(n16485), .A2(n16692), .ZN(n16475) );
  NOR2_X1 U19726 ( .A1(n17450), .A2(n16475), .ZN(n16474) );
  NOR2_X1 U19727 ( .A1(n16474), .A2(n16692), .ZN(n16464) );
  NOR2_X1 U19728 ( .A1(n17433), .A2(n16464), .ZN(n16463) );
  NOR2_X1 U19729 ( .A1(n16463), .A2(n16692), .ZN(n16455) );
  NOR2_X1 U19730 ( .A1(n16456), .A2(n16455), .ZN(n16454) );
  NOR2_X1 U19731 ( .A1(n16454), .A2(n16692), .ZN(n16440) );
  NOR2_X1 U19732 ( .A1(n16441), .A2(n16440), .ZN(n16439) );
  NOR2_X1 U19733 ( .A1(n16439), .A2(n16692), .ZN(n16430) );
  INV_X1 U19734 ( .A(n16764), .ZN(n18620) );
  NAND2_X1 U19735 ( .A1(n16749), .A2(n18620), .ZN(n16778) );
  NOR3_X1 U19736 ( .A1(n16431), .A2(n16430), .A3(n16778), .ZN(n16424) );
  NAND2_X1 U19737 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .ZN(n16420) );
  NAND2_X1 U19738 ( .A1(n16792), .A2(n16789), .ZN(n16791) );
  OAI21_X1 U19739 ( .B1(n16419), .B2(n16789), .A(n16792), .ZN(n16452) );
  AOI221_X1 U19740 ( .B1(n16420), .B2(n16791), .C1(n18695), .C2(n16791), .A(
        n16452), .ZN(n16450) );
  NOR2_X1 U19741 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16421), .ZN(n16434) );
  INV_X1 U19742 ( .A(n16434), .ZN(n16422) );
  AOI21_X1 U19743 ( .B1(n16450), .B2(n16422), .A(n18702), .ZN(n16423) );
  AOI211_X1 U19744 ( .C1(n16436), .C2(n16425), .A(n16424), .B(n16423), .ZN(
        n16426) );
  OAI211_X1 U19745 ( .C1(n16428), .C2(n16777), .A(n16427), .B(n16426), .ZN(
        P3_U2640) );
  NAND2_X1 U19746 ( .A1(n16790), .A2(n16429), .ZN(n16446) );
  XOR2_X1 U19747 ( .A(n16431), .B(n16430), .Z(n16435) );
  OAI22_X1 U19748 ( .A1(n16450), .A2(n18704), .B1(n16432), .B2(n16777), .ZN(
        n16433) );
  AOI211_X1 U19749 ( .C1(n16435), .C2(n18620), .A(n16434), .B(n16433), .ZN(
        n16438) );
  OAI21_X1 U19750 ( .B1(n16401), .B2(n16436), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16437) );
  INV_X1 U19751 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18699) );
  AOI211_X1 U19752 ( .C1(n16441), .C2(n16440), .A(n16439), .B(n16764), .ZN(
        n16445) );
  NAND2_X1 U19753 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16451), .ZN(n16443) );
  OAI22_X1 U19754 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16443), .B1(n16442), 
        .B2(n16777), .ZN(n16444) );
  AOI211_X1 U19755 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16758), .A(n16445), .B(
        n16444), .ZN(n16449) );
  INV_X1 U19756 ( .A(n16446), .ZN(n16447) );
  OAI21_X1 U19757 ( .B1(n16453), .B2(n16831), .A(n16447), .ZN(n16448) );
  OAI211_X1 U19758 ( .C1(n16450), .C2(n18699), .A(n16449), .B(n16448), .ZN(
        P3_U2642) );
  INV_X1 U19759 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16462) );
  INV_X1 U19760 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18698) );
  AOI22_X1 U19761 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16758), .B1(n16451), 
        .B2(n18698), .ZN(n16461) );
  INV_X1 U19762 ( .A(n16452), .ZN(n16481) );
  OAI21_X1 U19763 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16465), .A(n16481), 
        .ZN(n16459) );
  AOI211_X1 U19764 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16468), .A(n16453), .B(
        n16782), .ZN(n16458) );
  AOI211_X1 U19765 ( .C1(n16456), .C2(n16455), .A(n16454), .B(n16764), .ZN(
        n16457) );
  AOI211_X1 U19766 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16459), .A(n16458), 
        .B(n16457), .ZN(n16460) );
  OAI211_X1 U19767 ( .C1(n16462), .C2(n16777), .A(n16461), .B(n16460), .ZN(
        P3_U2643) );
  AOI211_X1 U19768 ( .C1(n17433), .C2(n16464), .A(n16463), .B(n16764), .ZN(
        n16467) );
  OAI22_X1 U19769 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16465), .B1(n17438), 
        .B2(n16777), .ZN(n16466) );
  AOI211_X1 U19770 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16758), .A(n16467), .B(
        n16466), .ZN(n16470) );
  OAI211_X1 U19771 ( .C1(n16472), .C2(n16840), .A(n16790), .B(n16468), .ZN(
        n16469) );
  OAI211_X1 U19772 ( .C1(n16481), .C2(n18695), .A(n16470), .B(n16469), .ZN(
        P3_U2644) );
  NOR2_X1 U19773 ( .A1(n16789), .A2(n16471), .ZN(n16490) );
  AOI21_X1 U19774 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n16490), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n16482) );
  AOI211_X1 U19775 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16473), .A(n16472), .B(
        n16782), .ZN(n16479) );
  AOI211_X1 U19776 ( .C1(n17450), .C2(n16475), .A(n16474), .B(n16764), .ZN(
        n16478) );
  INV_X1 U19777 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16844) );
  OAI22_X1 U19778 ( .A1(n16476), .A2(n16777), .B1(n16783), .B2(n16844), .ZN(
        n16477) );
  NOR3_X1 U19779 ( .A1(n16479), .A2(n16478), .A3(n16477), .ZN(n16480) );
  OAI21_X1 U19780 ( .B1(n16482), .B2(n16481), .A(n16480), .ZN(P3_U2645) );
  INV_X1 U19781 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18689) );
  OAI21_X1 U19782 ( .B1(n16495), .B2(n16789), .A(n16792), .ZN(n16509) );
  AOI21_X1 U19783 ( .B1(n16770), .B2(n18689), .A(n16509), .ZN(n16493) );
  AOI22_X1 U19784 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16761), .B1(
        n16758), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16492) );
  AOI211_X1 U19785 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n16484), .A(n16483), .B(
        n16782), .ZN(n16489) );
  AOI211_X1 U19786 ( .C1(n16487), .C2(n16486), .A(n16485), .B(n16764), .ZN(
        n16488) );
  AOI211_X1 U19787 ( .C1(n16490), .C2(n18691), .A(n16489), .B(n16488), .ZN(
        n16491) );
  OAI211_X1 U19788 ( .C1(n16493), .C2(n18691), .A(n16492), .B(n16491), .ZN(
        P3_U2646) );
  INV_X1 U19789 ( .A(n16509), .ZN(n16503) );
  NOR2_X1 U19790 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16789), .ZN(n16494) );
  AOI22_X1 U19791 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16761), .B1(
        n16495), .B2(n16494), .ZN(n16502) );
  AOI211_X1 U19792 ( .C1(n17469), .C2(n16497), .A(n16496), .B(n16764), .ZN(
        n16500) );
  AOI211_X1 U19793 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16511), .A(n16498), .B(
        n16782), .ZN(n16499) );
  AOI211_X1 U19794 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16758), .A(n16500), .B(
        n16499), .ZN(n16501) );
  OAI211_X1 U19795 ( .C1(n16503), .C2(n18689), .A(n16502), .B(n16501), .ZN(
        P3_U2647) );
  AOI22_X1 U19796 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16761), .B1(
        n16758), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n16514) );
  NAND3_X1 U19797 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_20__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .ZN(n16504) );
  NAND2_X1 U19798 ( .A1(n16770), .A2(n16571), .ZN(n16562) );
  NOR2_X1 U19799 ( .A1(n16504), .A2(n16562), .ZN(n16526) );
  NAND2_X1 U19800 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16526), .ZN(n16525) );
  NOR2_X1 U19801 ( .A1(n18685), .A2(n16525), .ZN(n16510) );
  AOI211_X1 U19802 ( .C1(n16507), .C2(n16506), .A(n16505), .B(n16764), .ZN(
        n16508) );
  AOI221_X1 U19803 ( .B1(n16510), .B2(n18687), .C1(n16509), .C2(
        P3_REIP_REG_23__SCAN_IN), .A(n16508), .ZN(n16513) );
  OAI211_X1 U19804 ( .C1(n16518), .C2(n16855), .A(n16790), .B(n16511), .ZN(
        n16512) );
  NAND3_X1 U19805 ( .A1(n16514), .A2(n16513), .A3(n16512), .ZN(P3_U2648) );
  OR2_X1 U19806 ( .A1(n16515), .A2(n16776), .ZN(n16542) );
  OAI21_X1 U19807 ( .B1(n18683), .B2(n16542), .A(n16791), .ZN(n16527) );
  AOI211_X1 U19808 ( .C1(n17496), .C2(n16517), .A(n16516), .B(n16764), .ZN(
        n16523) );
  AOI211_X1 U19809 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16534), .A(n16518), .B(
        n16782), .ZN(n16522) );
  OAI22_X1 U19810 ( .A1(n16520), .A2(n16777), .B1(n16783), .B2(n16519), .ZN(
        n16521) );
  NOR3_X1 U19811 ( .A1(n16523), .A2(n16522), .A3(n16521), .ZN(n16524) );
  OAI221_X1 U19812 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(n16525), .C1(n18685), 
        .C2(n16527), .A(n16524), .ZN(P3_U2649) );
  INV_X1 U19813 ( .A(n16526), .ZN(n16528) );
  AOI21_X1 U19814 ( .B1(n18683), .B2(n16528), .A(n16527), .ZN(n16533) );
  AOI211_X1 U19815 ( .C1(n16531), .C2(n16530), .A(n16529), .B(n16764), .ZN(
        n16532) );
  AOI211_X1 U19816 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n16758), .A(n16533), .B(
        n16532), .ZN(n16536) );
  OAI211_X1 U19817 ( .C1(n16540), .C2(n16887), .A(n16790), .B(n16534), .ZN(
        n16535) );
  OAI211_X1 U19818 ( .C1(n16777), .C2(n17509), .A(n16536), .B(n16535), .ZN(
        P3_U2650) );
  AOI211_X1 U19819 ( .C1(n17520), .C2(n16538), .A(n16537), .B(n16764), .ZN(
        n16539) );
  AOI21_X1 U19820 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16401), .A(n16539), .ZN(
        n16546) );
  AOI211_X1 U19821 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16553), .A(n16540), .B(
        n16782), .ZN(n16541) );
  AOI21_X1 U19822 ( .B1(n16761), .B2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16541), .ZN(n16545) );
  NAND3_X1 U19823 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16791), .A3(n16542), 
        .ZN(n16544) );
  INV_X1 U19824 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18677) );
  NOR2_X1 U19825 ( .A1(n18677), .A2(n16562), .ZN(n16552) );
  INV_X1 U19826 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18682) );
  NAND3_X1 U19827 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16552), .A3(n18682), 
        .ZN(n16543) );
  NAND4_X1 U19828 ( .A1(n16546), .A2(n16545), .A3(n16544), .A4(n16543), .ZN(
        P3_U2651) );
  INV_X1 U19829 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18680) );
  OAI221_X1 U19830 ( .B1(n16789), .B2(n16571), .C1(n16789), .C2(
        P3_REIP_REG_18__SCAN_IN), .A(n16792), .ZN(n16566) );
  AOI21_X1 U19831 ( .B1(n16556), .B2(n16557), .A(n17495), .ZN(n16547) );
  INV_X1 U19832 ( .A(n16547), .ZN(n17534) );
  INV_X1 U19833 ( .A(n16591), .ZN(n16548) );
  OAI21_X1 U19834 ( .B1(n16557), .B2(n16548), .A(n16749), .ZN(n16560) );
  AOI21_X1 U19835 ( .B1(n17534), .B2(n16560), .A(n16764), .ZN(n16549) );
  OAI21_X1 U19836 ( .B1(n17534), .B2(n16560), .A(n16549), .ZN(n16550) );
  OAI211_X1 U19837 ( .C1(n16783), .C2(n16902), .A(n17988), .B(n16550), .ZN(
        n16551) );
  AOI221_X1 U19838 ( .B1(n16552), .B2(n18680), .C1(n16566), .C2(
        P3_REIP_REG_19__SCAN_IN), .A(n16551), .ZN(n16555) );
  OAI211_X1 U19839 ( .C1(n16563), .C2(n16902), .A(n16790), .B(n16553), .ZN(
        n16554) );
  OAI211_X1 U19840 ( .C1(n16777), .C2(n16556), .A(n16555), .B(n16554), .ZN(
        P3_U2652) );
  INV_X1 U19841 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17543) );
  OAI21_X1 U19842 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17530), .A(
        n16557), .ZN(n17540) );
  NOR2_X1 U19843 ( .A1(n16764), .A2(n16749), .ZN(n16768) );
  INV_X1 U19844 ( .A(n16768), .ZN(n16559) );
  OAI221_X1 U19845 ( .B1(n17540), .B2(n16591), .C1(n17540), .C2(n17543), .A(
        n18620), .ZN(n16558) );
  AOI22_X1 U19846 ( .A1(n17540), .A2(n16560), .B1(n16559), .B2(n16558), .ZN(
        n16561) );
  AOI211_X1 U19847 ( .C1(n16758), .C2(P3_EBX_REG_18__SCAN_IN), .A(n9611), .B(
        n16561), .ZN(n16568) );
  INV_X1 U19848 ( .A(n16562), .ZN(n16565) );
  AOI211_X1 U19849 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16578), .A(n16563), .B(
        n16782), .ZN(n16564) );
  AOI221_X1 U19850 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16566), .C1(n16565), 
        .C2(n16566), .A(n16564), .ZN(n16567) );
  OAI211_X1 U19851 ( .C1(n17543), .C2(n16777), .A(n16568), .B(n16567), .ZN(
        P3_U2653) );
  AOI22_X1 U19852 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16761), .B1(
        n16758), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16581) );
  OAI21_X1 U19853 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16582), .A(
        n16569), .ZN(n17552) );
  AOI21_X1 U19854 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16591), .A(
        n16692), .ZN(n16570) );
  XNOR2_X1 U19855 ( .A(n17552), .B(n16570), .ZN(n16577) );
  NAND3_X1 U19856 ( .A1(n16770), .A2(P3_REIP_REG_14__SCAN_IN), .A3(n16608), 
        .ZN(n16605) );
  NOR2_X1 U19857 ( .A1(n16587), .A2(n16605), .ZN(n16575) );
  INV_X1 U19858 ( .A(n16571), .ZN(n16572) );
  AOI21_X1 U19859 ( .B1(n16770), .B2(n16572), .A(n16776), .ZN(n16573) );
  INV_X1 U19860 ( .A(n16573), .ZN(n16574) );
  MUX2_X1 U19861 ( .A(n16575), .B(n16574), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n16576) );
  AOI211_X1 U19862 ( .C1(n18620), .C2(n16577), .A(n9611), .B(n16576), .ZN(
        n16580) );
  OAI211_X1 U19863 ( .C1(n16585), .C2(n16930), .A(n16790), .B(n16578), .ZN(
        n16579) );
  NAND3_X1 U19864 ( .A1(n16581), .A2(n16580), .A3(n16579), .ZN(P3_U2654) );
  NOR2_X1 U19865 ( .A1(n16591), .A2(n16778), .ZN(n16603) );
  INV_X1 U19866 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16583) );
  AOI21_X1 U19867 ( .B1(n16583), .B2(n16595), .A(n16582), .ZN(n17564) );
  INV_X1 U19868 ( .A(n17564), .ZN(n16584) );
  AOI22_X1 U19869 ( .A1(n16758), .A2(P3_EBX_REG_16__SCAN_IN), .B1(n16603), 
        .B2(n16584), .ZN(n16594) );
  AOI211_X1 U19870 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16596), .A(n16585), .B(
        n16782), .ZN(n16590) );
  AOI21_X1 U19871 ( .B1(n16770), .B2(n16586), .A(n16776), .ZN(n16609) );
  INV_X1 U19872 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18673) );
  OAI21_X1 U19873 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(P3_REIP_REG_15__SCAN_IN), 
        .A(n16587), .ZN(n16588) );
  OAI22_X1 U19874 ( .A1(n16609), .A2(n18673), .B1(n16605), .B2(n16588), .ZN(
        n16589) );
  AOI211_X1 U19875 ( .C1(n16761), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16590), .B(n16589), .ZN(n16593) );
  OAI211_X1 U19876 ( .C1(n16591), .C2(n16692), .A(n18620), .B(n17564), .ZN(
        n16592) );
  NAND4_X1 U19877 ( .A1(n16594), .A2(n16593), .A3(n17988), .A4(n16592), .ZN(
        P3_U2655) );
  INV_X1 U19878 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18671) );
  OAI21_X1 U19879 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17563), .A(
        n16595), .ZN(n17574) );
  OAI211_X1 U19880 ( .C1(n16611), .C2(n16598), .A(n16790), .B(n16596), .ZN(
        n16597) );
  OAI21_X1 U19881 ( .B1(n16783), .B2(n16598), .A(n16597), .ZN(n16602) );
  INV_X1 U19882 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17577) );
  INV_X1 U19883 ( .A(n17574), .ZN(n16599) );
  AOI21_X1 U19884 ( .B1(n16749), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16764), .ZN(n16785) );
  OAI211_X1 U19885 ( .C1(n17577), .C2(n16692), .A(n16599), .B(n16785), .ZN(
        n16600) );
  OAI211_X1 U19886 ( .C1(n17577), .C2(n16777), .A(n17988), .B(n16600), .ZN(
        n16601) );
  AOI211_X1 U19887 ( .C1(n16603), .C2(n17574), .A(n16602), .B(n16601), .ZN(
        n16604) );
  OAI221_X1 U19888 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16605), .C1(n18671), 
        .C2(n16609), .A(n16604), .ZN(P3_U2656) );
  AND2_X1 U19889 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17589), .ZN(
        n16618) );
  OAI21_X1 U19890 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16618), .A(
        n16606), .ZN(n17590) );
  NAND2_X1 U19891 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17673), .ZN(
        n16645) );
  INV_X1 U19892 ( .A(n16645), .ZN(n16694) );
  NAND2_X1 U19893 ( .A1(n16607), .A2(n16694), .ZN(n17601) );
  OAI21_X1 U19894 ( .B1(n17601), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16749), .ZN(n16635) );
  INV_X1 U19895 ( .A(n16635), .ZN(n16634) );
  AOI21_X1 U19896 ( .B1(n16749), .B2(n17613), .A(n16634), .ZN(n16620) );
  XNOR2_X1 U19897 ( .A(n17590), .B(n16620), .ZN(n16617) );
  INV_X1 U19898 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18670) );
  NAND2_X1 U19899 ( .A1(n16770), .A2(n16608), .ZN(n16610) );
  AOI21_X1 U19900 ( .B1(n18670), .B2(n16610), .A(n16609), .ZN(n16615) );
  AOI211_X1 U19901 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16626), .A(n16611), .B(
        n16782), .ZN(n16614) );
  AOI22_X1 U19902 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16761), .B1(
        n16401), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n16612) );
  INV_X1 U19903 ( .A(n16612), .ZN(n16613) );
  NOR4_X1 U19904 ( .A1(n9611), .A2(n16615), .A3(n16614), .A4(n16613), .ZN(
        n16616) );
  OAI21_X1 U19905 ( .B1(n16617), .B2(n16764), .A(n16616), .ZN(P3_U2657) );
  INV_X1 U19906 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16622) );
  INV_X1 U19907 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17619) );
  NOR2_X1 U19908 ( .A1(n17619), .A2(n17601), .ZN(n16633) );
  INV_X1 U19909 ( .A(n16633), .ZN(n16619) );
  AOI21_X1 U19910 ( .B1(n16622), .B2(n16619), .A(n16618), .ZN(n17604) );
  NOR3_X1 U19911 ( .A1(n17604), .A2(n16620), .A3(n16764), .ZN(n16625) );
  NOR3_X1 U19912 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16789), .A3(n16621), 
        .ZN(n16624) );
  OAI22_X1 U19913 ( .A1(n16622), .A2(n16777), .B1(n16783), .B2(n16627), .ZN(
        n16623) );
  NOR4_X1 U19914 ( .A1(n9611), .A2(n16625), .A3(n16624), .A4(n16623), .ZN(
        n16631) );
  OAI21_X1 U19915 ( .B1(n16642), .B2(n16789), .A(n16792), .ZN(n16651) );
  NOR2_X1 U19916 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16789), .ZN(n16641) );
  OAI21_X1 U19917 ( .B1(n16651), .B2(n16641), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16630) );
  OAI211_X1 U19918 ( .C1(n16632), .C2(n16627), .A(n16790), .B(n16626), .ZN(
        n16629) );
  OAI211_X1 U19919 ( .C1(n16633), .C2(n16768), .A(n17604), .B(n16785), .ZN(
        n16628) );
  NAND4_X1 U19920 ( .A1(n16631), .A2(n16630), .A3(n16629), .A4(n16628), .ZN(
        P3_U2658) );
  AOI211_X1 U19921 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16653), .A(n16632), .B(
        n16782), .ZN(n16640) );
  AOI21_X1 U19922 ( .B1(n17619), .B2(n17601), .A(n16633), .ZN(n16636) );
  INV_X1 U19923 ( .A(n16636), .ZN(n17630) );
  AOI221_X1 U19924 ( .B1(n16636), .B2(n16635), .C1(n17630), .C2(n16634), .A(
        n9611), .ZN(n16637) );
  OAI22_X1 U19925 ( .A1(n16638), .A2(n16637), .B1(n17619), .B2(n16777), .ZN(
        n16639) );
  AOI211_X1 U19926 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16758), .A(n16640), .B(
        n16639), .ZN(n16644) );
  AOI22_X1 U19927 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16651), .B1(n16642), 
        .B2(n16641), .ZN(n16643) );
  NAND2_X1 U19928 ( .A1(n16644), .A2(n16643), .ZN(P3_U2659) );
  AOI22_X1 U19929 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16761), .B1(
        n16758), .B2(P3_EBX_REG_11__SCAN_IN), .ZN(n16656) );
  OR2_X1 U19930 ( .A1(n16647), .A2(n16645), .ZN(n16659) );
  INV_X1 U19931 ( .A(n17601), .ZN(n16646) );
  AOI21_X1 U19932 ( .B1(n17638), .B2(n16659), .A(n16646), .ZN(n17632) );
  INV_X1 U19933 ( .A(n17699), .ZN(n17703) );
  NOR2_X1 U19934 ( .A1(n17763), .A2(n17703), .ZN(n16722) );
  NAND2_X1 U19935 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16722), .ZN(
        n16712) );
  NOR2_X1 U19936 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16712), .ZN(
        n16693) );
  AOI21_X1 U19937 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16693), .A(
        n16692), .ZN(n16682) );
  AOI21_X1 U19938 ( .B1(n16749), .B2(n16647), .A(n16682), .ZN(n16648) );
  XNOR2_X1 U19939 ( .A(n17632), .B(n16648), .ZN(n16652) );
  OAI21_X1 U19940 ( .B1(n16789), .B2(n16649), .A(n18663), .ZN(n16650) );
  AOI22_X1 U19941 ( .A1(n18620), .A2(n16652), .B1(n16651), .B2(n16650), .ZN(
        n16655) );
  OAI211_X1 U19942 ( .C1(n16657), .C2(n16961), .A(n16790), .B(n16653), .ZN(
        n16654) );
  NAND4_X1 U19943 ( .A1(n16656), .A2(n16655), .A3(n17988), .A4(n16654), .ZN(
        P3_U2660) );
  AOI211_X1 U19944 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16658), .A(n16657), .B(
        n16782), .ZN(n16663) );
  INV_X1 U19945 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17657) );
  NAND2_X1 U19946 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17672) );
  OR2_X1 U19947 ( .A1(n17672), .A2(n16712), .ZN(n16680) );
  NOR2_X1 U19948 ( .A1(n17657), .A2(n16680), .ZN(n16669) );
  OAI21_X1 U19949 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16669), .A(
        n16659), .ZN(n16660) );
  INV_X1 U19950 ( .A(n16660), .ZN(n17645) );
  INV_X1 U19951 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16779) );
  AOI21_X1 U19952 ( .B1(n16669), .B2(n16779), .A(n16692), .ZN(n16670) );
  XNOR2_X1 U19953 ( .A(n17645), .B(n16670), .ZN(n16661) );
  OAI22_X1 U19954 ( .A1(n16783), .A2(n17067), .B1(n16764), .B2(n16661), .ZN(
        n16662) );
  AOI211_X1 U19955 ( .C1(n16761), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16663), .B(n16662), .ZN(n16668) );
  NOR3_X1 U19956 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16789), .A3(n16664), .ZN(
        n16674) );
  NAND2_X1 U19957 ( .A1(n16770), .A2(n16664), .ZN(n16690) );
  NAND2_X1 U19958 ( .A1(n16792), .A2(n16690), .ZN(n16687) );
  OAI21_X1 U19959 ( .B1(n16674), .B2(n16687), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16667) );
  INV_X1 U19960 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18661) );
  NAND3_X1 U19961 ( .A1(n16770), .A2(n16665), .A3(n18661), .ZN(n16666) );
  NAND4_X1 U19962 ( .A1(n16668), .A2(n17988), .A3(n16667), .A4(n16666), .ZN(
        P3_U2661) );
  INV_X1 U19963 ( .A(n16687), .ZN(n16678) );
  OR2_X1 U19964 ( .A1(n16782), .A2(n16675), .ZN(n16685) );
  AOI21_X1 U19965 ( .B1(n17657), .B2(n16680), .A(n16669), .ZN(n17660) );
  AOI221_X1 U19966 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17660), .C1(
        n16680), .C2(n17660), .A(n16764), .ZN(n16671) );
  OAI22_X1 U19967 ( .A1(n16768), .A2(n16671), .B1(n17660), .B2(n16670), .ZN(
        n16672) );
  OAI211_X1 U19968 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n16685), .A(n17988), .B(
        n16672), .ZN(n16673) );
  AOI211_X1 U19969 ( .C1(n16761), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16674), .B(n16673), .ZN(n16677) );
  OAI221_X1 U19970 ( .B1(n16758), .B2(n16790), .C1(n16758), .C2(n16675), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n16676) );
  OAI211_X1 U19971 ( .C1(n16678), .C2(n18659), .A(n16677), .B(n16676), .ZN(
        P3_U2662) );
  INV_X1 U19972 ( .A(n16679), .ZN(n16691) );
  AOI22_X1 U19973 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16761), .B1(
        n16758), .B2(P3_EBX_REG_8__SCAN_IN), .ZN(n16689) );
  OAI21_X1 U19974 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16694), .A(
        n16680), .ZN(n17675) );
  INV_X1 U19975 ( .A(n17675), .ZN(n16683) );
  INV_X1 U19976 ( .A(n16682), .ZN(n16681) );
  OAI221_X1 U19977 ( .B1(n16683), .B2(n16682), .C1(n17675), .C2(n16681), .A(
        n18620), .ZN(n16684) );
  OAI221_X1 U19978 ( .B1(n16685), .B2(P3_EBX_REG_8__SCAN_IN), .C1(n16685), 
        .C2(n16702), .A(n16684), .ZN(n16686) );
  AOI211_X1 U19979 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n16687), .A(n9611), .B(
        n16686), .ZN(n16688) );
  OAI211_X1 U19980 ( .C1(n16691), .C2(n16690), .A(n16689), .B(n16688), .ZN(
        P3_U2663) );
  NOR2_X1 U19981 ( .A1(n16693), .A2(n16692), .ZN(n16713) );
  AOI21_X1 U19982 ( .B1(n17685), .B2(n16712), .A(n16694), .ZN(n17693) );
  XNOR2_X1 U19983 ( .A(n16713), .B(n17693), .ZN(n16695) );
  OAI21_X1 U19984 ( .B1(n16695), .B2(n16764), .A(n17988), .ZN(n16701) );
  NOR2_X1 U19985 ( .A1(n16789), .A2(n16696), .ZN(n16718) );
  INV_X1 U19986 ( .A(n16718), .ZN(n16741) );
  NOR2_X1 U19987 ( .A1(n16697), .A2(n16741), .ZN(n16699) );
  AOI21_X1 U19988 ( .B1(n16696), .B2(n16770), .A(n16776), .ZN(n16760) );
  INV_X1 U19989 ( .A(n16760), .ZN(n16720) );
  AOI21_X1 U19990 ( .B1(n16697), .B2(n16791), .A(n16720), .ZN(n16709) );
  INV_X1 U19991 ( .A(n16709), .ZN(n16698) );
  MUX2_X1 U19992 ( .A(n16699), .B(n16698), .S(P3_REIP_REG_7__SCAN_IN), .Z(
        n16700) );
  AOI211_X1 U19993 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16758), .A(n16701), .B(
        n16700), .ZN(n16705) );
  OAI211_X1 U19994 ( .C1(n16706), .C2(n16703), .A(n16790), .B(n16702), .ZN(
        n16704) );
  OAI211_X1 U19995 ( .C1(n16777), .C2(n17685), .A(n16705), .B(n16704), .ZN(
        P3_U2664) );
  AOI211_X1 U19996 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16727), .A(n16706), .B(
        n16782), .ZN(n16711) );
  INV_X1 U19997 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18651) );
  INV_X1 U19998 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18649) );
  NOR2_X1 U19999 ( .A1(n18651), .A2(n18649), .ZN(n16719) );
  AOI21_X1 U20000 ( .B1(n16719), .B2(n16718), .A(P3_REIP_REG_6__SCAN_IN), .ZN(
        n16708) );
  OAI22_X1 U20001 ( .A1(n16709), .A2(n16708), .B1(n16707), .B2(n16783), .ZN(
        n16710) );
  AOI211_X1 U20002 ( .C1(n16761), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16711), .B(n16710), .ZN(n16717) );
  OAI21_X1 U20003 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16722), .A(
        n16712), .ZN(n17705) );
  NAND3_X1 U20004 ( .A1(n18620), .A2(n16713), .A3(n17705), .ZN(n16716) );
  INV_X1 U20005 ( .A(n17705), .ZN(n16714) );
  OAI211_X1 U20006 ( .C1(n16722), .C2(n16768), .A(n16714), .B(n16785), .ZN(
        n16715) );
  NAND4_X1 U20007 ( .A1(n16717), .A2(n17988), .A3(n16716), .A4(n16715), .ZN(
        P3_U2665) );
  AOI21_X1 U20008 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16718), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n16725) );
  INV_X1 U20009 ( .A(n16719), .ZN(n16721) );
  AOI21_X1 U20010 ( .B1(n16721), .B2(n16791), .A(n16720), .ZN(n16724) );
  NAND3_X1 U20011 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17729), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16732) );
  AOI21_X1 U20012 ( .B1(n17720), .B2(n16732), .A(n16722), .ZN(n17722) );
  OAI21_X1 U20013 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16732), .A(
        n16749), .ZN(n16734) );
  XOR2_X1 U20014 ( .A(n17722), .B(n16734), .Z(n16723) );
  OAI22_X1 U20015 ( .A1(n16725), .A2(n16724), .B1(n16764), .B2(n16723), .ZN(
        n16726) );
  AOI211_X1 U20016 ( .C1(n16758), .C2(P3_EBX_REG_5__SCAN_IN), .A(n9611), .B(
        n16726), .ZN(n16730) );
  OAI211_X1 U20017 ( .C1(n16731), .C2(n16728), .A(n16790), .B(n16727), .ZN(
        n16729) );
  OAI211_X1 U20018 ( .C1(n16777), .C2(n17720), .A(n16730), .B(n16729), .ZN(
        P3_U2666) );
  INV_X1 U20019 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16746) );
  AOI211_X1 U20020 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16752), .A(n16731), .B(
        n16782), .ZN(n16743) );
  NAND2_X1 U20021 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17729), .ZN(
        n16747) );
  INV_X1 U20022 ( .A(n16747), .ZN(n16733) );
  OAI21_X1 U20023 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16733), .A(
        n16732), .ZN(n17731) );
  INV_X1 U20024 ( .A(n17731), .ZN(n16735) );
  OAI221_X1 U20025 ( .B1(n16735), .B2(n16734), .C1(n17731), .C2(n16749), .A(
        n17988), .ZN(n16739) );
  NOR2_X1 U20026 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16736), .ZN(
        n17727) );
  NAND2_X1 U20027 ( .A1(n16779), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16765) );
  INV_X1 U20028 ( .A(n16765), .ZN(n16738) );
  OAI221_X1 U20029 ( .B1(n16739), .B2(n17727), .C1(n16739), .C2(n16738), .A(
        n16737), .ZN(n16740) );
  OAI221_X1 U20030 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16741), .C1(n18649), 
        .C2(n16760), .A(n16740), .ZN(n16742) );
  AOI211_X1 U20031 ( .C1(n16761), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16743), .B(n16742), .ZN(n16745) );
  NOR2_X1 U20032 ( .A1(n18125), .A2(n18769), .ZN(n18784) );
  OAI21_X1 U20033 ( .B1(n9600), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n18784), .ZN(n16744) );
  OAI211_X1 U20034 ( .C1(n16746), .C2(n16783), .A(n16745), .B(n16744), .ZN(
        P3_U2667) );
  INV_X1 U20035 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18648) );
  NAND2_X1 U20036 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16769) );
  NOR3_X1 U20037 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n16789), .A3(n16769), .ZN(
        n16757) );
  INV_X1 U20038 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16755) );
  AOI21_X1 U20039 ( .B1(n18722), .B2(n18563), .A(n9600), .ZN(n18720) );
  INV_X1 U20040 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17756) );
  NOR2_X1 U20041 ( .A1(n17763), .A2(n17756), .ZN(n16748) );
  OAI21_X1 U20042 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16748), .A(
        n16747), .ZN(n17741) );
  OAI21_X1 U20043 ( .B1(n17756), .B2(n16765), .A(n16749), .ZN(n16763) );
  OAI21_X1 U20044 ( .B1(n17741), .B2(n16763), .A(n18620), .ZN(n16750) );
  AOI21_X1 U20045 ( .B1(n17741), .B2(n16763), .A(n16750), .ZN(n16751) );
  AOI21_X1 U20046 ( .B1(n18784), .B2(n18720), .A(n16751), .ZN(n16754) );
  OAI211_X1 U20047 ( .C1(n16762), .C2(n17132), .A(n16790), .B(n16752), .ZN(
        n16753) );
  OAI211_X1 U20048 ( .C1(n16777), .C2(n16755), .A(n16754), .B(n16753), .ZN(
        n16756) );
  AOI211_X1 U20049 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n16758), .A(n16757), .B(
        n16756), .ZN(n16759) );
  OAI21_X1 U20050 ( .B1(n18648), .B2(n16760), .A(n16759), .ZN(P3_U2668) );
  NAND2_X1 U20051 ( .A1(n18734), .A2(n18568), .ZN(n18561) );
  NAND2_X1 U20052 ( .A1(n18563), .A2(n18561), .ZN(n18580) );
  INV_X1 U20053 ( .A(n18580), .ZN(n18732) );
  AOI22_X1 U20054 ( .A1(n16776), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n18732), 
        .B2(n18784), .ZN(n16774) );
  AOI22_X1 U20055 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16761), .B1(
        n16758), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n16773) );
  OAI22_X1 U20056 ( .A1(n17763), .A2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n17756), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17749) );
  INV_X1 U20057 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n16795) );
  INV_X1 U20058 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17144) );
  NAND2_X1 U20059 ( .A1(n16795), .A2(n17144), .ZN(n16781) );
  AOI211_X1 U20060 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16781), .A(n16762), .B(
        n16782), .ZN(n16767) );
  AOI211_X1 U20061 ( .C1(n17749), .C2(n16765), .A(n16764), .B(n16763), .ZN(
        n16766) );
  AOI211_X1 U20062 ( .C1(n16768), .C2(n17749), .A(n16767), .B(n16766), .ZN(
        n16772) );
  OAI211_X1 U20063 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16770), .B(n16769), .ZN(n16771) );
  NAND4_X1 U20064 ( .A1(n16774), .A2(n16773), .A3(n16772), .A4(n16771), .ZN(
        P3_U2669) );
  NAND2_X1 U20065 ( .A1(n18568), .A2(n16775), .ZN(n18587) );
  INV_X1 U20066 ( .A(n18587), .ZN(n18737) );
  AOI22_X1 U20067 ( .A1(n16776), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18737), 
        .B2(n18784), .ZN(n16788) );
  OAI211_X1 U20068 ( .C1(n16779), .C2(n16778), .A(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B(n16777), .ZN(n16786) );
  NAND2_X1 U20069 ( .A1(n16781), .A2(n16780), .ZN(n17145) );
  OAI22_X1 U20070 ( .A1(n16783), .A2(n17144), .B1(n16782), .B2(n17145), .ZN(
        n16784) );
  AOI221_X1 U20071 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16786), .C1(
        n16785), .C2(n16786), .A(n16784), .ZN(n16787) );
  OAI211_X1 U20072 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n16789), .A(n16788), .B(
        n16787), .ZN(P3_U2670) );
  NOR2_X1 U20073 ( .A1(n16401), .A2(n16790), .ZN(n16796) );
  AOI22_X1 U20074 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16791), .B1(n18784), 
        .B2(n18749), .ZN(n16794) );
  NAND3_X1 U20075 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18729), .A3(
        n16792), .ZN(n16793) );
  OAI211_X1 U20076 ( .C1(n16796), .C2(n16795), .A(n16794), .B(n16793), .ZN(
        P3_U2671) );
  NAND2_X1 U20077 ( .A1(n16833), .A2(n16832), .ZN(n16797) );
  NOR3_X1 U20078 ( .A1(n16831), .A2(n16873), .A3(n16797), .ZN(n16825) );
  NAND2_X1 U20079 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16825), .ZN(n16824) );
  INV_X1 U20080 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16799) );
  INV_X1 U20081 ( .A(n16824), .ZN(n16798) );
  OAI33_X1 U20082 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18158), .A3(n16824), 
        .B1(n16799), .B2(n17147), .B3(n16798), .ZN(P3_U2672) );
  OAI22_X1 U20083 ( .A1(n16986), .A2(n16801), .B1(n12454), .B2(n16800), .ZN(
        n16811) );
  AOI22_X1 U20084 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16809) );
  AOI22_X1 U20085 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12442), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16808) );
  AOI22_X1 U20086 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16802) );
  OAI21_X1 U20087 ( .B1(n17077), .B2(n16985), .A(n16802), .ZN(n16806) );
  AOI22_X1 U20088 ( .A1(n17096), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16804) );
  AOI22_X1 U20089 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16972), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16803) );
  OAI211_X1 U20090 ( .C1(n17106), .C2(n16862), .A(n16804), .B(n16803), .ZN(
        n16805) );
  AOI211_X1 U20091 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n16806), .B(n16805), .ZN(n16807) );
  NAND3_X1 U20092 ( .A1(n16809), .A2(n16808), .A3(n16807), .ZN(n16810) );
  AOI211_X1 U20093 ( .C1(n16812), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n16811), .B(n16810), .ZN(n16829) );
  NOR2_X1 U20094 ( .A1(n16829), .A2(n16828), .ZN(n16827) );
  AOI22_X1 U20095 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17078), .B1(
        n17070), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16822) );
  AOI22_X1 U20096 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17115), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16821) );
  AOI22_X1 U20097 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n12486), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16820) );
  OAI22_X1 U20098 ( .A1(n16969), .A2(n17038), .B1(n16968), .B2(n17077), .ZN(
        n16818) );
  AOI22_X1 U20099 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17095), .ZN(n16816) );
  AOI22_X1 U20100 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n16972), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16815) );
  AOI22_X1 U20101 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12405), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17096), .ZN(n16814) );
  NAND2_X1 U20102 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n16813) );
  NAND4_X1 U20103 ( .A1(n16816), .A2(n16815), .A3(n16814), .A4(n16813), .ZN(
        n16817) );
  AOI211_X1 U20104 ( .C1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .C2(n16949), .A(
        n16818), .B(n16817), .ZN(n16819) );
  NAND4_X1 U20105 ( .A1(n16822), .A2(n16821), .A3(n16820), .A4(n16819), .ZN(
        n16823) );
  XNOR2_X1 U20106 ( .A(n16827), .B(n16823), .ZN(n17157) );
  OAI211_X1 U20107 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16825), .A(n16824), .B(
        n17139), .ZN(n16826) );
  OAI21_X1 U20108 ( .B1(n17157), .B2(n17139), .A(n16826), .ZN(P3_U2673) );
  AOI21_X1 U20109 ( .B1(n16829), .B2(n16828), .A(n16827), .ZN(n17161) );
  AOI22_X1 U20110 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16830), .B1(n17147), 
        .B2(n17161), .ZN(n16835) );
  NAND4_X1 U20111 ( .A1(n16885), .A2(n16833), .A3(n16832), .A4(n16831), .ZN(
        n16834) );
  NAND2_X1 U20112 ( .A1(n16835), .A2(n16834), .ZN(P3_U2674) );
  AOI21_X1 U20113 ( .B1(n16837), .B2(n17175), .A(n16836), .ZN(n17170) );
  AOI22_X1 U20114 ( .A1(n17170), .A2(n17147), .B1(n16838), .B2(n16840), .ZN(
        n16839) );
  OAI21_X1 U20115 ( .B1(n16840), .B2(n16843), .A(n16839), .ZN(P3_U2676) );
  NAND2_X1 U20116 ( .A1(n16885), .A2(n16841), .ZN(n16857) );
  OAI211_X1 U20117 ( .C1(n17177), .C2(n17176), .A(n17147), .B(n17175), .ZN(
        n16842) );
  XNOR2_X1 U20118 ( .A(n16845), .B(n16848), .ZN(n17186) );
  OAI211_X1 U20119 ( .C1(n16851), .C2(P3_EBX_REG_25__SCAN_IN), .A(n17139), .B(
        n9669), .ZN(n16846) );
  OAI21_X1 U20120 ( .B1(n17186), .B2(n17139), .A(n16846), .ZN(P3_U2678) );
  AOI21_X1 U20121 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17139), .A(n16847), .ZN(
        n16850) );
  OAI21_X1 U20122 ( .B1(n16852), .B2(n16849), .A(n16848), .ZN(n17192) );
  OAI22_X1 U20123 ( .A1(n16851), .A2(n16850), .B1(n17139), .B2(n17192), .ZN(
        P3_U2679) );
  AOI21_X1 U20124 ( .B1(n16854), .B2(n16853), .A(n16852), .ZN(n17193) );
  NAND3_X1 U20125 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n16885), .ZN(n16859) );
  OAI21_X1 U20126 ( .B1(n17147), .B2(n16855), .A(n16859), .ZN(n16856) );
  AOI22_X1 U20127 ( .A1(n17147), .A2(n17193), .B1(n16857), .B2(n16856), .ZN(
        n16858) );
  INV_X1 U20128 ( .A(n16858), .ZN(P3_U2680) );
  INV_X1 U20129 ( .A(n16859), .ZN(n16872) );
  AOI22_X1 U20130 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17139), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n16885), .ZN(n16871) );
  AOI22_X1 U20131 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16860) );
  OAI21_X1 U20132 ( .B1(n16986), .B2(n12420), .A(n16860), .ZN(n16870) );
  AOI22_X1 U20133 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17115), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16868) );
  AOI22_X1 U20134 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16861) );
  OAI21_X1 U20135 ( .B1(n17038), .B2(n16862), .A(n16861), .ZN(n16866) );
  AOI22_X1 U20136 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16864) );
  AOI22_X1 U20137 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16863) );
  OAI211_X1 U20138 ( .C1(n17106), .C2(n16985), .A(n16864), .B(n16863), .ZN(
        n16865) );
  AOI211_X1 U20139 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n16866), .B(n16865), .ZN(n16867) );
  OAI211_X1 U20140 ( .C1(n17077), .C2(n17124), .A(n16868), .B(n16867), .ZN(
        n16869) );
  AOI211_X1 U20141 ( .C1(n17102), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n16870), .B(n16869), .ZN(n17201) );
  OAI22_X1 U20142 ( .A1(n16872), .A2(n16871), .B1(n17201), .B2(n17139), .ZN(
        P3_U2681) );
  NAND2_X1 U20143 ( .A1(n17139), .A2(n16873), .ZN(n16899) );
  AOI22_X1 U20144 ( .A1(n16949), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16884) );
  INV_X1 U20145 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16876) );
  AOI22_X1 U20146 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16875) );
  AOI22_X1 U20147 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16874) );
  OAI211_X1 U20148 ( .C1(n17005), .C2(n16876), .A(n16875), .B(n16874), .ZN(
        n16882) );
  AOI22_X1 U20149 ( .A1(n17101), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16880) );
  AOI22_X1 U20150 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16906), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16879) );
  AOI22_X1 U20151 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17115), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16878) );
  NAND2_X1 U20152 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n16877) );
  NAND4_X1 U20153 ( .A1(n16880), .A2(n16879), .A3(n16878), .A4(n16877), .ZN(
        n16881) );
  AOI211_X1 U20154 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n16882), .B(n16881), .ZN(n16883) );
  OAI211_X1 U20155 ( .C1(n17077), .C2(n17128), .A(n16884), .B(n16883), .ZN(
        n17207) );
  AOI22_X1 U20156 ( .A1(n17147), .A2(n17207), .B1(n16885), .B2(n16887), .ZN(
        n16886) );
  OAI21_X1 U20157 ( .B1(n16887), .B2(n16899), .A(n16886), .ZN(P3_U2682) );
  NOR2_X1 U20158 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16917), .ZN(n16900) );
  AOI22_X1 U20159 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16888) );
  OAI21_X1 U20160 ( .B1(n10169), .B2(n17018), .A(n16888), .ZN(n16898) );
  AOI22_X1 U20161 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12486), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16896) );
  OAI22_X1 U20162 ( .A1(n17053), .A2(n16889), .B1(n12445), .B2(n17019), .ZN(
        n16894) );
  AOI22_X1 U20163 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16892) );
  AOI22_X1 U20164 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16906), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16891) );
  AOI22_X1 U20165 ( .A1(n16949), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16890) );
  NAND3_X1 U20166 ( .A1(n16892), .A2(n16891), .A3(n16890), .ZN(n16893) );
  AOI211_X1 U20167 ( .C1(n17074), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n16894), .B(n16893), .ZN(n16895) );
  OAI211_X1 U20168 ( .C1(n17077), .C2(n17131), .A(n16896), .B(n16895), .ZN(
        n16897) );
  AOI211_X1 U20169 ( .C1(n17101), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n16898), .B(n16897), .ZN(n17216) );
  OAI22_X1 U20170 ( .A1(n16900), .A2(n16899), .B1(n17216), .B2(n17139), .ZN(
        P3_U2683) );
  AOI21_X1 U20171 ( .B1(n16902), .B2(n16901), .A(n17147), .ZN(n16903) );
  INV_X1 U20172 ( .A(n16903), .ZN(n16916) );
  INV_X1 U20173 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16905) );
  AOI22_X1 U20174 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16904) );
  OAI21_X1 U20175 ( .B1(n17073), .B2(n16905), .A(n16904), .ZN(n16915) );
  AOI22_X1 U20176 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16906), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20177 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16907) );
  OAI21_X1 U20178 ( .B1(n17106), .B2(n17037), .A(n16907), .ZN(n16911) );
  AOI22_X1 U20179 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16909) );
  AOI22_X1 U20180 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16972), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16908) );
  OAI211_X1 U20181 ( .C1(n17038), .C2(n17035), .A(n16909), .B(n16908), .ZN(
        n16910) );
  AOI211_X1 U20182 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n16911), .B(n16910), .ZN(n16912) );
  OAI211_X1 U20183 ( .C1(n17077), .C2(n17134), .A(n16913), .B(n16912), .ZN(
        n16914) );
  AOI211_X1 U20184 ( .C1(n17070), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n16915), .B(n16914), .ZN(n17221) );
  OAI22_X1 U20185 ( .A1(n16917), .A2(n16916), .B1(n17221), .B2(n17139), .ZN(
        P3_U2684) );
  INV_X1 U20186 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17141) );
  OAI22_X1 U20187 ( .A1(n16918), .A2(n17087), .B1(n17077), .B2(n17141), .ZN(
        n16929) );
  AOI22_X1 U20188 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16927) );
  AOI22_X1 U20189 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16926) );
  OAI22_X1 U20190 ( .A1(n17100), .A2(n17052), .B1(n12454), .B2(n16919), .ZN(
        n16924) );
  AOI22_X1 U20191 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n17095), .B1(
        n17101), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16922) );
  AOI22_X1 U20192 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16921) );
  AOI22_X1 U20193 ( .A1(n16949), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16920) );
  NAND3_X1 U20194 ( .A1(n16922), .A2(n16921), .A3(n16920), .ZN(n16923) );
  AOI211_X1 U20195 ( .C1(n12486), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n16924), .B(n16923), .ZN(n16925) );
  NAND3_X1 U20196 ( .A1(n16927), .A2(n16926), .A3(n16925), .ZN(n16928) );
  AOI211_X1 U20197 ( .C1(n17096), .C2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n16929), .B(n16928), .ZN(n17225) );
  NOR2_X1 U20198 ( .A1(n17147), .A2(n9701), .ZN(n16945) );
  NOR4_X1 U20199 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18158), .A3(n16930), .A4(
        n16944), .ZN(n16931) );
  AOI21_X1 U20200 ( .B1(n16945), .B2(P3_EBX_REG_18__SCAN_IN), .A(n16931), .ZN(
        n16932) );
  OAI21_X1 U20201 ( .B1(n17225), .B2(n17139), .A(n16932), .ZN(P3_U2685) );
  AOI22_X1 U20202 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16933) );
  OAI21_X1 U20203 ( .B1(n10165), .B2(n17072), .A(n16933), .ZN(n16943) );
  AOI22_X1 U20204 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16941) );
  AOI22_X1 U20205 ( .A1(n17074), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16949), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16934) );
  OAI21_X1 U20206 ( .B1(n17005), .B2(n16935), .A(n16934), .ZN(n16939) );
  INV_X1 U20207 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20208 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17096), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16937) );
  AOI22_X1 U20209 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16936) );
  OAI211_X1 U20210 ( .C1(n17038), .C2(n17086), .A(n16937), .B(n16936), .ZN(
        n16938) );
  AOI211_X1 U20211 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n16939), .B(n16938), .ZN(n16940) );
  OAI211_X1 U20212 ( .C1(n17077), .C2(n17142), .A(n16941), .B(n16940), .ZN(
        n16942) );
  AOI211_X1 U20213 ( .C1(n17102), .C2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n16943), .B(n16942), .ZN(n17232) );
  INV_X1 U20214 ( .A(n16944), .ZN(n16946) );
  OAI21_X1 U20215 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16946), .A(n16945), .ZN(
        n16947) );
  OAI21_X1 U20216 ( .B1(n17232), .B2(n17139), .A(n16947), .ZN(P3_U2686) );
  AOI22_X1 U20217 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16972), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16948) );
  OAI21_X1 U20218 ( .B1(n12430), .B2(n17094), .A(n16948), .ZN(n16959) );
  INV_X1 U20219 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20220 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16956) );
  OAI22_X1 U20221 ( .A1(n17077), .A2(n17105), .B1(n12420), .B2(n17112), .ZN(
        n16954) );
  AOI22_X1 U20222 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16952) );
  AOI22_X1 U20223 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n17075), .B1(
        n12405), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16951) );
  AOI22_X1 U20224 ( .A1(n16949), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16950) );
  NAND3_X1 U20225 ( .A1(n16952), .A2(n16951), .A3(n16950), .ZN(n16953) );
  AOI211_X1 U20226 ( .C1(n17070), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n16954), .B(n16953), .ZN(n16955) );
  OAI211_X1 U20227 ( .C1(n17100), .C2(n16957), .A(n16956), .B(n16955), .ZN(
        n16958) );
  AOI211_X1 U20228 ( .C1(n17102), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n16959), .B(n16958), .ZN(n17239) );
  NOR2_X1 U20229 ( .A1(n17147), .A2(n16960), .ZN(n16982) );
  NOR2_X1 U20230 ( .A1(n18158), .A2(n17129), .ZN(n17122) );
  NAND2_X1 U20231 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n16965) );
  NAND2_X1 U20232 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .ZN(n16964) );
  NAND4_X1 U20233 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(P3_EBX_REG_7__SCAN_IN), .ZN(n16963) );
  OR4_X1 U20234 ( .A1(n16999), .A2(n16961), .A3(n17067), .A4(
        P3_EBX_REG_16__SCAN_IN), .ZN(n16962) );
  NOR4_X1 U20235 ( .A1(n16965), .A2(n16964), .A3(n16963), .A4(n16962), .ZN(
        n16966) );
  AOI22_X1 U20236 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16982), .B1(n17122), 
        .B2(n16966), .ZN(n16967) );
  OAI21_X1 U20237 ( .B1(n17239), .B2(n17139), .A(n16967), .ZN(P3_U2687) );
  OAI22_X1 U20238 ( .A1(n16969), .A2(n17100), .B1(n16968), .B2(n17038), .ZN(
        n16981) );
  AOI22_X1 U20239 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17078), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17096), .ZN(n16979) );
  AOI22_X1 U20240 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17075), .ZN(n16978) );
  AOI22_X1 U20241 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17074), .ZN(n16970) );
  OAI21_X1 U20242 ( .B1(n17087), .B2(n16971), .A(n16970), .ZN(n16976) );
  AOI22_X1 U20243 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n16972), .B1(
        n17102), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20244 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n16812), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17095), .ZN(n16973) );
  OAI211_X1 U20245 ( .C1(n17119), .C2(n17106), .A(n16974), .B(n16973), .ZN(
        n16975) );
  AOI211_X1 U20246 ( .C1(n12486), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n16976), .B(n16975), .ZN(n16977) );
  NAND3_X1 U20247 ( .A1(n16979), .A2(n16978), .A3(n16977), .ZN(n16980) );
  AOI211_X1 U20248 ( .C1(n17097), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n16981), .B(n16980), .ZN(n17243) );
  OAI21_X1 U20249 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n16983), .A(n16982), .ZN(
        n16984) );
  OAI21_X1 U20250 ( .B1(n17243), .B2(n17139), .A(n16984), .ZN(P3_U2688) );
  AOI22_X1 U20251 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16997) );
  AOI22_X1 U20252 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17096), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16996) );
  OAI22_X1 U20253 ( .A1(n16986), .A2(n12454), .B1(n17038), .B2(n16985), .ZN(
        n16994) );
  AOI22_X1 U20254 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16991) );
  AOI22_X1 U20255 ( .A1(n17115), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16972), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20256 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16987) );
  OAI211_X1 U20257 ( .C1(n17106), .C2(n17124), .A(n16988), .B(n16987), .ZN(
        n16989) );
  AOI21_X1 U20258 ( .B1(n12486), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n16989), .ZN(n16990) );
  OAI211_X1 U20259 ( .C1(n17077), .C2(n16992), .A(n16991), .B(n16990), .ZN(
        n16993) );
  AOI211_X1 U20260 ( .C1(n17060), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n16994), .B(n16993), .ZN(n16995) );
  NAND3_X1 U20261 ( .A1(n16997), .A2(n16996), .A3(n16995), .ZN(n17244) );
  INV_X1 U20262 ( .A(n17016), .ZN(n16998) );
  OAI33_X1 U20263 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17016), .A3(n18158), 
        .B1(n16999), .B2(n17147), .B3(n16998), .ZN(n17000) );
  AOI21_X1 U20264 ( .B1(n17147), .B2(n17244), .A(n17000), .ZN(n17001) );
  INV_X1 U20265 ( .A(n17001), .ZN(P3_U2689) );
  AOI22_X1 U20266 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17096), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17002) );
  OAI21_X1 U20267 ( .B1(n17073), .B2(n17003), .A(n17002), .ZN(n17015) );
  AOI22_X1 U20268 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17115), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17012) );
  OAI22_X1 U20269 ( .A1(n17005), .A2(n17004), .B1(n17106), .B2(n17128), .ZN(
        n17010) );
  AOI22_X1 U20270 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20271 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17007) );
  AOI22_X1 U20272 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17006) );
  NAND3_X1 U20273 ( .A1(n17008), .A2(n17007), .A3(n17006), .ZN(n17009) );
  AOI211_X1 U20274 ( .C1(n17074), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n17010), .B(n17009), .ZN(n17011) );
  OAI211_X1 U20275 ( .C1(n17077), .C2(n17013), .A(n17012), .B(n17011), .ZN(
        n17014) );
  AOI211_X1 U20276 ( .C1(n17070), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n17015), .B(n17014), .ZN(n17249) );
  AND2_X1 U20277 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17031), .ZN(n17033) );
  OAI211_X1 U20278 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n17033), .A(n17016), .B(
        n17139), .ZN(n17017) );
  OAI21_X1 U20279 ( .B1(n17249), .B2(n17139), .A(n17017), .ZN(P3_U2690) );
  OAI22_X1 U20280 ( .A1(n17077), .A2(n17019), .B1(n12445), .B2(n17018), .ZN(
        n17030) );
  AOI22_X1 U20281 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20282 ( .A1(n17096), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17027) );
  INV_X1 U20283 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17021) );
  AOI22_X1 U20284 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17020) );
  OAI21_X1 U20285 ( .B1(n17100), .B2(n17021), .A(n17020), .ZN(n17025) );
  AOI22_X1 U20286 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20287 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17022) );
  OAI211_X1 U20288 ( .C1(n17106), .C2(n17131), .A(n17023), .B(n17022), .ZN(
        n17024) );
  NAND3_X1 U20289 ( .A1(n17028), .A2(n17027), .A3(n17026), .ZN(n17029) );
  AOI211_X1 U20290 ( .C1(n12442), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n17030), .B(n17029), .ZN(n17254) );
  OAI21_X1 U20291 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17031), .A(n17139), .ZN(
        n17032) );
  OAI22_X1 U20292 ( .A1(n17254), .A2(n17139), .B1(n17033), .B2(n17032), .ZN(
        P3_U2691) );
  AOI22_X1 U20293 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17034) );
  OAI21_X1 U20294 ( .B1(n17087), .B2(n17035), .A(n17034), .ZN(n17048) );
  AOI22_X1 U20295 ( .A1(n17096), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20296 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17036) );
  OAI21_X1 U20297 ( .B1(n17038), .B2(n17037), .A(n17036), .ZN(n17043) );
  AOI22_X1 U20298 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20299 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12405), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17040) );
  OAI211_X1 U20300 ( .C1(n17106), .C2(n17134), .A(n17041), .B(n17040), .ZN(
        n17042) );
  AOI211_X1 U20301 ( .C1(n12486), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n17043), .B(n17042), .ZN(n17044) );
  OAI211_X1 U20302 ( .C1(n17077), .C2(n17046), .A(n17045), .B(n17044), .ZN(
        n17047) );
  AOI211_X1 U20303 ( .C1(n17102), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n17048), .B(n17047), .ZN(n17257) );
  OAI21_X1 U20304 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n9728), .A(n17049), .ZN(
        n17050) );
  AOI22_X1 U20305 ( .A1(n17147), .A2(n17257), .B1(n17050), .B2(n17139), .ZN(
        P3_U2692) );
  AOI22_X1 U20306 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17051) );
  OAI21_X1 U20307 ( .B1(n17053), .B2(n17052), .A(n17051), .ZN(n17065) );
  AOI22_X1 U20308 ( .A1(n12442), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17062) );
  OAI22_X1 U20309 ( .A1(n17077), .A2(n17054), .B1(n17106), .B2(n17141), .ZN(
        n17059) );
  AOI22_X1 U20310 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20311 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20312 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17055) );
  NAND3_X1 U20313 ( .A1(n17057), .A2(n17056), .A3(n17055), .ZN(n17058) );
  AOI211_X1 U20314 ( .C1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .C2(n17060), .A(
        n17059), .B(n17058), .ZN(n17061) );
  OAI211_X1 U20315 ( .C1(n10165), .C2(n17063), .A(n17062), .B(n17061), .ZN(
        n17064) );
  AOI211_X1 U20316 ( .C1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .C2(n17096), .A(
        n17065), .B(n17064), .ZN(n17264) );
  INV_X1 U20317 ( .A(n17090), .ZN(n17066) );
  OAI33_X1 U20318 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18158), .A3(n17090), 
        .B1(n17067), .B2(n17147), .B3(n17066), .ZN(n17068) );
  INV_X1 U20319 ( .A(n17068), .ZN(n17069) );
  OAI21_X1 U20320 ( .B1(n17264), .B2(n17139), .A(n17069), .ZN(P3_U2693) );
  AOI22_X1 U20321 ( .A1(n17070), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17071) );
  OAI21_X1 U20322 ( .B1(n17073), .B2(n17072), .A(n17071), .ZN(n17089) );
  AOI22_X1 U20323 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17074), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17085) );
  OAI22_X1 U20324 ( .A1(n17077), .A2(n17076), .B1(n17106), .B2(n17142), .ZN(
        n17083) );
  AOI22_X1 U20325 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17096), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17081) );
  AOI22_X1 U20326 ( .A1(n17078), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17080) );
  AOI22_X1 U20327 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17079) );
  NAND3_X1 U20328 ( .A1(n17081), .A2(n17080), .A3(n17079), .ZN(n17082) );
  AOI211_X1 U20329 ( .C1(n12486), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n17083), .B(n17082), .ZN(n17084) );
  OAI211_X1 U20330 ( .C1(n17087), .C2(n17086), .A(n17085), .B(n17084), .ZN(
        n17088) );
  AOI211_X1 U20331 ( .C1(n17102), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n17089), .B(n17088), .ZN(n17266) );
  OAI211_X1 U20332 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n17117), .A(n17090), .B(
        n17139), .ZN(n17091) );
  OAI21_X1 U20333 ( .B1(n17266), .B2(n17139), .A(n17091), .ZN(P3_U2694) );
  OAI21_X1 U20334 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17121), .A(n17139), .ZN(
        n17116) );
  AOI22_X1 U20335 ( .A1(n16972), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17092), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17093) );
  OAI21_X1 U20336 ( .B1(n10169), .B2(n17094), .A(n17093), .ZN(n17114) );
  AOI22_X1 U20337 ( .A1(n17096), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17095), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20338 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12486), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17098) );
  OAI21_X1 U20339 ( .B1(n17100), .B2(n17099), .A(n17098), .ZN(n17108) );
  AOI22_X1 U20340 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n17101), .B1(
        n16812), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U20341 ( .A1(n17102), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17078), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17103) );
  OAI211_X1 U20342 ( .C1(n17106), .C2(n17105), .A(n17104), .B(n17103), .ZN(
        n17107) );
  OAI211_X1 U20343 ( .C1(n12454), .C2(n17112), .A(n17111), .B(n17110), .ZN(
        n17113) );
  AOI211_X1 U20344 ( .C1(n17115), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17114), .B(n17113), .ZN(n17273) );
  OAI22_X1 U20345 ( .A1(n17117), .A2(n17116), .B1(n17273), .B2(n17139), .ZN(
        P3_U2695) );
  AOI22_X1 U20346 ( .A1(n17199), .A2(n17118), .B1(P3_EBX_REG_7__SCAN_IN), .B2(
        n17139), .ZN(n17120) );
  OAI22_X1 U20347 ( .A1(n17121), .A2(n17120), .B1(n17119), .B2(n17139), .ZN(
        P3_U2696) );
  NAND2_X1 U20348 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17122), .ZN(n17125) );
  NAND3_X1 U20349 ( .A1(n17125), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17139), .ZN(
        n17123) );
  OAI221_X1 U20350 ( .B1(n17125), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17139), 
        .C2(n17124), .A(n17123), .ZN(P3_U2697) );
  INV_X1 U20351 ( .A(n17129), .ZN(n17126) );
  OAI211_X1 U20352 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17126), .A(n17125), .B(
        n17139), .ZN(n17127) );
  OAI21_X1 U20353 ( .B1(n17139), .B2(n17128), .A(n17127), .ZN(P3_U2698) );
  OAI21_X1 U20354 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17136), .A(n17129), .ZN(
        n17130) );
  AOI22_X1 U20355 ( .A1(n17147), .A2(n17131), .B1(n17130), .B2(n17139), .ZN(
        P3_U2699) );
  AOI21_X1 U20356 ( .B1(n17132), .B2(n17137), .A(n17147), .ZN(n17133) );
  INV_X1 U20357 ( .A(n17133), .ZN(n17135) );
  OAI22_X1 U20358 ( .A1(n17136), .A2(n17135), .B1(n17134), .B2(n17139), .ZN(
        P3_U2700) );
  OAI21_X1 U20359 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n17138), .A(n17137), .ZN(
        n17140) );
  AOI22_X1 U20360 ( .A1(n17147), .A2(n17141), .B1(n17140), .B2(n17139), .ZN(
        P3_U2701) );
  OAI222_X1 U20361 ( .A1(n17145), .A2(n17149), .B1(n17144), .B2(n17143), .C1(
        n17142), .C2(n17139), .ZN(P3_U2702) );
  AOI22_X1 U20362 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17147), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17146), .ZN(n17148) );
  OAI21_X1 U20363 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17149), .A(n17148), .ZN(
        P3_U2703) );
  NAND2_X1 U20364 ( .A1(n18158), .A2(n17150), .ZN(n17296) );
  INV_X1 U20365 ( .A(n17234), .ZN(n17200) );
  INV_X1 U20366 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17372) );
  INV_X1 U20367 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17368) );
  INV_X1 U20368 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17366) );
  INV_X1 U20369 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17364) );
  INV_X1 U20370 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17350) );
  INV_X1 U20371 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17383) );
  INV_X1 U20372 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17395) );
  NAND2_X1 U20373 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n17275) );
  NOR4_X1 U20374 ( .A1(n17385), .A2(n17395), .A3(n17381), .A4(n17275), .ZN(
        n17153) );
  INV_X1 U20375 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17403) );
  NAND2_X1 U20376 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n17245), .ZN(n17240) );
  NOR2_X2 U20377 ( .A1(n17350), .A2(n17240), .ZN(n17235) );
  INV_X1 U20378 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17356) );
  INV_X1 U20379 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17360) );
  INV_X1 U20380 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17358) );
  INV_X1 U20381 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17354) );
  NOR4_X1 U20382 ( .A1(n17356), .A2(n17360), .A3(n17358), .A4(n17354), .ZN(
        n17204) );
  NAND4_X1 U20383 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(n17235), .A4(n17204), .ZN(n17195) );
  NAND2_X1 U20384 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17171), .ZN(n17166) );
  NAND2_X1 U20385 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17163), .ZN(n17162) );
  NOR2_X1 U20386 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17162), .ZN(n17155) );
  INV_X1 U20387 ( .A(n17301), .ZN(n17274) );
  NAND2_X1 U20388 ( .A1(n17296), .A2(n17162), .ZN(n17160) );
  OAI21_X1 U20389 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17274), .A(n17160), .ZN(
        n17154) );
  AOI22_X1 U20390 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17155), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17154), .ZN(n17156) );
  OAI21_X1 U20391 ( .B1(n18162), .B2(n17200), .A(n17156), .ZN(P3_U2704) );
  INV_X1 U20392 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17378) );
  NOR2_X2 U20393 ( .A1(n18148), .A2(n17296), .ZN(n17233) );
  OAI22_X1 U20394 ( .A1(n17157), .A2(n17308), .B1(n19185), .B2(n17200), .ZN(
        n17158) );
  AOI21_X1 U20395 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17233), .A(n17158), .ZN(
        n17159) );
  OAI221_X1 U20396 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17162), .C1(n17378), 
        .C2(n17160), .A(n17159), .ZN(P3_U2705) );
  INV_X1 U20397 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18150) );
  AOI22_X1 U20398 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17233), .B1(n17283), .B2(
        n17161), .ZN(n17165) );
  OAI211_X1 U20399 ( .C1(n17163), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17296), .B(
        n17162), .ZN(n17164) );
  OAI211_X1 U20400 ( .C1(n17200), .C2(n18150), .A(n17165), .B(n17164), .ZN(
        P3_U2706) );
  AOI22_X1 U20401 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17234), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n17233), .ZN(n17168) );
  OAI211_X1 U20402 ( .C1(n17171), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17296), .B(
        n17166), .ZN(n17167) );
  OAI211_X1 U20403 ( .C1(n17169), .C2(n17308), .A(n17168), .B(n17167), .ZN(
        P3_U2707) );
  INV_X1 U20404 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18138) );
  AOI22_X1 U20405 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17233), .B1(n17283), .B2(
        n17170), .ZN(n17174) );
  AOI211_X1 U20406 ( .C1(n17372), .C2(n17178), .A(n17171), .B(n17285), .ZN(
        n17172) );
  INV_X1 U20407 ( .A(n17172), .ZN(n17173) );
  OAI211_X1 U20408 ( .C1(n17200), .C2(n18138), .A(n17174), .B(n17173), .ZN(
        P3_U2708) );
  OAI21_X1 U20409 ( .B1(n17177), .B2(n17176), .A(n17175), .ZN(n17181) );
  AOI22_X1 U20410 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n17234), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n17233), .ZN(n17180) );
  OAI211_X1 U20411 ( .C1(n17182), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17296), .B(
        n17178), .ZN(n17179) );
  OAI211_X1 U20412 ( .C1(n17181), .C2(n17308), .A(n17180), .B(n17179), .ZN(
        P3_U2709) );
  AOI22_X1 U20413 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n17234), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n17233), .ZN(n17185) );
  AOI211_X1 U20414 ( .C1(n17368), .C2(n17188), .A(n17182), .B(n17285), .ZN(
        n17183) );
  INV_X1 U20415 ( .A(n17183), .ZN(n17184) );
  OAI211_X1 U20416 ( .C1(n17186), .C2(n17308), .A(n17185), .B(n17184), .ZN(
        P3_U2710) );
  AOI22_X1 U20417 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17234), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17233), .ZN(n17191) );
  OAI21_X1 U20418 ( .B1(n17366), .B2(n17285), .A(n17187), .ZN(n17189) );
  NAND2_X1 U20419 ( .A1(n17189), .A2(n17188), .ZN(n17190) );
  OAI211_X1 U20420 ( .C1(n17192), .C2(n17308), .A(n17191), .B(n17190), .ZN(
        P3_U2711) );
  AOI22_X1 U20421 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n17234), .B1(n17283), .B2(
        n17193), .ZN(n17198) );
  AOI211_X1 U20422 ( .C1(n17364), .C2(n17195), .A(n17285), .B(n17194), .ZN(
        n17196) );
  AOI21_X1 U20423 ( .B1(n17233), .B2(BUF2_REG_7__SCAN_IN), .A(n17196), .ZN(
        n17197) );
  NAND2_X1 U20424 ( .A1(n17198), .A2(n17197), .ZN(P3_U2712) );
  INV_X1 U20425 ( .A(n17233), .ZN(n17209) );
  INV_X1 U20426 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18154) );
  INV_X1 U20427 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17352) );
  NAND2_X1 U20428 ( .A1(n17199), .A2(n17235), .ZN(n17226) );
  NAND2_X1 U20429 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17227), .ZN(n17222) );
  NAND2_X1 U20430 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17217), .ZN(n17213) );
  NAND2_X1 U20431 ( .A1(n17296), .A2(n17213), .ZN(n17208) );
  OAI21_X1 U20432 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17274), .A(n17208), .ZN(
        n17203) );
  INV_X1 U20433 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18155) );
  OAI22_X1 U20434 ( .A1(n17201), .A2(n17308), .B1(n18155), .B2(n17200), .ZN(
        n17202) );
  AOI21_X1 U20435 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(n17203), .A(n17202), .ZN(
        n17206) );
  INV_X1 U20436 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17362) );
  NAND3_X1 U20437 ( .A1(n17204), .A2(n17227), .A3(n17362), .ZN(n17205) );
  OAI211_X1 U20438 ( .C1(n17209), .C2(n18154), .A(n17206), .B(n17205), .ZN(
        P3_U2713) );
  AOI22_X1 U20439 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17234), .B1(n17283), .B2(
        n17207), .ZN(n17212) );
  INV_X1 U20440 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18149) );
  OAI22_X1 U20441 ( .A1(n18149), .A2(n17209), .B1(n17360), .B2(n17208), .ZN(
        n17210) );
  INV_X1 U20442 ( .A(n17210), .ZN(n17211) );
  OAI211_X1 U20443 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n17213), .A(n17212), .B(
        n17211), .ZN(P3_U2714) );
  AOI22_X1 U20444 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17234), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n17233), .ZN(n17215) );
  OAI211_X1 U20445 ( .C1(n17217), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17296), .B(
        n17213), .ZN(n17214) );
  OAI211_X1 U20446 ( .C1(n17216), .C2(n17308), .A(n17215), .B(n17214), .ZN(
        P3_U2715) );
  AOI22_X1 U20447 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n17234), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n17233), .ZN(n17220) );
  AOI211_X1 U20448 ( .C1(n17356), .C2(n17222), .A(n17217), .B(n17285), .ZN(
        n17218) );
  INV_X1 U20449 ( .A(n17218), .ZN(n17219) );
  OAI211_X1 U20450 ( .C1(n17221), .C2(n17308), .A(n17220), .B(n17219), .ZN(
        P3_U2716) );
  AOI22_X1 U20451 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17234), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n17233), .ZN(n17224) );
  OAI211_X1 U20452 ( .C1(n17227), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17296), .B(
        n17222), .ZN(n17223) );
  OAI211_X1 U20453 ( .C1(n17225), .C2(n17308), .A(n17224), .B(n17223), .ZN(
        P3_U2717) );
  AOI22_X1 U20454 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n17234), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17233), .ZN(n17231) );
  OAI21_X1 U20455 ( .B1(n17352), .B2(n17285), .A(n17226), .ZN(n17229) );
  INV_X1 U20456 ( .A(n17227), .ZN(n17228) );
  NAND2_X1 U20457 ( .A1(n17229), .A2(n17228), .ZN(n17230) );
  OAI211_X1 U20458 ( .C1(n17232), .C2(n17308), .A(n17231), .B(n17230), .ZN(
        P3_U2718) );
  AOI22_X1 U20459 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n17234), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n17233), .ZN(n17238) );
  AOI211_X1 U20460 ( .C1(n17350), .C2(n17240), .A(n17285), .B(n17235), .ZN(
        n17236) );
  INV_X1 U20461 ( .A(n17236), .ZN(n17237) );
  OAI211_X1 U20462 ( .C1(n17239), .C2(n17308), .A(n17238), .B(n17237), .ZN(
        P3_U2719) );
  OAI211_X1 U20463 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17245), .A(n17296), .B(
        n17240), .ZN(n17242) );
  NAND2_X1 U20464 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17306), .ZN(n17241) );
  OAI211_X1 U20465 ( .C1(n17243), .C2(n17308), .A(n17242), .B(n17241), .ZN(
        P3_U2720) );
  INV_X1 U20466 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17406) );
  NOR2_X1 U20467 ( .A1(n18158), .A2(n17270), .ZN(n17278) );
  NAND2_X1 U20468 ( .A1(n9739), .A2(n17278), .ZN(n17265) );
  NAND2_X1 U20469 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17261), .ZN(n17253) );
  NOR2_X1 U20470 ( .A1(n17406), .A2(n17253), .ZN(n17256) );
  NAND2_X1 U20471 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17256), .ZN(n17248) );
  AOI22_X1 U20472 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17306), .B1(n17283), .B2(
        n17244), .ZN(n17247) );
  INV_X1 U20473 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17410) );
  OR3_X1 U20474 ( .A1(n17410), .A2(n17285), .A3(n17245), .ZN(n17246) );
  OAI211_X1 U20475 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17248), .A(n17247), .B(
        n17246), .ZN(P3_U2721) );
  INV_X1 U20476 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17252) );
  INV_X1 U20477 ( .A(n17248), .ZN(n17251) );
  AOI21_X1 U20478 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17296), .A(n17256), .ZN(
        n17250) );
  OAI222_X1 U20479 ( .A1(n17300), .A2(n17252), .B1(n17251), .B2(n17250), .C1(
        n17308), .C2(n17249), .ZN(P3_U2722) );
  INV_X1 U20480 ( .A(n17253), .ZN(n17259) );
  AOI21_X1 U20481 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17296), .A(n17259), .ZN(
        n17255) );
  OAI222_X1 U20482 ( .A1(n17300), .A2(n12737), .B1(n17256), .B2(n17255), .C1(
        n17308), .C2(n17254), .ZN(P3_U2723) );
  INV_X1 U20483 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17260) );
  AOI21_X1 U20484 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17296), .A(n17261), .ZN(
        n17258) );
  OAI222_X1 U20485 ( .A1(n17300), .A2(n17260), .B1(n17259), .B2(n17258), .C1(
        n17308), .C2(n17257), .ZN(P3_U2724) );
  AOI211_X1 U20486 ( .C1(n17401), .C2(n17265), .A(n17261), .B(n17285), .ZN(
        n17262) );
  AOI21_X1 U20487 ( .B1(n17306), .B2(BUF2_REG_10__SCAN_IN), .A(n17262), .ZN(
        n17263) );
  OAI21_X1 U20488 ( .B1(n17264), .B2(n17308), .A(n17263), .ZN(P3_U2725) );
  INV_X1 U20489 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17269) );
  INV_X1 U20490 ( .A(n17265), .ZN(n17268) );
  AOI22_X1 U20491 ( .A1(n17278), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17296), .ZN(n17267) );
  OAI222_X1 U20492 ( .A1(n17300), .A2(n17269), .B1(n17268), .B2(n17267), .C1(
        n17308), .C2(n17266), .ZN(P3_U2726) );
  INV_X1 U20493 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U20494 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17306), .B1(n17278), .B2(
        n17397), .ZN(n17272) );
  NAND3_X1 U20495 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17296), .A3(n17270), .ZN(
        n17271) );
  OAI211_X1 U20496 ( .C1(n17273), .C2(n17308), .A(n17272), .B(n17271), .ZN(
        P3_U2727) );
  INV_X1 U20497 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18160) );
  INV_X1 U20498 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17387) );
  NOR3_X1 U20499 ( .A1(n17383), .A2(n17381), .A3(n17274), .ZN(n17295) );
  NAND2_X1 U20500 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17295), .ZN(n17291) );
  NOR2_X1 U20501 ( .A1(n17387), .A2(n17291), .ZN(n17294) );
  NAND2_X1 U20502 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17294), .ZN(n17287) );
  NOR2_X1 U20503 ( .A1(n17275), .A2(n17287), .ZN(n17281) );
  AOI21_X1 U20504 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17296), .A(n17281), .ZN(
        n17277) );
  OAI222_X1 U20505 ( .A1(n17300), .A2(n18160), .B1(n17278), .B2(n17277), .C1(
        n17308), .C2(n17276), .ZN(P3_U2728) );
  INV_X1 U20506 ( .A(n17287), .ZN(n17290) );
  AOI22_X1 U20507 ( .A1(n17290), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n17296), .ZN(n17280) );
  OAI222_X1 U20508 ( .A1(n18154), .A2(n17300), .B1(n17281), .B2(n17280), .C1(
        n17308), .C2(n17279), .ZN(P3_U2729) );
  NAND2_X1 U20509 ( .A1(n17287), .A2(P3_EAX_REG_5__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20510 ( .A1(n17306), .A2(BUF2_REG_5__SCAN_IN), .B1(n17283), .B2(
        n17282), .ZN(n17284) );
  OAI221_X1 U20511 ( .B1(n17287), .B2(P3_EAX_REG_5__SCAN_IN), .C1(n17286), 
        .C2(n17285), .A(n17284), .ZN(P3_U2730) );
  INV_X1 U20512 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18144) );
  AOI21_X1 U20513 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17296), .A(n17294), .ZN(
        n17289) );
  OAI222_X1 U20514 ( .A1(n18144), .A2(n17300), .B1(n17290), .B2(n17289), .C1(
        n17308), .C2(n17288), .ZN(P3_U2731) );
  INV_X1 U20515 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18139) );
  INV_X1 U20516 ( .A(n17291), .ZN(n17299) );
  AOI21_X1 U20517 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17296), .A(n17299), .ZN(
        n17293) );
  OAI222_X1 U20518 ( .A1(n18139), .A2(n17300), .B1(n17294), .B2(n17293), .C1(
        n17308), .C2(n17292), .ZN(P3_U2732) );
  INV_X1 U20519 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18134) );
  AOI21_X1 U20520 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17296), .A(n17295), .ZN(
        n17298) );
  OAI222_X1 U20521 ( .A1(n18134), .A2(n17300), .B1(n17299), .B2(n17298), .C1(
        n17308), .C2(n17297), .ZN(P3_U2733) );
  NAND2_X1 U20522 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17301), .ZN(n17302) );
  AOI22_X1 U20523 ( .A1(n17304), .A2(n17303), .B1(n17383), .B2(n17302), .ZN(
        n17305) );
  AOI21_X1 U20524 ( .B1(n17306), .B2(BUF2_REG_1__SCAN_IN), .A(n17305), .ZN(
        n17307) );
  OAI21_X1 U20525 ( .B1(n12501), .B2(n17308), .A(n17307), .ZN(P3_U2734) );
  NOR2_X2 U20526 ( .A1(n18726), .A2(n17771), .ZN(n18774) );
  NOR2_X4 U20527 ( .A1(n18774), .A2(n17326), .ZN(n17336) );
  AND2_X1 U20528 ( .A1(n17336), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  AOI22_X1 U20529 ( .A1(n18774), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17310) );
  OAI21_X1 U20530 ( .B1(n17378), .B2(n17325), .A(n17310), .ZN(P3_U2737) );
  INV_X1 U20531 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17376) );
  AOI22_X1 U20532 ( .A1(n18774), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17311) );
  OAI21_X1 U20533 ( .B1(n17376), .B2(n17325), .A(n17311), .ZN(P3_U2738) );
  INV_X1 U20534 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17374) );
  AOI22_X1 U20535 ( .A1(n18774), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17312) );
  OAI21_X1 U20536 ( .B1(n17374), .B2(n17325), .A(n17312), .ZN(P3_U2739) );
  AOI22_X1 U20537 ( .A1(n18774), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17313) );
  OAI21_X1 U20538 ( .B1(n17372), .B2(n17325), .A(n17313), .ZN(P3_U2740) );
  INV_X1 U20539 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17370) );
  AOI22_X1 U20540 ( .A1(n18774), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17314) );
  OAI21_X1 U20541 ( .B1(n17370), .B2(n17325), .A(n17314), .ZN(P3_U2741) );
  AOI22_X1 U20542 ( .A1(n18774), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17315) );
  OAI21_X1 U20543 ( .B1(n17368), .B2(n17325), .A(n17315), .ZN(P3_U2742) );
  AOI22_X1 U20544 ( .A1(P3_UWORD_REG_8__SCAN_IN), .A2(n18774), .B1(n17336), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17316) );
  OAI21_X1 U20545 ( .B1(n17366), .B2(n17325), .A(n17316), .ZN(P3_U2743) );
  AOI22_X1 U20546 ( .A1(n18774), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17317) );
  OAI21_X1 U20547 ( .B1(n17364), .B2(n17325), .A(n17317), .ZN(P3_U2744) );
  CLKBUF_X1 U20548 ( .A(n18774), .Z(n18609) );
  AOI22_X1 U20549 ( .A1(n18609), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17318) );
  OAI21_X1 U20550 ( .B1(n17362), .B2(n17325), .A(n17318), .ZN(P3_U2745) );
  AOI22_X1 U20551 ( .A1(n18609), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17319) );
  OAI21_X1 U20552 ( .B1(n17360), .B2(n17325), .A(n17319), .ZN(P3_U2746) );
  AOI22_X1 U20553 ( .A1(n18609), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17320) );
  OAI21_X1 U20554 ( .B1(n17358), .B2(n17325), .A(n17320), .ZN(P3_U2747) );
  AOI22_X1 U20555 ( .A1(n18609), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17321) );
  OAI21_X1 U20556 ( .B1(n17356), .B2(n17325), .A(n17321), .ZN(P3_U2748) );
  AOI22_X1 U20557 ( .A1(n18609), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17322) );
  OAI21_X1 U20558 ( .B1(n17354), .B2(n17325), .A(n17322), .ZN(P3_U2749) );
  AOI22_X1 U20559 ( .A1(n18609), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17323) );
  OAI21_X1 U20560 ( .B1(n17352), .B2(n17325), .A(n17323), .ZN(P3_U2750) );
  AOI22_X1 U20561 ( .A1(n18609), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17324) );
  OAI21_X1 U20562 ( .B1(n17350), .B2(n17325), .A(n17324), .ZN(P3_U2751) );
  INV_X1 U20563 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17415) );
  AOI22_X1 U20564 ( .A1(n18609), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17327) );
  OAI21_X1 U20565 ( .B1(n17415), .B2(n17344), .A(n17327), .ZN(P3_U2752) );
  AOI22_X1 U20566 ( .A1(n18609), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17328) );
  OAI21_X1 U20567 ( .B1(n17410), .B2(n17344), .A(n17328), .ZN(P3_U2753) );
  INV_X1 U20568 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U20569 ( .A1(n18609), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17329) );
  OAI21_X1 U20570 ( .B1(n17408), .B2(n17344), .A(n17329), .ZN(P3_U2754) );
  AOI22_X1 U20571 ( .A1(n18609), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17330) );
  OAI21_X1 U20572 ( .B1(n17406), .B2(n17344), .A(n17330), .ZN(P3_U2755) );
  AOI22_X1 U20573 ( .A1(n18609), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17331) );
  OAI21_X1 U20574 ( .B1(n17403), .B2(n17344), .A(n17331), .ZN(P3_U2756) );
  AOI22_X1 U20575 ( .A1(n18609), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17332) );
  OAI21_X1 U20576 ( .B1(n17401), .B2(n17344), .A(n17332), .ZN(P3_U2757) );
  INV_X1 U20577 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U20578 ( .A1(n18609), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17333) );
  OAI21_X1 U20579 ( .B1(n17399), .B2(n17344), .A(n17333), .ZN(P3_U2758) );
  AOI22_X1 U20580 ( .A1(n18609), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17334) );
  OAI21_X1 U20581 ( .B1(n17397), .B2(n17344), .A(n17334), .ZN(P3_U2759) );
  AOI22_X1 U20582 ( .A1(n18609), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17335) );
  OAI21_X1 U20583 ( .B1(n17395), .B2(n17344), .A(n17335), .ZN(P3_U2760) );
  INV_X1 U20584 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17393) );
  AOI22_X1 U20585 ( .A1(n18609), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17337) );
  OAI21_X1 U20586 ( .B1(n17393), .B2(n17344), .A(n17337), .ZN(P3_U2761) );
  INV_X1 U20587 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17391) );
  AOI22_X1 U20588 ( .A1(n18609), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17338) );
  OAI21_X1 U20589 ( .B1(n17391), .B2(n17344), .A(n17338), .ZN(P3_U2762) );
  INV_X1 U20590 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17389) );
  AOI22_X1 U20591 ( .A1(n18609), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17339) );
  OAI21_X1 U20592 ( .B1(n17389), .B2(n17344), .A(n17339), .ZN(P3_U2763) );
  AOI22_X1 U20593 ( .A1(n18609), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17340) );
  OAI21_X1 U20594 ( .B1(n17387), .B2(n17344), .A(n17340), .ZN(P3_U2764) );
  AOI22_X1 U20595 ( .A1(n18609), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17341) );
  OAI21_X1 U20596 ( .B1(n17385), .B2(n17344), .A(n17341), .ZN(P3_U2765) );
  AOI22_X1 U20597 ( .A1(n18609), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17342) );
  OAI21_X1 U20598 ( .B1(n17383), .B2(n17344), .A(n17342), .ZN(P3_U2766) );
  AOI22_X1 U20599 ( .A1(n18609), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17336), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17343) );
  OAI21_X1 U20600 ( .B1(n17381), .B2(n17344), .A(n17343), .ZN(P3_U2767) );
  AOI22_X1 U20601 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17412), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17411), .ZN(n17349) );
  OAI21_X1 U20602 ( .B1(n17350), .B2(n17414), .A(n17349), .ZN(P3_U2768) );
  AOI22_X1 U20603 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17412), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17411), .ZN(n17351) );
  OAI21_X1 U20604 ( .B1(n17352), .B2(n17414), .A(n17351), .ZN(P3_U2769) );
  AOI22_X1 U20605 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17412), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17411), .ZN(n17353) );
  OAI21_X1 U20606 ( .B1(n17354), .B2(n17414), .A(n17353), .ZN(P3_U2770) );
  AOI22_X1 U20607 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17404), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17411), .ZN(n17355) );
  OAI21_X1 U20608 ( .B1(n17356), .B2(n17414), .A(n17355), .ZN(P3_U2771) );
  AOI22_X1 U20609 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17412), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17379), .ZN(n17357) );
  OAI21_X1 U20610 ( .B1(n17358), .B2(n17414), .A(n17357), .ZN(P3_U2772) );
  AOI22_X1 U20611 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17404), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17411), .ZN(n17359) );
  OAI21_X1 U20612 ( .B1(n17360), .B2(n17414), .A(n17359), .ZN(P3_U2773) );
  AOI22_X1 U20613 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17412), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17379), .ZN(n17361) );
  OAI21_X1 U20614 ( .B1(n17362), .B2(n17414), .A(n17361), .ZN(P3_U2774) );
  AOI22_X1 U20615 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17412), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17379), .ZN(n17363) );
  OAI21_X1 U20616 ( .B1(n17364), .B2(n17414), .A(n17363), .ZN(P3_U2775) );
  AOI22_X1 U20617 ( .A1(P3_UWORD_REG_8__SCAN_IN), .A2(n17411), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17412), .ZN(n17365) );
  OAI21_X1 U20618 ( .B1(n17366), .B2(n17414), .A(n17365), .ZN(P3_U2776) );
  AOI22_X1 U20619 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17412), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17379), .ZN(n17367) );
  OAI21_X1 U20620 ( .B1(n17368), .B2(n17414), .A(n17367), .ZN(P3_U2777) );
  AOI22_X1 U20621 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17412), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17379), .ZN(n17369) );
  OAI21_X1 U20622 ( .B1(n17370), .B2(n17414), .A(n17369), .ZN(P3_U2778) );
  AOI22_X1 U20623 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17412), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17379), .ZN(n17371) );
  OAI21_X1 U20624 ( .B1(n17372), .B2(n17414), .A(n17371), .ZN(P3_U2779) );
  AOI22_X1 U20625 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17412), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17379), .ZN(n17373) );
  OAI21_X1 U20626 ( .B1(n17374), .B2(n17414), .A(n17373), .ZN(P3_U2780) );
  AOI22_X1 U20627 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17412), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17379), .ZN(n17375) );
  OAI21_X1 U20628 ( .B1(n17376), .B2(n17414), .A(n17375), .ZN(P3_U2781) );
  AOI22_X1 U20629 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17412), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17379), .ZN(n17377) );
  OAI21_X1 U20630 ( .B1(n17378), .B2(n17414), .A(n17377), .ZN(P3_U2782) );
  AOI22_X1 U20631 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17412), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17379), .ZN(n17380) );
  OAI21_X1 U20632 ( .B1(n17381), .B2(n17414), .A(n17380), .ZN(P3_U2783) );
  AOI22_X1 U20633 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17412), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17411), .ZN(n17382) );
  OAI21_X1 U20634 ( .B1(n17383), .B2(n17414), .A(n17382), .ZN(P3_U2784) );
  AOI22_X1 U20635 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17412), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17411), .ZN(n17384) );
  OAI21_X1 U20636 ( .B1(n17385), .B2(n17414), .A(n17384), .ZN(P3_U2785) );
  AOI22_X1 U20637 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17412), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17411), .ZN(n17386) );
  OAI21_X1 U20638 ( .B1(n17387), .B2(n17414), .A(n17386), .ZN(P3_U2786) );
  AOI22_X1 U20639 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17404), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17411), .ZN(n17388) );
  OAI21_X1 U20640 ( .B1(n17389), .B2(n17414), .A(n17388), .ZN(P3_U2787) );
  AOI22_X1 U20641 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17404), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17411), .ZN(n17390) );
  OAI21_X1 U20642 ( .B1(n17391), .B2(n17414), .A(n17390), .ZN(P3_U2788) );
  AOI22_X1 U20643 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17404), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17411), .ZN(n17392) );
  OAI21_X1 U20644 ( .B1(n17393), .B2(n17414), .A(n17392), .ZN(P3_U2789) );
  AOI22_X1 U20645 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17404), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17411), .ZN(n17394) );
  OAI21_X1 U20646 ( .B1(n17395), .B2(n17414), .A(n17394), .ZN(P3_U2790) );
  AOI22_X1 U20647 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17404), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17411), .ZN(n17396) );
  OAI21_X1 U20648 ( .B1(n17397), .B2(n17414), .A(n17396), .ZN(P3_U2791) );
  AOI22_X1 U20649 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17404), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17411), .ZN(n17398) );
  OAI21_X1 U20650 ( .B1(n17399), .B2(n17414), .A(n17398), .ZN(P3_U2792) );
  AOI22_X1 U20651 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17404), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17411), .ZN(n17400) );
  OAI21_X1 U20652 ( .B1(n17401), .B2(n17414), .A(n17400), .ZN(P3_U2793) );
  AOI22_X1 U20653 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17404), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17411), .ZN(n17402) );
  OAI21_X1 U20654 ( .B1(n17403), .B2(n17414), .A(n17402), .ZN(P3_U2794) );
  AOI22_X1 U20655 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17404), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17411), .ZN(n17405) );
  OAI21_X1 U20656 ( .B1(n17406), .B2(n17414), .A(n17405), .ZN(P3_U2795) );
  AOI22_X1 U20657 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17412), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17411), .ZN(n17407) );
  OAI21_X1 U20658 ( .B1(n17408), .B2(n17414), .A(n17407), .ZN(P3_U2796) );
  AOI22_X1 U20659 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17412), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17411), .ZN(n17409) );
  OAI21_X1 U20660 ( .B1(n17410), .B2(n17414), .A(n17409), .ZN(P3_U2797) );
  AOI22_X1 U20661 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17412), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17411), .ZN(n17413) );
  OAI21_X1 U20662 ( .B1(n17415), .B2(n17414), .A(n17413), .ZN(P3_U2798) );
  INV_X1 U20663 ( .A(n17573), .ZN(n17512) );
  NAND2_X1 U20664 ( .A1(n17898), .A2(n17512), .ZN(n17550) );
  OAI21_X1 U20665 ( .B1(n17416), .B2(n17771), .A(n17770), .ZN(n17417) );
  AOI21_X1 U20666 ( .B1(n17600), .B2(n17420), .A(n17417), .ZN(n17448) );
  OAI21_X1 U20667 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17516), .A(
        n17448), .ZN(n17434) );
  NOR2_X1 U20668 ( .A1(n17607), .A2(n17762), .ZN(n17521) );
  OAI22_X1 U20669 ( .A1(n17783), .A2(n17678), .B1(n17782), .B2(n17775), .ZN(
        n17452) );
  NOR2_X1 U20670 ( .A1(n17792), .A2(n17452), .ZN(n17419) );
  NOR3_X1 U20671 ( .A1(n17521), .A2(n17419), .A3(n17418), .ZN(n17426) );
  NOR2_X1 U20672 ( .A1(n17612), .A2(n17420), .ZN(n17439) );
  OAI211_X1 U20673 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17439), .B(n17421), .ZN(n17422) );
  OAI211_X1 U20674 ( .C1(n17631), .C2(n17424), .A(n17423), .B(n17422), .ZN(
        n17425) );
  AOI211_X1 U20675 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17434), .A(
        n17426), .B(n17425), .ZN(n17431) );
  OAI211_X1 U20676 ( .C1(n17429), .C2(n17428), .A(n9608), .B(n17427), .ZN(
        n17430) );
  OAI211_X1 U20677 ( .C1(n17550), .C2(n17432), .A(n17431), .B(n17430), .ZN(
        P3_U2802) );
  AOI22_X1 U20678 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17434), .B1(
        n17605), .B2(n17433), .ZN(n17443) );
  NAND2_X1 U20679 ( .A1(n17436), .A2(n17435), .ZN(n17437) );
  XOR2_X1 U20680 ( .A(n17662), .B(n17437), .Z(n17789) );
  AOI22_X1 U20681 ( .A1(n17664), .A2(n17789), .B1(n17439), .B2(n17438), .ZN(
        n17442) );
  AOI22_X1 U20682 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17452), .B1(
        n17440), .B2(n17792), .ZN(n17441) );
  NAND2_X1 U20683 ( .A1(n9611), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17790) );
  NAND4_X1 U20684 ( .A1(n17443), .A2(n17442), .A3(n17441), .A4(n17790), .ZN(
        P3_U2803) );
  AOI21_X1 U20685 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17445), .A(
        n17444), .ZN(n17799) );
  AOI21_X1 U20686 ( .B1(n17446), .B2(n18493), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17447) );
  OAI22_X1 U20687 ( .A1(n17448), .A2(n17447), .B1(n17988), .B2(n18693), .ZN(
        n17449) );
  AOI221_X1 U20688 ( .B1(n17605), .B2(n17450), .C1(n12648), .C2(n17450), .A(
        n17449), .ZN(n17454) );
  INV_X1 U20689 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17794) );
  NAND3_X1 U20690 ( .A1(n17794), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17793) );
  INV_X1 U20691 ( .A(n17793), .ZN(n17451) );
  INV_X1 U20692 ( .A(n17550), .ZN(n17536) );
  AND3_X1 U20693 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17803), .A3(
        n17536), .ZN(n17476) );
  AOI22_X1 U20694 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17452), .B1(
        n17451), .B2(n17476), .ZN(n17453) );
  OAI211_X1 U20695 ( .C1(n17799), .C2(n17682), .A(n17454), .B(n17453), .ZN(
        P3_U2804) );
  NAND2_X1 U20696 ( .A1(n17845), .A2(n17801), .ZN(n17819) );
  NOR2_X1 U20697 ( .A1(n17819), .A2(n17825), .ZN(n17455) );
  XOR2_X1 U20698 ( .A(n17455), .B(n17810), .Z(n17817) );
  OAI21_X1 U20699 ( .B1(n17456), .B2(n17771), .A(n17770), .ZN(n17457) );
  AOI21_X1 U20700 ( .B1(n18493), .B2(n17458), .A(n17457), .ZN(n17484) );
  OAI21_X1 U20701 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17516), .A(
        n17484), .ZN(n17470) );
  NOR2_X1 U20702 ( .A1(n17612), .A2(n17458), .ZN(n17472) );
  OAI211_X1 U20703 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17472), .B(n17459), .ZN(n17460) );
  NAND2_X1 U20704 ( .A1(n9611), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17809) );
  OAI211_X1 U20705 ( .C1(n17631), .C2(n17461), .A(n17460), .B(n17809), .ZN(
        n17467) );
  NAND2_X1 U20706 ( .A1(n17847), .A2(n17801), .ZN(n17818) );
  NOR2_X1 U20707 ( .A1(n17818), .A2(n17825), .ZN(n17462) );
  XOR2_X1 U20708 ( .A(n17462), .B(n17810), .Z(n17812) );
  OAI21_X1 U20709 ( .B1(n17670), .B2(n17464), .A(n17463), .ZN(n17465) );
  XOR2_X1 U20710 ( .A(n17465), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17811) );
  OAI22_X1 U20711 ( .A1(n17812), .A2(n17678), .B1(n17682), .B2(n17811), .ZN(
        n17466) );
  AOI211_X1 U20712 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17470), .A(
        n17467), .B(n17466), .ZN(n17468) );
  OAI21_X1 U20713 ( .B1(n17817), .B2(n17775), .A(n17468), .ZN(P3_U2805) );
  INV_X1 U20714 ( .A(n17469), .ZN(n17479) );
  NOR2_X1 U20715 ( .A1(n17988), .A2(n18689), .ZN(n17830) );
  AOI221_X1 U20716 ( .B1(n17472), .B2(n17471), .C1(n17470), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17830), .ZN(n17478) );
  AOI22_X1 U20717 ( .A1(n17607), .A2(n17818), .B1(n17762), .B2(n17819), .ZN(
        n17488) );
  AOI21_X1 U20718 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17474), .A(
        n17473), .ZN(n17832) );
  OAI22_X1 U20719 ( .A1(n17488), .A2(n17825), .B1(n17832), .B2(n17682), .ZN(
        n17475) );
  AOI21_X1 U20720 ( .B1(n17476), .B2(n17825), .A(n17475), .ZN(n17477) );
  OAI211_X1 U20721 ( .C1(n17631), .C2(n17479), .A(n17478), .B(n17477), .ZN(
        P3_U2806) );
  NAND2_X1 U20722 ( .A1(n17803), .A2(n17536), .ZN(n17490) );
  AOI22_X1 U20723 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17670), .B1(
        n17480), .B2(n17492), .ZN(n17481) );
  NAND2_X1 U20724 ( .A1(n17522), .A2(n17481), .ZN(n17482) );
  XOR2_X1 U20725 ( .A(n17482), .B(n17489), .Z(n17836) );
  NOR2_X1 U20726 ( .A1(n17988), .A2(n18687), .ZN(n17835) );
  AOI21_X1 U20727 ( .B1(n9737), .B2(n18493), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17483) );
  OAI22_X1 U20728 ( .A1(n17754), .A2(n17485), .B1(n17484), .B2(n17483), .ZN(
        n17486) );
  AOI211_X1 U20729 ( .C1(n17836), .C2(n9608), .A(n17835), .B(n17486), .ZN(
        n17487) );
  OAI221_X1 U20730 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17490), 
        .C1(n17489), .C2(n17488), .A(n17487), .ZN(P3_U2807) );
  INV_X1 U20731 ( .A(n17851), .ZN(n17494) );
  INV_X1 U20732 ( .A(n17522), .ZN(n17491) );
  AOI221_X1 U20733 ( .B1(n12528), .B2(n17492), .C1(n17494), .C2(n17492), .A(
        n17491), .ZN(n17493) );
  XOR2_X1 U20734 ( .A(n17500), .B(n17493), .Z(n17857) );
  NOR2_X1 U20735 ( .A1(n9613), .A2(n17494), .ZN(n17501) );
  AOI22_X1 U20736 ( .A1(n17607), .A2(n17923), .B1(n17762), .B2(n17920), .ZN(
        n17571) );
  OAI21_X1 U20737 ( .B1(n17851), .B2(n17521), .A(n17571), .ZN(n17513) );
  OAI21_X1 U20738 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17516), .A(
        n9624), .ZN(n17508) );
  NOR2_X1 U20739 ( .A1(n17612), .A2(n17497), .ZN(n17510) );
  OAI211_X1 U20740 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17510), .B(n17498), .ZN(n17499) );
  NOR3_X1 U20741 ( .A1(n17670), .A2(n17897), .A3(n17502), .ZN(n17528) );
  INV_X1 U20742 ( .A(n17503), .ZN(n17546) );
  AOI22_X1 U20743 ( .A1(n17860), .A2(n17528), .B1(n17546), .B2(n17504), .ZN(
        n17505) );
  XOR2_X1 U20744 ( .A(n17505), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(
        n17867) );
  OAI22_X1 U20745 ( .A1(n18683), .A2(n17988), .B1(n17631), .B2(n17506), .ZN(
        n17507) );
  AOI221_X1 U20746 ( .B1(n17510), .B2(n17509), .C1(n17508), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17507), .ZN(n17515) );
  INV_X1 U20747 ( .A(n17860), .ZN(n17511) );
  NOR3_X1 U20748 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17862), .A3(
        n17511), .ZN(n17858) );
  AOI22_X1 U20749 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17513), .B1(
        n17858), .B2(n17512), .ZN(n17514) );
  OAI211_X1 U20750 ( .C1(n17867), .C2(n17682), .A(n17515), .B(n17514), .ZN(
        P3_U2809) );
  NOR2_X1 U20751 ( .A1(n17862), .A2(n17523), .ZN(n17872) );
  NAND2_X1 U20752 ( .A1(n17872), .A2(n17525), .ZN(n17877) );
  AOI21_X1 U20753 ( .B1(n17517), .B2(n18493), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17518) );
  OAI22_X1 U20754 ( .A1(n9624), .A2(n17518), .B1(n17988), .B2(n18682), .ZN(
        n17519) );
  AOI221_X1 U20755 ( .B1(n17605), .B2(n17520), .C1(n12648), .C2(n17520), .A(
        n17519), .ZN(n17527) );
  OAI21_X1 U20756 ( .B1(n17521), .B2(n17872), .A(n17571), .ZN(n17537) );
  OAI221_X1 U20757 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17545), 
        .C1(n17523), .C2(n17528), .A(n17522), .ZN(n17524) );
  XOR2_X1 U20758 ( .A(n17525), .B(n17524), .Z(n17868) );
  AOI22_X1 U20759 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17537), .B1(
        n9608), .B2(n17868), .ZN(n17526) );
  OAI211_X1 U20760 ( .C1(n9613), .C2(n17877), .A(n17527), .B(n17526), .ZN(
        P3_U2810) );
  AOI21_X1 U20761 ( .B1(n17546), .B2(n17545), .A(n17528), .ZN(n17529) );
  XOR2_X1 U20762 ( .A(n17529), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n17883) );
  AOI21_X1 U20763 ( .B1(n17600), .B2(n17531), .A(n17757), .ZN(n17553) );
  OAI21_X1 U20764 ( .B1(n17530), .B2(n17771), .A(n17553), .ZN(n17542) );
  NOR2_X1 U20765 ( .A1(n17612), .A2(n17531), .ZN(n17544) );
  OAI211_X1 U20766 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17544), .B(n17532), .ZN(n17533) );
  NAND2_X1 U20767 ( .A1(n9611), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17881) );
  OAI211_X1 U20768 ( .C1(n17631), .C2(n17534), .A(n17533), .B(n17881), .ZN(
        n17535) );
  AOI21_X1 U20769 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17542), .A(
        n17535), .ZN(n17539) );
  NOR2_X1 U20770 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17897), .ZN(
        n17878) );
  AOI22_X1 U20771 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17537), .B1(
        n17536), .B2(n17878), .ZN(n17538) );
  OAI211_X1 U20772 ( .C1(n17883), .C2(n17682), .A(n17539), .B(n17538), .ZN(
        P3_U2811) );
  OAI22_X1 U20773 ( .A1(n17988), .A2(n18677), .B1(n17631), .B2(n17540), .ZN(
        n17541) );
  AOI221_X1 U20774 ( .B1(n17544), .B2(n17543), .C1(n17542), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17541), .ZN(n17549) );
  OAI21_X1 U20775 ( .B1(n17898), .B2(n9613), .A(n17571), .ZN(n17558) );
  AOI21_X1 U20776 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17662), .A(
        n17545), .ZN(n17547) );
  XOR2_X1 U20777 ( .A(n17547), .B(n17546), .Z(n17890) );
  AOI22_X1 U20778 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17558), .B1(
        n9608), .B2(n17890), .ZN(n17548) );
  OAI211_X1 U20779 ( .C1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n17550), .A(
        n17549), .B(n17548), .ZN(P3_U2812) );
  NAND2_X1 U20780 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17902), .ZN(
        n17908) );
  AOI21_X1 U20781 ( .B1(n17551), .B2(n18493), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17554) );
  OAI22_X1 U20782 ( .A1(n17554), .A2(n17553), .B1(n17754), .B2(n17552), .ZN(
        n17555) );
  AOI21_X1 U20783 ( .B1(n9611), .B2(P3_REIP_REG_17__SCAN_IN), .A(n17555), .ZN(
        n17560) );
  OAI21_X1 U20784 ( .B1(n17557), .B2(n17902), .A(n17556), .ZN(n17906) );
  AOI22_X1 U20785 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17558), .B1(
        n17664), .B2(n17906), .ZN(n17559) );
  OAI211_X1 U20786 ( .C1(n9613), .C2(n17908), .A(n17560), .B(n17559), .ZN(
        P3_U2813) );
  AOI21_X1 U20787 ( .B1(n17662), .B2(n12528), .A(n17561), .ZN(n17562) );
  XOR2_X1 U20788 ( .A(n17562), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(
        n17915) );
  AOI21_X1 U20789 ( .B1(n17600), .B2(n17565), .A(n17757), .ZN(n17592) );
  OAI21_X1 U20790 ( .B1(n17563), .B2(n17771), .A(n17592), .ZN(n17576) );
  AOI22_X1 U20791 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17576), .B1(
        n17605), .B2(n17564), .ZN(n17568) );
  NAND2_X1 U20792 ( .A1(n9611), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17917) );
  NOR2_X1 U20793 ( .A1(n17612), .A2(n17565), .ZN(n17578) );
  OAI211_X1 U20794 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17578), .B(n17566), .ZN(n17567) );
  NAND3_X1 U20795 ( .A1(n17568), .A2(n17917), .A3(n17567), .ZN(n17569) );
  AOI21_X1 U20796 ( .B1(n17664), .B2(n17915), .A(n17569), .ZN(n17570) );
  OAI221_X1 U20797 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n9613), .C1(
        n17572), .C2(n17571), .A(n17570), .ZN(P3_U2814) );
  INV_X1 U20798 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17942) );
  NOR3_X1 U20799 ( .A1(n17960), .A2(n17942), .A3(n17955), .ZN(n17594) );
  NOR2_X1 U20800 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17594), .ZN(
        n17933) );
  NAND2_X1 U20801 ( .A1(n17762), .A2(n17920), .ZN(n17587) );
  OAI22_X1 U20802 ( .A1(n17988), .A2(n18671), .B1(n17631), .B2(n17574), .ZN(
        n17575) );
  AOI221_X1 U20803 ( .B1(n17578), .B2(n17577), .C1(n17576), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17575), .ZN(n17586) );
  NAND2_X1 U20804 ( .A1(n17974), .A2(n17942), .ZN(n17581) );
  NOR2_X1 U20805 ( .A1(n17670), .A2(n17974), .ZN(n17608) );
  INV_X1 U20806 ( .A(n17608), .ZN(n17580) );
  NOR3_X1 U20807 ( .A1(n17662), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n12524), .ZN(n17646) );
  INV_X1 U20808 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17997) );
  NAND2_X1 U20809 ( .A1(n17646), .A2(n17997), .ZN(n17633) );
  NOR2_X1 U20810 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17633), .ZN(
        n17621) );
  NAND2_X1 U20811 ( .A1(n17621), .A2(n17960), .ZN(n17596) );
  AOI22_X1 U20812 ( .A1(n17581), .A2(n17580), .B1(n17579), .B2(n17596), .ZN(
        n17582) );
  XOR2_X1 U20813 ( .A(n17582), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n17928) );
  NOR2_X1 U20814 ( .A1(n17847), .A2(n17678), .ZN(n17584) );
  INV_X1 U20815 ( .A(n17975), .ZN(n17637) );
  NOR2_X1 U20816 ( .A1(n17595), .A2(n17942), .ZN(n17921) );
  AOI21_X1 U20817 ( .B1(n17637), .B2(n17921), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17925) );
  INV_X1 U20818 ( .A(n17925), .ZN(n17583) );
  AOI22_X1 U20819 ( .A1(n9608), .A2(n17928), .B1(n17584), .B2(n17583), .ZN(
        n17585) );
  OAI211_X1 U20820 ( .C1(n17933), .C2(n17587), .A(n17586), .B(n17585), .ZN(
        P3_U2815) );
  INV_X1 U20821 ( .A(n17921), .ZN(n17913) );
  OAI22_X1 U20822 ( .A1(n17588), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n17975), .B2(n17913), .ZN(n17949) );
  AOI21_X1 U20823 ( .B1(n17589), .B2(n18493), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17591) );
  OAI22_X1 U20824 ( .A1(n17592), .A2(n17591), .B1(n17754), .B2(n17590), .ZN(
        n17593) );
  AOI21_X1 U20825 ( .B1(n9611), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17593), .ZN(
        n17599) );
  INV_X1 U20826 ( .A(n17636), .ZN(n17977) );
  AOI221_X1 U20827 ( .B1(n17977), .B2(n17942), .C1(n17595), .C2(n17942), .A(
        n17594), .ZN(n17946) );
  NOR2_X1 U20828 ( .A1(n17670), .A2(n17975), .ZN(n17647) );
  INV_X1 U20829 ( .A(n17647), .ZN(n17661) );
  OAI22_X1 U20830 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17596), .B1(
        n17661), .B2(n17595), .ZN(n17597) );
  XOR2_X1 U20831 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17597), .Z(
        n17945) );
  AOI22_X1 U20832 ( .A1(n17762), .A2(n17946), .B1(n9608), .B2(n17945), .ZN(
        n17598) );
  OAI211_X1 U20833 ( .C1(n17678), .C2(n17949), .A(n17599), .B(n17598), .ZN(
        P3_U2816) );
  AOI22_X1 U20834 ( .A1(n17602), .A2(n17601), .B1(n17600), .B2(n17640), .ZN(
        n17603) );
  NAND2_X1 U20835 ( .A1(n17603), .A2(n17770), .ZN(n17618) );
  AOI22_X1 U20836 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17618), .B1(
        n17605), .B2(n17604), .ZN(n17616) );
  NOR2_X1 U20837 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17936), .ZN(
        n17963) );
  AOI22_X1 U20838 ( .A1(n17636), .A2(n17762), .B1(n17607), .B2(n17637), .ZN(
        n17668) );
  INV_X1 U20839 ( .A(n17668), .ZN(n17635) );
  NAND2_X1 U20840 ( .A1(n17637), .A2(n17606), .ZN(n17954) );
  AOI22_X1 U20841 ( .A1(n17607), .A2(n17954), .B1(n17762), .B2(n17955), .ZN(
        n17624) );
  OAI22_X1 U20842 ( .A1(n17609), .A2(n17974), .B1(n17608), .B2(n17621), .ZN(
        n17610) );
  XOR2_X1 U20843 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17610), .Z(
        n17966) );
  OAI22_X1 U20844 ( .A1(n17624), .A2(n17960), .B1(n17682), .B2(n17966), .ZN(
        n17611) );
  AOI21_X1 U20845 ( .B1(n17963), .B2(n17635), .A(n17611), .ZN(n17615) );
  NAND2_X1 U20846 ( .A1(n9611), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17964) );
  NOR2_X1 U20847 ( .A1(n17612), .A2(n17640), .ZN(n17620) );
  OAI211_X1 U20848 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17620), .B(n17613), .ZN(n17614) );
  NAND4_X1 U20849 ( .A1(n17616), .A2(n17615), .A3(n17964), .A4(n17614), .ZN(
        P3_U2817) );
  INV_X1 U20850 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18665) );
  NOR2_X1 U20851 ( .A1(n17988), .A2(n18665), .ZN(n17617) );
  AOI221_X1 U20852 ( .B1(n17620), .B2(n17619), .C1(n17618), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17617), .ZN(n17629) );
  INV_X1 U20853 ( .A(n17621), .ZN(n17622) );
  OAI21_X1 U20854 ( .B1(n17968), .B2(n17661), .A(n17622), .ZN(n17623) );
  XOR2_X1 U20855 ( .A(n17623), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n17967) );
  NOR2_X1 U20856 ( .A1(n17668), .A2(n17968), .ZN(n17626) );
  INV_X1 U20857 ( .A(n17624), .ZN(n17625) );
  MUX2_X1 U20858 ( .A(n17626), .B(n17625), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n17627) );
  AOI21_X1 U20859 ( .B1(n9608), .B2(n17967), .A(n17627), .ZN(n17628) );
  OAI211_X1 U20860 ( .C1(n17631), .C2(n17630), .A(n17629), .B(n17628), .ZN(
        P3_U2818) );
  AOI22_X1 U20861 ( .A1(n9611), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17632), 
        .B2(n17764), .ZN(n17644) );
  OAI21_X1 U20862 ( .B1(n17982), .B2(n17661), .A(n17633), .ZN(n17634) );
  XOR2_X1 U20863 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17634), .Z(
        n17986) );
  NOR2_X1 U20864 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17982), .ZN(
        n17985) );
  AOI22_X1 U20865 ( .A1(n17664), .A2(n17986), .B1(n17985), .B2(n17635), .ZN(
        n17643) );
  NOR2_X1 U20866 ( .A1(n17952), .A2(n17668), .ZN(n17649) );
  OAI22_X1 U20867 ( .A1(n17637), .A2(n17678), .B1(n17775), .B2(n17636), .ZN(
        n17665) );
  OAI21_X1 U20868 ( .B1(n17649), .B2(n17665), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17642) );
  NOR2_X1 U20869 ( .A1(n17671), .A2(n18456), .ZN(n17686) );
  NAND3_X1 U20870 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(n17686), .ZN(n17658) );
  NOR2_X1 U20871 ( .A1(n17657), .A2(n17658), .ZN(n17655) );
  NAND2_X1 U20872 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17655), .ZN(
        n17650) );
  OAI21_X1 U20873 ( .B1(n17656), .B2(n17638), .A(n17650), .ZN(n17639) );
  OAI21_X1 U20874 ( .B1(n18456), .B2(n17640), .A(n17639), .ZN(n17641) );
  NAND4_X1 U20875 ( .A1(n17644), .A2(n17643), .A3(n17642), .A4(n17641), .ZN(
        P3_U2819) );
  AOI22_X1 U20876 ( .A1(n9611), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17645), 
        .B2(n17764), .ZN(n17654) );
  AOI21_X1 U20877 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17647), .A(
        n17646), .ZN(n17648) );
  XOR2_X1 U20878 ( .A(n17997), .B(n17648), .Z(n17990) );
  AOI22_X1 U20879 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17665), .B1(
        n9608), .B2(n17990), .ZN(n17653) );
  OAI21_X1 U20880 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17649), .ZN(n17652) );
  OAI211_X1 U20881 ( .C1(n17655), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17765), .B(n17650), .ZN(n17651) );
  NAND4_X1 U20882 ( .A1(n17654), .A2(n17653), .A3(n17652), .A4(n17651), .ZN(
        P3_U2820) );
  AOI211_X1 U20883 ( .C1(n17658), .C2(n17657), .A(n17656), .B(n17655), .ZN(
        n17659) );
  NOR2_X1 U20884 ( .A1(n17988), .A2(n18659), .ZN(n18007) );
  AOI211_X1 U20885 ( .C1(n17660), .C2(n17764), .A(n17659), .B(n18007), .ZN(
        n17667) );
  OAI21_X1 U20886 ( .B1(n12524), .B2(n17662), .A(n17661), .ZN(n17663) );
  XOR2_X1 U20887 ( .A(n17663), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18008) );
  AOI22_X1 U20888 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17665), .B1(
        n17664), .B2(n18008), .ZN(n17666) );
  OAI211_X1 U20889 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17668), .A(
        n17667), .B(n17666), .ZN(P3_U2821) );
  AOI21_X1 U20890 ( .B1(n17670), .B2(n18028), .A(n17669), .ZN(n18022) );
  OAI21_X1 U20891 ( .B1(n9886), .B2(n17728), .A(n17770), .ZN(n17687) );
  OAI211_X1 U20892 ( .C1(n17673), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n18493), .B(n17672), .ZN(n17674) );
  NAND2_X1 U20893 ( .A1(n9611), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18018) );
  OAI211_X1 U20894 ( .C1(n17754), .C2(n17675), .A(n17674), .B(n18018), .ZN(
        n17680) );
  OAI21_X1 U20895 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17677), .A(
        n17676), .ZN(n18020) );
  OAI22_X1 U20896 ( .A1(n17678), .A2(n18028), .B1(n17775), .B2(n18020), .ZN(
        n17679) );
  AOI211_X1 U20897 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17687), .A(
        n17680), .B(n17679), .ZN(n17681) );
  OAI21_X1 U20898 ( .B1(n18022), .B2(n17682), .A(n17681), .ZN(P3_U2822) );
  OAI21_X1 U20899 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17684), .A(
        n17683), .ZN(n18031) );
  NOR2_X1 U20900 ( .A1(n17988), .A2(n18655), .ZN(n18030) );
  AOI221_X1 U20901 ( .B1(n17687), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n17686), .C2(n17685), .A(n18030), .ZN(n17695) );
  AOI21_X1 U20902 ( .B1(n17690), .B2(n17689), .A(n17688), .ZN(n17692) );
  XNOR2_X1 U20903 ( .A(n17692), .B(n17691), .ZN(n18033) );
  AOI22_X1 U20904 ( .A1(n17762), .A2(n18033), .B1(n17693), .B2(n17764), .ZN(
        n17694) );
  OAI211_X1 U20905 ( .C1(n17774), .C2(n18031), .A(n17695), .B(n17694), .ZN(
        P3_U2823) );
  OAI21_X1 U20906 ( .B1(n17698), .B2(n17697), .A(n17696), .ZN(n18039) );
  NAND2_X1 U20907 ( .A1(n17699), .A2(n18493), .ZN(n17702) );
  OAI21_X1 U20908 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17701), .A(
        n17700), .ZN(n18044) );
  OAI22_X1 U20909 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17702), .B1(
        n17775), .B2(n18044), .ZN(n17707) );
  INV_X1 U20910 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17704) );
  OAI21_X1 U20911 ( .B1(n18456), .B2(n17703), .A(n17765), .ZN(n17718) );
  OAI22_X1 U20912 ( .A1(n17754), .A2(n17705), .B1(n17704), .B2(n17718), .ZN(
        n17706) );
  AOI211_X1 U20913 ( .C1(n9611), .C2(P3_REIP_REG_6__SCAN_IN), .A(n17707), .B(
        n17706), .ZN(n17708) );
  OAI21_X1 U20914 ( .B1(n17774), .B2(n18039), .A(n17708), .ZN(P3_U2824) );
  OAI21_X1 U20915 ( .B1(n17711), .B2(n17710), .A(n17709), .ZN(n18053) );
  OAI21_X1 U20916 ( .B1(n17714), .B2(n17713), .A(n17712), .ZN(n17716) );
  XOR2_X1 U20917 ( .A(n17716), .B(n17715), .Z(n18049) );
  AOI22_X1 U20918 ( .A1(n17717), .A2(n18049), .B1(n9611), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17724) );
  AOI221_X1 U20919 ( .B1(n17757), .B2(n17720), .C1(n17719), .C2(n17720), .A(
        n17718), .ZN(n17721) );
  AOI21_X1 U20920 ( .B1(n17722), .B2(n17764), .A(n17721), .ZN(n17723) );
  OAI211_X1 U20921 ( .C1(n17775), .C2(n18053), .A(n17724), .B(n17723), .ZN(
        P3_U2825) );
  OAI21_X1 U20922 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17726), .A(
        n17725), .ZN(n18056) );
  AOI22_X1 U20923 ( .A1(n9611), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18493), .B2(
        n17727), .ZN(n17734) );
  OAI21_X1 U20924 ( .B1(n17729), .B2(n17728), .A(n17770), .ZN(n17744) );
  OAI22_X1 U20925 ( .A1(n17754), .A2(n17731), .B1(n17774), .B2(n18062), .ZN(
        n17732) );
  AOI21_X1 U20926 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17744), .A(
        n17732), .ZN(n17733) );
  OAI211_X1 U20927 ( .C1(n17775), .C2(n18056), .A(n17734), .B(n17733), .ZN(
        P3_U2826) );
  OAI21_X1 U20928 ( .B1(n17737), .B2(n17736), .A(n17735), .ZN(n18064) );
  NOR2_X1 U20929 ( .A1(n17757), .A2(n17756), .ZN(n17743) );
  OAI21_X1 U20930 ( .B1(n17740), .B2(n17739), .A(n17738), .ZN(n18071) );
  OAI22_X1 U20931 ( .A1(n17754), .A2(n17741), .B1(n17774), .B2(n18071), .ZN(
        n17742) );
  AOI221_X1 U20932 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17744), .C1(
        n17743), .C2(n17744), .A(n17742), .ZN(n17745) );
  NAND2_X1 U20933 ( .A1(n9611), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18069) );
  OAI211_X1 U20934 ( .C1(n17775), .C2(n18064), .A(n17745), .B(n18069), .ZN(
        P3_U2827) );
  OAI21_X1 U20935 ( .B1(n17748), .B2(n17747), .A(n17746), .ZN(n18082) );
  INV_X1 U20936 ( .A(n17749), .ZN(n17753) );
  OAI21_X1 U20937 ( .B1(n17752), .B2(n17751), .A(n17750), .ZN(n18081) );
  OAI22_X1 U20938 ( .A1(n17754), .A2(n17753), .B1(n17774), .B2(n18081), .ZN(
        n17755) );
  AOI221_X1 U20939 ( .B1(n17757), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18493), .C2(n17756), .A(n17755), .ZN(n17758) );
  NAND2_X1 U20940 ( .A1(n9611), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18086) );
  OAI211_X1 U20941 ( .C1(n17775), .C2(n18082), .A(n17758), .B(n18086), .ZN(
        P3_U2828) );
  OAI21_X1 U20942 ( .B1(n17768), .B2(n17760), .A(n17759), .ZN(n18100) );
  NAND2_X1 U20943 ( .A1(n18725), .A2(n17769), .ZN(n17761) );
  XNOR2_X1 U20944 ( .A(n17761), .B(n17760), .ZN(n18096) );
  AOI22_X1 U20945 ( .A1(n17762), .A2(n18096), .B1(n9611), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17767) );
  AOI22_X1 U20946 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17765), .B1(
        n17764), .B2(n17763), .ZN(n17766) );
  OAI211_X1 U20947 ( .C1(n17774), .C2(n18100), .A(n17767), .B(n17766), .ZN(
        P3_U2829) );
  AOI21_X1 U20948 ( .B1(n17769), .B2(n18725), .A(n17768), .ZN(n18111) );
  INV_X1 U20949 ( .A(n18111), .ZN(n18109) );
  NAND3_X1 U20950 ( .A1(n18726), .A2(n17771), .A3(n17770), .ZN(n17772) );
  AOI22_X1 U20951 ( .A1(n9611), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17772), .ZN(n17773) );
  OAI221_X1 U20952 ( .B1(n18111), .B2(n17775), .C1(n18109), .C2(n17774), .A(
        n17773), .ZN(P3_U2830) );
  AOI21_X1 U20953 ( .B1(n17792), .B2(n17776), .A(n18016), .ZN(n17788) );
  INV_X1 U20954 ( .A(n18583), .ZN(n18572) );
  AOI21_X1 U20955 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18572), .A(
        n17777), .ZN(n17848) );
  NAND2_X1 U20956 ( .A1(n17851), .A2(n17884), .ZN(n17778) );
  OAI21_X1 U20957 ( .B1(n17848), .B2(n17778), .A(n18077), .ZN(n17820) );
  OAI21_X1 U20958 ( .B1(n17889), .B2(n17779), .A(n17820), .ZN(n17804) );
  INV_X1 U20959 ( .A(n17780), .ZN(n17781) );
  OAI22_X1 U20960 ( .A1(n18585), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18572), .B2(n17781), .ZN(n17785) );
  OAI22_X1 U20961 ( .A1(n17783), .A2(n17846), .B1(n17782), .B2(n17844), .ZN(
        n17784) );
  NOR4_X1 U20962 ( .A1(n17786), .A2(n17804), .A3(n17785), .A4(n17784), .ZN(
        n17795) );
  OAI211_X1 U20963 ( .C1(n18585), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17795), .ZN(n17787) );
  AOI22_X1 U20964 ( .A1(n18009), .A2(n17789), .B1(n17788), .B2(n17787), .ZN(
        n17791) );
  OAI211_X1 U20965 ( .C1(n18089), .C2(n17792), .A(n17791), .B(n17790), .ZN(
        P3_U2835) );
  NAND3_X1 U20966 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17833), .A3(
        n17850), .ZN(n17827) );
  OAI22_X1 U20967 ( .A1(n17795), .A2(n17794), .B1(n17793), .B2(n17827), .ZN(
        n17796) );
  AOI22_X1 U20968 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18092), .B1(
        n18101), .B2(n17796), .ZN(n17798) );
  NAND2_X1 U20969 ( .A1(n9611), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17797) );
  OAI211_X1 U20970 ( .C1(n17799), .C2(n18021), .A(n17798), .B(n17797), .ZN(
        P3_U2836) );
  NOR2_X1 U20971 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17825), .ZN(
        n17800) );
  NAND2_X1 U20972 ( .A1(n17801), .A2(n17800), .ZN(n17807) );
  AOI21_X1 U20973 ( .B1(n17898), .B2(n17840), .A(n9932), .ZN(n17802) );
  INV_X1 U20974 ( .A(n17802), .ZN(n17885) );
  OAI21_X1 U20975 ( .B1(n17803), .B2(n9932), .A(n17885), .ZN(n17822) );
  AOI211_X1 U20976 ( .C1(n18581), .C2(n17805), .A(n17804), .B(n17822), .ZN(
        n17806) );
  OAI22_X1 U20977 ( .A1(n17808), .A2(n17807), .B1(n17806), .B2(n17810), .ZN(
        n17815) );
  OAI21_X1 U20978 ( .B1(n18089), .B2(n17810), .A(n17809), .ZN(n17814) );
  OAI22_X1 U20979 ( .A1(n17812), .A2(n18027), .B1(n18021), .B2(n17811), .ZN(
        n17813) );
  AOI211_X1 U20980 ( .C1(n18101), .C2(n17815), .A(n17814), .B(n17813), .ZN(
        n17816) );
  OAI21_X1 U20981 ( .B1(n17817), .B2(n18110), .A(n17816), .ZN(P3_U2837) );
  AOI22_X1 U20982 ( .A1(n18549), .A2(n17819), .B1(n17976), .B2(n17818), .ZN(
        n17821) );
  AND3_X1 U20983 ( .A1(n17821), .A2(n18089), .A3(n17820), .ZN(n17826) );
  INV_X1 U20984 ( .A(n17822), .ZN(n17823) );
  NAND3_X1 U20985 ( .A1(n17823), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17826), .ZN(n17824) );
  NAND2_X1 U20986 ( .A1(n17988), .A2(n17824), .ZN(n17838) );
  AOI211_X1 U20987 ( .C1(n9622), .C2(n17826), .A(n17825), .B(n17838), .ZN(
        n17829) );
  NOR3_X1 U20988 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18016), .A3(
        n17827), .ZN(n17828) );
  NOR3_X1 U20989 ( .A1(n17830), .A2(n17829), .A3(n17828), .ZN(n17831) );
  OAI21_X1 U20990 ( .B1(n17832), .B2(n18021), .A(n17831), .ZN(P3_U2838) );
  AND2_X1 U20991 ( .A1(n17850), .A2(n17833), .ZN(n17834) );
  AOI21_X1 U20992 ( .B1(n17834), .B2(n18089), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17839) );
  AOI21_X1 U20993 ( .B1(n17836), .B2(n18009), .A(n17835), .ZN(n17837) );
  OAI21_X1 U20994 ( .B1(n17839), .B2(n17838), .A(n17837), .ZN(P3_U2839) );
  NOR2_X1 U20995 ( .A1(n17988), .A2(n18685), .ZN(n17855) );
  INV_X1 U20996 ( .A(n17840), .ZN(n17841) );
  OAI21_X1 U20997 ( .B1(n17862), .B2(n17841), .A(n18581), .ZN(n17842) );
  OAI221_X1 U20998 ( .B1(n18585), .B2(n17884), .C1(n18585), .C2(n17872), .A(
        n17842), .ZN(n17870) );
  NAND2_X1 U20999 ( .A1(n17844), .A2(n17846), .ZN(n17981) );
  INV_X1 U21000 ( .A(n17981), .ZN(n17886) );
  OAI22_X1 U21001 ( .A1(n18585), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17851), .B2(n17886), .ZN(n17843) );
  NOR2_X1 U21002 ( .A1(n17870), .A2(n17843), .ZN(n17859) );
  OAI22_X1 U21003 ( .A1(n17847), .A2(n17846), .B1(n17845), .B2(n17844), .ZN(
        n17861) );
  AOI211_X1 U21004 ( .C1(n17849), .C2(n17959), .A(n17848), .B(n17861), .ZN(
        n17853) );
  AOI21_X1 U21005 ( .B1(n17851), .B2(n17850), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17852) );
  AOI211_X1 U21006 ( .C1(n17859), .C2(n17853), .A(n17852), .B(n18016), .ZN(
        n17854) );
  AOI211_X1 U21007 ( .C1(n18092), .C2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n17855), .B(n17854), .ZN(n17856) );
  OAI21_X1 U21008 ( .B1(n18021), .B2(n17857), .A(n17856), .ZN(P3_U2840) );
  INV_X1 U21009 ( .A(n17876), .ZN(n17879) );
  AOI22_X1 U21010 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n9611), .B1(n17879), 
        .B2(n17858), .ZN(n17866) );
  OAI21_X1 U21011 ( .B1(n17860), .B2(n17938), .A(n17859), .ZN(n17864) );
  NOR2_X1 U21012 ( .A1(n18016), .A2(n17861), .ZN(n17914) );
  OAI21_X1 U21013 ( .B1(n17862), .B2(n17909), .A(n18583), .ZN(n17863) );
  NAND2_X1 U21014 ( .A1(n17914), .A2(n17863), .ZN(n17869) );
  OAI211_X1 U21015 ( .C1(n17864), .C2(n17869), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17988), .ZN(n17865) );
  OAI211_X1 U21016 ( .C1(n17867), .C2(n18021), .A(n17866), .B(n17865), .ZN(
        P3_U2841) );
  AOI22_X1 U21017 ( .A1(n9611), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18009), 
        .B2(n17868), .ZN(n17875) );
  NOR2_X1 U21018 ( .A1(n17870), .A2(n17869), .ZN(n17871) );
  AOI221_X1 U21019 ( .B1(n17872), .B2(n17871), .C1(n17886), .C2(n17871), .A(
        n9611), .ZN(n17880) );
  NOR3_X1 U21020 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17938), .A3(
        n18779), .ZN(n17873) );
  OAI21_X1 U21021 ( .B1(n17880), .B2(n17873), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17874) );
  OAI211_X1 U21022 ( .C1(n17877), .C2(n17876), .A(n17875), .B(n17874), .ZN(
        P3_U2842) );
  AOI22_X1 U21023 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17880), .B1(
        n17879), .B2(n17878), .ZN(n17882) );
  OAI211_X1 U21024 ( .C1(n17883), .C2(n18021), .A(n17882), .B(n17881), .ZN(
        P3_U2843) );
  NAND2_X1 U21025 ( .A1(n18583), .A2(n18725), .ZN(n18074) );
  NAND3_X1 U21026 ( .A1(n17884), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18074), .ZN(n17888) );
  OAI211_X1 U21027 ( .C1(n17898), .C2(n17886), .A(n17914), .B(n17885), .ZN(
        n17887) );
  AOI21_X1 U21028 ( .B1(n18077), .B2(n17888), .A(n17887), .ZN(n17903) );
  AOI221_X1 U21029 ( .B1(n17889), .B2(n17903), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17903), .A(n9611), .ZN(
        n17891) );
  AOI22_X1 U21030 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17891), .B1(
        n18009), .B2(n17890), .ZN(n17900) );
  NAND2_X1 U21031 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18054) );
  OAI22_X1 U21032 ( .A1(n17892), .A2(n9932), .B1(n18073), .B2(n18054), .ZN(
        n18067) );
  NAND2_X1 U21033 ( .A1(n17893), .A2(n18067), .ZN(n17950) );
  NOR2_X1 U21034 ( .A1(n17951), .A2(n17950), .ZN(n17922) );
  NAND2_X1 U21035 ( .A1(n17894), .A2(n17922), .ZN(n17941) );
  AOI211_X1 U21036 ( .C1(n17896), .C2(n17941), .A(n17895), .B(n18016), .ZN(
        n17901) );
  NAND3_X1 U21037 ( .A1(n17898), .A2(n17901), .A3(n17897), .ZN(n17899) );
  OAI211_X1 U21038 ( .C1(n18677), .C2(n17988), .A(n17900), .B(n17899), .ZN(
        P3_U2844) );
  INV_X1 U21039 ( .A(n17901), .ZN(n17919) );
  NOR2_X1 U21040 ( .A1(n17988), .A2(n18676), .ZN(n17905) );
  NOR3_X1 U21041 ( .A1(n9611), .A2(n17903), .A3(n17902), .ZN(n17904) );
  AOI211_X1 U21042 ( .C1(n18009), .C2(n17906), .A(n17905), .B(n17904), .ZN(
        n17907) );
  OAI21_X1 U21043 ( .B1(n17919), .B2(n17908), .A(n17907), .ZN(P3_U2845) );
  OAI21_X1 U21044 ( .B1(n17910), .B2(n18583), .A(n17909), .ZN(n17911) );
  INV_X1 U21045 ( .A(n17911), .ZN(n17912) );
  OAI22_X1 U21046 ( .A1(n18585), .A2(n17991), .B1(n17956), .B2(n9932), .ZN(
        n18001) );
  AOI211_X1 U21047 ( .C1(n17959), .C2(n17913), .A(n17912), .B(n18001), .ZN(
        n17927) );
  AOI221_X1 U21048 ( .B1(n9622), .B2(n17914), .C1(n17927), .C2(n17914), .A(
        n9611), .ZN(n17916) );
  AOI22_X1 U21049 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17916), .B1(
        n18009), .B2(n17915), .ZN(n17918) );
  OAI211_X1 U21050 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17919), .A(
        n17918), .B(n17917), .ZN(P3_U2846) );
  AOI22_X1 U21051 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18092), .B1(
        n18097), .B2(n17920), .ZN(n17932) );
  AOI21_X1 U21052 ( .B1(n17922), .B2(n17921), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17926) );
  NAND2_X1 U21053 ( .A1(n17976), .A2(n17923), .ZN(n17924) );
  OAI22_X1 U21054 ( .A1(n17927), .A2(n17926), .B1(n17925), .B2(n17924), .ZN(
        n17929) );
  AOI22_X1 U21055 ( .A1(n18101), .A2(n17929), .B1(n18009), .B2(n17928), .ZN(
        n17931) );
  NAND2_X1 U21056 ( .A1(n9611), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17930) );
  OAI211_X1 U21057 ( .C1(n17933), .C2(n17932), .A(n17931), .B(n17930), .ZN(
        P3_U2847) );
  NOR2_X1 U21058 ( .A1(n17988), .A2(n18670), .ZN(n17944) );
  AOI22_X1 U21059 ( .A1(n18581), .A2(n17935), .B1(n18559), .B2(n17934), .ZN(
        n17937) );
  NAND2_X1 U21060 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17991), .ZN(
        n18002) );
  OAI21_X1 U21061 ( .B1(n17936), .B2(n18002), .A(n18583), .ZN(n17957) );
  NAND3_X1 U21062 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17937), .A3(
        n17957), .ZN(n17939) );
  NOR2_X1 U21063 ( .A1(n17938), .A2(n18016), .ZN(n18102) );
  AOI22_X1 U21064 ( .A1(n18101), .A2(n17939), .B1(n18102), .B2(n17960), .ZN(
        n17940) );
  AOI21_X1 U21065 ( .B1(n17942), .B2(n17941), .A(n17940), .ZN(n17943) );
  AOI211_X1 U21066 ( .C1(n18092), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17944), .B(n17943), .ZN(n17948) );
  AOI22_X1 U21067 ( .A1(n18097), .A2(n17946), .B1(n18009), .B2(n17945), .ZN(
        n17947) );
  OAI211_X1 U21068 ( .C1(n18027), .C2(n17949), .A(n17948), .B(n17947), .ZN(
        P3_U2848) );
  INV_X1 U21069 ( .A(n17950), .ZN(n18029) );
  NAND2_X1 U21070 ( .A1(n18101), .A2(n18029), .ZN(n18040) );
  OAI222_X1 U21071 ( .A1(n18040), .A2(n17951), .B1(n18110), .B2(n17977), .C1(
        n17975), .C2(n18027), .ZN(n17996) );
  OAI21_X1 U21072 ( .B1(n18585), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17971) );
  AOI21_X1 U21073 ( .B1(n17952), .B2(n17991), .A(n18585), .ZN(n17953) );
  AOI21_X1 U21074 ( .B1(n18581), .B2(n17968), .A(n17953), .ZN(n17983) );
  AOI22_X1 U21075 ( .A1(n18549), .A2(n17955), .B1(n17976), .B2(n17954), .ZN(
        n17958) );
  OR2_X1 U21076 ( .A1(n17956), .A2(n9932), .ZN(n17979) );
  NAND4_X1 U21077 ( .A1(n17983), .A2(n17958), .A3(n17979), .A4(n17957), .ZN(
        n17970) );
  AOI211_X1 U21078 ( .C1(n17959), .C2(n17971), .A(n18016), .B(n17970), .ZN(
        n17961) );
  NOR3_X1 U21079 ( .A1(n9611), .A2(n17961), .A3(n17960), .ZN(n17962) );
  AOI21_X1 U21080 ( .B1(n17963), .B2(n17996), .A(n17962), .ZN(n17965) );
  OAI211_X1 U21081 ( .C1(n17966), .C2(n18021), .A(n17965), .B(n17964), .ZN(
        P3_U2849) );
  AOI22_X1 U21082 ( .A1(n9611), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n18009), 
        .B2(n17967), .ZN(n17973) );
  INV_X1 U21083 ( .A(n17996), .ZN(n18011) );
  OAI22_X1 U21084 ( .A1(n18011), .A2(n17968), .B1(n17974), .B2(n18016), .ZN(
        n17969) );
  OAI21_X1 U21085 ( .B1(n17971), .B2(n17970), .A(n17969), .ZN(n17972) );
  OAI211_X1 U21086 ( .C1(n18089), .C2(n17974), .A(n17973), .B(n17972), .ZN(
        P3_U2850) );
  AOI22_X1 U21087 ( .A1(n18549), .A2(n17977), .B1(n17976), .B2(n17975), .ZN(
        n18005) );
  INV_X1 U21088 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18003) );
  OAI21_X1 U21089 ( .B1(n18003), .B2(n18002), .A(n18583), .ZN(n17978) );
  NAND4_X1 U21090 ( .A1(n18101), .A2(n18005), .A3(n17979), .A4(n17978), .ZN(
        n17980) );
  AOI21_X1 U21091 ( .B1(n17982), .B2(n17981), .A(n17980), .ZN(n17992) );
  OAI211_X1 U21092 ( .C1(n18572), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17983), .B(n17992), .ZN(n17984) );
  NAND2_X1 U21093 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17984), .ZN(
        n17989) );
  AOI22_X1 U21094 ( .A1(n18009), .A2(n17986), .B1(n17985), .B2(n17996), .ZN(
        n17987) );
  OAI221_X1 U21095 ( .B1(n9611), .B2(n17989), .C1(n17988), .C2(n18663), .A(
        n17987), .ZN(P3_U2851) );
  AOI22_X1 U21096 ( .A1(n9611), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18009), 
        .B2(n17990), .ZN(n18000) );
  NOR2_X1 U21097 ( .A1(n18585), .A2(n17991), .ZN(n17995) );
  OAI21_X1 U21098 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17993), .A(
        n17992), .ZN(n17994) );
  OAI211_X1 U21099 ( .C1(n17995), .C2(n17994), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n17988), .ZN(n17999) );
  NAND3_X1 U21100 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17997), .A3(
        n17996), .ZN(n17998) );
  NAND3_X1 U21101 ( .A1(n18000), .A2(n17999), .A3(n17998), .ZN(P3_U2852) );
  AOI211_X1 U21102 ( .C1(n18583), .C2(n18002), .A(n18092), .B(n18001), .ZN(
        n18004) );
  AOI211_X1 U21103 ( .C1(n18005), .C2(n18004), .A(n9611), .B(n18003), .ZN(
        n18006) );
  AOI211_X1 U21104 ( .C1(n18009), .C2(n18008), .A(n18007), .B(n18006), .ZN(
        n18010) );
  OAI21_X1 U21105 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18011), .A(
        n18010), .ZN(P3_U2853) );
  NAND2_X1 U21106 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18012) );
  NOR3_X1 U21107 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18012), .A3(
        n18040), .ZN(n18025) );
  INV_X1 U21108 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18019) );
  AOI22_X1 U21109 ( .A1(n18581), .A2(n18014), .B1(n18077), .B2(n18013), .ZN(
        n18015) );
  AOI21_X1 U21110 ( .B1(n18015), .B2(n18074), .A(n18016), .ZN(n18038) );
  AOI211_X1 U21111 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n9622), .B(n18016), .ZN(n18017)
         );
  NOR2_X1 U21112 ( .A1(n18038), .A2(n18017), .ZN(n18037) );
  OAI221_X1 U21113 ( .B1(n18019), .B2(n18037), .C1(n18019), .C2(n18089), .A(
        n18018), .ZN(n18024) );
  OAI22_X1 U21114 ( .A1(n18022), .A2(n18021), .B1(n18110), .B2(n18020), .ZN(
        n18023) );
  NOR3_X1 U21115 ( .A1(n18025), .A2(n18024), .A3(n18023), .ZN(n18026) );
  OAI21_X1 U21116 ( .B1(n18028), .B2(n18027), .A(n18026), .ZN(P3_U2854) );
  AOI21_X1 U21117 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18029), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18036) );
  AOI21_X1 U21118 ( .B1(n18092), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18030), .ZN(n18035) );
  INV_X1 U21119 ( .A(n18031), .ZN(n18032) );
  AOI22_X1 U21120 ( .A1(n18097), .A2(n18033), .B1(n18050), .B2(n18032), .ZN(
        n18034) );
  OAI211_X1 U21121 ( .C1(n18037), .C2(n18036), .A(n18035), .B(n18034), .ZN(
        P3_U2855) );
  OR2_X1 U21122 ( .A1(n18092), .A2(n18038), .ZN(n18046) );
  INV_X1 U21123 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18653) );
  NOR2_X1 U21124 ( .A1(n17988), .A2(n18653), .ZN(n18042) );
  OAI22_X1 U21125 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18040), .B1(
        n18039), .B2(n18108), .ZN(n18041) );
  AOI211_X1 U21126 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18046), .A(
        n18042), .B(n18041), .ZN(n18043) );
  OAI21_X1 U21127 ( .B1(n18110), .B2(n18044), .A(n18043), .ZN(P3_U2856) );
  NAND3_X1 U21128 ( .A1(n18101), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18067), .ZN(n18057) );
  NOR2_X1 U21129 ( .A1(n18045), .A2(n18057), .ZN(n18047) );
  MUX2_X1 U21130 ( .A(n18047), .B(n18046), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18048) );
  AOI21_X1 U21131 ( .B1(n18050), .B2(n18049), .A(n18048), .ZN(n18052) );
  NAND2_X1 U21132 ( .A1(n9611), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18051) );
  OAI211_X1 U21133 ( .C1(n18053), .C2(n18110), .A(n18052), .B(n18051), .ZN(
        P3_U2857) );
  OAI211_X1 U21134 ( .C1(n9932), .C2(n18072), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18074), .ZN(n18055) );
  OAI221_X1 U21135 ( .B1(n18055), .B2(n18077), .C1(n18055), .C2(n18054), .A(
        n18101), .ZN(n18063) );
  OAI21_X1 U21136 ( .B1(n9622), .B2(n18063), .A(n18089), .ZN(n18059) );
  OAI22_X1 U21137 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18057), .B1(
        n18056), .B2(n18110), .ZN(n18058) );
  AOI21_X1 U21138 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18059), .A(
        n18058), .ZN(n18061) );
  NAND2_X1 U21139 ( .A1(n9611), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18060) );
  OAI211_X1 U21140 ( .C1(n18062), .C2(n18108), .A(n18061), .B(n18060), .ZN(
        P3_U2858) );
  INV_X1 U21141 ( .A(n18063), .ZN(n18068) );
  OAI22_X1 U21142 ( .A1(n18065), .A2(n18089), .B1(n18110), .B2(n18064), .ZN(
        n18066) );
  AOI221_X1 U21143 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18068), .C1(
        n18067), .C2(n18068), .A(n18066), .ZN(n18070) );
  OAI211_X1 U21144 ( .C1(n18071), .C2(n18108), .A(n18070), .B(n18069), .ZN(
        P3_U2859) );
  NOR2_X1 U21145 ( .A1(n9932), .A2(n18072), .ZN(n18085) );
  NOR2_X1 U21146 ( .A1(n18728), .A2(n18073), .ZN(n18080) );
  NAND2_X1 U21147 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18075) );
  OAI21_X1 U21148 ( .B1(n18075), .B2(n9932), .A(n18074), .ZN(n18076) );
  AOI21_X1 U21149 ( .B1(n18077), .B2(n18728), .A(n18076), .ZN(n18078) );
  INV_X1 U21150 ( .A(n18078), .ZN(n18079) );
  MUX2_X1 U21151 ( .A(n18080), .B(n18079), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18084) );
  OAI22_X1 U21152 ( .A1(n18110), .A2(n18082), .B1(n18108), .B2(n18081), .ZN(
        n18083) );
  AOI221_X1 U21153 ( .B1(n18085), .B2(n18101), .C1(n18084), .C2(n18101), .A(
        n18083), .ZN(n18087) );
  OAI211_X1 U21154 ( .C1(n18089), .C2(n18088), .A(n18087), .B(n18086), .ZN(
        P3_U2860) );
  NOR2_X1 U21155 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18559), .ZN(
        n18091) );
  NOR2_X1 U21156 ( .A1(n18091), .A2(n18090), .ZN(n18094) );
  AOI21_X1 U21157 ( .B1(n18102), .B2(n18725), .A(n18092), .ZN(n18105) );
  INV_X1 U21158 ( .A(n18105), .ZN(n18093) );
  MUX2_X1 U21159 ( .A(n18094), .B(n18093), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n18095) );
  AOI21_X1 U21160 ( .B1(n18097), .B2(n18096), .A(n18095), .ZN(n18099) );
  NAND2_X1 U21161 ( .A1(n9611), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18098) );
  OAI211_X1 U21162 ( .C1(n18100), .C2(n18108), .A(n18099), .B(n18098), .ZN(
        P3_U2861) );
  NAND2_X1 U21163 ( .A1(n18101), .A2(n18559), .ZN(n18104) );
  INV_X1 U21164 ( .A(n18102), .ZN(n18103) );
  AOI22_X1 U21165 ( .A1(n18105), .A2(n18104), .B1(n18725), .B2(n18103), .ZN(
        n18106) );
  AOI21_X1 U21166 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n9611), .A(n18106), .ZN(
        n18107) );
  OAI221_X1 U21167 ( .B1(n18111), .B2(n18110), .C1(n18109), .C2(n18108), .A(
        n18107), .ZN(P3_U2862) );
  AOI21_X1 U21168 ( .B1(n18114), .B2(n18113), .A(n18112), .ZN(n18614) );
  OAI21_X1 U21169 ( .B1(n18614), .B2(n18386), .A(n18119), .ZN(n18115) );
  OAI221_X1 U21170 ( .B1(n18589), .B2(n18770), .C1(n18589), .C2(n18119), .A(
        n18115), .ZN(P3_U2863) );
  INV_X1 U21171 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18599) );
  NAND2_X1 U21172 ( .A1(n18596), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18361) );
  INV_X1 U21173 ( .A(n18361), .ZN(n18387) );
  NAND2_X1 U21174 ( .A1(n18599), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18249) );
  INV_X1 U21175 ( .A(n18249), .ZN(n18297) );
  NOR2_X1 U21176 ( .A1(n18387), .A2(n18297), .ZN(n18117) );
  OAI22_X1 U21177 ( .A1(n18118), .A2(n18599), .B1(n18117), .B2(n18116), .ZN(
        P3_U2866) );
  NOR2_X1 U21178 ( .A1(n18600), .A2(n18119), .ZN(P3_U2867) );
  NOR2_X1 U21179 ( .A1(n18120), .A2(n18456), .ZN(n18489) );
  INV_X1 U21180 ( .A(n18489), .ZN(n18463) );
  NAND2_X1 U21181 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18433) );
  INV_X1 U21182 ( .A(n18433), .ZN(n18435) );
  NOR2_X1 U21183 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18589), .ZN(
        n18340) );
  NAND2_X1 U21184 ( .A1(n18435), .A2(n18340), .ZN(n18516) );
  AND2_X1 U21185 ( .A1(n18410), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18488) );
  NOR2_X1 U21186 ( .A1(n18599), .A2(n18272), .ZN(n18491) );
  NAND2_X1 U21187 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18491), .ZN(
        n18545) );
  NOR2_X1 U21188 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18226) );
  NOR2_X1 U21189 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18205) );
  NAND2_X1 U21190 ( .A1(n18226), .A2(n18205), .ZN(n18214) );
  NAND2_X1 U21191 ( .A1(n18545), .A2(n18214), .ZN(n18121) );
  INV_X1 U21192 ( .A(n18121), .ZN(n18185) );
  NOR2_X1 U21193 ( .A1(n18487), .A2(n18185), .ZN(n18161) );
  INV_X1 U21194 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19100) );
  NOR2_X2 U21195 ( .A1(n18456), .A2(n19100), .ZN(n18494) );
  NAND2_X1 U21196 ( .A1(n18589), .A2(n18491), .ZN(n18485) );
  INV_X1 U21197 ( .A(n18485), .ZN(n18469) );
  AOI22_X1 U21198 ( .A1(n18488), .A2(n18161), .B1(n18494), .B2(n18469), .ZN(
        n18127) );
  AOI21_X1 U21199 ( .B1(n18516), .B2(n18485), .A(n18385), .ZN(n18459) );
  AOI21_X1 U21200 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18385), .ZN(n18122) );
  AOI22_X1 U21201 ( .A1(n18123), .A2(n18459), .B1(n18122), .B2(n18121), .ZN(
        n18163) );
  NAND2_X1 U21202 ( .A1(n18125), .A2(n18159), .ZN(n18497) );
  INV_X1 U21203 ( .A(n18497), .ZN(n18460) );
  INV_X1 U21204 ( .A(n18214), .ZN(n18222) );
  AOI22_X1 U21205 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18163), .B1(
        n18460), .B2(n18222), .ZN(n18126) );
  OAI211_X1 U21206 ( .C1(n18463), .C2(n18516), .A(n18127), .B(n18126), .ZN(
        P3_U2868) );
  NAND2_X1 U21207 ( .A1(n18159), .A2(n18128), .ZN(n18503) );
  AND2_X1 U21208 ( .A1(n18410), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18498) );
  NOR2_X2 U21209 ( .A1(n18129), .A2(n18456), .ZN(n18499) );
  INV_X1 U21210 ( .A(n18516), .ZN(n18540) );
  AOI22_X1 U21211 ( .A1(n18498), .A2(n18161), .B1(n18499), .B2(n18540), .ZN(
        n18131) );
  NOR2_X2 U21212 ( .A1(n18456), .A2(n14757), .ZN(n18500) );
  AOI22_X1 U21213 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18163), .B1(
        n18500), .B2(n18469), .ZN(n18130) );
  OAI211_X1 U21214 ( .C1(n18503), .C2(n18214), .A(n18131), .B(n18130), .ZN(
        P3_U2869) );
  NAND2_X1 U21215 ( .A1(n18159), .A2(n18132), .ZN(n18509) );
  NOR2_X2 U21216 ( .A1(n18133), .A2(n18456), .ZN(n18506) );
  NOR2_X2 U21217 ( .A1(n18385), .A2(n18134), .ZN(n18504) );
  AOI22_X1 U21218 ( .A1(n18506), .A2(n18540), .B1(n18504), .B2(n18161), .ZN(
        n18137) );
  NOR2_X2 U21219 ( .A1(n18456), .A2(n18135), .ZN(n18505) );
  AOI22_X1 U21220 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18163), .B1(
        n18505), .B2(n18469), .ZN(n18136) );
  OAI211_X1 U21221 ( .C1(n18509), .C2(n18214), .A(n18137), .B(n18136), .ZN(
        P3_U2870) );
  NAND2_X1 U21222 ( .A1(n18493), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18517) );
  NOR2_X1 U21223 ( .A1(n18138), .A2(n18456), .ZN(n18511) );
  NOR2_X2 U21224 ( .A1(n18385), .A2(n18139), .ZN(n18510) );
  AOI22_X1 U21225 ( .A1(n18511), .A2(n18540), .B1(n18510), .B2(n18161), .ZN(
        n18142) );
  AND2_X1 U21226 ( .A1(n18140), .A2(n18159), .ZN(n18513) );
  AOI22_X1 U21227 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18163), .B1(
        n18513), .B2(n18222), .ZN(n18141) );
  OAI211_X1 U21228 ( .C1(n18517), .C2(n18485), .A(n18142), .B(n18141), .ZN(
        P3_U2871) );
  NAND2_X1 U21229 ( .A1(n18159), .A2(n18143), .ZN(n18523) );
  NOR2_X2 U21230 ( .A1(n18385), .A2(n18144), .ZN(n18518) );
  AND2_X1 U21231 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18493), .ZN(n18520) );
  AOI22_X1 U21232 ( .A1(n18518), .A2(n18161), .B1(n18520), .B2(n18540), .ZN(
        n18147) );
  NOR2_X2 U21233 ( .A1(n18456), .A2(n18145), .ZN(n18519) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18163), .B1(
        n18519), .B2(n18469), .ZN(n18146) );
  OAI211_X1 U21235 ( .C1(n18523), .C2(n18214), .A(n18147), .B(n18146), .ZN(
        P3_U2872) );
  NAND2_X1 U21236 ( .A1(n18159), .A2(n18148), .ZN(n18529) );
  AND2_X1 U21237 ( .A1(n18493), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18525) );
  NOR2_X2 U21238 ( .A1(n18385), .A2(n18149), .ZN(n18524) );
  AOI22_X1 U21239 ( .A1(n18525), .A2(n18469), .B1(n18524), .B2(n18161), .ZN(
        n18152) );
  NOR2_X2 U21240 ( .A1(n18150), .A2(n18456), .ZN(n18526) );
  AOI22_X1 U21241 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18163), .B1(
        n18526), .B2(n18540), .ZN(n18151) );
  OAI211_X1 U21242 ( .C1(n18529), .C2(n18214), .A(n18152), .B(n18151), .ZN(
        P3_U2873) );
  NAND2_X1 U21243 ( .A1(n18159), .A2(n18153), .ZN(n18535) );
  NOR2_X2 U21244 ( .A1(n19185), .A2(n18456), .ZN(n18532) );
  NOR2_X2 U21245 ( .A1(n18385), .A2(n18154), .ZN(n18530) );
  AOI22_X1 U21246 ( .A1(n18532), .A2(n18540), .B1(n18530), .B2(n18161), .ZN(
        n18157) );
  NOR2_X2 U21247 ( .A1(n18456), .A2(n18155), .ZN(n18531) );
  AOI22_X1 U21248 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18163), .B1(
        n18531), .B2(n18469), .ZN(n18156) );
  OAI211_X1 U21249 ( .C1(n18535), .C2(n18214), .A(n18157), .B(n18156), .ZN(
        P3_U2874) );
  NAND2_X1 U21250 ( .A1(n18159), .A2(n18158), .ZN(n18546) );
  AND2_X1 U21251 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18493), .ZN(n18541) );
  NOR2_X2 U21252 ( .A1(n18160), .A2(n18385), .ZN(n18537) );
  AOI22_X1 U21253 ( .A1(n18541), .A2(n18469), .B1(n18537), .B2(n18161), .ZN(
        n18165) );
  NOR2_X2 U21254 ( .A1(n18456), .A2(n18162), .ZN(n18538) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18163), .B1(
        n18538), .B2(n18540), .ZN(n18164) );
  OAI211_X1 U21256 ( .C1(n18546), .C2(n18214), .A(n18165), .B(n18164), .ZN(
        P3_U2875) );
  NAND2_X1 U21257 ( .A1(n18340), .A2(n18205), .ZN(n18237) );
  INV_X1 U21258 ( .A(n18205), .ZN(n18184) );
  NAND2_X1 U21259 ( .A1(n18591), .A2(n18613), .ZN(n18432) );
  NOR2_X1 U21260 ( .A1(n18184), .A2(n18432), .ZN(n18180) );
  AOI22_X1 U21261 ( .A1(n18489), .A2(n18469), .B1(n18488), .B2(n18180), .ZN(
        n18167) );
  NOR3_X1 U21262 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18386), .A3(
        n18385), .ZN(n18434) );
  AOI22_X1 U21263 ( .A1(n18493), .A2(n18491), .B1(n18205), .B2(n18434), .ZN(
        n18181) );
  INV_X1 U21264 ( .A(n18545), .ZN(n18512) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18181), .B1(
        n18494), .B2(n18512), .ZN(n18166) );
  OAI211_X1 U21266 ( .C1(n18497), .C2(n18237), .A(n18167), .B(n18166), .ZN(
        P3_U2876) );
  AOI22_X1 U21267 ( .A1(n18498), .A2(n18180), .B1(n18499), .B2(n18469), .ZN(
        n18169) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18181), .B1(
        n18500), .B2(n18512), .ZN(n18168) );
  OAI211_X1 U21269 ( .C1(n18503), .C2(n18237), .A(n18169), .B(n18168), .ZN(
        P3_U2877) );
  AOI22_X1 U21270 ( .A1(n18505), .A2(n18512), .B1(n18504), .B2(n18180), .ZN(
        n18171) );
  AOI22_X1 U21271 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18181), .B1(
        n18506), .B2(n18469), .ZN(n18170) );
  OAI211_X1 U21272 ( .C1(n18509), .C2(n18237), .A(n18171), .B(n18170), .ZN(
        P3_U2878) );
  INV_X1 U21273 ( .A(n18511), .ZN(n18472) );
  INV_X1 U21274 ( .A(n18517), .ZN(n18468) );
  AOI22_X1 U21275 ( .A1(n18468), .A2(n18512), .B1(n18510), .B2(n18180), .ZN(
        n18173) );
  INV_X1 U21276 ( .A(n18237), .ZN(n18244) );
  AOI22_X1 U21277 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18181), .B1(
        n18513), .B2(n18244), .ZN(n18172) );
  OAI211_X1 U21278 ( .C1(n18472), .C2(n18485), .A(n18173), .B(n18172), .ZN(
        P3_U2879) );
  AOI22_X1 U21279 ( .A1(n18519), .A2(n18512), .B1(n18518), .B2(n18180), .ZN(
        n18175) );
  AOI22_X1 U21280 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18181), .B1(
        n18520), .B2(n18469), .ZN(n18174) );
  OAI211_X1 U21281 ( .C1(n18523), .C2(n18237), .A(n18175), .B(n18174), .ZN(
        P3_U2880) );
  AOI22_X1 U21282 ( .A1(n18525), .A2(n18512), .B1(n18524), .B2(n18180), .ZN(
        n18177) );
  AOI22_X1 U21283 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18181), .B1(
        n18526), .B2(n18469), .ZN(n18176) );
  OAI211_X1 U21284 ( .C1(n18529), .C2(n18237), .A(n18177), .B(n18176), .ZN(
        P3_U2881) );
  AOI22_X1 U21285 ( .A1(n18532), .A2(n18469), .B1(n18530), .B2(n18180), .ZN(
        n18179) );
  AOI22_X1 U21286 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18181), .B1(
        n18531), .B2(n18512), .ZN(n18178) );
  OAI211_X1 U21287 ( .C1(n18535), .C2(n18237), .A(n18179), .B(n18178), .ZN(
        P3_U2882) );
  AOI22_X1 U21288 ( .A1(n18541), .A2(n18512), .B1(n18537), .B2(n18180), .ZN(
        n18183) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18181), .B1(
        n18538), .B2(n18469), .ZN(n18182) );
  OAI211_X1 U21290 ( .C1(n18546), .C2(n18237), .A(n18183), .B(n18182), .ZN(
        P3_U2883) );
  NOR2_X1 U21291 ( .A1(n18591), .A2(n18184), .ZN(n18250) );
  NAND2_X1 U21292 ( .A1(n18250), .A2(n18589), .ZN(n18259) );
  NOR2_X1 U21293 ( .A1(n18244), .A2(n18267), .ZN(n18227) );
  NOR2_X1 U21294 ( .A1(n18487), .A2(n18227), .ZN(n18201) );
  AOI22_X1 U21295 ( .A1(n18489), .A2(n18512), .B1(n18488), .B2(n18201), .ZN(
        n18188) );
  OAI21_X1 U21296 ( .B1(n18185), .B2(n18408), .A(n18227), .ZN(n18186) );
  OAI211_X1 U21297 ( .C1(n18267), .C2(n18743), .A(n18410), .B(n18186), .ZN(
        n18202) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18202), .B1(
        n18494), .B2(n18222), .ZN(n18187) );
  OAI211_X1 U21299 ( .C1(n18497), .C2(n18259), .A(n18188), .B(n18187), .ZN(
        P3_U2884) );
  AOI22_X1 U21300 ( .A1(n18500), .A2(n18222), .B1(n18498), .B2(n18201), .ZN(
        n18190) );
  AOI22_X1 U21301 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18202), .B1(
        n18499), .B2(n18512), .ZN(n18189) );
  OAI211_X1 U21302 ( .C1(n18503), .C2(n18259), .A(n18190), .B(n18189), .ZN(
        P3_U2885) );
  AOI22_X1 U21303 ( .A1(n18506), .A2(n18512), .B1(n18504), .B2(n18201), .ZN(
        n18192) );
  AOI22_X1 U21304 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18202), .B1(
        n18505), .B2(n18222), .ZN(n18191) );
  OAI211_X1 U21305 ( .C1(n18509), .C2(n18259), .A(n18192), .B(n18191), .ZN(
        P3_U2886) );
  AOI22_X1 U21306 ( .A1(n18511), .A2(n18512), .B1(n18510), .B2(n18201), .ZN(
        n18194) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18202), .B1(
        n18513), .B2(n18267), .ZN(n18193) );
  OAI211_X1 U21308 ( .C1(n18517), .C2(n18214), .A(n18194), .B(n18193), .ZN(
        P3_U2887) );
  AOI22_X1 U21309 ( .A1(n18518), .A2(n18201), .B1(n18520), .B2(n18512), .ZN(
        n18196) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18202), .B1(
        n18519), .B2(n18222), .ZN(n18195) );
  OAI211_X1 U21311 ( .C1(n18523), .C2(n18259), .A(n18196), .B(n18195), .ZN(
        P3_U2888) );
  AOI22_X1 U21312 ( .A1(n18525), .A2(n18222), .B1(n18524), .B2(n18201), .ZN(
        n18198) );
  AOI22_X1 U21313 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18202), .B1(
        n18526), .B2(n18512), .ZN(n18197) );
  OAI211_X1 U21314 ( .C1(n18529), .C2(n18259), .A(n18198), .B(n18197), .ZN(
        P3_U2889) );
  AOI22_X1 U21315 ( .A1(n18532), .A2(n18512), .B1(n18530), .B2(n18201), .ZN(
        n18200) );
  AOI22_X1 U21316 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18202), .B1(
        n18531), .B2(n18222), .ZN(n18199) );
  OAI211_X1 U21317 ( .C1(n18535), .C2(n18259), .A(n18200), .B(n18199), .ZN(
        P3_U2890) );
  AOI22_X1 U21318 ( .A1(n18541), .A2(n18222), .B1(n18537), .B2(n18201), .ZN(
        n18204) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18202), .B1(
        n18538), .B2(n18512), .ZN(n18203) );
  OAI211_X1 U21320 ( .C1(n18546), .C2(n18259), .A(n18204), .B(n18203), .ZN(
        P3_U2891) );
  NAND2_X1 U21321 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18250), .ZN(
        n18277) );
  AOI21_X1 U21322 ( .B1(n18591), .B2(n18408), .A(n18385), .ZN(n18296) );
  OAI211_X1 U21323 ( .C1(n18291), .C2(n18743), .A(n18205), .B(n18296), .ZN(
        n18223) );
  AND2_X1 U21324 ( .A1(n18613), .A2(n18250), .ZN(n18221) );
  AOI22_X1 U21325 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18223), .B1(
        n18488), .B2(n18221), .ZN(n18207) );
  AOI22_X1 U21326 ( .A1(n18489), .A2(n18222), .B1(n18494), .B2(n18244), .ZN(
        n18206) );
  OAI211_X1 U21327 ( .C1(n18497), .C2(n18277), .A(n18207), .B(n18206), .ZN(
        P3_U2892) );
  AOI22_X1 U21328 ( .A1(n18498), .A2(n18221), .B1(n18499), .B2(n18222), .ZN(
        n18209) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18223), .B1(
        n18500), .B2(n18244), .ZN(n18208) );
  OAI211_X1 U21330 ( .C1(n18503), .C2(n18277), .A(n18209), .B(n18208), .ZN(
        P3_U2893) );
  AOI22_X1 U21331 ( .A1(n18505), .A2(n18244), .B1(n18504), .B2(n18221), .ZN(
        n18211) );
  AOI22_X1 U21332 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18223), .B1(
        n18506), .B2(n18222), .ZN(n18210) );
  OAI211_X1 U21333 ( .C1(n18509), .C2(n18277), .A(n18211), .B(n18210), .ZN(
        P3_U2894) );
  AOI22_X1 U21334 ( .A1(n18468), .A2(n18244), .B1(n18510), .B2(n18221), .ZN(
        n18213) );
  AOI22_X1 U21335 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18223), .B1(
        n18513), .B2(n18291), .ZN(n18212) );
  OAI211_X1 U21336 ( .C1(n18472), .C2(n18214), .A(n18213), .B(n18212), .ZN(
        P3_U2895) );
  AOI22_X1 U21337 ( .A1(n18518), .A2(n18221), .B1(n18520), .B2(n18222), .ZN(
        n18216) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18223), .B1(
        n18519), .B2(n18244), .ZN(n18215) );
  OAI211_X1 U21339 ( .C1(n18523), .C2(n18277), .A(n18216), .B(n18215), .ZN(
        P3_U2896) );
  AOI22_X1 U21340 ( .A1(n18525), .A2(n18244), .B1(n18524), .B2(n18221), .ZN(
        n18218) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18223), .B1(
        n18526), .B2(n18222), .ZN(n18217) );
  OAI211_X1 U21342 ( .C1(n18529), .C2(n18277), .A(n18218), .B(n18217), .ZN(
        P3_U2897) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18223), .B1(
        n18530), .B2(n18221), .ZN(n18220) );
  AOI22_X1 U21344 ( .A1(n18531), .A2(n18244), .B1(n18532), .B2(n18222), .ZN(
        n18219) );
  OAI211_X1 U21345 ( .C1(n18535), .C2(n18277), .A(n18220), .B(n18219), .ZN(
        P3_U2898) );
  AOI22_X1 U21346 ( .A1(n18541), .A2(n18244), .B1(n18537), .B2(n18221), .ZN(
        n18225) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18223), .B1(
        n18538), .B2(n18222), .ZN(n18224) );
  OAI211_X1 U21348 ( .C1(n18546), .C2(n18277), .A(n18225), .B(n18224), .ZN(
        P3_U2899) );
  INV_X1 U21349 ( .A(n18226), .ZN(n18592) );
  NOR2_X2 U21350 ( .A1(n18592), .A2(n18249), .ZN(n18314) );
  INV_X1 U21351 ( .A(n18314), .ZN(n18306) );
  NOR2_X1 U21352 ( .A1(n18291), .A2(n18314), .ZN(n18273) );
  NOR2_X1 U21353 ( .A1(n18487), .A2(n18273), .ZN(n18245) );
  AOI22_X1 U21354 ( .A1(n18489), .A2(n18244), .B1(n18488), .B2(n18245), .ZN(
        n18230) );
  OAI21_X1 U21355 ( .B1(n18227), .B2(n18408), .A(n18273), .ZN(n18228) );
  OAI211_X1 U21356 ( .C1(n18314), .C2(n18743), .A(n18410), .B(n18228), .ZN(
        n18246) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18246), .B1(
        n18494), .B2(n18267), .ZN(n18229) );
  OAI211_X1 U21358 ( .C1(n18497), .C2(n18306), .A(n18230), .B(n18229), .ZN(
        P3_U2900) );
  AOI22_X1 U21359 ( .A1(n18500), .A2(n18267), .B1(n18498), .B2(n18245), .ZN(
        n18232) );
  AOI22_X1 U21360 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18246), .B1(
        n18499), .B2(n18244), .ZN(n18231) );
  OAI211_X1 U21361 ( .C1(n18503), .C2(n18306), .A(n18232), .B(n18231), .ZN(
        P3_U2901) );
  AOI22_X1 U21362 ( .A1(n18505), .A2(n18267), .B1(n18504), .B2(n18245), .ZN(
        n18234) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18246), .B1(
        n18506), .B2(n18244), .ZN(n18233) );
  OAI211_X1 U21364 ( .C1(n18509), .C2(n18306), .A(n18234), .B(n18233), .ZN(
        P3_U2902) );
  AOI22_X1 U21365 ( .A1(n18468), .A2(n18267), .B1(n18510), .B2(n18245), .ZN(
        n18236) );
  AOI22_X1 U21366 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18246), .B1(
        n18513), .B2(n18314), .ZN(n18235) );
  OAI211_X1 U21367 ( .C1(n18472), .C2(n18237), .A(n18236), .B(n18235), .ZN(
        P3_U2903) );
  AOI22_X1 U21368 ( .A1(n18518), .A2(n18245), .B1(n18520), .B2(n18244), .ZN(
        n18239) );
  AOI22_X1 U21369 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18246), .B1(
        n18519), .B2(n18267), .ZN(n18238) );
  OAI211_X1 U21370 ( .C1(n18523), .C2(n18306), .A(n18239), .B(n18238), .ZN(
        P3_U2904) );
  AOI22_X1 U21371 ( .A1(n18524), .A2(n18245), .B1(n18526), .B2(n18244), .ZN(
        n18241) );
  AOI22_X1 U21372 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18246), .B1(
        n18525), .B2(n18267), .ZN(n18240) );
  OAI211_X1 U21373 ( .C1(n18529), .C2(n18306), .A(n18241), .B(n18240), .ZN(
        P3_U2905) );
  AOI22_X1 U21374 ( .A1(n18531), .A2(n18267), .B1(n18530), .B2(n18245), .ZN(
        n18243) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18246), .B1(
        n18532), .B2(n18244), .ZN(n18242) );
  OAI211_X1 U21376 ( .C1(n18535), .C2(n18306), .A(n18243), .B(n18242), .ZN(
        P3_U2906) );
  AOI22_X1 U21377 ( .A1(n18537), .A2(n18245), .B1(n18538), .B2(n18244), .ZN(
        n18248) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18246), .B1(
        n18541), .B2(n18267), .ZN(n18247) );
  OAI211_X1 U21379 ( .C1(n18546), .C2(n18306), .A(n18248), .B(n18247), .ZN(
        P3_U2907) );
  NAND2_X1 U21380 ( .A1(n18297), .A2(n18340), .ZN(n18271) );
  NOR2_X1 U21381 ( .A1(n18249), .A2(n18432), .ZN(n18266) );
  AOI22_X1 U21382 ( .A1(n18489), .A2(n18267), .B1(n18488), .B2(n18266), .ZN(
        n18252) );
  AOI22_X1 U21383 ( .A1(n18493), .A2(n18250), .B1(n18297), .B2(n18434), .ZN(
        n18268) );
  AOI22_X1 U21384 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18268), .B1(
        n18494), .B2(n18291), .ZN(n18251) );
  OAI211_X1 U21385 ( .C1(n18497), .C2(n18271), .A(n18252), .B(n18251), .ZN(
        P3_U2908) );
  AOI22_X1 U21386 ( .A1(n18498), .A2(n18266), .B1(n18499), .B2(n18267), .ZN(
        n18254) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18268), .B1(
        n18500), .B2(n18291), .ZN(n18253) );
  OAI211_X1 U21388 ( .C1(n18503), .C2(n18271), .A(n18254), .B(n18253), .ZN(
        P3_U2909) );
  AOI22_X1 U21389 ( .A1(n18506), .A2(n18267), .B1(n18504), .B2(n18266), .ZN(
        n18256) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18268), .B1(
        n18505), .B2(n18291), .ZN(n18255) );
  OAI211_X1 U21391 ( .C1(n18509), .C2(n18271), .A(n18256), .B(n18255), .ZN(
        P3_U2910) );
  AOI22_X1 U21392 ( .A1(n18468), .A2(n18291), .B1(n18510), .B2(n18266), .ZN(
        n18258) );
  INV_X1 U21393 ( .A(n18271), .ZN(n18335) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18268), .B1(
        n18513), .B2(n18335), .ZN(n18257) );
  OAI211_X1 U21395 ( .C1(n18472), .C2(n18259), .A(n18258), .B(n18257), .ZN(
        P3_U2911) );
  AOI22_X1 U21396 ( .A1(n18518), .A2(n18266), .B1(n18520), .B2(n18267), .ZN(
        n18261) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18268), .B1(
        n18519), .B2(n18291), .ZN(n18260) );
  OAI211_X1 U21398 ( .C1(n18523), .C2(n18271), .A(n18261), .B(n18260), .ZN(
        P3_U2912) );
  AOI22_X1 U21399 ( .A1(n18524), .A2(n18266), .B1(n18526), .B2(n18267), .ZN(
        n18263) );
  AOI22_X1 U21400 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18268), .B1(
        n18525), .B2(n18291), .ZN(n18262) );
  OAI211_X1 U21401 ( .C1(n18529), .C2(n18271), .A(n18263), .B(n18262), .ZN(
        P3_U2913) );
  AOI22_X1 U21402 ( .A1(n18532), .A2(n18267), .B1(n18530), .B2(n18266), .ZN(
        n18265) );
  AOI22_X1 U21403 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18268), .B1(
        n18531), .B2(n18291), .ZN(n18264) );
  OAI211_X1 U21404 ( .C1(n18535), .C2(n18271), .A(n18265), .B(n18264), .ZN(
        P3_U2914) );
  AOI22_X1 U21405 ( .A1(n18541), .A2(n18291), .B1(n18537), .B2(n18266), .ZN(
        n18270) );
  AOI22_X1 U21406 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18268), .B1(
        n18538), .B2(n18267), .ZN(n18269) );
  OAI211_X1 U21407 ( .C1(n18546), .C2(n18271), .A(n18270), .B(n18269), .ZN(
        P3_U2915) );
  NOR2_X1 U21408 ( .A1(n18272), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18339) );
  NAND2_X1 U21409 ( .A1(n18589), .A2(n18339), .ZN(n18343) );
  INV_X1 U21410 ( .A(n18343), .ZN(n18357) );
  NOR2_X1 U21411 ( .A1(n18335), .A2(n18357), .ZN(n18318) );
  NOR2_X1 U21412 ( .A1(n18487), .A2(n18318), .ZN(n18290) );
  AOI22_X1 U21413 ( .A1(n18488), .A2(n18290), .B1(n18494), .B2(n18314), .ZN(
        n18276) );
  OAI22_X1 U21414 ( .A1(n18273), .A2(n18456), .B1(n18318), .B2(n18385), .ZN(
        n18274) );
  OAI21_X1 U21415 ( .B1(n18357), .B2(n18743), .A(n18274), .ZN(n18292) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18292), .B1(
        n18460), .B2(n18357), .ZN(n18275) );
  OAI211_X1 U21417 ( .C1(n18463), .C2(n18277), .A(n18276), .B(n18275), .ZN(
        P3_U2916) );
  AOI22_X1 U21418 ( .A1(n18498), .A2(n18290), .B1(n18499), .B2(n18291), .ZN(
        n18279) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18292), .B1(
        n18500), .B2(n18314), .ZN(n18278) );
  OAI211_X1 U21420 ( .C1(n18503), .C2(n18343), .A(n18279), .B(n18278), .ZN(
        P3_U2917) );
  AOI22_X1 U21421 ( .A1(n18506), .A2(n18291), .B1(n18504), .B2(n18290), .ZN(
        n18281) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18292), .B1(
        n18505), .B2(n18314), .ZN(n18280) );
  OAI211_X1 U21423 ( .C1(n18509), .C2(n18343), .A(n18281), .B(n18280), .ZN(
        P3_U2918) );
  AOI22_X1 U21424 ( .A1(n18511), .A2(n18291), .B1(n18510), .B2(n18290), .ZN(
        n18283) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18292), .B1(
        n18513), .B2(n18357), .ZN(n18282) );
  OAI211_X1 U21426 ( .C1(n18517), .C2(n18306), .A(n18283), .B(n18282), .ZN(
        P3_U2919) );
  AOI22_X1 U21427 ( .A1(n18519), .A2(n18314), .B1(n18518), .B2(n18290), .ZN(
        n18285) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18292), .B1(
        n18520), .B2(n18291), .ZN(n18284) );
  OAI211_X1 U21429 ( .C1(n18523), .C2(n18343), .A(n18285), .B(n18284), .ZN(
        P3_U2920) );
  AOI22_X1 U21430 ( .A1(n18524), .A2(n18290), .B1(n18526), .B2(n18291), .ZN(
        n18287) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18292), .B1(
        n18525), .B2(n18314), .ZN(n18286) );
  OAI211_X1 U21432 ( .C1(n18529), .C2(n18343), .A(n18287), .B(n18286), .ZN(
        P3_U2921) );
  AOI22_X1 U21433 ( .A1(n18532), .A2(n18291), .B1(n18530), .B2(n18290), .ZN(
        n18289) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18292), .B1(
        n18531), .B2(n18314), .ZN(n18288) );
  OAI211_X1 U21435 ( .C1(n18535), .C2(n18343), .A(n18289), .B(n18288), .ZN(
        P3_U2922) );
  AOI22_X1 U21436 ( .A1(n18541), .A2(n18314), .B1(n18537), .B2(n18290), .ZN(
        n18294) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18292), .B1(
        n18538), .B2(n18291), .ZN(n18293) );
  OAI211_X1 U21438 ( .C1(n18546), .C2(n18343), .A(n18294), .B(n18293), .ZN(
        P3_U2923) );
  INV_X1 U21439 ( .A(n18339), .ZN(n18295) );
  NOR2_X2 U21440 ( .A1(n18589), .A2(n18295), .ZN(n18379) );
  INV_X1 U21441 ( .A(n18379), .ZN(n18372) );
  NOR2_X1 U21442 ( .A1(n18487), .A2(n18295), .ZN(n18313) );
  AOI22_X1 U21443 ( .A1(n18489), .A2(n18314), .B1(n18488), .B2(n18313), .ZN(
        n18299) );
  OAI211_X1 U21444 ( .C1(n18379), .C2(n18743), .A(n18297), .B(n18296), .ZN(
        n18315) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18315), .B1(
        n18494), .B2(n18335), .ZN(n18298) );
  OAI211_X1 U21446 ( .C1(n18497), .C2(n18372), .A(n18299), .B(n18298), .ZN(
        P3_U2924) );
  AOI22_X1 U21447 ( .A1(n18500), .A2(n18335), .B1(n18498), .B2(n18313), .ZN(
        n18301) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18315), .B1(
        n18499), .B2(n18314), .ZN(n18300) );
  OAI211_X1 U21449 ( .C1(n18503), .C2(n18372), .A(n18301), .B(n18300), .ZN(
        P3_U2925) );
  AOI22_X1 U21450 ( .A1(n18505), .A2(n18335), .B1(n18504), .B2(n18313), .ZN(
        n18303) );
  AOI22_X1 U21451 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18315), .B1(
        n18506), .B2(n18314), .ZN(n18302) );
  OAI211_X1 U21452 ( .C1(n18509), .C2(n18372), .A(n18303), .B(n18302), .ZN(
        P3_U2926) );
  AOI22_X1 U21453 ( .A1(n18468), .A2(n18335), .B1(n18510), .B2(n18313), .ZN(
        n18305) );
  AOI22_X1 U21454 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18315), .B1(
        n18513), .B2(n18379), .ZN(n18304) );
  OAI211_X1 U21455 ( .C1(n18472), .C2(n18306), .A(n18305), .B(n18304), .ZN(
        P3_U2927) );
  AOI22_X1 U21456 ( .A1(n18519), .A2(n18335), .B1(n18518), .B2(n18313), .ZN(
        n18308) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18315), .B1(
        n18520), .B2(n18314), .ZN(n18307) );
  OAI211_X1 U21458 ( .C1(n18523), .C2(n18372), .A(n18308), .B(n18307), .ZN(
        P3_U2928) );
  AOI22_X1 U21459 ( .A1(n18524), .A2(n18313), .B1(n18526), .B2(n18314), .ZN(
        n18310) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18315), .B1(
        n18525), .B2(n18335), .ZN(n18309) );
  OAI211_X1 U21461 ( .C1(n18529), .C2(n18372), .A(n18310), .B(n18309), .ZN(
        P3_U2929) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18315), .B1(
        n18530), .B2(n18313), .ZN(n18312) );
  AOI22_X1 U21463 ( .A1(n18531), .A2(n18335), .B1(n18532), .B2(n18314), .ZN(
        n18311) );
  OAI211_X1 U21464 ( .C1(n18535), .C2(n18372), .A(n18312), .B(n18311), .ZN(
        P3_U2930) );
  AOI22_X1 U21465 ( .A1(n18541), .A2(n18335), .B1(n18537), .B2(n18313), .ZN(
        n18317) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18315), .B1(
        n18538), .B2(n18314), .ZN(n18316) );
  OAI211_X1 U21467 ( .C1(n18546), .C2(n18372), .A(n18317), .B(n18316), .ZN(
        P3_U2931) );
  NOR2_X2 U21468 ( .A1(n18592), .A2(n18361), .ZN(n18403) );
  INV_X1 U21469 ( .A(n18403), .ZN(n18396) );
  NOR2_X1 U21470 ( .A1(n18379), .A2(n18403), .ZN(n18362) );
  NOR2_X1 U21471 ( .A1(n18487), .A2(n18362), .ZN(n18334) );
  AOI22_X1 U21472 ( .A1(n18488), .A2(n18334), .B1(n18494), .B2(n18357), .ZN(
        n18321) );
  OAI21_X1 U21473 ( .B1(n18318), .B2(n18408), .A(n18362), .ZN(n18319) );
  OAI211_X1 U21474 ( .C1(n18403), .C2(n18743), .A(n18410), .B(n18319), .ZN(
        n18336) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18336), .B1(
        n18489), .B2(n18335), .ZN(n18320) );
  OAI211_X1 U21476 ( .C1(n18497), .C2(n18396), .A(n18321), .B(n18320), .ZN(
        P3_U2932) );
  AOI22_X1 U21477 ( .A1(n18500), .A2(n18357), .B1(n18498), .B2(n18334), .ZN(
        n18323) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18336), .B1(
        n18499), .B2(n18335), .ZN(n18322) );
  OAI211_X1 U21479 ( .C1(n18503), .C2(n18396), .A(n18323), .B(n18322), .ZN(
        P3_U2933) );
  AOI22_X1 U21480 ( .A1(n18505), .A2(n18357), .B1(n18504), .B2(n18334), .ZN(
        n18325) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18336), .B1(
        n18506), .B2(n18335), .ZN(n18324) );
  OAI211_X1 U21482 ( .C1(n18509), .C2(n18396), .A(n18325), .B(n18324), .ZN(
        P3_U2934) );
  AOI22_X1 U21483 ( .A1(n18511), .A2(n18335), .B1(n18510), .B2(n18334), .ZN(
        n18327) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18336), .B1(
        n18513), .B2(n18403), .ZN(n18326) );
  OAI211_X1 U21485 ( .C1(n18517), .C2(n18343), .A(n18327), .B(n18326), .ZN(
        P3_U2935) );
  AOI22_X1 U21486 ( .A1(n18518), .A2(n18334), .B1(n18520), .B2(n18335), .ZN(
        n18329) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18336), .B1(
        n18519), .B2(n18357), .ZN(n18328) );
  OAI211_X1 U21488 ( .C1(n18523), .C2(n18396), .A(n18329), .B(n18328), .ZN(
        P3_U2936) );
  AOI22_X1 U21489 ( .A1(n18524), .A2(n18334), .B1(n18526), .B2(n18335), .ZN(
        n18331) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18336), .B1(
        n18525), .B2(n18357), .ZN(n18330) );
  OAI211_X1 U21491 ( .C1(n18529), .C2(n18396), .A(n18331), .B(n18330), .ZN(
        P3_U2937) );
  AOI22_X1 U21492 ( .A1(n18531), .A2(n18357), .B1(n18530), .B2(n18334), .ZN(
        n18333) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18336), .B1(
        n18532), .B2(n18335), .ZN(n18332) );
  OAI211_X1 U21494 ( .C1(n18535), .C2(n18396), .A(n18333), .B(n18332), .ZN(
        P3_U2938) );
  AOI22_X1 U21495 ( .A1(n18541), .A2(n18357), .B1(n18537), .B2(n18334), .ZN(
        n18338) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18336), .B1(
        n18538), .B2(n18335), .ZN(n18337) );
  OAI211_X1 U21497 ( .C1(n18546), .C2(n18396), .A(n18338), .B(n18337), .ZN(
        P3_U2939) );
  NOR2_X1 U21498 ( .A1(n18361), .A2(n18432), .ZN(n18356) );
  AOI22_X1 U21499 ( .A1(n18488), .A2(n18356), .B1(n18494), .B2(n18379), .ZN(
        n18342) );
  AOI22_X1 U21500 ( .A1(n18493), .A2(n18339), .B1(n18387), .B2(n18434), .ZN(
        n18358) );
  NAND2_X1 U21501 ( .A1(n18387), .A2(n18340), .ZN(n18420) );
  INV_X1 U21502 ( .A(n18420), .ZN(n18428) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18358), .B1(
        n18428), .B2(n18460), .ZN(n18341) );
  OAI211_X1 U21504 ( .C1(n18463), .C2(n18343), .A(n18342), .B(n18341), .ZN(
        P3_U2940) );
  AOI22_X1 U21505 ( .A1(n18500), .A2(n18379), .B1(n18498), .B2(n18356), .ZN(
        n18345) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18358), .B1(
        n18499), .B2(n18357), .ZN(n18344) );
  OAI211_X1 U21507 ( .C1(n18420), .C2(n18503), .A(n18345), .B(n18344), .ZN(
        P3_U2941) );
  AOI22_X1 U21508 ( .A1(n18506), .A2(n18357), .B1(n18504), .B2(n18356), .ZN(
        n18347) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18358), .B1(
        n18505), .B2(n18379), .ZN(n18346) );
  OAI211_X1 U21510 ( .C1(n18420), .C2(n18509), .A(n18347), .B(n18346), .ZN(
        P3_U2942) );
  AOI22_X1 U21511 ( .A1(n18511), .A2(n18357), .B1(n18510), .B2(n18356), .ZN(
        n18349) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18358), .B1(
        n18428), .B2(n18513), .ZN(n18348) );
  OAI211_X1 U21513 ( .C1(n18517), .C2(n18372), .A(n18349), .B(n18348), .ZN(
        P3_U2943) );
  AOI22_X1 U21514 ( .A1(n18518), .A2(n18356), .B1(n18520), .B2(n18357), .ZN(
        n18351) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18358), .B1(
        n18519), .B2(n18379), .ZN(n18350) );
  OAI211_X1 U21516 ( .C1(n18420), .C2(n18523), .A(n18351), .B(n18350), .ZN(
        P3_U2944) );
  AOI22_X1 U21517 ( .A1(n18525), .A2(n18379), .B1(n18524), .B2(n18356), .ZN(
        n18353) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18358), .B1(
        n18526), .B2(n18357), .ZN(n18352) );
  OAI211_X1 U21519 ( .C1(n18420), .C2(n18529), .A(n18353), .B(n18352), .ZN(
        P3_U2945) );
  AOI22_X1 U21520 ( .A1(n18531), .A2(n18379), .B1(n18530), .B2(n18356), .ZN(
        n18355) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18358), .B1(
        n18532), .B2(n18357), .ZN(n18354) );
  OAI211_X1 U21522 ( .C1(n18420), .C2(n18535), .A(n18355), .B(n18354), .ZN(
        P3_U2946) );
  AOI22_X1 U21523 ( .A1(n18541), .A2(n18379), .B1(n18537), .B2(n18356), .ZN(
        n18360) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18358), .B1(
        n18538), .B2(n18357), .ZN(n18359) );
  OAI211_X1 U21525 ( .C1(n18420), .C2(n18546), .A(n18360), .B(n18359), .ZN(
        P3_U2947) );
  NOR2_X1 U21526 ( .A1(n18591), .A2(n18361), .ZN(n18436) );
  NAND2_X1 U21527 ( .A1(n18589), .A2(n18436), .ZN(n18445) );
  NOR2_X1 U21528 ( .A1(n18452), .A2(n18428), .ZN(n18409) );
  NOR2_X1 U21529 ( .A1(n18487), .A2(n18409), .ZN(n18380) );
  AOI22_X1 U21530 ( .A1(n18488), .A2(n18380), .B1(n18494), .B2(n18403), .ZN(
        n18365) );
  OAI21_X1 U21531 ( .B1(n18362), .B2(n18408), .A(n18409), .ZN(n18363) );
  OAI211_X1 U21532 ( .C1(n18452), .C2(n18743), .A(n18410), .B(n18363), .ZN(
        n18381) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18381), .B1(
        n18452), .B2(n18460), .ZN(n18364) );
  OAI211_X1 U21534 ( .C1(n18463), .C2(n18372), .A(n18365), .B(n18364), .ZN(
        P3_U2948) );
  AOI22_X1 U21535 ( .A1(n18500), .A2(n18403), .B1(n18498), .B2(n18380), .ZN(
        n18367) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18381), .B1(
        n18499), .B2(n18379), .ZN(n18366) );
  OAI211_X1 U21537 ( .C1(n18445), .C2(n18503), .A(n18367), .B(n18366), .ZN(
        P3_U2949) );
  AOI22_X1 U21538 ( .A1(n18506), .A2(n18379), .B1(n18504), .B2(n18380), .ZN(
        n18369) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18381), .B1(
        n18505), .B2(n18403), .ZN(n18368) );
  OAI211_X1 U21540 ( .C1(n18445), .C2(n18509), .A(n18369), .B(n18368), .ZN(
        P3_U2950) );
  AOI22_X1 U21541 ( .A1(n18468), .A2(n18403), .B1(n18510), .B2(n18380), .ZN(
        n18371) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18381), .B1(
        n18452), .B2(n18513), .ZN(n18370) );
  OAI211_X1 U21543 ( .C1(n18472), .C2(n18372), .A(n18371), .B(n18370), .ZN(
        P3_U2951) );
  AOI22_X1 U21544 ( .A1(n18518), .A2(n18380), .B1(n18520), .B2(n18379), .ZN(
        n18374) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18381), .B1(
        n18519), .B2(n18403), .ZN(n18373) );
  OAI211_X1 U21546 ( .C1(n18445), .C2(n18523), .A(n18374), .B(n18373), .ZN(
        P3_U2952) );
  AOI22_X1 U21547 ( .A1(n18525), .A2(n18403), .B1(n18524), .B2(n18380), .ZN(
        n18376) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18381), .B1(
        n18526), .B2(n18379), .ZN(n18375) );
  OAI211_X1 U21549 ( .C1(n18445), .C2(n18529), .A(n18376), .B(n18375), .ZN(
        P3_U2953) );
  AOI22_X1 U21550 ( .A1(n18532), .A2(n18379), .B1(n18530), .B2(n18380), .ZN(
        n18378) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18381), .B1(
        n18531), .B2(n18403), .ZN(n18377) );
  OAI211_X1 U21552 ( .C1(n18445), .C2(n18535), .A(n18378), .B(n18377), .ZN(
        P3_U2954) );
  AOI22_X1 U21553 ( .A1(n18537), .A2(n18380), .B1(n18538), .B2(n18379), .ZN(
        n18383) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18381), .B1(
        n18541), .B2(n18403), .ZN(n18382) );
  OAI211_X1 U21555 ( .C1(n18445), .C2(n18546), .A(n18383), .B(n18382), .ZN(
        P3_U2955) );
  INV_X1 U21556 ( .A(n18436), .ZN(n18384) );
  NOR2_X2 U21557 ( .A1(n18589), .A2(n18384), .ZN(n18481) );
  NOR2_X1 U21558 ( .A1(n18487), .A2(n18384), .ZN(n18404) );
  AOI22_X1 U21559 ( .A1(n18489), .A2(n18403), .B1(n18488), .B2(n18404), .ZN(
        n18389) );
  NOR2_X1 U21560 ( .A1(n18386), .A2(n18385), .ZN(n18490) );
  AOI22_X1 U21561 ( .A1(n18493), .A2(n18387), .B1(n18436), .B2(n18490), .ZN(
        n18405) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18405), .B1(
        n18428), .B2(n18494), .ZN(n18388) );
  OAI211_X1 U21563 ( .C1(n18473), .C2(n18497), .A(n18389), .B(n18388), .ZN(
        P3_U2956) );
  AOI22_X1 U21564 ( .A1(n18498), .A2(n18404), .B1(n18499), .B2(n18403), .ZN(
        n18391) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18405), .B1(
        n18428), .B2(n18500), .ZN(n18390) );
  OAI211_X1 U21566 ( .C1(n18473), .C2(n18503), .A(n18391), .B(n18390), .ZN(
        P3_U2957) );
  AOI22_X1 U21567 ( .A1(n18428), .A2(n18505), .B1(n18504), .B2(n18404), .ZN(
        n18393) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18405), .B1(
        n18506), .B2(n18403), .ZN(n18392) );
  OAI211_X1 U21569 ( .C1(n18473), .C2(n18509), .A(n18393), .B(n18392), .ZN(
        P3_U2958) );
  AOI22_X1 U21570 ( .A1(n18428), .A2(n18468), .B1(n18510), .B2(n18404), .ZN(
        n18395) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18405), .B1(
        n18481), .B2(n18513), .ZN(n18394) );
  OAI211_X1 U21572 ( .C1(n18472), .C2(n18396), .A(n18395), .B(n18394), .ZN(
        P3_U2959) );
  AOI22_X1 U21573 ( .A1(n18518), .A2(n18404), .B1(n18520), .B2(n18403), .ZN(
        n18398) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18405), .B1(
        n18428), .B2(n18519), .ZN(n18397) );
  OAI211_X1 U21575 ( .C1(n18473), .C2(n18523), .A(n18398), .B(n18397), .ZN(
        P3_U2960) );
  AOI22_X1 U21576 ( .A1(n18524), .A2(n18404), .B1(n18526), .B2(n18403), .ZN(
        n18400) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18405), .B1(
        n18428), .B2(n18525), .ZN(n18399) );
  OAI211_X1 U21578 ( .C1(n18473), .C2(n18529), .A(n18400), .B(n18399), .ZN(
        P3_U2961) );
  AOI22_X1 U21579 ( .A1(n18532), .A2(n18403), .B1(n18530), .B2(n18404), .ZN(
        n18402) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18405), .B1(
        n18428), .B2(n18531), .ZN(n18401) );
  OAI211_X1 U21581 ( .C1(n18473), .C2(n18535), .A(n18402), .B(n18401), .ZN(
        P3_U2962) );
  AOI22_X1 U21582 ( .A1(n18537), .A2(n18404), .B1(n18538), .B2(n18403), .ZN(
        n18407) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18405), .B1(
        n18428), .B2(n18541), .ZN(n18406) );
  OAI211_X1 U21584 ( .C1(n18473), .C2(n18546), .A(n18407), .B(n18406), .ZN(
        P3_U2963) );
  NOR2_X2 U21585 ( .A1(n18592), .A2(n18433), .ZN(n18539) );
  INV_X1 U21586 ( .A(n18539), .ZN(n18457) );
  AOI21_X1 U21587 ( .B1(n18457), .B2(n18473), .A(n18487), .ZN(n18427) );
  AOI22_X1 U21588 ( .A1(n18452), .A2(n18494), .B1(n18488), .B2(n18427), .ZN(
        n18413) );
  AOI221_X1 U21589 ( .B1(n18409), .B2(n18473), .C1(n18408), .C2(n18473), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18411) );
  OAI21_X1 U21590 ( .B1(n18539), .B2(n18411), .A(n18410), .ZN(n18429) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18429), .B1(
        n18539), .B2(n18460), .ZN(n18412) );
  OAI211_X1 U21592 ( .C1(n18420), .C2(n18463), .A(n18413), .B(n18412), .ZN(
        P3_U2964) );
  AOI22_X1 U21593 ( .A1(n18428), .A2(n18499), .B1(n18427), .B2(n18498), .ZN(
        n18415) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18429), .B1(
        n18452), .B2(n18500), .ZN(n18414) );
  OAI211_X1 U21595 ( .C1(n18457), .C2(n18503), .A(n18415), .B(n18414), .ZN(
        P3_U2965) );
  AOI22_X1 U21596 ( .A1(n18428), .A2(n18506), .B1(n18427), .B2(n18504), .ZN(
        n18417) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18429), .B1(
        n18452), .B2(n18505), .ZN(n18416) );
  OAI211_X1 U21598 ( .C1(n18457), .C2(n18509), .A(n18417), .B(n18416), .ZN(
        P3_U2966) );
  AOI22_X1 U21599 ( .A1(n18452), .A2(n18468), .B1(n18427), .B2(n18510), .ZN(
        n18419) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18429), .B1(
        n18539), .B2(n18513), .ZN(n18418) );
  OAI211_X1 U21601 ( .C1(n18420), .C2(n18472), .A(n18419), .B(n18418), .ZN(
        P3_U2967) );
  AOI22_X1 U21602 ( .A1(n18428), .A2(n18520), .B1(n18427), .B2(n18518), .ZN(
        n18422) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18429), .B1(
        n18452), .B2(n18519), .ZN(n18421) );
  OAI211_X1 U21604 ( .C1(n18457), .C2(n18523), .A(n18422), .B(n18421), .ZN(
        P3_U2968) );
  AOI22_X1 U21605 ( .A1(n18428), .A2(n18526), .B1(n18427), .B2(n18524), .ZN(
        n18424) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18429), .B1(
        n18452), .B2(n18525), .ZN(n18423) );
  OAI211_X1 U21607 ( .C1(n18457), .C2(n18529), .A(n18424), .B(n18423), .ZN(
        P3_U2969) );
  AOI22_X1 U21608 ( .A1(n18428), .A2(n18532), .B1(n18427), .B2(n18530), .ZN(
        n18426) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18429), .B1(
        n18452), .B2(n18531), .ZN(n18425) );
  OAI211_X1 U21610 ( .C1(n18457), .C2(n18535), .A(n18426), .B(n18425), .ZN(
        P3_U2970) );
  AOI22_X1 U21611 ( .A1(n18428), .A2(n18538), .B1(n18427), .B2(n18537), .ZN(
        n18431) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18429), .B1(
        n18452), .B2(n18541), .ZN(n18430) );
  OAI211_X1 U21613 ( .C1(n18457), .C2(n18546), .A(n18431), .B(n18430), .ZN(
        P3_U2971) );
  NOR2_X1 U21614 ( .A1(n18433), .A2(n18432), .ZN(n18492) );
  AOI22_X1 U21615 ( .A1(n18452), .A2(n18489), .B1(n18488), .B2(n18492), .ZN(
        n18438) );
  AOI22_X1 U21616 ( .A1(n18493), .A2(n18436), .B1(n18435), .B2(n18434), .ZN(
        n18453) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18453), .B1(
        n18481), .B2(n18494), .ZN(n18437) );
  OAI211_X1 U21618 ( .C1(n18497), .C2(n18516), .A(n18438), .B(n18437), .ZN(
        P3_U2972) );
  AOI22_X1 U21619 ( .A1(n18452), .A2(n18499), .B1(n18498), .B2(n18492), .ZN(
        n18440) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18453), .B1(
        n18481), .B2(n18500), .ZN(n18439) );
  OAI211_X1 U21621 ( .C1(n18503), .C2(n18516), .A(n18440), .B(n18439), .ZN(
        P3_U2973) );
  AOI22_X1 U21622 ( .A1(n18452), .A2(n18506), .B1(n18504), .B2(n18492), .ZN(
        n18442) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18453), .B1(
        n18481), .B2(n18505), .ZN(n18441) );
  OAI211_X1 U21624 ( .C1(n18509), .C2(n18516), .A(n18442), .B(n18441), .ZN(
        P3_U2974) );
  AOI22_X1 U21625 ( .A1(n18481), .A2(n18468), .B1(n18510), .B2(n18492), .ZN(
        n18444) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18453), .B1(
        n18513), .B2(n18540), .ZN(n18443) );
  OAI211_X1 U21627 ( .C1(n18445), .C2(n18472), .A(n18444), .B(n18443), .ZN(
        P3_U2975) );
  AOI22_X1 U21628 ( .A1(n18452), .A2(n18520), .B1(n18518), .B2(n18492), .ZN(
        n18447) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18453), .B1(
        n18481), .B2(n18519), .ZN(n18446) );
  OAI211_X1 U21630 ( .C1(n18523), .C2(n18516), .A(n18447), .B(n18446), .ZN(
        P3_U2976) );
  AOI22_X1 U21631 ( .A1(n18452), .A2(n18526), .B1(n18524), .B2(n18492), .ZN(
        n18449) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18453), .B1(
        n18481), .B2(n18525), .ZN(n18448) );
  OAI211_X1 U21633 ( .C1(n18529), .C2(n18516), .A(n18449), .B(n18448), .ZN(
        P3_U2977) );
  AOI22_X1 U21634 ( .A1(n18481), .A2(n18531), .B1(n18530), .B2(n18492), .ZN(
        n18451) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18453), .B1(
        n18452), .B2(n18532), .ZN(n18450) );
  OAI211_X1 U21636 ( .C1(n18535), .C2(n18516), .A(n18451), .B(n18450), .ZN(
        P3_U2978) );
  AOI22_X1 U21637 ( .A1(n18481), .A2(n18541), .B1(n18537), .B2(n18492), .ZN(
        n18455) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18453), .B1(
        n18452), .B2(n18538), .ZN(n18454) );
  OAI211_X1 U21639 ( .C1(n18546), .C2(n18516), .A(n18455), .B(n18454), .ZN(
        P3_U2979) );
  AOI21_X1 U21640 ( .B1(n18516), .B2(n18485), .A(n18487), .ZN(n18480) );
  AOI22_X1 U21641 ( .A1(n18539), .A2(n18494), .B1(n18488), .B2(n18480), .ZN(
        n18462) );
  AOI21_X1 U21642 ( .B1(n18457), .B2(n18473), .A(n18456), .ZN(n18458) );
  OAI22_X1 U21643 ( .A1(n18469), .A2(n18743), .B1(n18459), .B2(n18458), .ZN(
        n18482) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18482), .B1(
        n18460), .B2(n18469), .ZN(n18461) );
  OAI211_X1 U21645 ( .C1(n18473), .C2(n18463), .A(n18462), .B(n18461), .ZN(
        P3_U2980) );
  AOI22_X1 U21646 ( .A1(n18539), .A2(n18500), .B1(n18498), .B2(n18480), .ZN(
        n18465) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18482), .B1(
        n18481), .B2(n18499), .ZN(n18464) );
  OAI211_X1 U21648 ( .C1(n18503), .C2(n18485), .A(n18465), .B(n18464), .ZN(
        P3_U2981) );
  AOI22_X1 U21649 ( .A1(n18481), .A2(n18506), .B1(n18504), .B2(n18480), .ZN(
        n18467) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18482), .B1(
        n18539), .B2(n18505), .ZN(n18466) );
  OAI211_X1 U21651 ( .C1(n18509), .C2(n18485), .A(n18467), .B(n18466), .ZN(
        P3_U2982) );
  AOI22_X1 U21652 ( .A1(n18539), .A2(n18468), .B1(n18510), .B2(n18480), .ZN(
        n18471) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18482), .B1(
        n18513), .B2(n18469), .ZN(n18470) );
  OAI211_X1 U21654 ( .C1(n18473), .C2(n18472), .A(n18471), .B(n18470), .ZN(
        P3_U2983) );
  AOI22_X1 U21655 ( .A1(n18481), .A2(n18520), .B1(n18518), .B2(n18480), .ZN(
        n18475) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18482), .B1(
        n18539), .B2(n18519), .ZN(n18474) );
  OAI211_X1 U21657 ( .C1(n18523), .C2(n18485), .A(n18475), .B(n18474), .ZN(
        P3_U2984) );
  AOI22_X1 U21658 ( .A1(n18539), .A2(n18525), .B1(n18524), .B2(n18480), .ZN(
        n18477) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18482), .B1(
        n18481), .B2(n18526), .ZN(n18476) );
  OAI211_X1 U21660 ( .C1(n18529), .C2(n18485), .A(n18477), .B(n18476), .ZN(
        P3_U2985) );
  AOI22_X1 U21661 ( .A1(n18481), .A2(n18532), .B1(n18530), .B2(n18480), .ZN(
        n18479) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18482), .B1(
        n18539), .B2(n18531), .ZN(n18478) );
  OAI211_X1 U21663 ( .C1(n18535), .C2(n18485), .A(n18479), .B(n18478), .ZN(
        P3_U2986) );
  AOI22_X1 U21664 ( .A1(n18481), .A2(n18538), .B1(n18537), .B2(n18480), .ZN(
        n18484) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18482), .B1(
        n18539), .B2(n18541), .ZN(n18483) );
  OAI211_X1 U21666 ( .C1(n18546), .C2(n18485), .A(n18484), .B(n18483), .ZN(
        P3_U2987) );
  INV_X1 U21667 ( .A(n18491), .ZN(n18486) );
  NOR2_X1 U21668 ( .A1(n18487), .A2(n18486), .ZN(n18536) );
  AOI22_X1 U21669 ( .A1(n18539), .A2(n18489), .B1(n18488), .B2(n18536), .ZN(
        n18496) );
  AOI22_X1 U21670 ( .A1(n18493), .A2(n18492), .B1(n18491), .B2(n18490), .ZN(
        n18542) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18542), .B1(
        n18494), .B2(n18540), .ZN(n18495) );
  OAI211_X1 U21672 ( .C1(n18497), .C2(n18545), .A(n18496), .B(n18495), .ZN(
        P3_U2988) );
  AOI22_X1 U21673 ( .A1(n18539), .A2(n18499), .B1(n18498), .B2(n18536), .ZN(
        n18502) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18542), .B1(
        n18500), .B2(n18540), .ZN(n18501) );
  OAI211_X1 U21675 ( .C1(n18503), .C2(n18545), .A(n18502), .B(n18501), .ZN(
        P3_U2989) );
  AOI22_X1 U21676 ( .A1(n18505), .A2(n18540), .B1(n18504), .B2(n18536), .ZN(
        n18508) );
  AOI22_X1 U21677 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18542), .B1(
        n18539), .B2(n18506), .ZN(n18507) );
  OAI211_X1 U21678 ( .C1(n18509), .C2(n18545), .A(n18508), .B(n18507), .ZN(
        P3_U2990) );
  AOI22_X1 U21679 ( .A1(n18539), .A2(n18511), .B1(n18510), .B2(n18536), .ZN(
        n18515) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18542), .B1(
        n18513), .B2(n18512), .ZN(n18514) );
  OAI211_X1 U21681 ( .C1(n18517), .C2(n18516), .A(n18515), .B(n18514), .ZN(
        P3_U2991) );
  AOI22_X1 U21682 ( .A1(n18519), .A2(n18540), .B1(n18518), .B2(n18536), .ZN(
        n18522) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18542), .B1(
        n18539), .B2(n18520), .ZN(n18521) );
  OAI211_X1 U21684 ( .C1(n18523), .C2(n18545), .A(n18522), .B(n18521), .ZN(
        P3_U2992) );
  AOI22_X1 U21685 ( .A1(n18525), .A2(n18540), .B1(n18524), .B2(n18536), .ZN(
        n18528) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18542), .B1(
        n18539), .B2(n18526), .ZN(n18527) );
  OAI211_X1 U21687 ( .C1(n18529), .C2(n18545), .A(n18528), .B(n18527), .ZN(
        P3_U2993) );
  AOI22_X1 U21688 ( .A1(n18531), .A2(n18540), .B1(n18530), .B2(n18536), .ZN(
        n18534) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18542), .B1(
        n18539), .B2(n18532), .ZN(n18533) );
  OAI211_X1 U21690 ( .C1(n18535), .C2(n18545), .A(n18534), .B(n18533), .ZN(
        P3_U2994) );
  AOI22_X1 U21691 ( .A1(n18539), .A2(n18538), .B1(n18537), .B2(n18536), .ZN(
        n18544) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18540), .ZN(n18543) );
  OAI211_X1 U21693 ( .C1(n18546), .C2(n18545), .A(n18544), .B(n18543), .ZN(
        P3_U2995) );
  INV_X1 U21694 ( .A(n18547), .ZN(n18554) );
  INV_X1 U21695 ( .A(n18548), .ZN(n18553) );
  NOR2_X1 U21696 ( .A1(n18581), .A2(n18549), .ZN(n18552) );
  OAI222_X1 U21697 ( .A1(n18555), .A2(n18554), .B1(n18553), .B2(n18552), .C1(
        n18551), .C2(n18550), .ZN(n18761) );
  OAI21_X1 U21698 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18556), .ZN(n18558) );
  OAI211_X1 U21699 ( .C1(n18582), .C2(n18607), .A(n18558), .B(n18557), .ZN(
        n18605) );
  NOR2_X1 U21700 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18559), .ZN(
        n18586) );
  INV_X1 U21701 ( .A(n18586), .ZN(n18560) );
  AOI22_X1 U21702 ( .A1(n18569), .A2(n18560), .B1(n18581), .B2(n18561), .ZN(
        n18718) );
  NOR2_X1 U21703 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18718), .ZN(
        n18566) );
  INV_X1 U21704 ( .A(n18582), .ZN(n18594) );
  INV_X1 U21705 ( .A(n18561), .ZN(n18562) );
  AOI21_X1 U21706 ( .B1(n18563), .B2(n18567), .A(n18562), .ZN(n18564) );
  OAI21_X1 U21707 ( .B1(n18569), .B2(n18585), .A(n18564), .ZN(n18721) );
  OR2_X1 U21708 ( .A1(n18594), .A2(n18721), .ZN(n18565) );
  AOI22_X1 U21709 ( .A1(n18582), .A2(n18566), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18565), .ZN(n18603) );
  AOI21_X1 U21710 ( .B1(n18741), .B2(n18573), .A(n18567), .ZN(n18578) );
  NAND2_X1 U21711 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18568), .ZN(
        n18577) );
  INV_X1 U21712 ( .A(n18569), .ZN(n18570) );
  OAI211_X1 U21713 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18571), .B(n18570), .ZN(
        n18576) );
  NOR2_X1 U21714 ( .A1(n18572), .A2(n18749), .ZN(n18574) );
  OAI211_X1 U21715 ( .C1(n18574), .C2(n18573), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n18734), .ZN(n18575) );
  OAI211_X1 U21716 ( .C1(n18578), .C2(n18577), .A(n18576), .B(n18575), .ZN(
        n18579) );
  AOI21_X1 U21717 ( .B1(n18581), .B2(n18580), .A(n18579), .ZN(n18730) );
  AOI22_X1 U21718 ( .A1(n18594), .A2(n18734), .B1(n18730), .B2(n18582), .ZN(
        n18598) );
  NOR2_X1 U21719 ( .A1(n18584), .A2(n18583), .ZN(n18588) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18585), .B1(
        n18588), .B2(n18749), .ZN(n18744) );
  OAI22_X1 U21721 ( .A1(n18588), .A2(n18587), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18586), .ZN(n18738) );
  OR3_X1 U21722 ( .A1(n18744), .A2(n18591), .A3(n18589), .ZN(n18590) );
  AOI22_X1 U21723 ( .A1(n18744), .A2(n18591), .B1(n18738), .B2(n18590), .ZN(
        n18593) );
  OAI21_X1 U21724 ( .B1(n18594), .B2(n18593), .A(n18592), .ZN(n18597) );
  AND2_X1 U21725 ( .A1(n18598), .A2(n18597), .ZN(n18595) );
  OAI221_X1 U21726 ( .B1(n18598), .B2(n18597), .C1(n18596), .C2(n18595), .A(
        n18600), .ZN(n18602) );
  AOI21_X1 U21727 ( .B1(n18600), .B2(n18599), .A(n18598), .ZN(n18601) );
  AOI222_X1 U21728 ( .A1(n18603), .A2(n18602), .B1(n18603), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18602), .C2(n18601), .ZN(
        n18604) );
  NOR4_X1 U21729 ( .A1(n18606), .A2(n18761), .A3(n18605), .A4(n18604), .ZN(
        n18618) );
  NOR2_X1 U21730 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18613), .ZN(n18608) );
  AOI22_X1 U21731 ( .A1(n18609), .A2(n18764), .B1(n18608), .B2(n18607), .ZN(
        n18615) );
  OAI211_X1 U21732 ( .C1(n18611), .C2(n18610), .A(n18771), .B(n18618), .ZN(
        n18612) );
  NAND2_X1 U21733 ( .A1(n18764), .A2(n18779), .ZN(n18619) );
  OAI211_X1 U21734 ( .C1(P3_STATE2_REG_1__SCAN_IN), .C2(n18613), .A(n18717), 
        .B(n18619), .ZN(n18622) );
  OAI22_X1 U21735 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18615), .B1(n18614), 
        .B2(n18622), .ZN(n18616) );
  OAI21_X1 U21736 ( .B1(n18618), .B2(n18617), .A(n18616), .ZN(P3_U2996) );
  NOR3_X1 U21737 ( .A1(n18726), .A2(n18767), .A3(n18619), .ZN(n18624) );
  AOI211_X1 U21738 ( .C1(n18764), .C2(n18774), .A(n18620), .B(n18624), .ZN(
        n18621) );
  OAI21_X1 U21739 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18622), .A(n18621), 
        .ZN(P3_U2997) );
  NOR4_X1 U21740 ( .A1(n18626), .A2(n18625), .A3(n18624), .A4(n18623), .ZN(
        P3_U2998) );
  INV_X1 U21741 ( .A(n18715), .ZN(n18712) );
  AND2_X1 U21742 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18712), .ZN(
        P3_U2999) );
  AND2_X1 U21743 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18712), .ZN(
        P3_U3000) );
  AND2_X1 U21744 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18712), .ZN(
        P3_U3001) );
  AND2_X1 U21745 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18712), .ZN(
        P3_U3002) );
  AND2_X1 U21746 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18712), .ZN(
        P3_U3003) );
  AND2_X1 U21747 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18712), .ZN(
        P3_U3004) );
  AND2_X1 U21748 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18712), .ZN(
        P3_U3005) );
  AND2_X1 U21749 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18712), .ZN(
        P3_U3006) );
  AND2_X1 U21750 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18712), .ZN(
        P3_U3007) );
  AND2_X1 U21751 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18712), .ZN(
        P3_U3008) );
  AND2_X1 U21752 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18712), .ZN(
        P3_U3009) );
  AND2_X1 U21753 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18712), .ZN(
        P3_U3010) );
  AND2_X1 U21754 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18712), .ZN(
        P3_U3011) );
  AND2_X1 U21755 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18712), .ZN(
        P3_U3012) );
  AND2_X1 U21756 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18712), .ZN(
        P3_U3013) );
  AND2_X1 U21757 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18712), .ZN(
        P3_U3014) );
  AND2_X1 U21758 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18712), .ZN(
        P3_U3015) );
  AND2_X1 U21759 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18712), .ZN(
        P3_U3016) );
  AND2_X1 U21760 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18712), .ZN(
        P3_U3017) );
  AND2_X1 U21761 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18712), .ZN(
        P3_U3018) );
  AND2_X1 U21762 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18712), .ZN(
        P3_U3019) );
  AND2_X1 U21763 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18712), .ZN(
        P3_U3020) );
  AND2_X1 U21764 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18712), .ZN(P3_U3021) );
  AND2_X1 U21765 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18712), .ZN(P3_U3022) );
  AND2_X1 U21766 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18712), .ZN(P3_U3023) );
  AND2_X1 U21767 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18712), .ZN(P3_U3024) );
  AND2_X1 U21768 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18712), .ZN(P3_U3025) );
  AND2_X1 U21769 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18712), .ZN(P3_U3026) );
  AND2_X1 U21770 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18712), .ZN(P3_U3027) );
  AND2_X1 U21771 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18712), .ZN(P3_U3028) );
  INV_X1 U21772 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18633) );
  AOI21_X1 U21773 ( .B1(HOLD), .B2(n18627), .A(n18633), .ZN(n18630) );
  AOI21_X1 U21774 ( .B1(n18764), .B2(P3_STATE_REG_1__SCAN_IN), .A(n18628), 
        .ZN(n18642) );
  AOI21_X1 U21775 ( .B1(n18629), .B2(NA), .A(n18643), .ZN(n18637) );
  OAI22_X1 U21776 ( .A1(n18758), .A2(n18630), .B1(n18642), .B2(n18637), .ZN(
        P3_U3029) );
  NAND3_X1 U21777 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(HOLD), .A3(n18643), .ZN(
        n18631) );
  OAI221_X1 U21778 ( .B1(n18633), .B2(HOLD), .C1(n18633), .C2(n18632), .A(
        n18631), .ZN(n18634) );
  AOI22_X1 U21779 ( .A1(n18764), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18634), .ZN(n18636) );
  NAND2_X1 U21780 ( .A1(n18636), .A2(n18635), .ZN(P3_U3030) );
  INV_X1 U21781 ( .A(n18637), .ZN(n18641) );
  NAND2_X1 U21782 ( .A1(n18764), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18638) );
  OAI222_X1 U21783 ( .A1(n18643), .A2(n20761), .B1(P3_STATE_REG_1__SCAN_IN), 
        .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(n18638), .C2(NA), .ZN(n18639)
         );
  OAI211_X1 U21784 ( .C1(P3_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .B(n18639), .ZN(n18640) );
  OAI21_X1 U21785 ( .B1(n18642), .B2(n18641), .A(n18640), .ZN(P3_U3031) );
  INV_X1 U21786 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18645) );
  OAI222_X1 U21787 ( .A1(n18750), .A2(n18705), .B1(n18644), .B2(n18758), .C1(
        n18645), .C2(n18701), .ZN(P3_U3032) );
  OAI222_X1 U21788 ( .A1(n18701), .A2(n18648), .B1(n18646), .B2(n18758), .C1(
        n18645), .C2(n18705), .ZN(P3_U3033) );
  OAI222_X1 U21789 ( .A1(n18648), .A2(n18705), .B1(n18647), .B2(n18758), .C1(
        n18649), .C2(n18701), .ZN(P3_U3034) );
  OAI222_X1 U21790 ( .A1(n18701), .A2(n18651), .B1(n18650), .B2(n18758), .C1(
        n18649), .C2(n18705), .ZN(P3_U3035) );
  OAI222_X1 U21791 ( .A1(n18701), .A2(n18653), .B1(n18652), .B2(n18758), .C1(
        n18651), .C2(n18705), .ZN(P3_U3036) );
  OAI222_X1 U21792 ( .A1(n18701), .A2(n18655), .B1(n18654), .B2(n18758), .C1(
        n18653), .C2(n18705), .ZN(P3_U3037) );
  INV_X1 U21793 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18657) );
  OAI222_X1 U21794 ( .A1(n18701), .A2(n18657), .B1(n18656), .B2(n18758), .C1(
        n18655), .C2(n18705), .ZN(P3_U3038) );
  OAI222_X1 U21795 ( .A1(n18701), .A2(n18659), .B1(n18658), .B2(n18758), .C1(
        n18657), .C2(n18705), .ZN(P3_U3039) );
  OAI222_X1 U21796 ( .A1(n18701), .A2(n18661), .B1(n18660), .B2(n18758), .C1(
        n18659), .C2(n18705), .ZN(P3_U3040) );
  OAI222_X1 U21797 ( .A1(n18701), .A2(n18663), .B1(n18662), .B2(n18758), .C1(
        n18661), .C2(n18705), .ZN(P3_U3041) );
  OAI222_X1 U21798 ( .A1(n18701), .A2(n18665), .B1(n18664), .B2(n18758), .C1(
        n18663), .C2(n18705), .ZN(P3_U3042) );
  OAI222_X1 U21799 ( .A1(n18701), .A2(n18667), .B1(n18666), .B2(n18758), .C1(
        n18665), .C2(n18705), .ZN(P3_U3043) );
  OAI222_X1 U21800 ( .A1(n18701), .A2(n18670), .B1(n18668), .B2(n18758), .C1(
        n18667), .C2(n18705), .ZN(P3_U3044) );
  OAI222_X1 U21801 ( .A1(n18670), .A2(n18705), .B1(n18669), .B2(n18758), .C1(
        n18671), .C2(n18701), .ZN(P3_U3045) );
  OAI222_X1 U21802 ( .A1(n18701), .A2(n18673), .B1(n18672), .B2(n18758), .C1(
        n18671), .C2(n18705), .ZN(P3_U3046) );
  OAI222_X1 U21803 ( .A1(n18701), .A2(n18676), .B1(n18674), .B2(n18758), .C1(
        n18673), .C2(n18705), .ZN(P3_U3047) );
  OAI222_X1 U21804 ( .A1(n18676), .A2(n18705), .B1(n18675), .B2(n18758), .C1(
        n18677), .C2(n18701), .ZN(P3_U3048) );
  OAI222_X1 U21805 ( .A1(n18701), .A2(n18680), .B1(n18678), .B2(n18758), .C1(
        n18677), .C2(n18705), .ZN(P3_U3049) );
  OAI222_X1 U21806 ( .A1(n18680), .A2(n18705), .B1(n18679), .B2(n18758), .C1(
        n18682), .C2(n18701), .ZN(P3_U3050) );
  OAI222_X1 U21807 ( .A1(n18705), .A2(n18682), .B1(n18681), .B2(n18758), .C1(
        n18683), .C2(n18701), .ZN(P3_U3051) );
  OAI222_X1 U21808 ( .A1(n18701), .A2(n18685), .B1(n18684), .B2(n18758), .C1(
        n18683), .C2(n18705), .ZN(P3_U3052) );
  OAI222_X1 U21809 ( .A1(n18701), .A2(n18687), .B1(n18686), .B2(n18758), .C1(
        n18685), .C2(n18705), .ZN(P3_U3053) );
  OAI222_X1 U21810 ( .A1(n18701), .A2(n18689), .B1(n18688), .B2(n18758), .C1(
        n18687), .C2(n18705), .ZN(P3_U3054) );
  OAI222_X1 U21811 ( .A1(n18701), .A2(n18691), .B1(n18690), .B2(n18758), .C1(
        n18689), .C2(n18705), .ZN(P3_U3055) );
  OAI222_X1 U21812 ( .A1(n18701), .A2(n18693), .B1(n18692), .B2(n18758), .C1(
        n18691), .C2(n18705), .ZN(P3_U3056) );
  OAI222_X1 U21813 ( .A1(n18701), .A2(n18695), .B1(n18694), .B2(n18758), .C1(
        n18693), .C2(n18705), .ZN(P3_U3057) );
  OAI222_X1 U21814 ( .A1(n18701), .A2(n18698), .B1(n18696), .B2(n18758), .C1(
        n18695), .C2(n18705), .ZN(P3_U3058) );
  OAI222_X1 U21815 ( .A1(n18698), .A2(n18705), .B1(n18697), .B2(n18758), .C1(
        n18699), .C2(n18701), .ZN(P3_U3059) );
  OAI222_X1 U21816 ( .A1(n18701), .A2(n18704), .B1(n18700), .B2(n18758), .C1(
        n18699), .C2(n18705), .ZN(P3_U3060) );
  OAI222_X1 U21817 ( .A1(n18705), .A2(n18704), .B1(n18703), .B2(n18758), .C1(
        n18702), .C2(n18701), .ZN(P3_U3061) );
  OAI22_X1 U21818 ( .A1(n18777), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18758), .ZN(n18706) );
  INV_X1 U21819 ( .A(n18706), .ZN(P3_U3274) );
  OAI22_X1 U21820 ( .A1(n18777), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18758), .ZN(n18707) );
  INV_X1 U21821 ( .A(n18707), .ZN(P3_U3275) );
  OAI22_X1 U21822 ( .A1(n18777), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18758), .ZN(n18708) );
  INV_X1 U21823 ( .A(n18708), .ZN(P3_U3276) );
  OAI22_X1 U21824 ( .A1(n18777), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18758), .ZN(n18709) );
  INV_X1 U21825 ( .A(n18709), .ZN(P3_U3277) );
  INV_X1 U21826 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18711) );
  INV_X1 U21827 ( .A(n18713), .ZN(n18710) );
  AOI21_X1 U21828 ( .B1(n18712), .B2(n18711), .A(n18710), .ZN(P3_U3280) );
  OAI21_X1 U21829 ( .B1(n18715), .B2(n18714), .A(n18713), .ZN(P3_U3281) );
  OAI21_X1 U21830 ( .B1(n18717), .B2(n18743), .A(n18716), .ZN(P3_U3282) );
  NOR3_X1 U21831 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18718), .A3(
        n18729), .ZN(n18719) );
  AOI21_X1 U21832 ( .B1(n18720), .B2(n18745), .A(n18719), .ZN(n18724) );
  AOI21_X1 U21833 ( .B1(n18780), .B2(n18721), .A(n18748), .ZN(n18723) );
  OAI22_X1 U21834 ( .A1(n18748), .A2(n18724), .B1(n18723), .B2(n18722), .ZN(
        P3_U3285) );
  NOR2_X1 U21835 ( .A1(n18726), .A2(n18725), .ZN(n18735) );
  INV_X1 U21836 ( .A(n18735), .ZN(n18742) );
  AOI22_X1 U21837 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18728), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18727), .ZN(n18736) );
  OAI22_X1 U21838 ( .A1(n18730), .A2(n18729), .B1(n18742), .B2(n18736), .ZN(
        n18731) );
  AOI21_X1 U21839 ( .B1(n18745), .B2(n18732), .A(n18731), .ZN(n18733) );
  INV_X1 U21840 ( .A(n18748), .ZN(n18739) );
  AOI22_X1 U21841 ( .A1(n18748), .A2(n18734), .B1(n18733), .B2(n18739), .ZN(
        P3_U3288) );
  AOI222_X1 U21842 ( .A1(n18738), .A2(n18780), .B1(n18745), .B2(n18737), .C1(
        n18736), .C2(n18735), .ZN(n18740) );
  AOI22_X1 U21843 ( .A1(n18748), .A2(n18741), .B1(n18740), .B2(n18739), .ZN(
        P3_U3289) );
  OAI221_X1 U21844 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18744), .C1(
        P3_STATE2_REG_1__SCAN_IN), .C2(n18743), .A(n18742), .ZN(n18747) );
  AOI21_X1 U21845 ( .B1(n18749), .B2(n18745), .A(n18748), .ZN(n18746) );
  AOI22_X1 U21846 ( .A1(n18749), .A2(n18748), .B1(n18747), .B2(n18746), .ZN(
        P3_U3290) );
  AOI21_X1 U21847 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18751) );
  AOI22_X1 U21848 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18751), .B2(n18750), .ZN(n18754) );
  INV_X1 U21849 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18753) );
  AOI22_X1 U21850 ( .A1(n18757), .A2(n18754), .B1(n18753), .B2(n18752), .ZN(
        P3_U3292) );
  INV_X1 U21851 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18756) );
  OAI21_X1 U21852 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18757), .ZN(n18755) );
  OAI21_X1 U21853 ( .B1(n18757), .B2(n18756), .A(n18755), .ZN(P3_U3293) );
  INV_X1 U21854 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18783) );
  OAI22_X1 U21855 ( .A1(n18777), .A2(n18783), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18758), .ZN(n18759) );
  INV_X1 U21856 ( .A(n18759), .ZN(P3_U3294) );
  MUX2_X1 U21857 ( .A(P3_MORE_REG_SCAN_IN), .B(n18761), .S(n18760), .Z(
        P3_U3295) );
  OAI21_X1 U21858 ( .B1(n18763), .B2(P3_STATEBS16_REG_SCAN_IN), .A(n18762), 
        .ZN(n18765) );
  AOI211_X1 U21859 ( .C1(n18781), .C2(n18765), .A(n18764), .B(n18779), .ZN(
        n18768) );
  OAI21_X1 U21860 ( .B1(n18768), .B2(n18767), .A(n18766), .ZN(n18776) );
  OAI21_X1 U21861 ( .B1(n18771), .B2(n18770), .A(n18769), .ZN(n18772) );
  AOI21_X1 U21862 ( .B1(n18774), .B2(n18773), .A(n18772), .ZN(n18775) );
  MUX2_X1 U21863 ( .A(n18776), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n18775), 
        .Z(P3_U3296) );
  OAI22_X1 U21864 ( .A1(n18777), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18758), .ZN(n18778) );
  INV_X1 U21865 ( .A(n18778), .ZN(P3_U3297) );
  AOI21_X1 U21866 ( .B1(n18780), .B2(n18779), .A(n18782), .ZN(n18786) );
  AOI22_X1 U21867 ( .A1(n18786), .A2(n18783), .B1(n18782), .B2(n18781), .ZN(
        P3_U3298) );
  INV_X1 U21868 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18785) );
  AOI21_X1 U21869 ( .B1(n18786), .B2(n18785), .A(n18784), .ZN(P3_U3299) );
  INV_X1 U21870 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19729) );
  AND2_X1 U21871 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19729), .ZN(n19719) );
  NOR2_X1 U21872 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19712) );
  AOI21_X1 U21873 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19719), .A(n19712), 
        .ZN(n19711) );
  INV_X1 U21874 ( .A(n19711), .ZN(n19787) );
  AOI21_X1 U21875 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19787), .ZN(n18787) );
  INV_X1 U21876 ( .A(n18787), .ZN(P2_U2815) );
  INV_X1 U21877 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18789) );
  OAI22_X1 U21878 ( .A1(n19846), .A2(n18789), .B1(n19855), .B2(n18788), .ZN(
        P2_U2816) );
  AOI21_X1 U21879 ( .B1(n19717), .B2(n19729), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18790) );
  AOI22_X1 U21880 ( .A1(n19867), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18790), 
        .B2(n19864), .ZN(P2_U2817) );
  OAI21_X1 U21881 ( .B1(n19713), .B2(BS16), .A(n19787), .ZN(n19785) );
  OAI21_X1 U21882 ( .B1(n19787), .B2(n19797), .A(n19785), .ZN(P2_U2818) );
  NOR2_X1 U21883 ( .A1(n18791), .A2(n19849), .ZN(n19841) );
  OAI21_X1 U21884 ( .B1(n19841), .B2(n10339), .A(n18792), .ZN(P2_U2819) );
  NOR4_X1 U21885 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18802) );
  NOR4_X1 U21886 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n18801) );
  NOR4_X1 U21887 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18793) );
  INV_X1 U21888 ( .A(P2_DATAWIDTH_REG_24__SCAN_IN), .ZN(n19708) );
  NAND3_X1 U21889 ( .A1(n18793), .A2(n19709), .A3(n19708), .ZN(n18799) );
  NOR4_X1 U21890 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18797) );
  NOR4_X1 U21891 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18796) );
  NOR4_X1 U21892 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18795) );
  NOR4_X1 U21893 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18794) );
  NAND4_X1 U21894 ( .A1(n18797), .A2(n18796), .A3(n18795), .A4(n18794), .ZN(
        n18798) );
  AOI211_X1 U21895 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n18799), .B(n18798), .ZN(n18800) );
  NAND3_X1 U21896 ( .A1(n18802), .A2(n18801), .A3(n18800), .ZN(n18810) );
  NOR2_X1 U21897 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18810), .ZN(n18805) );
  INV_X1 U21898 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18803) );
  AOI22_X1 U21899 ( .A1(n18805), .A2(n19024), .B1(n18810), .B2(n18803), .ZN(
        P2_U2820) );
  OR3_X1 U21900 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18809) );
  INV_X1 U21901 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18804) );
  AOI22_X1 U21902 ( .A1(n18805), .A2(n18809), .B1(n18810), .B2(n18804), .ZN(
        P2_U2821) );
  INV_X1 U21903 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19786) );
  NAND2_X1 U21904 ( .A1(n18805), .A2(n19786), .ZN(n18808) );
  INV_X1 U21905 ( .A(n18810), .ZN(n18812) );
  OAI21_X1 U21906 ( .B1(n19024), .B2(n19731), .A(n18812), .ZN(n18806) );
  OAI21_X1 U21907 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18812), .A(n18806), 
        .ZN(n18807) );
  OAI221_X1 U21908 ( .B1(n18808), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18808), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18807), .ZN(P2_U2822) );
  INV_X1 U21909 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18811) );
  OAI221_X1 U21910 ( .B1(n18812), .B2(n18811), .C1(n18810), .C2(n18809), .A(
        n18808), .ZN(P2_U2823) );
  OAI22_X1 U21911 ( .A1(n19760), .A2(n19004), .B1(n18813), .B2(n18850), .ZN(
        n18816) );
  OAI22_X1 U21912 ( .A1(n19006), .A2(n12041), .B1(n18814), .B2(n18989), .ZN(
        n18815) );
  AOI211_X1 U21913 ( .C1(n18817), .C2(n18998), .A(n18816), .B(n18815), .ZN(
        n18822) );
  OAI211_X1 U21914 ( .C1(n18820), .C2(n18819), .A(n19000), .B(n18818), .ZN(
        n18821) );
  OAI211_X1 U21915 ( .C1(n19032), .C2(n18823), .A(n18822), .B(n18821), .ZN(
        P2_U2834) );
  INV_X1 U21916 ( .A(n18824), .ZN(n18829) );
  AOI22_X1 U21917 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19038), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19027), .ZN(n18825) );
  INV_X1 U21918 ( .A(n18825), .ZN(n18828) );
  OAI22_X1 U21919 ( .A1(n19006), .A2(n9997), .B1(n18826), .B2(n18989), .ZN(
        n18827) );
  AOI211_X1 U21920 ( .C1(n18829), .C2(n19008), .A(n18828), .B(n18827), .ZN(
        n18834) );
  OAI211_X1 U21921 ( .C1(n18832), .C2(n18831), .A(n19000), .B(n18830), .ZN(
        n18833) );
  OAI211_X1 U21922 ( .C1(n19022), .C2(n18835), .A(n18834), .B(n18833), .ZN(
        P2_U2835) );
  AOI22_X1 U21923 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n19028), .B1(n18836), 
        .B2(n19026), .ZN(n18837) );
  OAI211_X1 U21924 ( .C1(n19756), .C2(n19004), .A(n18837), .B(n18966), .ZN(
        n18838) );
  AOI21_X1 U21925 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19038), .A(
        n18838), .ZN(n18846) );
  AOI22_X1 U21926 ( .A1(n18840), .A2(n18998), .B1(n18839), .B2(n19008), .ZN(
        n18845) );
  OAI211_X1 U21927 ( .C1(n18843), .C2(n18842), .A(n19000), .B(n18841), .ZN(
        n18844) );
  NAND3_X1 U21928 ( .A1(n18846), .A2(n18845), .A3(n18844), .ZN(P2_U2836) );
  AOI21_X1 U21929 ( .B1(P2_REIP_REG_18__SCAN_IN), .B2(n19027), .A(n18992), 
        .ZN(n18849) );
  AOI22_X1 U21930 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n19028), .B1(n18847), 
        .B2(n19026), .ZN(n18848) );
  OAI211_X1 U21931 ( .C1(n10032), .C2(n18850), .A(n18849), .B(n18848), .ZN(
        n18851) );
  AOI21_X1 U21932 ( .B1(n18852), .B2(n19008), .A(n18851), .ZN(n18857) );
  OAI211_X1 U21933 ( .C1(n18855), .C2(n18854), .A(n19000), .B(n18853), .ZN(
        n18856) );
  OAI211_X1 U21934 ( .C1(n19022), .C2(n18858), .A(n18857), .B(n18856), .ZN(
        P2_U2837) );
  AOI21_X1 U21935 ( .B1(P2_REIP_REG_17__SCAN_IN), .B2(n19027), .A(n18992), 
        .ZN(n18860) );
  AOI22_X1 U21936 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19038), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n19028), .ZN(n18859) );
  OAI211_X1 U21937 ( .C1(n18861), .C2(n18989), .A(n18860), .B(n18859), .ZN(
        n18862) );
  AOI21_X1 U21938 ( .B1(n18863), .B2(n18998), .A(n18862), .ZN(n18868) );
  OAI211_X1 U21939 ( .C1(n18866), .C2(n18865), .A(n19000), .B(n18864), .ZN(
        n18867) );
  OAI211_X1 U21940 ( .C1(n19032), .C2(n18869), .A(n18868), .B(n18867), .ZN(
        P2_U2838) );
  AOI21_X1 U21941 ( .B1(P2_REIP_REG_16__SCAN_IN), .B2(n19027), .A(n18992), 
        .ZN(n18871) );
  AOI22_X1 U21942 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19038), .B1(
        P2_EBX_REG_16__SCAN_IN), .B2(n19028), .ZN(n18870) );
  OAI211_X1 U21943 ( .C1(n18872), .C2(n18989), .A(n18871), .B(n18870), .ZN(
        n18873) );
  AOI21_X1 U21944 ( .B1(n19097), .B2(n19008), .A(n18873), .ZN(n18878) );
  OAI211_X1 U21945 ( .C1(n18876), .C2(n18875), .A(n19000), .B(n18874), .ZN(
        n18877) );
  OAI211_X1 U21946 ( .C1(n19022), .C2(n19047), .A(n18878), .B(n18877), .ZN(
        P2_U2839) );
  OAI21_X1 U21947 ( .B1(n19750), .B2(n19004), .A(n18974), .ZN(n18881) );
  OAI22_X1 U21948 ( .A1(n19006), .A2(n11010), .B1(n18879), .B2(n18989), .ZN(
        n18880) );
  AOI211_X1 U21949 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18979), .A(
        n18881), .B(n18880), .ZN(n18888) );
  NAND2_X1 U21950 ( .A1(n18994), .A2(n18882), .ZN(n18883) );
  XNOR2_X1 U21951 ( .A(n18884), .B(n18883), .ZN(n18885) );
  AOI22_X1 U21952 ( .A1(n18886), .A2(n18998), .B1(n19000), .B2(n18885), .ZN(
        n18887) );
  OAI211_X1 U21953 ( .C1(n18889), .C2(n19032), .A(n18888), .B(n18887), .ZN(
        P2_U2840) );
  AOI22_X1 U21954 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19038), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19028), .ZN(n18890) );
  OAI21_X1 U21955 ( .B1(n18891), .B2(n18989), .A(n18890), .ZN(n18892) );
  AOI211_X1 U21956 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19027), .A(n18992), 
        .B(n18892), .ZN(n18898) );
  NOR2_X1 U21957 ( .A1(n19016), .A2(n18899), .ZN(n18894) );
  XNOR2_X1 U21958 ( .A(n18894), .B(n18893), .ZN(n18896) );
  AOI22_X1 U21959 ( .A1(n19000), .A2(n18896), .B1(n19008), .B2(n18895), .ZN(
        n18897) );
  OAI211_X1 U21960 ( .C1(n19022), .C2(n19052), .A(n18898), .B(n18897), .ZN(
        P2_U2841) );
  NAND2_X1 U21961 ( .A1(n19000), .A2(n18994), .ZN(n19041) );
  AOI211_X1 U21962 ( .C1(n18906), .C2(n18900), .A(n18899), .B(n19041), .ZN(
        n18903) );
  AOI22_X1 U21963 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19038), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n19028), .ZN(n18901) );
  OAI211_X1 U21964 ( .C1(n14957), .C2(n19004), .A(n18901), .B(n18974), .ZN(
        n18902) );
  AOI211_X1 U21965 ( .C1(n19026), .C2(n18904), .A(n18903), .B(n18902), .ZN(
        n18908) );
  AOI22_X1 U21966 ( .A1(n18906), .A2(n19037), .B1(n18998), .B2(n18905), .ZN(
        n18907) );
  OAI211_X1 U21967 ( .C1(n19032), .C2(n18909), .A(n18908), .B(n18907), .ZN(
        P2_U2842) );
  OR2_X1 U21968 ( .A1(n19016), .A2(n18910), .ZN(n18924) );
  XNOR2_X1 U21969 ( .A(n18924), .B(n18911), .ZN(n18918) );
  INV_X1 U21970 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n19058) );
  AOI22_X1 U21971 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19038), .B1(
        n18912), .B2(n19026), .ZN(n18913) );
  OAI21_X1 U21972 ( .B1(n19006), .B2(n19058), .A(n18913), .ZN(n18914) );
  AOI211_X1 U21973 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19027), .A(n18992), 
        .B(n18914), .ZN(n18917) );
  AOI22_X1 U21974 ( .A1(n19008), .A2(n18915), .B1(n18998), .B2(n19055), .ZN(
        n18916) );
  OAI211_X1 U21975 ( .C1(n19705), .C2(n18918), .A(n18917), .B(n18916), .ZN(
        P2_U2843) );
  AOI22_X1 U21976 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19038), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n19028), .ZN(n18919) );
  OAI211_X1 U21977 ( .C1(n19745), .C2(n19004), .A(n18919), .B(n18974), .ZN(
        n18923) );
  OAI22_X1 U21978 ( .A1(n18921), .A2(n18989), .B1(n19032), .B2(n18920), .ZN(
        n18922) );
  AOI211_X1 U21979 ( .C1(n10153), .C2(n19037), .A(n18923), .B(n18922), .ZN(
        n18928) );
  AOI211_X1 U21980 ( .C1(n18925), .C2(n10153), .A(n19705), .B(n18924), .ZN(
        n18926) );
  INV_X1 U21981 ( .A(n18926), .ZN(n18927) );
  OAI211_X1 U21982 ( .C1(n18929), .C2(n19022), .A(n18928), .B(n18927), .ZN(
        P2_U2844) );
  NOR2_X1 U21983 ( .A1(n19016), .A2(n18930), .ZN(n18931) );
  XOR2_X1 U21984 ( .A(n18932), .B(n18931), .Z(n18940) );
  INV_X1 U21985 ( .A(n18933), .ZN(n18934) );
  AOI22_X1 U21986 ( .A1(n18934), .A2(n19026), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n19028), .ZN(n18935) );
  OAI211_X1 U21987 ( .C1(n10895), .C2(n19004), .A(n18935), .B(n18966), .ZN(
        n18938) );
  OAI22_X1 U21988 ( .A1(n19032), .A2(n18936), .B1(n19022), .B2(n19059), .ZN(
        n18937) );
  AOI211_X1 U21989 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n18979), .A(
        n18938), .B(n18937), .ZN(n18939) );
  OAI21_X1 U21990 ( .B1(n19705), .B2(n18940), .A(n18939), .ZN(P2_U2845) );
  OAI21_X1 U21991 ( .B1(n19742), .B2(n19004), .A(n18974), .ZN(n18943) );
  OAI22_X1 U21992 ( .A1(n18941), .A2(n18989), .B1(n19006), .B2(n10988), .ZN(
        n18942) );
  AOI211_X1 U21993 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18979), .A(
        n18943), .B(n18942), .ZN(n18950) );
  NAND2_X1 U21994 ( .A1(n18994), .A2(n18944), .ZN(n18945) );
  XNOR2_X1 U21995 ( .A(n18946), .B(n18945), .ZN(n18948) );
  AOI22_X1 U21996 ( .A1(n19000), .A2(n18948), .B1(n18998), .B2(n18947), .ZN(
        n18949) );
  OAI211_X1 U21997 ( .C1(n19032), .C2(n18951), .A(n18950), .B(n18949), .ZN(
        P2_U2846) );
  AOI22_X1 U21998 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19038), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19028), .ZN(n18952) );
  OAI21_X1 U21999 ( .B1(n18953), .B2(n18989), .A(n18952), .ZN(n18954) );
  AOI211_X1 U22000 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19027), .A(n18992), .B(
        n18954), .ZN(n18961) );
  NOR2_X1 U22001 ( .A1(n19016), .A2(n18955), .ZN(n18957) );
  XNOR2_X1 U22002 ( .A(n18957), .B(n18956), .ZN(n18959) );
  AOI22_X1 U22003 ( .A1(n19000), .A2(n18959), .B1(n19008), .B2(n18958), .ZN(
        n18960) );
  OAI211_X1 U22004 ( .C1(n19022), .C2(n19079), .A(n18961), .B(n18960), .ZN(
        P2_U2847) );
  NAND2_X1 U22005 ( .A1(n18994), .A2(n18962), .ZN(n18964) );
  XOR2_X1 U22006 ( .A(n18964), .B(n18963), .Z(n18973) );
  AOI22_X1 U22007 ( .A1(P2_EBX_REG_7__SCAN_IN), .A2(n19028), .B1(n18965), .B2(
        n19026), .ZN(n18967) );
  OAI211_X1 U22008 ( .C1(n19739), .C2(n19004), .A(n18967), .B(n18966), .ZN(
        n18971) );
  OAI22_X1 U22009 ( .A1(n19032), .A2(n18969), .B1(n19022), .B2(n18968), .ZN(
        n18970) );
  AOI211_X1 U22010 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18979), .A(
        n18971), .B(n18970), .ZN(n18972) );
  OAI21_X1 U22011 ( .B1(n18973), .B2(n19705), .A(n18972), .ZN(P2_U2848) );
  OAI21_X1 U22012 ( .B1(n19737), .B2(n19004), .A(n18974), .ZN(n18978) );
  OAI22_X1 U22013 ( .A1(n19006), .A2(n18976), .B1(n18975), .B2(n18989), .ZN(
        n18977) );
  AOI211_X1 U22014 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18979), .A(
        n18978), .B(n18977), .ZN(n18986) );
  NOR2_X1 U22015 ( .A1(n19016), .A2(n18980), .ZN(n18982) );
  XNOR2_X1 U22016 ( .A(n18982), .B(n18981), .ZN(n18984) );
  AOI22_X1 U22017 ( .A1(n19000), .A2(n18984), .B1(n18998), .B2(n18983), .ZN(
        n18985) );
  OAI211_X1 U22018 ( .C1(n19032), .C2(n18987), .A(n18986), .B(n18985), .ZN(
        P2_U2849) );
  AOI22_X1 U22019 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19038), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n19028), .ZN(n18988) );
  OAI21_X1 U22020 ( .B1(n18990), .B2(n18989), .A(n18988), .ZN(n18991) );
  AOI211_X1 U22021 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19027), .A(n18992), .B(
        n18991), .ZN(n19002) );
  NAND2_X1 U22022 ( .A1(n18994), .A2(n18993), .ZN(n18995) );
  XNOR2_X1 U22023 ( .A(n18996), .B(n18995), .ZN(n18999) );
  AOI22_X1 U22024 ( .A1(n19000), .A2(n18999), .B1(n18998), .B2(n18997), .ZN(
        n19001) );
  OAI211_X1 U22025 ( .C1(n19032), .C2(n19110), .A(n19002), .B(n19001), .ZN(
        P2_U2850) );
  AOI22_X1 U22026 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19038), .B1(
        n19003), .B2(n19026), .ZN(n19011) );
  OAI22_X1 U22027 ( .A1(n19006), .A2(n19005), .B1(n10972), .B2(n19004), .ZN(
        n19007) );
  AOI211_X1 U22028 ( .C1(n19009), .C2(n19008), .A(n18992), .B(n19007), .ZN(
        n19010) );
  OAI211_X1 U22029 ( .C1(n19080), .C2(n19012), .A(n19011), .B(n19010), .ZN(
        n19013) );
  INV_X1 U22030 ( .A(n19013), .ZN(n19021) );
  INV_X1 U22031 ( .A(n19014), .ZN(n19019) );
  NOR2_X1 U22032 ( .A1(n19016), .A2(n19015), .ZN(n19018) );
  AOI21_X1 U22033 ( .B1(n19019), .B2(n19018), .A(n19705), .ZN(n19017) );
  OAI21_X1 U22034 ( .B1(n19019), .B2(n19018), .A(n19017), .ZN(n19020) );
  OAI211_X1 U22035 ( .C1(n19083), .C2(n19022), .A(n19021), .B(n19020), .ZN(
        P2_U2851) );
  NOR2_X1 U22036 ( .A1(n19023), .A2(n19022), .ZN(n19034) );
  AOI22_X1 U22037 ( .A1(n19027), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19026), 
        .B2(n19025), .ZN(n19030) );
  NAND2_X1 U22038 ( .A1(n19028), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n19029) );
  OAI211_X1 U22039 ( .C1(n19032), .C2(n19031), .A(n19030), .B(n19029), .ZN(
        n19033) );
  AOI211_X1 U22040 ( .C1(n19036), .C2(n19035), .A(n19034), .B(n19033), .ZN(
        n19040) );
  OAI21_X1 U22041 ( .B1(n19038), .B2(n19037), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19039) );
  OAI211_X1 U22042 ( .C1(n19042), .C2(n19041), .A(n19040), .B(n19039), .ZN(
        P2_U2855) );
  AOI21_X1 U22043 ( .B1(n19045), .B2(n19044), .A(n19043), .ZN(n19095) );
  AOI22_X1 U22044 ( .A1(n19095), .A2(n19081), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n19084), .ZN(n19046) );
  OAI21_X1 U22045 ( .B1(n19084), .B2(n19047), .A(n19046), .ZN(P2_U2871) );
  XOR2_X1 U22046 ( .A(n19049), .B(n19048), .Z(n19050) );
  AOI22_X1 U22047 ( .A1(n19050), .A2(n19081), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19084), .ZN(n19051) );
  OAI21_X1 U22048 ( .B1(n19052), .B2(n19084), .A(n19051), .ZN(P2_U2873) );
  XOR2_X1 U22049 ( .A(n19054), .B(n19053), .Z(n19056) );
  AOI22_X1 U22050 ( .A1(n19056), .A2(n19081), .B1(n19070), .B2(n19055), .ZN(
        n19057) );
  OAI21_X1 U22051 ( .B1(n19070), .B2(n19058), .A(n19057), .ZN(P2_U2875) );
  INV_X1 U22052 ( .A(n19059), .ZN(n19067) );
  INV_X1 U22053 ( .A(n19060), .ZN(n19074) );
  AOI21_X1 U22054 ( .B1(n19074), .B2(n19062), .A(n19061), .ZN(n19065) );
  INV_X1 U22055 ( .A(n19063), .ZN(n19064) );
  NOR3_X1 U22056 ( .A1(n19065), .A2(n19064), .A3(n19075), .ZN(n19066) );
  AOI21_X1 U22057 ( .B1(n19067), .B2(n19070), .A(n19066), .ZN(n19068) );
  OAI21_X1 U22058 ( .B1(n19070), .B2(n19069), .A(n19068), .ZN(P2_U2877) );
  INV_X1 U22059 ( .A(n19071), .ZN(n19076) );
  AOI211_X1 U22060 ( .C1(n19076), .C2(n9727), .A(n19075), .B(n19074), .ZN(
        n19077) );
  AOI21_X1 U22061 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19084), .A(n19077), .ZN(
        n19078) );
  OAI21_X1 U22062 ( .B1(n19079), .B2(n19084), .A(n19078), .ZN(P2_U2879) );
  INV_X1 U22063 ( .A(n19080), .ZN(n19106) );
  AOI22_X1 U22064 ( .A1(n19106), .A2(n19081), .B1(P2_EBX_REG_4__SCAN_IN), .B2(
        n19084), .ZN(n19082) );
  OAI21_X1 U22065 ( .B1(n19084), .B2(n19083), .A(n19082), .ZN(P2_U2883) );
  AOI22_X1 U22066 ( .A1(n19086), .A2(n19096), .B1(n19085), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19089) );
  AOI22_X1 U22067 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19102), .B1(n19087), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19088) );
  NAND2_X1 U22068 ( .A1(n19089), .A2(n19088), .ZN(P2_U2888) );
  OAI22_X1 U22069 ( .A1(n19093), .A2(n19092), .B1(n19091), .B2(n19090), .ZN(
        n19094) );
  AOI21_X1 U22070 ( .B1(P2_EAX_REG_16__SCAN_IN), .B2(n19102), .A(n19094), .ZN(
        n19099) );
  AOI22_X1 U22071 ( .A1(n19097), .A2(n19096), .B1(n19105), .B2(n19095), .ZN(
        n19098) );
  OAI211_X1 U22072 ( .C1(n19101), .C2(n19100), .A(n19099), .B(n19098), .ZN(
        P2_U2903) );
  AOI22_X1 U22073 ( .A1(n19104), .A2(n19103), .B1(n19102), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n19109) );
  NAND3_X1 U22074 ( .A1(n19107), .A2(n19106), .A3(n19105), .ZN(n19108) );
  OAI211_X1 U22075 ( .C1(n19111), .C2(n19110), .A(n19109), .B(n19108), .ZN(
        P2_U2914) );
  NOR2_X1 U22076 ( .A1(n19117), .A2(n19112), .ZN(P2_U2920) );
  INV_X1 U22077 ( .A(n19113), .ZN(n19114) );
  AOI22_X1 U22078 ( .A1(n19114), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_UWORD_REG_14__SCAN_IN), .B2(n19148), .ZN(n19115) );
  OAI21_X1 U22079 ( .B1(n19117), .B2(n19116), .A(n19115), .ZN(P2_U2921) );
  AOI22_X1 U22080 ( .A1(n19148), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19118) );
  OAI21_X1 U22081 ( .B1(n12722), .B2(n19150), .A(n19118), .ZN(P2_U2936) );
  AOI22_X1 U22082 ( .A1(n19148), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19119) );
  OAI21_X1 U22083 ( .B1(n19120), .B2(n19150), .A(n19119), .ZN(P2_U2937) );
  AOI22_X1 U22084 ( .A1(n19148), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19121) );
  OAI21_X1 U22085 ( .B1(n19122), .B2(n19150), .A(n19121), .ZN(P2_U2938) );
  AOI22_X1 U22086 ( .A1(n19148), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19123) );
  OAI21_X1 U22087 ( .B1(n19124), .B2(n19150), .A(n19123), .ZN(P2_U2939) );
  AOI22_X1 U22088 ( .A1(n19148), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19125) );
  OAI21_X1 U22089 ( .B1(n19126), .B2(n19150), .A(n19125), .ZN(P2_U2940) );
  AOI22_X1 U22090 ( .A1(n19148), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19127) );
  OAI21_X1 U22091 ( .B1(n19128), .B2(n19150), .A(n19127), .ZN(P2_U2941) );
  AOI22_X1 U22092 ( .A1(n19148), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19129) );
  OAI21_X1 U22093 ( .B1(n19130), .B2(n19150), .A(n19129), .ZN(P2_U2942) );
  AOI22_X1 U22094 ( .A1(n19148), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19131) );
  OAI21_X1 U22095 ( .B1(n19132), .B2(n19150), .A(n19131), .ZN(P2_U2943) );
  AOI22_X1 U22096 ( .A1(n19148), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19133) );
  OAI21_X1 U22097 ( .B1(n19134), .B2(n19150), .A(n19133), .ZN(P2_U2944) );
  AOI22_X1 U22098 ( .A1(n19148), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19135) );
  OAI21_X1 U22099 ( .B1(n19136), .B2(n19150), .A(n19135), .ZN(P2_U2945) );
  INV_X1 U22100 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19138) );
  AOI22_X1 U22101 ( .A1(n19148), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19137) );
  OAI21_X1 U22102 ( .B1(n19138), .B2(n19150), .A(n19137), .ZN(P2_U2946) );
  INV_X1 U22103 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19140) );
  AOI22_X1 U22104 ( .A1(n19148), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19139) );
  OAI21_X1 U22105 ( .B1(n19140), .B2(n19150), .A(n19139), .ZN(P2_U2947) );
  INV_X1 U22106 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19142) );
  AOI22_X1 U22107 ( .A1(n19148), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19141) );
  OAI21_X1 U22108 ( .B1(n19142), .B2(n19150), .A(n19141), .ZN(P2_U2948) );
  AOI22_X1 U22109 ( .A1(n19148), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19143) );
  OAI21_X1 U22110 ( .B1(n19144), .B2(n19150), .A(n19143), .ZN(P2_U2949) );
  INV_X1 U22111 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19146) );
  AOI22_X1 U22112 ( .A1(n19148), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19145) );
  OAI21_X1 U22113 ( .B1(n19146), .B2(n19150), .A(n19145), .ZN(P2_U2950) );
  INV_X1 U22114 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19151) );
  AOI22_X1 U22115 ( .A1(n19148), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19147), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19149) );
  OAI21_X1 U22116 ( .B1(n19151), .B2(n19150), .A(n19149), .ZN(P2_U2951) );
  AOI22_X1 U22117 ( .A1(n19153), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19152), .B2(n19819), .ZN(n19167) );
  INV_X1 U22118 ( .A(n19154), .ZN(n19156) );
  OAI22_X1 U22119 ( .A1(n19158), .A2(n19157), .B1(n19156), .B2(n19155), .ZN(
        n19159) );
  AOI211_X1 U22120 ( .C1(n19162), .C2(n19161), .A(n19160), .B(n19159), .ZN(
        n19166) );
  OAI211_X1 U22121 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n19164), .B(n19163), .ZN(n19165) );
  NAND3_X1 U22122 ( .A1(n19167), .A2(n19166), .A3(n19165), .ZN(P2_U3045) );
  AOI22_X1 U22123 ( .A1(n19693), .A2(n19629), .B1(n19190), .B2(n19628), .ZN(
        n19169) );
  AOI22_X1 U22124 ( .A1(n13567), .A2(n19195), .B1(n19194), .B2(n19630), .ZN(
        n19168) );
  OAI211_X1 U22125 ( .C1(n19199), .C2(n19170), .A(n19169), .B(n19168), .ZN(
        P2_U3050) );
  AOI22_X1 U22126 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19193), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19192), .ZN(n19607) );
  INV_X1 U22127 ( .A(n19607), .ZN(n19665) );
  NAND2_X1 U22128 ( .A1(n19172), .A2(n19171), .ZN(n19661) );
  INV_X1 U22129 ( .A(n19661), .ZN(n19634) );
  AOI22_X1 U22130 ( .A1(n19693), .A2(n19665), .B1(n19190), .B2(n19634), .ZN(
        n19175) );
  NOR2_X2 U22131 ( .A1(n19173), .A2(n19285), .ZN(n19659) );
  AOI22_X1 U22132 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19193), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19192), .ZN(n19533) );
  INV_X1 U22133 ( .A(n19533), .ZN(n19664) );
  AOI22_X1 U22134 ( .A1(n19659), .A2(n19195), .B1(n19194), .B2(n19664), .ZN(
        n19174) );
  OAI211_X1 U22135 ( .C1(n19199), .C2(n19176), .A(n19175), .B(n19174), .ZN(
        P2_U3051) );
  AOI22_X1 U22136 ( .A1(n19693), .A2(n19672), .B1(n19670), .B2(n19190), .ZN(
        n19178) );
  AOI22_X1 U22137 ( .A1(n19671), .A2(n19195), .B1(n19194), .B2(n19673), .ZN(
        n19177) );
  OAI211_X1 U22138 ( .C1(n19199), .C2(n19179), .A(n19178), .B(n19177), .ZN(
        P2_U3052) );
  AOI22_X1 U22139 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19192), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19193), .ZN(n19613) );
  INV_X1 U22140 ( .A(n19613), .ZN(n19679) );
  NOR2_X2 U22141 ( .A1(n19189), .A2(n10302), .ZN(n19676) );
  AOI22_X1 U22142 ( .A1(n19693), .A2(n19679), .B1(n19190), .B2(n19676), .ZN(
        n19183) );
  NOR2_X2 U22143 ( .A1(n19181), .A2(n19285), .ZN(n19677) );
  AOI22_X1 U22144 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19193), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19192), .ZN(n19539) );
  INV_X1 U22145 ( .A(n19539), .ZN(n19678) );
  AOI22_X1 U22146 ( .A1(n19677), .A2(n19195), .B1(n19194), .B2(n19678), .ZN(
        n19182) );
  OAI211_X1 U22147 ( .C1(n19199), .C2(n13121), .A(n19183), .B(n19182), .ZN(
        P2_U3053) );
  OAI22_X1 U22148 ( .A1(n19187), .A2(n19186), .B1(n19185), .B2(n19184), .ZN(
        n19684) );
  NOR2_X2 U22149 ( .A1(n19189), .A2(n19188), .ZN(n19682) );
  AOI22_X1 U22150 ( .A1(n19693), .A2(n19684), .B1(n19190), .B2(n19682), .ZN(
        n19197) );
  NOR2_X2 U22151 ( .A1(n19191), .A2(n19285), .ZN(n19683) );
  AOI22_X1 U22152 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19193), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19192), .ZN(n19542) );
  AOI22_X1 U22153 ( .A1(n19683), .A2(n19195), .B1(n19194), .B2(n19685), .ZN(
        n19196) );
  OAI211_X1 U22154 ( .C1(n19199), .C2(n19198), .A(n19197), .B(n19196), .ZN(
        P2_U3054) );
  OR2_X1 U22155 ( .A1(n19245), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19202) );
  NOR3_X2 U22156 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19830), .A3(
        n19245), .ZN(n19220) );
  INV_X1 U22157 ( .A(n19203), .ZN(n19201) );
  AOI211_X2 U22158 ( .C1(n19202), .C2(n19843), .A(n19378), .B(n19201), .ZN(
        n19221) );
  AOI22_X1 U22159 ( .A1(n19221), .A2(n13539), .B1(n19586), .B2(n19220), .ZN(
        n19207) );
  NOR4_X1 U22160 ( .A1(n19803), .A2(n19442), .A3(P2_STATE2_REG_3__SCAN_IN), 
        .A4(n19797), .ZN(n19205) );
  NOR2_X1 U22161 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19587), .ZN(
        n19827) );
  NOR3_X1 U22162 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19827), .A3(
        n19245), .ZN(n19204) );
  OAI211_X1 U22163 ( .C1(n19205), .C2(n19204), .A(n19593), .B(n19203), .ZN(
        n19222) );
  AOI22_X1 U22164 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19222), .B1(
        n19240), .B2(n19595), .ZN(n19206) );
  OAI211_X1 U22165 ( .C1(n19598), .C2(n19225), .A(n19207), .B(n19206), .ZN(
        P2_U3056) );
  INV_X1 U22166 ( .A(n19651), .ZN(n19624) );
  AOI22_X1 U22167 ( .A1(n19221), .A2(n15341), .B1(n19624), .B2(n19220), .ZN(
        n19209) );
  AOI22_X1 U22168 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19222), .B1(
        n19240), .B2(n19655), .ZN(n19208) );
  OAI211_X1 U22169 ( .C1(n19601), .C2(n19225), .A(n19209), .B(n19208), .ZN(
        P2_U3057) );
  AOI22_X1 U22170 ( .A1(n19221), .A2(n13567), .B1(n19628), .B2(n19220), .ZN(
        n19211) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19222), .B1(
        n19240), .B2(n19630), .ZN(n19210) );
  OAI211_X1 U22172 ( .C1(n19604), .C2(n19225), .A(n19211), .B(n19210), .ZN(
        P2_U3058) );
  AOI22_X1 U22173 ( .A1(n19221), .A2(n19659), .B1(n19634), .B2(n19220), .ZN(
        n19213) );
  AOI22_X1 U22174 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19222), .B1(
        n19240), .B2(n19664), .ZN(n19212) );
  OAI211_X1 U22175 ( .C1(n19607), .C2(n19225), .A(n19213), .B(n19212), .ZN(
        P2_U3059) );
  AOI22_X1 U22176 ( .A1(n19221), .A2(n19671), .B1(n19670), .B2(n19220), .ZN(
        n19215) );
  AOI22_X1 U22177 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19222), .B1(
        n19240), .B2(n19673), .ZN(n19214) );
  OAI211_X1 U22178 ( .C1(n19610), .C2(n19225), .A(n19215), .B(n19214), .ZN(
        P2_U3060) );
  AOI22_X1 U22179 ( .A1(n19221), .A2(n19677), .B1(n19676), .B2(n19220), .ZN(
        n19217) );
  AOI22_X1 U22180 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19222), .B1(
        n19240), .B2(n19678), .ZN(n19216) );
  OAI211_X1 U22181 ( .C1(n19613), .C2(n19225), .A(n19217), .B(n19216), .ZN(
        P2_U3061) );
  AOI22_X1 U22182 ( .A1(n19221), .A2(n19683), .B1(n19682), .B2(n19220), .ZN(
        n19219) );
  AOI22_X1 U22183 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19222), .B1(
        n19240), .B2(n19685), .ZN(n19218) );
  OAI211_X1 U22184 ( .C1(n19616), .C2(n19225), .A(n19219), .B(n19218), .ZN(
        P2_U3062) );
  AOI22_X1 U22185 ( .A1(n19221), .A2(n19690), .B1(n19688), .B2(n19220), .ZN(
        n19224) );
  AOI22_X1 U22186 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19222), .B1(
        n19240), .B2(n19692), .ZN(n19223) );
  OAI211_X1 U22187 ( .C1(n19623), .C2(n19225), .A(n19224), .B(n19223), .ZN(
        P2_U3063) );
  AOI22_X1 U22188 ( .A1(n19239), .A2(n13539), .B1(n19238), .B2(n19586), .ZN(
        n19227) );
  AOI22_X1 U22189 ( .A1(n19255), .A2(n19595), .B1(n19240), .B2(n19521), .ZN(
        n19226) );
  OAI211_X1 U22190 ( .C1(n19243), .C2(n19228), .A(n19227), .B(n19226), .ZN(
        P2_U3064) );
  AOI22_X1 U22191 ( .A1(n19239), .A2(n15341), .B1(n19238), .B2(n19624), .ZN(
        n19230) );
  AOI22_X1 U22192 ( .A1(n19255), .A2(n19655), .B1(n19240), .B2(n19654), .ZN(
        n19229) );
  OAI211_X1 U22193 ( .C1(n19243), .C2(n10507), .A(n19230), .B(n19229), .ZN(
        P2_U3065) );
  INV_X1 U22194 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n19233) );
  AOI22_X1 U22195 ( .A1(n19239), .A2(n13567), .B1(n19238), .B2(n19628), .ZN(
        n19232) );
  AOI22_X1 U22196 ( .A1(n19255), .A2(n19630), .B1(n19240), .B2(n19629), .ZN(
        n19231) );
  OAI211_X1 U22197 ( .C1(n19243), .C2(n19233), .A(n19232), .B(n19231), .ZN(
        P2_U3066) );
  AOI22_X1 U22198 ( .A1(n19239), .A2(n19659), .B1(n19238), .B2(n19634), .ZN(
        n19235) );
  AOI22_X1 U22199 ( .A1(n19240), .A2(n19665), .B1(n19255), .B2(n19664), .ZN(
        n19234) );
  OAI211_X1 U22200 ( .C1(n19243), .C2(n10480), .A(n19235), .B(n19234), .ZN(
        P2_U3067) );
  AOI22_X1 U22201 ( .A1(n19239), .A2(n19677), .B1(n19238), .B2(n19676), .ZN(
        n19237) );
  AOI22_X1 U22202 ( .A1(n19240), .A2(n19679), .B1(n19255), .B2(n19678), .ZN(
        n19236) );
  OAI211_X1 U22203 ( .C1(n19243), .C2(n10596), .A(n19237), .B(n19236), .ZN(
        P2_U3069) );
  AOI22_X1 U22204 ( .A1(n19239), .A2(n19683), .B1(n19238), .B2(n19682), .ZN(
        n19242) );
  AOI22_X1 U22205 ( .A1(n19255), .A2(n19685), .B1(n19240), .B2(n19684), .ZN(
        n19241) );
  OAI211_X1 U22206 ( .C1(n19243), .C2(n10632), .A(n19242), .B(n19241), .ZN(
        P2_U3070) );
  NOR2_X1 U22207 ( .A1(n19511), .A2(n19245), .ZN(n19270) );
  AOI22_X1 U22208 ( .A1(n19521), .A2(n19255), .B1(n19586), .B2(n19270), .ZN(
        n19254) );
  AOI21_X1 U22209 ( .B1(n19249), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19247) );
  NAND3_X1 U22210 ( .A1(n19791), .A2(n19482), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19244) );
  NAND2_X1 U22211 ( .A1(n19244), .A2(n19806), .ZN(n19252) );
  NOR2_X1 U22212 ( .A1(n19821), .A2(n19245), .ZN(n19248) );
  OR2_X1 U22213 ( .A1(n19252), .A2(n19248), .ZN(n19246) );
  OAI211_X1 U22214 ( .C1(n19270), .C2(n19247), .A(n19246), .B(n19593), .ZN(
        n19277) );
  INV_X1 U22215 ( .A(n19248), .ZN(n19251) );
  OAI21_X1 U22216 ( .B1(n9752), .B2(n19270), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19250) );
  OAI21_X1 U22217 ( .B1(n19252), .B2(n19251), .A(n19250), .ZN(n19276) );
  AOI22_X1 U22218 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19277), .B1(
        n13539), .B2(n19276), .ZN(n19253) );
  OAI211_X1 U22219 ( .C1(n19524), .C2(n19318), .A(n19254), .B(n19253), .ZN(
        P2_U3072) );
  AOI22_X1 U22220 ( .A1(n19654), .A2(n19255), .B1(n19624), .B2(n19270), .ZN(
        n19257) );
  AOI22_X1 U22221 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19277), .B1(
        n15341), .B2(n19276), .ZN(n19256) );
  OAI211_X1 U22222 ( .C1(n19527), .C2(n19318), .A(n19257), .B(n19256), .ZN(
        P2_U3073) );
  INV_X1 U22223 ( .A(n19270), .ZN(n19273) );
  INV_X1 U22224 ( .A(n19628), .ZN(n19333) );
  OAI22_X1 U22225 ( .A1(n19274), .A2(n19604), .B1(n19273), .B2(n19333), .ZN(
        n19258) );
  INV_X1 U22226 ( .A(n19258), .ZN(n19260) );
  AOI22_X1 U22227 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19277), .B1(
        n13567), .B2(n19276), .ZN(n19259) );
  OAI211_X1 U22228 ( .C1(n19530), .C2(n19318), .A(n19260), .B(n19259), .ZN(
        P2_U3074) );
  OAI22_X1 U22229 ( .A1(n19318), .A2(n19533), .B1(n19273), .B2(n19661), .ZN(
        n19261) );
  INV_X1 U22230 ( .A(n19261), .ZN(n19263) );
  AOI22_X1 U22231 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19277), .B1(
        n19659), .B2(n19276), .ZN(n19262) );
  OAI211_X1 U22232 ( .C1(n19607), .C2(n19274), .A(n19263), .B(n19262), .ZN(
        P2_U3075) );
  INV_X1 U22233 ( .A(n19670), .ZN(n19461) );
  OAI22_X1 U22234 ( .A1(n19274), .A2(n19610), .B1(n19461), .B2(n19273), .ZN(
        n19264) );
  INV_X1 U22235 ( .A(n19264), .ZN(n19266) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19277), .B1(
        n19671), .B2(n19276), .ZN(n19265) );
  OAI211_X1 U22237 ( .C1(n19536), .C2(n19318), .A(n19266), .B(n19265), .ZN(
        P2_U3076) );
  INV_X1 U22238 ( .A(n19676), .ZN(n19427) );
  OAI22_X1 U22239 ( .A1(n19274), .A2(n19613), .B1(n19273), .B2(n19427), .ZN(
        n19267) );
  INV_X1 U22240 ( .A(n19267), .ZN(n19269) );
  AOI22_X1 U22241 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19277), .B1(
        n19677), .B2(n19276), .ZN(n19268) );
  OAI211_X1 U22242 ( .C1(n19539), .C2(n19318), .A(n19269), .B(n19268), .ZN(
        P2_U3077) );
  INV_X1 U22243 ( .A(n19318), .ZN(n19281) );
  AOI22_X1 U22244 ( .A1(n19685), .A2(n19281), .B1(n19682), .B2(n19270), .ZN(
        n19272) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19277), .B1(
        n19683), .B2(n19276), .ZN(n19271) );
  OAI211_X1 U22246 ( .C1(n19616), .C2(n19274), .A(n19272), .B(n19271), .ZN(
        P2_U3078) );
  OAI22_X1 U22247 ( .A1(n19274), .A2(n19623), .B1(n19472), .B2(n19273), .ZN(
        n19275) );
  INV_X1 U22248 ( .A(n19275), .ZN(n19279) );
  AOI22_X1 U22249 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19277), .B1(
        n19690), .B2(n19276), .ZN(n19278) );
  OAI211_X1 U22250 ( .C1(n19549), .C2(n19318), .A(n19279), .B(n19278), .ZN(
        P2_U3079) );
  NOR2_X1 U22251 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19326), .ZN(
        n19309) );
  AOI22_X1 U22252 ( .A1(n19595), .A2(n19330), .B1(n19586), .B2(n19309), .ZN(
        n19294) );
  NOR2_X1 U22253 ( .A1(n19330), .A2(n19281), .ZN(n19282) );
  OAI21_X1 U22254 ( .B1(n19282), .B2(n19797), .A(n19806), .ZN(n19292) );
  NAND2_X1 U22255 ( .A1(n19284), .A2(n19283), .ZN(n19550) );
  NOR2_X1 U22256 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19550), .ZN(
        n19288) );
  OAI21_X1 U22257 ( .B1(n19289), .B2(n19843), .A(n19587), .ZN(n19286) );
  INV_X1 U22258 ( .A(n19309), .ZN(n19312) );
  AOI21_X1 U22259 ( .B1(n19286), .B2(n19312), .A(n19285), .ZN(n19287) );
  INV_X1 U22260 ( .A(n19288), .ZN(n19291) );
  OAI21_X1 U22261 ( .B1(n19289), .B2(n19309), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19290) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19315), .B1(
        n13539), .B2(n19314), .ZN(n19293) );
  OAI211_X1 U22263 ( .C1(n19598), .C2(n19318), .A(n19294), .B(n19293), .ZN(
        P2_U3080) );
  OAI22_X1 U22264 ( .A1(n19355), .A2(n19527), .B1(n19312), .B2(n19651), .ZN(
        n19295) );
  INV_X1 U22265 ( .A(n19295), .ZN(n19297) );
  AOI22_X1 U22266 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19315), .B1(
        n15341), .B2(n19314), .ZN(n19296) );
  OAI211_X1 U22267 ( .C1(n19601), .C2(n19318), .A(n19297), .B(n19296), .ZN(
        P2_U3081) );
  OAI22_X1 U22268 ( .A1(n19318), .A2(n19604), .B1(n19312), .B2(n19333), .ZN(
        n19298) );
  INV_X1 U22269 ( .A(n19298), .ZN(n19300) );
  AOI22_X1 U22270 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19315), .B1(
        n13567), .B2(n19314), .ZN(n19299) );
  OAI211_X1 U22271 ( .C1(n19530), .C2(n19355), .A(n19300), .B(n19299), .ZN(
        P2_U3082) );
  OAI22_X1 U22272 ( .A1(n19318), .A2(n19607), .B1(n19312), .B2(n19661), .ZN(
        n19301) );
  INV_X1 U22273 ( .A(n19301), .ZN(n19303) );
  AOI22_X1 U22274 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19315), .B1(
        n19659), .B2(n19314), .ZN(n19302) );
  OAI211_X1 U22275 ( .C1(n19533), .C2(n19355), .A(n19303), .B(n19302), .ZN(
        P2_U3083) );
  AOI22_X1 U22276 ( .A1(n19673), .A2(n19330), .B1(n19670), .B2(n19309), .ZN(
        n19305) );
  AOI22_X1 U22277 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19315), .B1(
        n19671), .B2(n19314), .ZN(n19304) );
  OAI211_X1 U22278 ( .C1(n19610), .C2(n19318), .A(n19305), .B(n19304), .ZN(
        P2_U3084) );
  OAI22_X1 U22279 ( .A1(n19355), .A2(n19539), .B1(n19312), .B2(n19427), .ZN(
        n19306) );
  INV_X1 U22280 ( .A(n19306), .ZN(n19308) );
  AOI22_X1 U22281 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19315), .B1(
        n19677), .B2(n19314), .ZN(n19307) );
  OAI211_X1 U22282 ( .C1(n19613), .C2(n19318), .A(n19308), .B(n19307), .ZN(
        P2_U3085) );
  AOI22_X1 U22283 ( .A1(n19685), .A2(n19330), .B1(n19309), .B2(n19682), .ZN(
        n19311) );
  AOI22_X1 U22284 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19315), .B1(
        n19683), .B2(n19314), .ZN(n19310) );
  OAI211_X1 U22285 ( .C1(n19616), .C2(n19318), .A(n19311), .B(n19310), .ZN(
        P2_U3086) );
  OAI22_X1 U22286 ( .A1(n19355), .A2(n19549), .B1(n19472), .B2(n19312), .ZN(
        n19313) );
  INV_X1 U22287 ( .A(n19313), .ZN(n19317) );
  AOI22_X1 U22288 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19315), .B1(
        n19690), .B2(n19314), .ZN(n19316) );
  OAI211_X1 U22289 ( .C1(n19623), .C2(n19318), .A(n19317), .B(n19316), .ZN(
        P2_U3087) );
  AOI22_X1 U22290 ( .A1(n19595), .A2(n19371), .B1(n19586), .B2(n19346), .ZN(
        n19329) );
  AOI21_X1 U22291 ( .B1(n19319), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19323) );
  NAND3_X1 U22292 ( .A1(n19791), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19588), 
        .ZN(n19320) );
  NAND2_X1 U22293 ( .A1(n19320), .A2(n19806), .ZN(n19327) );
  OR2_X1 U22294 ( .A1(n19327), .A2(n19321), .ZN(n19322) );
  OAI211_X1 U22295 ( .C1(n19346), .C2(n19323), .A(n19322), .B(n19593), .ZN(
        n19352) );
  OAI21_X1 U22296 ( .B1(n19324), .B2(n19346), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19325) );
  OAI21_X1 U22297 ( .B1(n19327), .B2(n19326), .A(n19325), .ZN(n19351) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19352), .B1(
        n13539), .B2(n19351), .ZN(n19328) );
  OAI211_X1 U22299 ( .C1(n19598), .C2(n19355), .A(n19329), .B(n19328), .ZN(
        P2_U3088) );
  AOI22_X1 U22300 ( .A1(n19654), .A2(n19330), .B1(n19624), .B2(n19346), .ZN(
        n19332) );
  AOI22_X1 U22301 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19352), .B1(
        n15341), .B2(n19351), .ZN(n19331) );
  OAI211_X1 U22302 ( .C1(n19527), .C2(n19368), .A(n19332), .B(n19331), .ZN(
        P2_U3089) );
  INV_X1 U22303 ( .A(n19346), .ZN(n19349) );
  OAI22_X1 U22304 ( .A1(n19355), .A2(n19604), .B1(n19349), .B2(n19333), .ZN(
        n19334) );
  INV_X1 U22305 ( .A(n19334), .ZN(n19336) );
  AOI22_X1 U22306 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19352), .B1(
        n13567), .B2(n19351), .ZN(n19335) );
  OAI211_X1 U22307 ( .C1(n19530), .C2(n19368), .A(n19336), .B(n19335), .ZN(
        P2_U3090) );
  OAI22_X1 U22308 ( .A1(n19368), .A2(n19533), .B1(n19349), .B2(n19661), .ZN(
        n19337) );
  INV_X1 U22309 ( .A(n19337), .ZN(n19339) );
  AOI22_X1 U22310 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19352), .B1(
        n19659), .B2(n19351), .ZN(n19338) );
  OAI211_X1 U22311 ( .C1(n19607), .C2(n19355), .A(n19339), .B(n19338), .ZN(
        P2_U3091) );
  OAI22_X1 U22312 ( .A1(n19355), .A2(n19610), .B1(n19461), .B2(n19349), .ZN(
        n19340) );
  INV_X1 U22313 ( .A(n19340), .ZN(n19342) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19352), .B1(
        n19671), .B2(n19351), .ZN(n19341) );
  OAI211_X1 U22315 ( .C1(n19536), .C2(n19368), .A(n19342), .B(n19341), .ZN(
        P2_U3092) );
  OAI22_X1 U22316 ( .A1(n19368), .A2(n19539), .B1(n19349), .B2(n19427), .ZN(
        n19343) );
  INV_X1 U22317 ( .A(n19343), .ZN(n19345) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19352), .B1(
        n19677), .B2(n19351), .ZN(n19344) );
  OAI211_X1 U22319 ( .C1(n19613), .C2(n19355), .A(n19345), .B(n19344), .ZN(
        P2_U3093) );
  AOI22_X1 U22320 ( .A1(n19685), .A2(n19371), .B1(n19346), .B2(n19682), .ZN(
        n19348) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19352), .B1(
        n19683), .B2(n19351), .ZN(n19347) );
  OAI211_X1 U22322 ( .C1(n19616), .C2(n19355), .A(n19348), .B(n19347), .ZN(
        P2_U3094) );
  OAI22_X1 U22323 ( .A1(n19368), .A2(n19549), .B1(n19472), .B2(n19349), .ZN(
        n19350) );
  INV_X1 U22324 ( .A(n19350), .ZN(n19354) );
  AOI22_X1 U22325 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19352), .B1(
        n19690), .B2(n19351), .ZN(n19353) );
  OAI211_X1 U22326 ( .C1(n19623), .C2(n19355), .A(n19354), .B(n19353), .ZN(
        P2_U3095) );
  AOI22_X1 U22327 ( .A1(n19370), .A2(n15341), .B1(n19369), .B2(n19624), .ZN(
        n19357) );
  AOI22_X1 U22328 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19372), .B1(
        n19401), .B2(n19655), .ZN(n19356) );
  OAI211_X1 U22329 ( .C1(n19601), .C2(n19368), .A(n19357), .B(n19356), .ZN(
        P2_U3097) );
  AOI22_X1 U22330 ( .A1(n19370), .A2(n13567), .B1(n19369), .B2(n19628), .ZN(
        n19359) );
  AOI22_X1 U22331 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19372), .B1(
        n19401), .B2(n19630), .ZN(n19358) );
  OAI211_X1 U22332 ( .C1(n19604), .C2(n19368), .A(n19359), .B(n19358), .ZN(
        P2_U3098) );
  AOI22_X1 U22333 ( .A1(n19370), .A2(n19659), .B1(n19369), .B2(n19634), .ZN(
        n19361) );
  AOI22_X1 U22334 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19372), .B1(
        n19401), .B2(n19664), .ZN(n19360) );
  OAI211_X1 U22335 ( .C1(n19607), .C2(n19368), .A(n19361), .B(n19360), .ZN(
        P2_U3099) );
  AOI22_X1 U22336 ( .A1(n19370), .A2(n19671), .B1(n19670), .B2(n19369), .ZN(
        n19363) );
  AOI22_X1 U22337 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19372), .B1(
        n19401), .B2(n19673), .ZN(n19362) );
  OAI211_X1 U22338 ( .C1(n19610), .C2(n19368), .A(n19363), .B(n19362), .ZN(
        P2_U3100) );
  AOI22_X1 U22339 ( .A1(n19370), .A2(n19677), .B1(n19369), .B2(n19676), .ZN(
        n19365) );
  AOI22_X1 U22340 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19372), .B1(
        n19371), .B2(n19679), .ZN(n19364) );
  OAI211_X1 U22341 ( .C1(n19539), .C2(n19397), .A(n19365), .B(n19364), .ZN(
        P2_U3101) );
  AOI22_X1 U22342 ( .A1(n19370), .A2(n19683), .B1(n19369), .B2(n19682), .ZN(
        n19367) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19372), .B1(
        n19401), .B2(n19685), .ZN(n19366) );
  OAI211_X1 U22344 ( .C1(n19616), .C2(n19368), .A(n19367), .B(n19366), .ZN(
        P2_U3102) );
  AOI22_X1 U22345 ( .A1(n19370), .A2(n19690), .B1(n19688), .B2(n19369), .ZN(
        n19374) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19372), .B1(
        n19371), .B2(n19694), .ZN(n19373) );
  OAI211_X1 U22347 ( .C1(n19549), .C2(n19397), .A(n19374), .B(n19373), .ZN(
        P2_U3103) );
  NOR2_X1 U22348 ( .A1(n19830), .A2(n19379), .ZN(n19411) );
  INV_X1 U22349 ( .A(n19411), .ZN(n19408) );
  AND2_X1 U22350 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19408), .ZN(n19376) );
  AOI211_X2 U22351 ( .C1(n19379), .C2(n19843), .A(n19378), .B(n19380), .ZN(
        n19400) );
  AOI22_X1 U22352 ( .A1(n19400), .A2(n13539), .B1(n19586), .B2(n19411), .ZN(
        n19385) );
  NOR3_X1 U22353 ( .A1(n19803), .A2(n19797), .A3(n19796), .ZN(n19801) );
  OAI21_X1 U22354 ( .B1(n19587), .B2(n19411), .A(n19593), .ZN(n19381) );
  NOR2_X1 U22355 ( .A1(n19381), .A2(n19380), .ZN(n19382) );
  OAI21_X1 U22356 ( .B1(n19383), .B2(n19801), .A(n19382), .ZN(n19402) );
  AOI22_X1 U22357 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19521), .ZN(n19384) );
  OAI211_X1 U22358 ( .C1(n19524), .C2(n19436), .A(n19385), .B(n19384), .ZN(
        P2_U3104) );
  AOI22_X1 U22359 ( .A1(n19400), .A2(n15341), .B1(n19624), .B2(n19411), .ZN(
        n19387) );
  INV_X1 U22360 ( .A(n19436), .ZN(n19394) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19402), .B1(
        n19394), .B2(n19655), .ZN(n19386) );
  OAI211_X1 U22362 ( .C1(n19601), .C2(n19397), .A(n19387), .B(n19386), .ZN(
        P2_U3105) );
  AOI22_X1 U22363 ( .A1(n19400), .A2(n13567), .B1(n19628), .B2(n19411), .ZN(
        n19389) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19402), .B1(
        n19394), .B2(n19630), .ZN(n19388) );
  OAI211_X1 U22365 ( .C1(n19604), .C2(n19397), .A(n19389), .B(n19388), .ZN(
        P2_U3106) );
  AOI22_X1 U22366 ( .A1(n19400), .A2(n19659), .B1(n19634), .B2(n19411), .ZN(
        n19391) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19665), .ZN(n19390) );
  OAI211_X1 U22368 ( .C1(n19533), .C2(n19436), .A(n19391), .B(n19390), .ZN(
        P2_U3107) );
  AOI22_X1 U22369 ( .A1(n19400), .A2(n19671), .B1(n19670), .B2(n19411), .ZN(
        n19393) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19672), .ZN(n19392) );
  OAI211_X1 U22371 ( .C1(n19536), .C2(n19436), .A(n19393), .B(n19392), .ZN(
        P2_U3108) );
  AOI22_X1 U22372 ( .A1(n19400), .A2(n19677), .B1(n19676), .B2(n19411), .ZN(
        n19396) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19402), .B1(
        n19394), .B2(n19678), .ZN(n19395) );
  OAI211_X1 U22374 ( .C1(n19613), .C2(n19397), .A(n19396), .B(n19395), .ZN(
        P2_U3109) );
  AOI22_X1 U22375 ( .A1(n19400), .A2(n19683), .B1(n19682), .B2(n19411), .ZN(
        n19399) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19684), .ZN(n19398) );
  OAI211_X1 U22377 ( .C1(n19542), .C2(n19436), .A(n19399), .B(n19398), .ZN(
        P2_U3110) );
  AOI22_X1 U22378 ( .A1(n19400), .A2(n19690), .B1(n19688), .B2(n19411), .ZN(
        n19404) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19694), .ZN(n19403) );
  OAI211_X1 U22380 ( .C1(n19549), .C2(n19436), .A(n19404), .B(n19403), .ZN(
        P2_U3111) );
  INV_X1 U22381 ( .A(n19442), .ZN(n19444) );
  INV_X1 U22382 ( .A(n19473), .ZN(n19432) );
  NAND2_X1 U22383 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19813), .ZN(
        n19517) );
  NOR2_X1 U22384 ( .A1(n19405), .A2(n19517), .ZN(n19431) );
  AOI22_X1 U22385 ( .A1(n19595), .A2(n19432), .B1(n19586), .B2(n19431), .ZN(
        n19416) );
  AOI21_X1 U22386 ( .B1(n19473), .B2(n19436), .A(n19797), .ZN(n19406) );
  INV_X1 U22387 ( .A(n19806), .ZN(n19556) );
  NOR2_X1 U22388 ( .A1(n19406), .A2(n19556), .ZN(n19410) );
  OAI21_X1 U22389 ( .B1(n19412), .B2(n19843), .A(n19587), .ZN(n19407) );
  AOI21_X1 U22390 ( .B1(n19410), .B2(n19408), .A(n19407), .ZN(n19409) );
  OAI21_X1 U22391 ( .B1(n19431), .B2(n19409), .A(n19593), .ZN(n19439) );
  OAI21_X1 U22392 ( .B1(n19431), .B2(n19411), .A(n19410), .ZN(n19414) );
  OAI21_X1 U22393 ( .B1(n19412), .B2(n19431), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19413) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19439), .B1(
        n13539), .B2(n19438), .ZN(n19415) );
  OAI211_X1 U22395 ( .C1(n19598), .C2(n19436), .A(n19416), .B(n19415), .ZN(
        P2_U3112) );
  INV_X1 U22396 ( .A(n19431), .ZN(n19435) );
  OAI22_X1 U22397 ( .A1(n19473), .A2(n19527), .B1(n19435), .B2(n19651), .ZN(
        n19417) );
  INV_X1 U22398 ( .A(n19417), .ZN(n19419) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19439), .B1(
        n15341), .B2(n19438), .ZN(n19418) );
  OAI211_X1 U22400 ( .C1(n19601), .C2(n19436), .A(n19419), .B(n19418), .ZN(
        P2_U3113) );
  AOI22_X1 U22401 ( .A1(n19630), .A2(n19432), .B1(n19628), .B2(n19431), .ZN(
        n19421) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19439), .B1(
        n13567), .B2(n19438), .ZN(n19420) );
  OAI211_X1 U22403 ( .C1(n19604), .C2(n19436), .A(n19421), .B(n19420), .ZN(
        P2_U3114) );
  OAI22_X1 U22404 ( .A1(n19436), .A2(n19607), .B1(n19435), .B2(n19661), .ZN(
        n19422) );
  INV_X1 U22405 ( .A(n19422), .ZN(n19424) );
  AOI22_X1 U22406 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19439), .B1(
        n19659), .B2(n19438), .ZN(n19423) );
  OAI211_X1 U22407 ( .C1(n19533), .C2(n19473), .A(n19424), .B(n19423), .ZN(
        P2_U3115) );
  AOI22_X1 U22408 ( .A1(n19673), .A2(n19432), .B1(n19670), .B2(n19431), .ZN(
        n19426) );
  AOI22_X1 U22409 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19439), .B1(
        n19671), .B2(n19438), .ZN(n19425) );
  OAI211_X1 U22410 ( .C1(n19610), .C2(n19436), .A(n19426), .B(n19425), .ZN(
        P2_U3116) );
  OAI22_X1 U22411 ( .A1(n19436), .A2(n19613), .B1(n19435), .B2(n19427), .ZN(
        n19428) );
  INV_X1 U22412 ( .A(n19428), .ZN(n19430) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19439), .B1(
        n19677), .B2(n19438), .ZN(n19429) );
  OAI211_X1 U22414 ( .C1(n19539), .C2(n19473), .A(n19430), .B(n19429), .ZN(
        P2_U3117) );
  AOI22_X1 U22415 ( .A1(n19685), .A2(n19432), .B1(n19682), .B2(n19431), .ZN(
        n19434) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19439), .B1(
        n19683), .B2(n19438), .ZN(n19433) );
  OAI211_X1 U22417 ( .C1(n19616), .C2(n19436), .A(n19434), .B(n19433), .ZN(
        P2_U3118) );
  OAI22_X1 U22418 ( .A1(n19436), .A2(n19623), .B1(n19472), .B2(n19435), .ZN(
        n19437) );
  INV_X1 U22419 ( .A(n19437), .ZN(n19441) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19439), .B1(
        n19690), .B2(n19438), .ZN(n19440) );
  OAI211_X1 U22421 ( .C1(n19549), .C2(n19473), .A(n19441), .B(n19440), .ZN(
        P2_U3119) );
  AOI22_X1 U22422 ( .A1(n19595), .A2(n19498), .B1(n19586), .B2(n19484), .ZN(
        n19453) );
  AOI21_X1 U22423 ( .B1(n19443), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19446) );
  AOI21_X1 U22424 ( .B1(n19516), .B2(n19444), .A(n19556), .ZN(n19447) );
  OR2_X1 U22425 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19517), .ZN(
        n19450) );
  NAND2_X1 U22426 ( .A1(n19447), .A2(n19450), .ZN(n19445) );
  OAI211_X1 U22427 ( .C1(n19484), .C2(n19446), .A(n19445), .B(n19593), .ZN(
        n19476) );
  INV_X1 U22428 ( .A(n19447), .ZN(n19451) );
  OAI21_X1 U22429 ( .B1(n19448), .B2(n19484), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19449) );
  OAI21_X1 U22430 ( .B1(n19451), .B2(n19450), .A(n19449), .ZN(n19475) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19476), .B1(
        n13539), .B2(n19475), .ZN(n19452) );
  OAI211_X1 U22432 ( .C1(n19598), .C2(n19473), .A(n19453), .B(n19452), .ZN(
        P2_U3120) );
  AOI22_X1 U22433 ( .A1(n19498), .A2(n19655), .B1(n19484), .B2(n19624), .ZN(
        n19455) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19476), .B1(
        n15341), .B2(n19475), .ZN(n19454) );
  OAI211_X1 U22435 ( .C1(n19601), .C2(n19473), .A(n19455), .B(n19454), .ZN(
        P2_U3121) );
  AOI22_X1 U22436 ( .A1(n19630), .A2(n19498), .B1(n19484), .B2(n19628), .ZN(
        n19457) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19476), .B1(
        n13567), .B2(n19475), .ZN(n19456) );
  OAI211_X1 U22438 ( .C1(n19604), .C2(n19473), .A(n19457), .B(n19456), .ZN(
        P2_U3122) );
  INV_X1 U22439 ( .A(n19484), .ZN(n19471) );
  OAI22_X1 U22440 ( .A1(n19473), .A2(n19607), .B1(n19471), .B2(n19661), .ZN(
        n19458) );
  INV_X1 U22441 ( .A(n19458), .ZN(n19460) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19476), .B1(
        n19659), .B2(n19475), .ZN(n19459) );
  OAI211_X1 U22443 ( .C1(n19533), .C2(n19509), .A(n19460), .B(n19459), .ZN(
        P2_U3123) );
  OAI22_X1 U22444 ( .A1(n19473), .A2(n19610), .B1(n19461), .B2(n19471), .ZN(
        n19462) );
  INV_X1 U22445 ( .A(n19462), .ZN(n19464) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19476), .B1(
        n19671), .B2(n19475), .ZN(n19463) );
  OAI211_X1 U22447 ( .C1(n19536), .C2(n19509), .A(n19464), .B(n19463), .ZN(
        P2_U3124) );
  AOI22_X1 U22448 ( .A1(n19498), .A2(n19678), .B1(n19484), .B2(n19676), .ZN(
        n19466) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19476), .B1(
        n19677), .B2(n19475), .ZN(n19465) );
  OAI211_X1 U22450 ( .C1(n19613), .C2(n19473), .A(n19466), .B(n19465), .ZN(
        P2_U3125) );
  INV_X1 U22451 ( .A(n19682), .ZN(n19467) );
  OAI22_X1 U22452 ( .A1(n19473), .A2(n19616), .B1(n19467), .B2(n19471), .ZN(
        n19468) );
  INV_X1 U22453 ( .A(n19468), .ZN(n19470) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19476), .B1(
        n19683), .B2(n19475), .ZN(n19469) );
  OAI211_X1 U22455 ( .C1(n19542), .C2(n19509), .A(n19470), .B(n19469), .ZN(
        P2_U3126) );
  OAI22_X1 U22456 ( .A1(n19473), .A2(n19623), .B1(n19472), .B2(n19471), .ZN(
        n19474) );
  INV_X1 U22457 ( .A(n19474), .ZN(n19478) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19476), .B1(
        n19690), .B2(n19475), .ZN(n19477) );
  OAI211_X1 U22459 ( .C1(n19549), .C2(n19509), .A(n19478), .B(n19477), .ZN(
        P2_U3127) );
  NOR3_X2 U22460 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19821), .A3(
        n19517), .ZN(n19504) );
  OAI21_X1 U22461 ( .B1(n19479), .B2(n19504), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19480) );
  OAI21_X1 U22462 ( .B1(n19517), .B2(n19481), .A(n19480), .ZN(n19505) );
  AOI22_X1 U22463 ( .A1(n19505), .A2(n13539), .B1(n19586), .B2(n19504), .ZN(
        n19489) );
  NAND2_X1 U22464 ( .A1(n19483), .A2(n19482), .ZN(n19501) );
  AOI221_X1 U22465 ( .B1(n19498), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19545), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19484), .ZN(n19485) );
  AOI211_X1 U22466 ( .C1(n19486), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19485), .ZN(n19487) );
  OAI21_X1 U22467 ( .B1(n19487), .B2(n19504), .A(n19593), .ZN(n19506) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19506), .B1(
        n19545), .B2(n19595), .ZN(n19488) );
  OAI211_X1 U22469 ( .C1(n19598), .C2(n19509), .A(n19489), .B(n19488), .ZN(
        P2_U3128) );
  AOI22_X1 U22470 ( .A1(n19505), .A2(n15341), .B1(n19624), .B2(n19504), .ZN(
        n19491) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19506), .B1(
        n19545), .B2(n19655), .ZN(n19490) );
  OAI211_X1 U22472 ( .C1(n19601), .C2(n19509), .A(n19491), .B(n19490), .ZN(
        P2_U3129) );
  AOI22_X1 U22473 ( .A1(n19505), .A2(n13567), .B1(n19628), .B2(n19504), .ZN(
        n19493) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19506), .B1(
        n19545), .B2(n19630), .ZN(n19492) );
  OAI211_X1 U22475 ( .C1(n19604), .C2(n19509), .A(n19493), .B(n19492), .ZN(
        P2_U3130) );
  AOI22_X1 U22476 ( .A1(n19505), .A2(n19659), .B1(n19634), .B2(n19504), .ZN(
        n19495) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19506), .B1(
        n19498), .B2(n19665), .ZN(n19494) );
  OAI211_X1 U22478 ( .C1(n19533), .C2(n19501), .A(n19495), .B(n19494), .ZN(
        P2_U3131) );
  AOI22_X1 U22479 ( .A1(n19505), .A2(n19671), .B1(n19670), .B2(n19504), .ZN(
        n19497) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19506), .B1(
        n19545), .B2(n19673), .ZN(n19496) );
  OAI211_X1 U22481 ( .C1(n19610), .C2(n19509), .A(n19497), .B(n19496), .ZN(
        P2_U3132) );
  AOI22_X1 U22482 ( .A1(n19505), .A2(n19677), .B1(n19676), .B2(n19504), .ZN(
        n19500) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19506), .B1(
        n19498), .B2(n19679), .ZN(n19499) );
  OAI211_X1 U22484 ( .C1(n19539), .C2(n19501), .A(n19500), .B(n19499), .ZN(
        P2_U3133) );
  AOI22_X1 U22485 ( .A1(n19505), .A2(n19683), .B1(n19682), .B2(n19504), .ZN(
        n19503) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19506), .B1(
        n19545), .B2(n19685), .ZN(n19502) );
  OAI211_X1 U22487 ( .C1(n19616), .C2(n19509), .A(n19503), .B(n19502), .ZN(
        P2_U3134) );
  AOI22_X1 U22488 ( .A1(n19505), .A2(n19690), .B1(n19688), .B2(n19504), .ZN(
        n19508) );
  AOI22_X1 U22489 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19506), .B1(
        n19545), .B2(n19692), .ZN(n19507) );
  OAI211_X1 U22490 ( .C1(n19623), .C2(n19509), .A(n19508), .B(n19507), .ZN(
        P2_U3135) );
  OR2_X1 U22491 ( .A1(n19821), .A2(n19517), .ZN(n19514) );
  NOR2_X1 U22492 ( .A1(n19511), .A2(n19517), .ZN(n19543) );
  OAI21_X1 U22493 ( .B1(n19512), .B2(n19543), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19513) );
  OAI21_X1 U22494 ( .B1(n19514), .B2(n19556), .A(n19513), .ZN(n19544) );
  AOI22_X1 U22495 ( .A1(n19544), .A2(n13539), .B1(n19586), .B2(n19543), .ZN(
        n19523) );
  AOI21_X1 U22496 ( .B1(n19515), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19520) );
  INV_X1 U22497 ( .A(n19516), .ZN(n19591) );
  OAI22_X1 U22498 ( .A1(n19591), .A2(n19518), .B1(n19517), .B2(n19821), .ZN(
        n19519) );
  OAI211_X1 U22499 ( .C1(n19543), .C2(n19520), .A(n19519), .B(n19593), .ZN(
        n19546) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19521), .ZN(n19522) );
  OAI211_X1 U22501 ( .C1(n19524), .C2(n19582), .A(n19523), .B(n19522), .ZN(
        P2_U3136) );
  AOI22_X1 U22502 ( .A1(n19544), .A2(n15341), .B1(n19624), .B2(n19543), .ZN(
        n19526) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19654), .ZN(n19525) );
  OAI211_X1 U22504 ( .C1(n19527), .C2(n19582), .A(n19526), .B(n19525), .ZN(
        P2_U3137) );
  AOI22_X1 U22505 ( .A1(n19544), .A2(n13567), .B1(n19628), .B2(n19543), .ZN(
        n19529) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19629), .ZN(n19528) );
  OAI211_X1 U22507 ( .C1(n19530), .C2(n19582), .A(n19529), .B(n19528), .ZN(
        P2_U3138) );
  AOI22_X1 U22508 ( .A1(n19544), .A2(n19659), .B1(n19634), .B2(n19543), .ZN(
        n19532) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19665), .ZN(n19531) );
  OAI211_X1 U22510 ( .C1(n19533), .C2(n19582), .A(n19532), .B(n19531), .ZN(
        P2_U3139) );
  AOI22_X1 U22511 ( .A1(n19544), .A2(n19671), .B1(n19670), .B2(n19543), .ZN(
        n19535) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19672), .ZN(n19534) );
  OAI211_X1 U22513 ( .C1(n19536), .C2(n19582), .A(n19535), .B(n19534), .ZN(
        P2_U3140) );
  AOI22_X1 U22514 ( .A1(n19544), .A2(n19677), .B1(n19676), .B2(n19543), .ZN(
        n19538) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19679), .ZN(n19537) );
  OAI211_X1 U22516 ( .C1(n19539), .C2(n19582), .A(n19538), .B(n19537), .ZN(
        P2_U3141) );
  AOI22_X1 U22517 ( .A1(n19544), .A2(n19683), .B1(n19682), .B2(n19543), .ZN(
        n19541) );
  AOI22_X1 U22518 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19684), .ZN(n19540) );
  OAI211_X1 U22519 ( .C1(n19542), .C2(n19582), .A(n19541), .B(n19540), .ZN(
        P2_U3142) );
  AOI22_X1 U22520 ( .A1(n19544), .A2(n19690), .B1(n19688), .B2(n19543), .ZN(
        n19548) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19694), .ZN(n19547) );
  OAI211_X1 U22522 ( .C1(n19549), .C2(n19582), .A(n19548), .B(n19547), .ZN(
        P2_U3143) );
  NOR2_X1 U22523 ( .A1(n19805), .A2(n19550), .ZN(n19560) );
  INV_X1 U22524 ( .A(n19560), .ZN(n19553) );
  NOR2_X1 U22525 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19589), .ZN(
        n19576) );
  OAI21_X1 U22526 ( .B1(n19551), .B2(n19576), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19552) );
  OAI21_X1 U22527 ( .B1(n19553), .B2(n19556), .A(n19552), .ZN(n19577) );
  AOI22_X1 U22528 ( .A1(n19577), .A2(n13539), .B1(n19586), .B2(n19576), .ZN(
        n19563) );
  AOI21_X1 U22529 ( .B1(n19622), .B2(n19582), .A(n19797), .ZN(n19561) );
  INV_X1 U22530 ( .A(n19576), .ZN(n19557) );
  OAI211_X1 U22531 ( .C1(n19558), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19557), 
        .B(n19556), .ZN(n19559) );
  OAI211_X1 U22532 ( .C1(n19561), .C2(n19560), .A(n19593), .B(n19559), .ZN(
        n19579) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19579), .B1(
        n19578), .B2(n19595), .ZN(n19562) );
  OAI211_X1 U22534 ( .C1(n19598), .C2(n19582), .A(n19563), .B(n19562), .ZN(
        P2_U3144) );
  AOI22_X1 U22535 ( .A1(n19577), .A2(n15341), .B1(n19624), .B2(n19576), .ZN(
        n19565) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19579), .B1(
        n19578), .B2(n19655), .ZN(n19564) );
  OAI211_X1 U22537 ( .C1(n19601), .C2(n19582), .A(n19565), .B(n19564), .ZN(
        P2_U3145) );
  AOI22_X1 U22538 ( .A1(n19577), .A2(n13567), .B1(n19628), .B2(n19576), .ZN(
        n19567) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19579), .B1(
        n19578), .B2(n19630), .ZN(n19566) );
  OAI211_X1 U22540 ( .C1(n19604), .C2(n19582), .A(n19567), .B(n19566), .ZN(
        P2_U3146) );
  AOI22_X1 U22541 ( .A1(n19577), .A2(n19659), .B1(n19634), .B2(n19576), .ZN(
        n19569) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19579), .B1(
        n19578), .B2(n19664), .ZN(n19568) );
  OAI211_X1 U22543 ( .C1(n19607), .C2(n19582), .A(n19569), .B(n19568), .ZN(
        P2_U3147) );
  AOI22_X1 U22544 ( .A1(n19577), .A2(n19671), .B1(n19670), .B2(n19576), .ZN(
        n19571) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19579), .B1(
        n19578), .B2(n19673), .ZN(n19570) );
  OAI211_X1 U22546 ( .C1(n19610), .C2(n19582), .A(n19571), .B(n19570), .ZN(
        P2_U3148) );
  AOI22_X1 U22547 ( .A1(n19577), .A2(n19677), .B1(n19676), .B2(n19576), .ZN(
        n19573) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19579), .B1(
        n19578), .B2(n19678), .ZN(n19572) );
  OAI211_X1 U22549 ( .C1(n19613), .C2(n19582), .A(n19573), .B(n19572), .ZN(
        P2_U3149) );
  AOI22_X1 U22550 ( .A1(n19577), .A2(n19683), .B1(n19682), .B2(n19576), .ZN(
        n19575) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19579), .B1(
        n19578), .B2(n19685), .ZN(n19574) );
  OAI211_X1 U22552 ( .C1(n19616), .C2(n19582), .A(n19575), .B(n19574), .ZN(
        P2_U3150) );
  AOI22_X1 U22553 ( .A1(n19577), .A2(n19690), .B1(n19688), .B2(n19576), .ZN(
        n19581) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19579), .B1(
        n19578), .B2(n19692), .ZN(n19580) );
  OAI211_X1 U22555 ( .C1(n19623), .C2(n19582), .A(n19581), .B(n19580), .ZN(
        P2_U3151) );
  INV_X1 U22556 ( .A(n19617), .ZN(n19583) );
  NAND3_X1 U22557 ( .A1(n19584), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19583), 
        .ZN(n19592) );
  OAI21_X1 U22558 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19589), .A(n19843), 
        .ZN(n19585) );
  AOI22_X1 U22559 ( .A1(n19618), .A2(n13539), .B1(n19586), .B2(n19617), .ZN(
        n19597) );
  NAND2_X1 U22560 ( .A1(n19588), .A2(n19587), .ZN(n19590) );
  OAI22_X1 U22561 ( .A1(n19591), .A2(n19590), .B1(n19827), .B2(n19589), .ZN(
        n19594) );
  NAND3_X1 U22562 ( .A1(n19594), .A2(n19593), .A3(n19592), .ZN(n19619) );
  AOI22_X1 U22563 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19619), .B1(
        n19645), .B2(n19595), .ZN(n19596) );
  OAI211_X1 U22564 ( .C1(n19598), .C2(n19622), .A(n19597), .B(n19596), .ZN(
        P2_U3152) );
  AOI22_X1 U22565 ( .A1(n19618), .A2(n15341), .B1(n19624), .B2(n19617), .ZN(
        n19600) );
  AOI22_X1 U22566 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19619), .B1(
        n19645), .B2(n19655), .ZN(n19599) );
  OAI211_X1 U22567 ( .C1(n19601), .C2(n19622), .A(n19600), .B(n19599), .ZN(
        P2_U3153) );
  AOI22_X1 U22568 ( .A1(n19618), .A2(n13567), .B1(n19628), .B2(n19617), .ZN(
        n19603) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19619), .B1(
        n19645), .B2(n19630), .ZN(n19602) );
  OAI211_X1 U22570 ( .C1(n19604), .C2(n19622), .A(n19603), .B(n19602), .ZN(
        P2_U3154) );
  AOI22_X1 U22571 ( .A1(n19618), .A2(n19659), .B1(n19634), .B2(n19617), .ZN(
        n19606) );
  AOI22_X1 U22572 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19619), .B1(
        n19645), .B2(n19664), .ZN(n19605) );
  OAI211_X1 U22573 ( .C1(n19607), .C2(n19622), .A(n19606), .B(n19605), .ZN(
        P2_U3155) );
  AOI22_X1 U22574 ( .A1(n19618), .A2(n19671), .B1(n19670), .B2(n19617), .ZN(
        n19609) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19619), .B1(
        n19645), .B2(n19673), .ZN(n19608) );
  OAI211_X1 U22576 ( .C1(n19610), .C2(n19622), .A(n19609), .B(n19608), .ZN(
        P2_U3156) );
  AOI22_X1 U22577 ( .A1(n19618), .A2(n19677), .B1(n19676), .B2(n19617), .ZN(
        n19612) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19619), .B1(
        n19645), .B2(n19678), .ZN(n19611) );
  OAI211_X1 U22579 ( .C1(n19613), .C2(n19622), .A(n19612), .B(n19611), .ZN(
        P2_U3157) );
  AOI22_X1 U22580 ( .A1(n19618), .A2(n19683), .B1(n19682), .B2(n19617), .ZN(
        n19615) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19619), .B1(
        n19645), .B2(n19685), .ZN(n19614) );
  OAI211_X1 U22582 ( .C1(n19616), .C2(n19622), .A(n19615), .B(n19614), .ZN(
        P2_U3158) );
  AOI22_X1 U22583 ( .A1(n19618), .A2(n19690), .B1(n19688), .B2(n19617), .ZN(
        n19621) );
  AOI22_X1 U22584 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19619), .B1(
        n19645), .B2(n19692), .ZN(n19620) );
  OAI211_X1 U22585 ( .C1(n19623), .C2(n19622), .A(n19621), .B(n19620), .ZN(
        P2_U3159) );
  AOI22_X1 U22586 ( .A1(n19695), .A2(n19655), .B1(n19644), .B2(n19624), .ZN(
        n19626) );
  AOI22_X1 U22587 ( .A1(n15341), .A2(n19646), .B1(n19645), .B2(n19654), .ZN(
        n19625) );
  OAI211_X1 U22588 ( .C1(n19650), .C2(n19627), .A(n19626), .B(n19625), .ZN(
        P2_U3161) );
  AOI22_X1 U22589 ( .A1(n19645), .A2(n19629), .B1(n19644), .B2(n19628), .ZN(
        n19632) );
  AOI22_X1 U22590 ( .A1(n13567), .A2(n19646), .B1(n19695), .B2(n19630), .ZN(
        n19631) );
  OAI211_X1 U22591 ( .C1(n19650), .C2(n19633), .A(n19632), .B(n19631), .ZN(
        P2_U3162) );
  INV_X1 U22592 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n19637) );
  AOI22_X1 U22593 ( .A1(n19695), .A2(n19664), .B1(n19644), .B2(n19634), .ZN(
        n19636) );
  AOI22_X1 U22594 ( .A1(n19659), .A2(n19646), .B1(n19645), .B2(n19665), .ZN(
        n19635) );
  OAI211_X1 U22595 ( .C1(n19650), .C2(n19637), .A(n19636), .B(n19635), .ZN(
        P2_U3163) );
  INV_X1 U22596 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19640) );
  AOI22_X1 U22597 ( .A1(n19645), .A2(n19672), .B1(n19670), .B2(n19644), .ZN(
        n19639) );
  AOI22_X1 U22598 ( .A1(n19671), .A2(n19646), .B1(n19695), .B2(n19673), .ZN(
        n19638) );
  OAI211_X1 U22599 ( .C1(n19650), .C2(n19640), .A(n19639), .B(n19638), .ZN(
        P2_U3164) );
  INV_X1 U22600 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n19643) );
  AOI22_X1 U22601 ( .A1(n19645), .A2(n19679), .B1(n19644), .B2(n19676), .ZN(
        n19642) );
  AOI22_X1 U22602 ( .A1(n19677), .A2(n19646), .B1(n19695), .B2(n19678), .ZN(
        n19641) );
  OAI211_X1 U22603 ( .C1(n19650), .C2(n19643), .A(n19642), .B(n19641), .ZN(
        P2_U3165) );
  INV_X1 U22604 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n19649) );
  AOI22_X1 U22605 ( .A1(n19645), .A2(n19684), .B1(n19644), .B2(n19682), .ZN(
        n19648) );
  AOI22_X1 U22606 ( .A1(n19683), .A2(n19646), .B1(n19695), .B2(n19685), .ZN(
        n19647) );
  OAI211_X1 U22607 ( .C1(n19650), .C2(n19649), .A(n19648), .B(n19647), .ZN(
        P2_U3166) );
  INV_X1 U22608 ( .A(n15341), .ZN(n19652) );
  OAI22_X1 U22609 ( .A1(n19669), .A2(n19652), .B1(n19651), .B2(n19660), .ZN(
        n19653) );
  INV_X1 U22610 ( .A(n19653), .ZN(n19657) );
  AOI22_X1 U22611 ( .A1(n19693), .A2(n19655), .B1(n19695), .B2(n19654), .ZN(
        n19656) );
  OAI211_X1 U22612 ( .C1(n19699), .C2(n19658), .A(n19657), .B(n19656), .ZN(
        P2_U3169) );
  INV_X1 U22613 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n19668) );
  INV_X1 U22614 ( .A(n19659), .ZN(n19662) );
  OAI22_X1 U22615 ( .A1(n19669), .A2(n19662), .B1(n19661), .B2(n19660), .ZN(
        n19663) );
  INV_X1 U22616 ( .A(n19663), .ZN(n19667) );
  AOI22_X1 U22617 ( .A1(n19695), .A2(n19665), .B1(n19693), .B2(n19664), .ZN(
        n19666) );
  OAI211_X1 U22618 ( .C1(n19699), .C2(n19668), .A(n19667), .B(n19666), .ZN(
        P2_U3171) );
  INV_X1 U22619 ( .A(n19669), .ZN(n19691) );
  AOI22_X1 U22620 ( .A1(n19691), .A2(n19671), .B1(n19689), .B2(n19670), .ZN(
        n19675) );
  AOI22_X1 U22621 ( .A1(n19693), .A2(n19673), .B1(n19695), .B2(n19672), .ZN(
        n19674) );
  OAI211_X1 U22622 ( .C1(n19699), .C2(n12308), .A(n19675), .B(n19674), .ZN(
        P2_U3172) );
  AOI22_X1 U22623 ( .A1(n19691), .A2(n19677), .B1(n19689), .B2(n19676), .ZN(
        n19681) );
  AOI22_X1 U22624 ( .A1(n19695), .A2(n19679), .B1(n19693), .B2(n19678), .ZN(
        n19680) );
  OAI211_X1 U22625 ( .C1(n19699), .C2(n12334), .A(n19681), .B(n19680), .ZN(
        P2_U3173) );
  AOI22_X1 U22626 ( .A1(n19691), .A2(n19683), .B1(n19689), .B2(n19682), .ZN(
        n19687) );
  AOI22_X1 U22627 ( .A1(n19693), .A2(n19685), .B1(n19695), .B2(n19684), .ZN(
        n19686) );
  OAI211_X1 U22628 ( .C1(n19699), .C2(n12355), .A(n19687), .B(n19686), .ZN(
        P2_U3174) );
  INV_X1 U22629 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19698) );
  AOI22_X1 U22630 ( .A1(n19691), .A2(n19690), .B1(n19689), .B2(n19688), .ZN(
        n19697) );
  AOI22_X1 U22631 ( .A1(n19695), .A2(n19694), .B1(n19693), .B2(n19692), .ZN(
        n19696) );
  OAI211_X1 U22632 ( .C1(n19699), .C2(n19698), .A(n19697), .B(n19696), .ZN(
        P2_U3175) );
  AOI21_X1 U22633 ( .B1(n19702), .B2(n19701), .A(n19700), .ZN(n19707) );
  OAI211_X1 U22634 ( .C1(n19703), .C2(n19706), .A(n19845), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19704) );
  OAI211_X1 U22635 ( .C1(n19707), .C2(n19706), .A(n19705), .B(n19704), .ZN(
        P2_U3177) );
  AND2_X1 U22636 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19711), .ZN(
        P2_U3179) );
  AND2_X1 U22637 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19711), .ZN(
        P2_U3180) );
  AND2_X1 U22638 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19711), .ZN(
        P2_U3181) );
  AND2_X1 U22639 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19711), .ZN(
        P2_U3182) );
  AND2_X1 U22640 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19711), .ZN(
        P2_U3183) );
  AND2_X1 U22641 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19711), .ZN(
        P2_U3184) );
  AND2_X1 U22642 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19711), .ZN(
        P2_U3185) );
  NOR2_X1 U22643 ( .A1(n19708), .A2(n19787), .ZN(P2_U3186) );
  AND2_X1 U22644 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19711), .ZN(
        P2_U3187) );
  AND2_X1 U22645 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19711), .ZN(
        P2_U3188) );
  AND2_X1 U22646 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19711), .ZN(
        P2_U3189) );
  INV_X1 U22647 ( .A(n19787), .ZN(n19710) );
  AND2_X1 U22648 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19710), .ZN(
        P2_U3190) );
  AND2_X1 U22649 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19710), .ZN(
        P2_U3191) );
  AND2_X1 U22650 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19710), .ZN(
        P2_U3192) );
  AND2_X1 U22651 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19710), .ZN(
        P2_U3193) );
  AND2_X1 U22652 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19710), .ZN(
        P2_U3194) );
  AND2_X1 U22653 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19710), .ZN(
        P2_U3195) );
  AND2_X1 U22654 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19710), .ZN(
        P2_U3196) );
  AND2_X1 U22655 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19710), .ZN(
        P2_U3197) );
  NOR2_X1 U22656 ( .A1(n19709), .A2(n19787), .ZN(P2_U3198) );
  AND2_X1 U22657 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19710), .ZN(
        P2_U3199) );
  AND2_X1 U22658 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19710), .ZN(
        P2_U3200) );
  AND2_X1 U22659 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19710), .ZN(P2_U3201) );
  AND2_X1 U22660 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19710), .ZN(P2_U3202) );
  AND2_X1 U22661 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19711), .ZN(P2_U3203) );
  AND2_X1 U22662 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19711), .ZN(P2_U3204) );
  AND2_X1 U22663 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19711), .ZN(P2_U3205) );
  AND2_X1 U22664 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19710), .ZN(P2_U3206) );
  AND2_X1 U22665 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19710), .ZN(P2_U3207) );
  AND2_X1 U22666 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19711), .ZN(P2_U3208) );
  INV_X1 U22667 ( .A(NA), .ZN(n20767) );
  INV_X1 U22668 ( .A(n19712), .ZN(n19718) );
  OAI21_X1 U22669 ( .B1(n20767), .B2(n19718), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19728) );
  NAND2_X1 U22670 ( .A1(n19845), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19726) );
  NAND3_X1 U22671 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19726), .ZN(n19715) );
  AOI211_X1 U22672 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20761), .A(
        n19867), .B(n19713), .ZN(n19714) );
  AOI21_X1 U22673 ( .B1(n19728), .B2(n19715), .A(n19714), .ZN(n19716) );
  INV_X1 U22674 ( .A(n19716), .ZN(P2_U3209) );
  NOR2_X1 U22675 ( .A1(HOLD), .A2(n19717), .ZN(n19727) );
  AOI21_X1 U22676 ( .B1(n19729), .B2(n19718), .A(n19727), .ZN(n19722) );
  INV_X1 U22677 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19721) );
  AOI21_X1 U22678 ( .B1(HOLD), .B2(n19719), .A(n19856), .ZN(n19720) );
  OAI211_X1 U22679 ( .C1(n19722), .C2(n19721), .A(n19720), .B(n19726), .ZN(
        P2_U3210) );
  OAI22_X1 U22680 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19723), .B1(NA), 
        .B2(n19726), .ZN(n19724) );
  OAI211_X1 U22681 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19724), .ZN(n19725) );
  OAI221_X1 U22682 ( .B1(n19728), .B2(n19727), .C1(n19728), .C2(n19726), .A(
        n19725), .ZN(P2_U3211) );
  OAI222_X1 U22683 ( .A1(n19776), .A2(n19731), .B1(n19730), .B2(n19867), .C1(
        n19733), .C2(n19780), .ZN(P2_U3212) );
  OAI222_X1 U22684 ( .A1(n19776), .A2(n19733), .B1(n19732), .B2(n19867), .C1(
        n13454), .C2(n19780), .ZN(P2_U3213) );
  OAI222_X1 U22685 ( .A1(n19776), .A2(n13454), .B1(n19734), .B2(n19867), .C1(
        n10972), .C2(n19780), .ZN(P2_U3214) );
  OAI222_X1 U22686 ( .A1(n19780), .A2(n15310), .B1(n19735), .B2(n19867), .C1(
        n10972), .C2(n19776), .ZN(P2_U3215) );
  OAI222_X1 U22687 ( .A1(n19780), .A2(n19737), .B1(n19736), .B2(n19867), .C1(
        n15310), .C2(n19776), .ZN(P2_U3216) );
  OAI222_X1 U22688 ( .A1(n19780), .A2(n19739), .B1(n19738), .B2(n19867), .C1(
        n19737), .C2(n19776), .ZN(P2_U3217) );
  OAI222_X1 U22689 ( .A1(n19780), .A2(n10868), .B1(n19740), .B2(n19867), .C1(
        n19739), .C2(n19776), .ZN(P2_U3218) );
  OAI222_X1 U22690 ( .A1(n19780), .A2(n19742), .B1(n19741), .B2(n19867), .C1(
        n10868), .C2(n19776), .ZN(P2_U3219) );
  OAI222_X1 U22691 ( .A1(n19780), .A2(n10895), .B1(n19743), .B2(n19867), .C1(
        n19742), .C2(n19776), .ZN(P2_U3220) );
  OAI222_X1 U22692 ( .A1(n19780), .A2(n19745), .B1(n19744), .B2(n19867), .C1(
        n10895), .C2(n19776), .ZN(P2_U3221) );
  OAI222_X1 U22693 ( .A1(n19780), .A2(n14973), .B1(n19746), .B2(n19867), .C1(
        n19745), .C2(n19776), .ZN(P2_U3222) );
  OAI222_X1 U22694 ( .A1(n19780), .A2(n14957), .B1(n19747), .B2(n19867), .C1(
        n14973), .C2(n19776), .ZN(P2_U3223) );
  OAI222_X1 U22695 ( .A1(n19780), .A2(n14945), .B1(n19748), .B2(n19867), .C1(
        n14957), .C2(n19776), .ZN(P2_U3224) );
  OAI222_X1 U22696 ( .A1(n19780), .A2(n19750), .B1(n19749), .B2(n19867), .C1(
        n14945), .C2(n19776), .ZN(P2_U3225) );
  OAI222_X1 U22697 ( .A1(n19780), .A2(n11014), .B1(n19751), .B2(n19867), .C1(
        n19750), .C2(n19776), .ZN(P2_U3226) );
  OAI222_X1 U22698 ( .A1(n19780), .A2(n19753), .B1(n19752), .B2(n19867), .C1(
        n11014), .C2(n19776), .ZN(P2_U3227) );
  OAI222_X1 U22699 ( .A1(n19780), .A2(n14904), .B1(n19754), .B2(n19867), .C1(
        n19753), .C2(n19776), .ZN(P2_U3228) );
  OAI222_X1 U22700 ( .A1(n19780), .A2(n19756), .B1(n19755), .B2(n19867), .C1(
        n14904), .C2(n19776), .ZN(P2_U3229) );
  OAI222_X1 U22701 ( .A1(n19780), .A2(n19758), .B1(n19757), .B2(n19867), .C1(
        n19756), .C2(n19776), .ZN(P2_U3230) );
  OAI222_X1 U22702 ( .A1(n19780), .A2(n19760), .B1(n19759), .B2(n19867), .C1(
        n19758), .C2(n19776), .ZN(P2_U3231) );
  OAI222_X1 U22703 ( .A1(n19780), .A2(n12045), .B1(n19761), .B2(n19867), .C1(
        n19760), .C2(n19776), .ZN(P2_U3232) );
  OAI222_X1 U22704 ( .A1(n19780), .A2(n19763), .B1(n19762), .B2(n19867), .C1(
        n12045), .C2(n19776), .ZN(P2_U3233) );
  OAI222_X1 U22705 ( .A1(n19780), .A2(n14832), .B1(n19764), .B2(n19867), .C1(
        n19763), .C2(n19776), .ZN(P2_U3234) );
  OAI222_X1 U22706 ( .A1(n19780), .A2(n19766), .B1(n19765), .B2(n19867), .C1(
        n14832), .C2(n19776), .ZN(P2_U3235) );
  OAI222_X1 U22707 ( .A1(n19780), .A2(n19768), .B1(n19767), .B2(n19867), .C1(
        n19766), .C2(n19776), .ZN(P2_U3236) );
  INV_X1 U22708 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19771) );
  OAI222_X1 U22709 ( .A1(n19780), .A2(n19771), .B1(n19769), .B2(n19867), .C1(
        n19768), .C2(n19776), .ZN(P2_U3237) );
  INV_X1 U22710 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19772) );
  OAI222_X1 U22711 ( .A1(n19776), .A2(n19771), .B1(n19770), .B2(n19867), .C1(
        n19772), .C2(n19780), .ZN(P2_U3238) );
  OAI222_X1 U22712 ( .A1(n19780), .A2(n19774), .B1(n19773), .B2(n19867), .C1(
        n19772), .C2(n19776), .ZN(P2_U3239) );
  OAI222_X1 U22713 ( .A1(n19780), .A2(n19777), .B1(n19775), .B2(n19867), .C1(
        n19774), .C2(n19776), .ZN(P2_U3240) );
  OAI222_X1 U22714 ( .A1(n19780), .A2(n19779), .B1(n19778), .B2(n19867), .C1(
        n19777), .C2(n19776), .ZN(P2_U3241) );
  OAI22_X1 U22715 ( .A1(n19864), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19867), .ZN(n19781) );
  INV_X1 U22716 ( .A(n19781), .ZN(P2_U3585) );
  MUX2_X1 U22717 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19864), .Z(P2_U3586) );
  OAI22_X1 U22718 ( .A1(n19864), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19867), .ZN(n19782) );
  INV_X1 U22719 ( .A(n19782), .ZN(P2_U3587) );
  OAI22_X1 U22720 ( .A1(n19864), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19867), .ZN(n19783) );
  INV_X1 U22721 ( .A(n19783), .ZN(P2_U3588) );
  OAI21_X1 U22722 ( .B1(n19787), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19785), 
        .ZN(n19784) );
  INV_X1 U22723 ( .A(n19784), .ZN(P2_U3591) );
  OAI21_X1 U22724 ( .B1(n19787), .B2(n19786), .A(n19785), .ZN(P2_U3592) );
  INV_X1 U22725 ( .A(n19788), .ZN(n19789) );
  OAI22_X1 U22726 ( .A1(n19791), .A2(n19790), .B1(n19799), .B2(n19789), .ZN(
        n19793) );
  OAI22_X1 U22727 ( .A1(n19794), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19793), .B2(n19792), .ZN(n19795) );
  INV_X1 U22728 ( .A(n19795), .ZN(P2_U3596) );
  INV_X1 U22729 ( .A(n19831), .ZN(n19822) );
  OR2_X1 U22730 ( .A1(n19797), .A2(n19796), .ZN(n19798) );
  NAND2_X1 U22731 ( .A1(n19806), .A2(n19798), .ZN(n19800) );
  NAND2_X1 U22732 ( .A1(n19800), .A2(n19799), .ZN(n19809) );
  AOI222_X1 U22733 ( .A1(n19809), .A2(n19803), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19802), .C1(n19806), .C2(n19801), .ZN(n19804) );
  AOI22_X1 U22734 ( .A1(n19822), .A2(n19805), .B1(n19804), .B2(n19831), .ZN(
        P2_U3602) );
  NAND2_X1 U22735 ( .A1(n19806), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19816) );
  OAI21_X1 U22736 ( .B1(n19808), .B2(n19816), .A(n19807), .ZN(n19810) );
  AOI22_X1 U22737 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19811), .B1(n19810), 
        .B2(n19809), .ZN(n19812) );
  AOI22_X1 U22738 ( .A1(n19822), .A2(n19813), .B1(n19812), .B2(n19831), .ZN(
        P2_U3603) );
  NAND3_X1 U22739 ( .A1(n19817), .A2(n19848), .A3(n19814), .ZN(n19815) );
  OAI21_X1 U22740 ( .B1(n19817), .B2(n19816), .A(n19815), .ZN(n19818) );
  AOI21_X1 U22741 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19819), .A(n19818), 
        .ZN(n19820) );
  AOI22_X1 U22742 ( .A1(n19822), .A2(n19821), .B1(n19820), .B2(n19831), .ZN(
        P2_U3604) );
  INV_X1 U22743 ( .A(n19848), .ZN(n19825) );
  NAND3_X1 U22744 ( .A1(n19823), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19824) );
  OAI21_X1 U22745 ( .B1(n19826), .B2(n19825), .A(n19824), .ZN(n19828) );
  OAI21_X1 U22746 ( .B1(n19828), .B2(n19827), .A(n19831), .ZN(n19829) );
  OAI21_X1 U22747 ( .B1(n19831), .B2(n19830), .A(n19829), .ZN(P2_U3605) );
  OAI22_X1 U22748 ( .A1(n19864), .A2(n19832), .B1(P2_W_R_N_REG_SCAN_IN), .B2(
        n19867), .ZN(n19833) );
  INV_X1 U22749 ( .A(n19833), .ZN(P2_U3608) );
  INV_X1 U22750 ( .A(n19834), .ZN(n19835) );
  AOI22_X1 U22751 ( .A1(n19838), .A2(n19837), .B1(n19836), .B2(n19835), .ZN(
        n19839) );
  NAND2_X1 U22752 ( .A1(n19840), .A2(n19839), .ZN(n19842) );
  MUX2_X1 U22753 ( .A(P2_MORE_REG_SCAN_IN), .B(n19842), .S(n19841), .Z(
        P2_U3609) );
  NOR4_X1 U22754 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19845), .A3(n19844), 
        .A4(n19843), .ZN(n19847) );
  AOI211_X1 U22755 ( .C1(n19849), .C2(n19848), .A(n19847), .B(n19846), .ZN(
        n19863) );
  NAND2_X1 U22756 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19850), .ZN(n19860) );
  INV_X1 U22757 ( .A(n19851), .ZN(n19853) );
  NOR3_X1 U22758 ( .A1(n19853), .A2(n19852), .A3(n19856), .ZN(n19858) );
  AOI211_X1 U22759 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n19856), .A(n19855), 
        .B(n19854), .ZN(n19857) );
  AOI211_X1 U22760 ( .C1(n19860), .C2(n19859), .A(n19858), .B(n19857), .ZN(
        n19862) );
  NAND2_X1 U22761 ( .A1(n19863), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19861) );
  OAI21_X1 U22762 ( .B1(n19863), .B2(n19862), .A(n19861), .ZN(P2_U3610) );
  AOI22_X1 U22763 ( .A1(n19867), .A2(n19866), .B1(n19865), .B2(n19864), .ZN(
        P2_U3611) );
  INV_X1 U22764 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20772) );
  AOI21_X1 U22765 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20775), .A(n20772), 
        .ZN(n19874) );
  INV_X1 U22766 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19868) );
  AND2_X1 U22767 ( .A1(n20772), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20861) );
  AOI21_X1 U22768 ( .B1(n19874), .B2(n19868), .A(n20861), .ZN(P1_U2802) );
  OAI21_X1 U22769 ( .B1(n19870), .B2(n19869), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19871) );
  OAI21_X1 U22770 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19872), .A(n19871), 
        .ZN(P1_U2803) );
  INV_X2 U22771 ( .A(n20861), .ZN(n20858) );
  NOR2_X1 U22772 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19875) );
  OAI21_X1 U22773 ( .B1(n19875), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20858), .ZN(
        n19873) );
  OAI21_X1 U22774 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20858), .A(n19873), 
        .ZN(P1_U2804) );
  NOR2_X1 U22775 ( .A1(n20861), .A2(n19874), .ZN(n20830) );
  OAI21_X1 U22776 ( .B1(BS16), .B2(n19875), .A(n20830), .ZN(n20828) );
  OAI21_X1 U22777 ( .B1(n20830), .B2(n14399), .A(n20828), .ZN(P1_U2805) );
  AOI21_X1 U22778 ( .B1(n19876), .B2(P1_FLUSH_REG_SCAN_IN), .A(n20071), .ZN(
        n19877) );
  INV_X1 U22779 ( .A(n19877), .ZN(P1_U2806) );
  NOR4_X1 U22780 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19881) );
  NOR4_X1 U22781 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19880) );
  NOR4_X1 U22782 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19879) );
  NOR4_X1 U22783 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19878) );
  NAND4_X1 U22784 ( .A1(n19881), .A2(n19880), .A3(n19879), .A4(n19878), .ZN(
        n19887) );
  NOR4_X1 U22785 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19885) );
  AOI211_X1 U22786 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_17__SCAN_IN), .B(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19884) );
  NOR4_X1 U22787 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A3(P1_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n19883) );
  NOR4_X1 U22788 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19882) );
  NAND4_X1 U22789 ( .A1(n19885), .A2(n19884), .A3(n19883), .A4(n19882), .ZN(
        n19886) );
  NOR2_X1 U22790 ( .A1(n19887), .A2(n19886), .ZN(n20842) );
  INV_X1 U22791 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20825) );
  NOR3_X1 U22792 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19889) );
  OAI21_X1 U22793 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19889), .A(n20842), .ZN(
        n19888) );
  OAI21_X1 U22794 ( .B1(n20842), .B2(n20825), .A(n19888), .ZN(P1_U2807) );
  INV_X1 U22795 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20829) );
  AOI21_X1 U22796 ( .B1(n20838), .B2(n20829), .A(n19889), .ZN(n19891) );
  INV_X1 U22797 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19890) );
  INV_X1 U22798 ( .A(n20842), .ZN(n20845) );
  AOI22_X1 U22799 ( .A1(n20842), .A2(n19891), .B1(n19890), .B2(n20845), .ZN(
        P1_U2808) );
  AOI22_X1 U22800 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n19955), .B1(
        n19926), .B2(n19964), .ZN(n19899) );
  AOI21_X1 U22801 ( .B1(n19937), .B2(P1_EBX_REG_9__SCAN_IN), .A(n19941), .ZN(
        n19898) );
  AOI22_X1 U22802 ( .A1(n19967), .A2(n19905), .B1(n19961), .B2(n19892), .ZN(
        n19897) );
  AND2_X1 U22803 ( .A1(n19925), .A2(n19893), .ZN(n19895) );
  OAI21_X1 U22804 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n19895), .A(n19894), .ZN(
        n19896) );
  NAND4_X1 U22805 ( .A1(n19899), .A2(n19898), .A3(n19897), .A4(n19896), .ZN(
        P1_U2831) );
  NAND2_X1 U22806 ( .A1(n19925), .A2(n19904), .ZN(n19902) );
  AOI22_X1 U22807 ( .A1(n19900), .A2(n19926), .B1(n19937), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n19901) );
  OAI21_X1 U22808 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n19902), .A(n19901), .ZN(
        n19903) );
  AOI211_X1 U22809 ( .C1(n19955), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19941), .B(n19903), .ZN(n19908) );
  OAI21_X1 U22810 ( .B1(n19958), .B2(n19904), .A(n19931), .ZN(n19922) );
  AOI22_X1 U22811 ( .A1(n19906), .A2(n19905), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n19922), .ZN(n19907) );
  OAI211_X1 U22812 ( .C1(n19909), .C2(n19948), .A(n19908), .B(n19907), .ZN(
        P1_U2833) );
  INV_X1 U22813 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19912) );
  NAND2_X1 U22814 ( .A1(n19937), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n19911) );
  OAI211_X1 U22815 ( .C1(n19913), .C2(n19912), .A(n19911), .B(n19910), .ZN(
        n19916) );
  NOR3_X1 U22816 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n19958), .A3(n19914), .ZN(
        n19915) );
  AOI211_X1 U22817 ( .C1(n19926), .C2(n19917), .A(n19916), .B(n19915), .ZN(
        n19918) );
  OAI21_X1 U22818 ( .B1(n19920), .B2(n19919), .A(n19918), .ZN(n19921) );
  AOI21_X1 U22819 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n19922), .A(n19921), .ZN(
        n19923) );
  OAI21_X1 U22820 ( .B1(n19924), .B2(n19948), .A(n19923), .ZN(P1_U2834) );
  NAND2_X1 U22821 ( .A1(n19925), .A2(n19932), .ZN(n19929) );
  AOI22_X1 U22822 ( .A1(n19927), .A2(n19926), .B1(n19937), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n19928) );
  OAI21_X1 U22823 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n19929), .A(n19928), .ZN(
        n19930) );
  AOI211_X1 U22824 ( .C1(n19955), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n19941), .B(n19930), .ZN(n19935) );
  INV_X1 U22825 ( .A(n19963), .ZN(n19945) );
  OAI21_X1 U22826 ( .B1(n19958), .B2(n19932), .A(n19931), .ZN(n19944) );
  AOI22_X1 U22827 ( .A1(n19933), .A2(n19945), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n19944), .ZN(n19934) );
  OAI211_X1 U22828 ( .C1(n19936), .C2(n19948), .A(n19935), .B(n19934), .ZN(
        P1_U2835) );
  AOI22_X1 U22829 ( .A1(n19938), .A2(n19953), .B1(n19937), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n19939) );
  OAI21_X1 U22830 ( .B1(n19952), .B2(n20094), .A(n19939), .ZN(n19940) );
  AOI211_X1 U22831 ( .C1(n19955), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19941), .B(n19940), .ZN(n19947) );
  OAI21_X1 U22832 ( .B1(n19958), .B2(n19942), .A(n20781), .ZN(n19943) );
  AOI22_X1 U22833 ( .A1(n20069), .A2(n19945), .B1(n19944), .B2(n19943), .ZN(
        n19946) );
  OAI211_X1 U22834 ( .C1(n20074), .C2(n19948), .A(n19947), .B(n19946), .ZN(
        P1_U2836) );
  INV_X1 U22835 ( .A(n20132), .ZN(n19951) );
  OAI22_X1 U22836 ( .A1(n19952), .A2(n19951), .B1(n19950), .B2(n19949), .ZN(
        n19960) );
  NAND2_X1 U22837 ( .A1(n20638), .A2(n19953), .ZN(n19957) );
  AOI22_X1 U22838 ( .A1(n19955), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19954), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n19956) );
  OAI211_X1 U22839 ( .C1(P1_REIP_REG_1__SCAN_IN), .C2(n19958), .A(n19957), .B(
        n19956), .ZN(n19959) );
  AOI211_X1 U22840 ( .C1(n19961), .C2(n20078), .A(n19960), .B(n19959), .ZN(
        n19962) );
  OAI21_X1 U22841 ( .B1(n19963), .B2(n20082), .A(n19962), .ZN(P1_U2839) );
  AOI22_X1 U22842 ( .A1(n19967), .A2(n19966), .B1(n19965), .B2(n19964), .ZN(
        n19968) );
  OAI21_X1 U22843 ( .B1(n19970), .B2(n19969), .A(n19968), .ZN(P1_U2863) );
  INV_X1 U22844 ( .A(n20159), .ZN(n19971) );
  INV_X1 U22845 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20034) );
  OAI222_X1 U22846 ( .A1(n20082), .A2(n19975), .B1(n19974), .B2(n19971), .C1(
        n20034), .C2(n19972), .ZN(P1_U2903) );
  INV_X1 U22847 ( .A(n20150), .ZN(n19973) );
  INV_X1 U22848 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20039) );
  OAI222_X1 U22849 ( .A1(n20083), .A2(n19975), .B1(n19974), .B2(n19973), .C1(
        n20039), .C2(n19972), .ZN(P1_U2904) );
  NAND2_X1 U22850 ( .A1(n20008), .A2(n19976), .ZN(n20004) );
  AOI22_X1 U22851 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n19977) );
  OAI21_X1 U22852 ( .B1(n14100), .B2(n20004), .A(n19977), .ZN(P1_U2906) );
  INV_X1 U22853 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n19979) );
  AOI22_X1 U22854 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n19978) );
  OAI21_X1 U22855 ( .B1(n19979), .B2(n20004), .A(n19978), .ZN(P1_U2907) );
  INV_X1 U22856 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n19981) );
  AOI22_X1 U22857 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20036), .B1(n20022), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n19980) );
  OAI21_X1 U22858 ( .B1(n19981), .B2(n20004), .A(n19980), .ZN(P1_U2908) );
  INV_X1 U22859 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n19983) );
  AOI22_X1 U22860 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20036), .B1(n20022), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n19982) );
  OAI21_X1 U22861 ( .B1(n19983), .B2(n20004), .A(n19982), .ZN(P1_U2909) );
  INV_X1 U22862 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n19985) );
  AOI22_X1 U22863 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20036), .B1(n20022), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n19984) );
  OAI21_X1 U22864 ( .B1(n19985), .B2(n20004), .A(n19984), .ZN(P1_U2910) );
  INV_X1 U22865 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n19987) );
  AOI22_X1 U22866 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20036), .B1(n20022), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n19986) );
  OAI21_X1 U22867 ( .B1(n19987), .B2(n20004), .A(n19986), .ZN(P1_U2911) );
  INV_X1 U22868 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n19989) );
  AOI22_X1 U22869 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20036), .B1(n20022), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n19988) );
  OAI21_X1 U22870 ( .B1(n19989), .B2(n20004), .A(n19988), .ZN(P1_U2912) );
  INV_X1 U22871 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n19991) );
  AOI22_X1 U22872 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n19990) );
  OAI21_X1 U22873 ( .B1(n19991), .B2(n20004), .A(n19990), .ZN(P1_U2913) );
  INV_X1 U22874 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n19993) );
  AOI22_X1 U22875 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n19992) );
  OAI21_X1 U22876 ( .B1(n19993), .B2(n20004), .A(n19992), .ZN(P1_U2914) );
  INV_X1 U22877 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n19995) );
  AOI22_X1 U22878 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n19994) );
  OAI21_X1 U22879 ( .B1(n19995), .B2(n20004), .A(n19994), .ZN(P1_U2915) );
  INV_X1 U22880 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n19997) );
  AOI22_X1 U22881 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n19996) );
  OAI21_X1 U22882 ( .B1(n19997), .B2(n20004), .A(n19996), .ZN(P1_U2916) );
  INV_X1 U22883 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n19999) );
  AOI22_X1 U22884 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n19998) );
  OAI21_X1 U22885 ( .B1(n19999), .B2(n20004), .A(n19998), .ZN(P1_U2917) );
  INV_X1 U22886 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n20001) );
  AOI22_X1 U22887 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n20000) );
  OAI21_X1 U22888 ( .B1(n20001), .B2(n20004), .A(n20000), .ZN(P1_U2918) );
  AOI22_X1 U22889 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n20002) );
  OAI21_X1 U22890 ( .B1(n11552), .B2(n20004), .A(n20002), .ZN(P1_U2919) );
  INV_X1 U22891 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n20005) );
  AOI22_X1 U22892 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n20003) );
  OAI21_X1 U22893 ( .B1(n20005), .B2(n20004), .A(n20003), .ZN(P1_U2920) );
  AOI22_X1 U22894 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20008), .B1(n20035), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20006) );
  OAI21_X1 U22895 ( .B1(n20007), .B2(n20850), .A(n20006), .ZN(P1_U2921) );
  AOI22_X1 U22896 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20009) );
  OAI21_X1 U22897 ( .B1(n13633), .B2(n20038), .A(n20009), .ZN(P1_U2922) );
  AOI22_X1 U22898 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20010) );
  OAI21_X1 U22899 ( .B1(n14159), .B2(n20038), .A(n20010), .ZN(P1_U2923) );
  AOI22_X1 U22900 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20035), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20036), .ZN(n20011) );
  OAI21_X1 U22901 ( .B1(n11488), .B2(n20038), .A(n20011), .ZN(P1_U2924) );
  INV_X1 U22902 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20013) );
  AOI22_X1 U22903 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20012) );
  OAI21_X1 U22904 ( .B1(n20013), .B2(n20038), .A(n20012), .ZN(P1_U2925) );
  INV_X1 U22905 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20015) );
  AOI22_X1 U22906 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20036), .B1(n20022), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20014) );
  OAI21_X1 U22907 ( .B1(n20015), .B2(n20038), .A(n20014), .ZN(P1_U2926) );
  INV_X1 U22908 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20017) );
  AOI22_X1 U22909 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20036), .B1(n20022), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20016) );
  OAI21_X1 U22910 ( .B1(n20017), .B2(n20038), .A(n20016), .ZN(P1_U2927) );
  AOI22_X1 U22911 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20036), .B1(n20022), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20018) );
  OAI21_X1 U22912 ( .B1(n20019), .B2(n20038), .A(n20018), .ZN(P1_U2928) );
  AOI22_X1 U22913 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20036), .B1(n20022), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20020) );
  OAI21_X1 U22914 ( .B1(n20021), .B2(n20038), .A(n20020), .ZN(P1_U2929) );
  AOI22_X1 U22915 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20036), .B1(n20022), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20023) );
  OAI21_X1 U22916 ( .B1(n20024), .B2(n20038), .A(n20023), .ZN(P1_U2930) );
  AOI22_X1 U22917 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20025) );
  OAI21_X1 U22918 ( .B1(n20026), .B2(n20038), .A(n20025), .ZN(P1_U2931) );
  AOI22_X1 U22919 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20027) );
  OAI21_X1 U22920 ( .B1(n20028), .B2(n20038), .A(n20027), .ZN(P1_U2932) );
  AOI22_X1 U22921 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20029) );
  OAI21_X1 U22922 ( .B1(n20030), .B2(n20038), .A(n20029), .ZN(P1_U2933) );
  AOI22_X1 U22923 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20035), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20036), .ZN(n20031) );
  OAI21_X1 U22924 ( .B1(n20032), .B2(n20038), .A(n20031), .ZN(P1_U2934) );
  AOI22_X1 U22925 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20033) );
  OAI21_X1 U22926 ( .B1(n20034), .B2(n20038), .A(n20033), .ZN(P1_U2935) );
  AOI22_X1 U22927 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20036), .B1(n20035), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20037) );
  OAI21_X1 U22928 ( .B1(n20039), .B2(n20038), .A(n20037), .ZN(P1_U2936) );
  AOI22_X1 U22929 ( .A1(n13133), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20064), .ZN(n20041) );
  NAND2_X1 U22930 ( .A1(n20052), .A2(n20040), .ZN(n20054) );
  NAND2_X1 U22931 ( .A1(n20041), .A2(n20054), .ZN(P1_U2946) );
  AOI22_X1 U22932 ( .A1(n13133), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20043) );
  NAND2_X1 U22933 ( .A1(n20052), .A2(n20042), .ZN(n20056) );
  NAND2_X1 U22934 ( .A1(n20043), .A2(n20056), .ZN(P1_U2947) );
  AOI22_X1 U22935 ( .A1(n13133), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20045) );
  NAND2_X1 U22936 ( .A1(n20052), .A2(n20044), .ZN(n20058) );
  NAND2_X1 U22937 ( .A1(n20045), .A2(n20058), .ZN(P1_U2948) );
  AOI22_X1 U22938 ( .A1(n13133), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20047) );
  NAND2_X1 U22939 ( .A1(n20052), .A2(n20046), .ZN(n20060) );
  NAND2_X1 U22940 ( .A1(n20047), .A2(n20060), .ZN(P1_U2949) );
  AOI22_X1 U22941 ( .A1(n13133), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20049) );
  NAND2_X1 U22942 ( .A1(n20052), .A2(n20048), .ZN(n20062) );
  NAND2_X1 U22943 ( .A1(n20049), .A2(n20062), .ZN(P1_U2950) );
  AOI22_X1 U22944 ( .A1(n13133), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20064), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20053) );
  INV_X1 U22945 ( .A(n20050), .ZN(n20051) );
  NAND2_X1 U22946 ( .A1(n20052), .A2(n20051), .ZN(n20065) );
  NAND2_X1 U22947 ( .A1(n20053), .A2(n20065), .ZN(P1_U2951) );
  AOI22_X1 U22948 ( .A1(n13133), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20064), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20055) );
  NAND2_X1 U22949 ( .A1(n20055), .A2(n20054), .ZN(P1_U2961) );
  AOI22_X1 U22950 ( .A1(n13133), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20064), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20057) );
  NAND2_X1 U22951 ( .A1(n20057), .A2(n20056), .ZN(P1_U2962) );
  AOI22_X1 U22952 ( .A1(n13133), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20064), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20059) );
  NAND2_X1 U22953 ( .A1(n20059), .A2(n20058), .ZN(P1_U2963) );
  AOI22_X1 U22954 ( .A1(n13133), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20064), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20061) );
  NAND2_X1 U22955 ( .A1(n20061), .A2(n20060), .ZN(P1_U2964) );
  AOI22_X1 U22956 ( .A1(n13133), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20064), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20063) );
  NAND2_X1 U22957 ( .A1(n20063), .A2(n20062), .ZN(P1_U2965) );
  AOI22_X1 U22958 ( .A1(n13133), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20064), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20066) );
  NAND2_X1 U22959 ( .A1(n20066), .A2(n20065), .ZN(P1_U2966) );
  AOI22_X1 U22960 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20073) );
  AOI21_X1 U22961 ( .B1(n20068), .B2(n20067), .A(n9699), .ZN(n20096) );
  AOI22_X1 U22962 ( .A1(n20096), .A2(n20071), .B1(n20070), .B2(n20069), .ZN(
        n20072) );
  OAI211_X1 U22963 ( .C1(n20075), .C2(n20074), .A(n20073), .B(n20072), .ZN(
        P1_U2995) );
  AOI22_X1 U22964 ( .A1(n20086), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20128), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n20081) );
  AOI21_X1 U22965 ( .B1(n20077), .B2(n20135), .A(n20076), .ZN(n20129) );
  AOI22_X1 U22966 ( .A1(n20071), .A2(n20129), .B1(n20079), .B2(n20078), .ZN(
        n20080) );
  OAI211_X1 U22967 ( .C1(n20149), .C2(n20082), .A(n20081), .B(n20080), .ZN(
        P1_U2998) );
  OAI22_X1 U22968 ( .A1(n20149), .A2(n20083), .B1(n20114), .B2(n20844), .ZN(
        n20084) );
  INV_X1 U22969 ( .A(n20084), .ZN(n20088) );
  OAI21_X1 U22970 ( .B1(n20086), .B2(n20085), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20087) );
  OAI211_X1 U22971 ( .C1(n20090), .C2(n20089), .A(n20088), .B(n20087), .ZN(
        P1_U2999) );
  AND2_X1 U22972 ( .A1(n20092), .A2(n20091), .ZN(n20118) );
  AOI211_X1 U22973 ( .C1(n20113), .C2(n20093), .A(n20118), .B(n20111), .ZN(
        n20108) );
  OAI22_X1 U22974 ( .A1(n20094), .A2(n20116), .B1(n20781), .B2(n20114), .ZN(
        n20095) );
  AOI21_X1 U22975 ( .B1(n20096), .B2(n20130), .A(n20095), .ZN(n20099) );
  OAI211_X1 U22976 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20103), .B(n20097), .ZN(n20098) );
  OAI211_X1 U22977 ( .C1(n20108), .C2(n20100), .A(n20099), .B(n20098), .ZN(
        P1_U3027) );
  AOI21_X1 U22978 ( .B1(n20102), .B2(n20131), .A(n20101), .ZN(n20106) );
  AOI22_X1 U22979 ( .A1(n20104), .A2(n20130), .B1(n20107), .B2(n20103), .ZN(
        n20105) );
  OAI211_X1 U22980 ( .C1(n20108), .C2(n20107), .A(n20106), .B(n20105), .ZN(
        P1_U3028) );
  NOR3_X1 U22981 ( .A1(n20110), .A2(n20135), .A3(n20109), .ZN(n20112) );
  AOI211_X1 U22982 ( .C1(n20135), .C2(n20113), .A(n20112), .B(n20111), .ZN(
        n20124) );
  INV_X1 U22983 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20778) );
  OAI22_X1 U22984 ( .A1(n20116), .A2(n20115), .B1(n20778), .B2(n20114), .ZN(
        n20117) );
  NOR2_X1 U22985 ( .A1(n20118), .A2(n20117), .ZN(n20119) );
  OAI21_X1 U22986 ( .B1(n20121), .B2(n20120), .A(n20119), .ZN(n20122) );
  INV_X1 U22987 ( .A(n20122), .ZN(n20123) );
  OAI221_X1 U22988 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20125), .C1(
        n11873), .C2(n20124), .A(n20123), .ZN(P1_U3029) );
  NAND2_X1 U22989 ( .A1(n20127), .A2(n20126), .ZN(n20136) );
  AOI222_X1 U22990 ( .A1(n20132), .A2(n20131), .B1(n20130), .B2(n20129), .C1(
        P1_REIP_REG_1__SCAN_IN), .C2(n20128), .ZN(n20133) );
  OAI221_X1 U22991 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20136), .C1(
        n20135), .C2(n20134), .A(n20133), .ZN(P1_U3030) );
  NOR2_X1 U22992 ( .A1(n20138), .A2(n20137), .ZN(P1_U3032) );
  OR2_X1 U22993 ( .A1(n20431), .A2(n20482), .ZN(n20307) );
  NAND2_X1 U22994 ( .A1(n20151), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20639) );
  NAND2_X1 U22995 ( .A1(n20197), .A2(n20639), .ZN(n20232) );
  OAI21_X1 U22996 ( .B1(n20228), .B2(n20170), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20142) );
  NAND2_X1 U22997 ( .A1(n20142), .A2(n20701), .ZN(n20153) );
  INV_X1 U22998 ( .A(n12991), .ZN(n20143) );
  NAND2_X1 U22999 ( .A1(n9719), .A2(n14385), .ZN(n20152) );
  INV_X1 U23000 ( .A(n20152), .ZN(n20144) );
  NAND2_X1 U23001 ( .A1(n20234), .A2(n20429), .ZN(n20268) );
  OR2_X1 U23002 ( .A1(n20564), .A2(n20268), .ZN(n20195) );
  INV_X1 U23003 ( .A(n20195), .ZN(n20171) );
  OAI22_X1 U23004 ( .A1(n20153), .A2(n20144), .B1(n20171), .B2(n20570), .ZN(
        n20145) );
  NOR2_X2 U23005 ( .A1(n20146), .A2(n20168), .ZN(n20691) );
  NOR2_X2 U23006 ( .A1(n14158), .A2(n20149), .ZN(n20199) );
  AOI22_X1 U23007 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20148), .B1(DATAI_24_), 
        .B2(n20199), .ZN(n20652) );
  INV_X1 U23008 ( .A(n20652), .ZN(n20702) );
  AOI22_X1 U23009 ( .A1(n20171), .A2(n20691), .B1(n20170), .B2(n20702), .ZN(
        n20155) );
  NAND2_X1 U23010 ( .A1(n20150), .A2(n20197), .ZN(n20493) );
  NOR2_X1 U23011 ( .A1(n20151), .A2(n11268), .ZN(n20483) );
  INV_X1 U23012 ( .A(n20483), .ZN(n20432) );
  OAI22_X1 U23013 ( .A1(n20153), .A2(n20152), .B1(n20432), .B2(n20307), .ZN(
        n20200) );
  AOI22_X1 U23014 ( .A1(DATAI_16_), .A2(n20199), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20148), .ZN(n20705) );
  INV_X1 U23015 ( .A(n20705), .ZN(n20649) );
  AOI22_X1 U23016 ( .A1(n20692), .A2(n20200), .B1(n20228), .B2(n20649), .ZN(
        n20154) );
  OAI211_X1 U23017 ( .C1(n20204), .C2(n20156), .A(n20155), .B(n20154), .ZN(
        P1_U3033) );
  NAND2_X1 U23018 ( .A1(n9614), .A2(n20194), .ZN(n20577) );
  OAI22_X1 U23019 ( .A1(n20751), .A2(n20656), .B1(n20195), .B2(n20577), .ZN(
        n20158) );
  INV_X1 U23020 ( .A(n20158), .ZN(n20161) );
  NAND2_X1 U23021 ( .A1(n20159), .A2(n20197), .ZN(n20497) );
  AOI22_X1 U23022 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20148), .B1(DATAI_17_), 
        .B2(n20199), .ZN(n20711) );
  INV_X1 U23023 ( .A(n20711), .ZN(n20653) );
  AOI22_X1 U23024 ( .A1(n20707), .A2(n20200), .B1(n20228), .B2(n20653), .ZN(
        n20160) );
  OAI211_X1 U23025 ( .C1(n20204), .C2(n11235), .A(n20161), .B(n20160), .ZN(
        P1_U3034) );
  AOI22_X1 U23026 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20148), .B1(DATAI_26_), 
        .B2(n20199), .ZN(n20660) );
  NAND2_X1 U23027 ( .A1(n20162), .A2(n20194), .ZN(n20581) );
  OAI22_X1 U23028 ( .A1(n20751), .A2(n20660), .B1(n20195), .B2(n20581), .ZN(
        n20163) );
  INV_X1 U23029 ( .A(n20163), .ZN(n20166) );
  NAND2_X1 U23030 ( .A1(n20164), .A2(n20197), .ZN(n20501) );
  AOI22_X1 U23031 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20148), .B1(DATAI_18_), 
        .B2(n20199), .ZN(n20717) );
  INV_X1 U23032 ( .A(n20717), .ZN(n20657) );
  AOI22_X1 U23033 ( .A1(n20713), .A2(n20200), .B1(n20228), .B2(n20657), .ZN(
        n20165) );
  OAI211_X1 U23034 ( .C1(n20204), .C2(n20167), .A(n20166), .B(n20165), .ZN(
        P1_U3035) );
  INV_X1 U23035 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20175) );
  NOR2_X2 U23036 ( .A1(n20169), .A2(n20168), .ZN(n20718) );
  AOI22_X1 U23037 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20148), .B1(DATAI_27_), 
        .B2(n20199), .ZN(n20664) );
  INV_X1 U23038 ( .A(n20664), .ZN(n20720) );
  AOI22_X1 U23039 ( .A1(n20171), .A2(n20718), .B1(n20170), .B2(n20720), .ZN(
        n20174) );
  NAND2_X1 U23040 ( .A1(n20172), .A2(n20197), .ZN(n20505) );
  AOI22_X1 U23041 ( .A1(DATAI_19_), .A2(n20199), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20148), .ZN(n20723) );
  INV_X1 U23042 ( .A(n20723), .ZN(n20661) );
  AOI22_X1 U23043 ( .A1(n20719), .A2(n20200), .B1(n20228), .B2(n20661), .ZN(
        n20173) );
  OAI211_X1 U23044 ( .C1(n20204), .C2(n20175), .A(n20174), .B(n20173), .ZN(
        P1_U3036) );
  INV_X1 U23045 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20181) );
  AOI22_X1 U23046 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20148), .B1(DATAI_28_), 
        .B2(n20199), .ZN(n20668) );
  NAND2_X1 U23047 ( .A1(n20176), .A2(n20194), .ZN(n20588) );
  OAI22_X1 U23048 ( .A1(n20751), .A2(n20668), .B1(n20195), .B2(n20588), .ZN(
        n20177) );
  INV_X1 U23049 ( .A(n20177), .ZN(n20180) );
  NAND2_X1 U23050 ( .A1(n20178), .A2(n20197), .ZN(n20509) );
  AOI22_X1 U23051 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20148), .B1(DATAI_20_), 
        .B2(n20199), .ZN(n20729) );
  INV_X1 U23052 ( .A(n20729), .ZN(n20665) );
  AOI22_X1 U23053 ( .A1(n20725), .A2(n20200), .B1(n20228), .B2(n20665), .ZN(
        n20179) );
  OAI211_X1 U23054 ( .C1(n20204), .C2(n20181), .A(n20180), .B(n20179), .ZN(
        P1_U3037) );
  INV_X1 U23055 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20187) );
  NAND2_X1 U23056 ( .A1(n20182), .A2(n20194), .ZN(n20592) );
  OAI22_X1 U23057 ( .A1(n20751), .A2(n20672), .B1(n20195), .B2(n20592), .ZN(
        n20183) );
  INV_X1 U23058 ( .A(n20183), .ZN(n20186) );
  NAND2_X1 U23059 ( .A1(n20184), .A2(n20197), .ZN(n20514) );
  AOI22_X1 U23060 ( .A1(DATAI_21_), .A2(n20199), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20148), .ZN(n20735) );
  INV_X1 U23061 ( .A(n20735), .ZN(n20669) );
  AOI22_X1 U23062 ( .A1(n20731), .A2(n20200), .B1(n20228), .B2(n20669), .ZN(
        n20185) );
  OAI211_X1 U23063 ( .C1(n20204), .C2(n20187), .A(n20186), .B(n20185), .ZN(
        P1_U3038) );
  AOI22_X1 U23064 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20148), .B1(DATAI_30_), 
        .B2(n20199), .ZN(n20676) );
  NAND2_X1 U23065 ( .A1(n20188), .A2(n20194), .ZN(n20596) );
  OAI22_X1 U23066 ( .A1(n20751), .A2(n20676), .B1(n20195), .B2(n20596), .ZN(
        n20189) );
  INV_X1 U23067 ( .A(n20189), .ZN(n20192) );
  NAND2_X1 U23068 ( .A1(n20190), .A2(n20197), .ZN(n20518) );
  AOI22_X1 U23069 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20148), .B1(DATAI_22_), 
        .B2(n20199), .ZN(n20741) );
  INV_X1 U23070 ( .A(n20741), .ZN(n20673) );
  AOI22_X1 U23071 ( .A1(n20737), .A2(n20200), .B1(n20228), .B2(n20673), .ZN(
        n20191) );
  OAI211_X1 U23072 ( .C1(n20204), .C2(n20193), .A(n20192), .B(n20191), .ZN(
        P1_U3039) );
  AOI22_X1 U23073 ( .A1(DATAI_31_), .A2(n20199), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20148), .ZN(n20684) );
  NAND2_X1 U23074 ( .A1(n11154), .A2(n20194), .ZN(n20601) );
  OAI22_X1 U23075 ( .A1(n20751), .A2(n20684), .B1(n20195), .B2(n20601), .ZN(
        n20196) );
  INV_X1 U23076 ( .A(n20196), .ZN(n20202) );
  NAND2_X1 U23077 ( .A1(n20198), .A2(n20197), .ZN(n20525) );
  AOI22_X1 U23078 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20148), .B1(DATAI_23_), 
        .B2(n20199), .ZN(n20752) );
  INV_X1 U23079 ( .A(n20752), .ZN(n20679) );
  AOI22_X1 U23080 ( .A1(n20744), .A2(n20200), .B1(n20228), .B2(n20679), .ZN(
        n20201) );
  OAI211_X1 U23081 ( .C1(n20204), .C2(n20203), .A(n20202), .B(n20201), .ZN(
        P1_U3040) );
  INV_X1 U23082 ( .A(n20205), .ZN(n20612) );
  NOR2_X1 U23083 ( .A1(n20268), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20209) );
  INV_X1 U23084 ( .A(n20209), .ZN(n20206) );
  NOR2_X1 U23085 ( .A1(n20611), .A2(n20206), .ZN(n20226) );
  AOI21_X1 U23086 ( .B1(n9719), .B2(n20612), .A(n20226), .ZN(n20207) );
  OAI22_X1 U23087 ( .A1(n20207), .A2(n20693), .B1(n20206), .B2(n11268), .ZN(
        n20227) );
  AOI22_X1 U23088 ( .A1(n20692), .A2(n20227), .B1(n20691), .B2(n20226), .ZN(
        n20211) );
  OAI211_X1 U23089 ( .C1(n20276), .C2(n14399), .A(n20701), .B(n20207), .ZN(
        n20208) );
  OAI211_X1 U23090 ( .C1(n20617), .C2(n20209), .A(n20699), .B(n20208), .ZN(
        n20229) );
  AOI22_X1 U23091 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20229), .B1(
        n20222), .B2(n20649), .ZN(n20210) );
  OAI211_X1 U23092 ( .C1(n20652), .C2(n20225), .A(n20211), .B(n20210), .ZN(
        P1_U3041) );
  AOI22_X1 U23093 ( .A1(n20227), .A2(n20707), .B1(n20706), .B2(n20226), .ZN(
        n20213) );
  AOI22_X1 U23094 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20229), .B1(
        n20222), .B2(n20653), .ZN(n20212) );
  OAI211_X1 U23095 ( .C1(n20656), .C2(n20225), .A(n20213), .B(n20212), .ZN(
        P1_U3042) );
  AOI22_X1 U23096 ( .A1(n20227), .A2(n20713), .B1(n20712), .B2(n20226), .ZN(
        n20215) );
  INV_X1 U23097 ( .A(n20660), .ZN(n20714) );
  AOI22_X1 U23098 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20229), .B1(
        n20228), .B2(n20714), .ZN(n20214) );
  OAI211_X1 U23099 ( .C1(n20717), .C2(n20260), .A(n20215), .B(n20214), .ZN(
        P1_U3043) );
  AOI22_X1 U23100 ( .A1(n20719), .A2(n20227), .B1(n20718), .B2(n20226), .ZN(
        n20217) );
  AOI22_X1 U23101 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20229), .B1(
        n20222), .B2(n20661), .ZN(n20216) );
  OAI211_X1 U23102 ( .C1(n20664), .C2(n20225), .A(n20217), .B(n20216), .ZN(
        P1_U3044) );
  AOI22_X1 U23103 ( .A1(n20227), .A2(n20725), .B1(n20724), .B2(n20226), .ZN(
        n20219) );
  AOI22_X1 U23104 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20229), .B1(
        n20222), .B2(n20665), .ZN(n20218) );
  OAI211_X1 U23105 ( .C1(n20668), .C2(n20225), .A(n20219), .B(n20218), .ZN(
        P1_U3045) );
  AOI22_X1 U23106 ( .A1(n20227), .A2(n20731), .B1(n20730), .B2(n20226), .ZN(
        n20221) );
  AOI22_X1 U23107 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20229), .B1(
        n20222), .B2(n20669), .ZN(n20220) );
  OAI211_X1 U23108 ( .C1(n20672), .C2(n20225), .A(n20221), .B(n20220), .ZN(
        P1_U3046) );
  AOI22_X1 U23109 ( .A1(n20227), .A2(n20737), .B1(n20736), .B2(n20226), .ZN(
        n20224) );
  AOI22_X1 U23110 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20229), .B1(
        n20222), .B2(n20673), .ZN(n20223) );
  OAI211_X1 U23111 ( .C1(n20676), .C2(n20225), .A(n20224), .B(n20223), .ZN(
        P1_U3047) );
  AOI22_X1 U23112 ( .A1(n20227), .A2(n20744), .B1(n20743), .B2(n20226), .ZN(
        n20231) );
  INV_X1 U23113 ( .A(n20684), .ZN(n20746) );
  AOI22_X1 U23114 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20229), .B1(
        n20228), .B2(n20746), .ZN(n20230) );
  OAI211_X1 U23115 ( .C1(n20752), .C2(n20260), .A(n20231), .B(n20230), .ZN(
        P1_U3048) );
  NOR2_X1 U23116 ( .A1(n20689), .A2(n20268), .ZN(n20271) );
  NAND2_X1 U23117 ( .A1(n20611), .A2(n20271), .ZN(n20259) );
  INV_X1 U23118 ( .A(n20259), .ZN(n20247) );
  AOI22_X1 U23119 ( .A1(n20247), .A2(n20691), .B1(n20300), .B2(n20649), .ZN(
        n20240) );
  AOI21_X1 U23120 ( .B1(n20291), .B2(n20260), .A(n14399), .ZN(n20233) );
  NOR2_X1 U23121 ( .A1(n20233), .A2(n20693), .ZN(n20236) );
  NAND2_X1 U23122 ( .A1(n9719), .A2(n20638), .ZN(n20237) );
  AOI22_X1 U23123 ( .A1(n20236), .A2(n20237), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20259), .ZN(n20235) );
  NAND2_X1 U23124 ( .A1(n20482), .A2(n20234), .ZN(n20360) );
  NAND2_X1 U23125 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20360), .ZN(n20367) );
  NAND3_X1 U23126 ( .A1(n20490), .A2(n20235), .A3(n20367), .ZN(n20263) );
  INV_X1 U23127 ( .A(n20236), .ZN(n20238) );
  OAI22_X1 U23128 ( .A1(n20238), .A2(n20237), .B1(n20432), .B2(n20360), .ZN(
        n20262) );
  AOI22_X1 U23129 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20263), .B1(
        n20692), .B2(n20262), .ZN(n20239) );
  OAI211_X1 U23130 ( .C1(n20652), .C2(n20260), .A(n20240), .B(n20239), .ZN(
        P1_U3049) );
  OAI22_X1 U23131 ( .A1(n20291), .A2(n20711), .B1(n20577), .B2(n20259), .ZN(
        n20241) );
  INV_X1 U23132 ( .A(n20241), .ZN(n20243) );
  AOI22_X1 U23133 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20263), .B1(
        n20707), .B2(n20262), .ZN(n20242) );
  OAI211_X1 U23134 ( .C1(n20656), .C2(n20260), .A(n20243), .B(n20242), .ZN(
        P1_U3050) );
  OAI22_X1 U23135 ( .A1(n20260), .A2(n20660), .B1(n20581), .B2(n20259), .ZN(
        n20244) );
  INV_X1 U23136 ( .A(n20244), .ZN(n20246) );
  AOI22_X1 U23137 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20263), .B1(
        n20713), .B2(n20262), .ZN(n20245) );
  OAI211_X1 U23138 ( .C1(n20717), .C2(n20291), .A(n20246), .B(n20245), .ZN(
        P1_U3051) );
  AOI22_X1 U23139 ( .A1(n20247), .A2(n20718), .B1(n20300), .B2(n20661), .ZN(
        n20249) );
  AOI22_X1 U23140 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20263), .B1(
        n20719), .B2(n20262), .ZN(n20248) );
  OAI211_X1 U23141 ( .C1(n20664), .C2(n20260), .A(n20249), .B(n20248), .ZN(
        P1_U3052) );
  OAI22_X1 U23142 ( .A1(n20260), .A2(n20668), .B1(n20588), .B2(n20259), .ZN(
        n20250) );
  INV_X1 U23143 ( .A(n20250), .ZN(n20252) );
  AOI22_X1 U23144 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20263), .B1(
        n20725), .B2(n20262), .ZN(n20251) );
  OAI211_X1 U23145 ( .C1(n20729), .C2(n20291), .A(n20252), .B(n20251), .ZN(
        P1_U3053) );
  OAI22_X1 U23146 ( .A1(n20291), .A2(n20735), .B1(n20592), .B2(n20259), .ZN(
        n20253) );
  INV_X1 U23147 ( .A(n20253), .ZN(n20255) );
  AOI22_X1 U23148 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20263), .B1(
        n20731), .B2(n20262), .ZN(n20254) );
  OAI211_X1 U23149 ( .C1(n20672), .C2(n20260), .A(n20255), .B(n20254), .ZN(
        P1_U3054) );
  OAI22_X1 U23150 ( .A1(n20260), .A2(n20676), .B1(n20596), .B2(n20259), .ZN(
        n20256) );
  INV_X1 U23151 ( .A(n20256), .ZN(n20258) );
  AOI22_X1 U23152 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20263), .B1(
        n20737), .B2(n20262), .ZN(n20257) );
  OAI211_X1 U23153 ( .C1(n20741), .C2(n20291), .A(n20258), .B(n20257), .ZN(
        P1_U3055) );
  OAI22_X1 U23154 ( .A1(n20260), .A2(n20684), .B1(n20601), .B2(n20259), .ZN(
        n20261) );
  INV_X1 U23155 ( .A(n20261), .ZN(n20265) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20263), .B1(
        n20744), .B2(n20262), .ZN(n20264) );
  OAI211_X1 U23157 ( .C1(n20752), .C2(n20291), .A(n20265), .B(n20264), .ZN(
        P1_U3056) );
  INV_X1 U23158 ( .A(n20276), .ZN(n20266) );
  OAI21_X1 U23159 ( .B1(n20266), .B2(n20693), .A(n20538), .ZN(n20274) );
  AND2_X1 U23160 ( .A1(n20267), .A2(n11289), .ZN(n20686) );
  INV_X1 U23161 ( .A(n20268), .ZN(n20269) );
  AND2_X1 U23162 ( .A1(n20529), .A2(n20269), .ZN(n20285) );
  AOI21_X1 U23163 ( .B1(n9719), .B2(n20686), .A(n20285), .ZN(n20273) );
  INV_X1 U23164 ( .A(n20273), .ZN(n20270) );
  AOI22_X1 U23165 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20271), .B1(n20274), 
        .B2(n20270), .ZN(n20304) );
  AOI22_X1 U23166 ( .A1(n20285), .A2(n20691), .B1(n20300), .B2(n20702), .ZN(
        n20278) );
  OAI21_X1 U23167 ( .B1(n20701), .B2(n20271), .A(n20699), .ZN(n20272) );
  AOI21_X1 U23168 ( .B1(n20274), .B2(n20273), .A(n20272), .ZN(n20275) );
  AOI22_X1 U23169 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20301), .B1(
        n20329), .B2(n20649), .ZN(n20277) );
  OAI211_X1 U23170 ( .C1(n20304), .C2(n20493), .A(n20278), .B(n20277), .ZN(
        P1_U3057) );
  INV_X1 U23171 ( .A(n20285), .ZN(n20298) );
  OAI22_X1 U23172 ( .A1(n20325), .A2(n20711), .B1(n20577), .B2(n20298), .ZN(
        n20279) );
  INV_X1 U23173 ( .A(n20279), .ZN(n20281) );
  INV_X1 U23174 ( .A(n20656), .ZN(n20708) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20301), .B1(
        n20300), .B2(n20708), .ZN(n20280) );
  OAI211_X1 U23176 ( .C1(n20304), .C2(n20497), .A(n20281), .B(n20280), .ZN(
        P1_U3058) );
  OAI22_X1 U23177 ( .A1(n20325), .A2(n20717), .B1(n20581), .B2(n20298), .ZN(
        n20282) );
  INV_X1 U23178 ( .A(n20282), .ZN(n20284) );
  AOI22_X1 U23179 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20301), .B1(
        n20300), .B2(n20714), .ZN(n20283) );
  OAI211_X1 U23180 ( .C1(n20304), .C2(n20501), .A(n20284), .B(n20283), .ZN(
        P1_U3059) );
  AOI22_X1 U23181 ( .A1(n20285), .A2(n20718), .B1(n20329), .B2(n20661), .ZN(
        n20287) );
  AOI22_X1 U23182 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20301), .B1(
        n20300), .B2(n20720), .ZN(n20286) );
  OAI211_X1 U23183 ( .C1(n20304), .C2(n20505), .A(n20287), .B(n20286), .ZN(
        P1_U3060) );
  OAI22_X1 U23184 ( .A1(n20325), .A2(n20729), .B1(n20588), .B2(n20298), .ZN(
        n20288) );
  INV_X1 U23185 ( .A(n20288), .ZN(n20290) );
  INV_X1 U23186 ( .A(n20668), .ZN(n20726) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20301), .B1(
        n20300), .B2(n20726), .ZN(n20289) );
  OAI211_X1 U23188 ( .C1(n20304), .C2(n20509), .A(n20290), .B(n20289), .ZN(
        P1_U3061) );
  OAI22_X1 U23189 ( .A1(n20291), .A2(n20672), .B1(n20592), .B2(n20298), .ZN(
        n20292) );
  INV_X1 U23190 ( .A(n20292), .ZN(n20294) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20301), .B1(
        n20329), .B2(n20669), .ZN(n20293) );
  OAI211_X1 U23192 ( .C1(n20304), .C2(n20514), .A(n20294), .B(n20293), .ZN(
        P1_U3062) );
  OAI22_X1 U23193 ( .A1(n20325), .A2(n20741), .B1(n20596), .B2(n20298), .ZN(
        n20295) );
  INV_X1 U23194 ( .A(n20295), .ZN(n20297) );
  INV_X1 U23195 ( .A(n20676), .ZN(n20738) );
  AOI22_X1 U23196 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20301), .B1(
        n20300), .B2(n20738), .ZN(n20296) );
  OAI211_X1 U23197 ( .C1(n20304), .C2(n20518), .A(n20297), .B(n20296), .ZN(
        P1_U3063) );
  OAI22_X1 U23198 ( .A1(n20325), .A2(n20752), .B1(n20601), .B2(n20298), .ZN(
        n20299) );
  INV_X1 U23199 ( .A(n20299), .ZN(n20303) );
  AOI22_X1 U23200 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20301), .B1(
        n20300), .B2(n20746), .ZN(n20302) );
  OAI211_X1 U23201 ( .C1(n20304), .C2(n20525), .A(n20303), .B(n20302), .ZN(
        P1_U3064) );
  OR2_X1 U23202 ( .A1(n12991), .A2(n20305), .ZN(n20401) );
  INV_X1 U23203 ( .A(n20401), .ZN(n20334) );
  NAND3_X1 U23204 ( .A1(n20334), .A2(n20701), .A3(n14385), .ZN(n20306) );
  OAI21_X1 U23205 ( .B1(n20639), .B2(n20307), .A(n20306), .ZN(n20328) );
  AOI22_X1 U23206 ( .A1(n20692), .A2(n20328), .B1(n20691), .B2(n10159), .ZN(
        n20313) );
  NAND2_X1 U23207 ( .A1(n20325), .A2(n20358), .ZN(n20308) );
  AOI22_X1 U23208 ( .A1(n20308), .A2(P1_STATEBS16_REG_SCAN_IN), .B1(n20334), 
        .B2(n14385), .ZN(n20309) );
  NOR2_X1 U23209 ( .A1(n20309), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20311) );
  INV_X1 U23210 ( .A(n20358), .ZN(n20322) );
  AOI22_X1 U23211 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20330), .B1(
        n20322), .B2(n20649), .ZN(n20312) );
  OAI211_X1 U23212 ( .C1(n20652), .C2(n20325), .A(n20313), .B(n20312), .ZN(
        P1_U3065) );
  AOI22_X1 U23213 ( .A1(n20328), .A2(n20707), .B1(n20706), .B2(n10159), .ZN(
        n20315) );
  AOI22_X1 U23214 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20330), .B1(
        n20322), .B2(n20653), .ZN(n20314) );
  OAI211_X1 U23215 ( .C1(n20656), .C2(n20325), .A(n20315), .B(n20314), .ZN(
        P1_U3066) );
  AOI22_X1 U23216 ( .A1(n20328), .A2(n20713), .B1(n20712), .B2(n10159), .ZN(
        n20317) );
  AOI22_X1 U23217 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20330), .B1(
        n20329), .B2(n20714), .ZN(n20316) );
  OAI211_X1 U23218 ( .C1(n20717), .C2(n20358), .A(n20317), .B(n20316), .ZN(
        P1_U3067) );
  AOI22_X1 U23219 ( .A1(n20719), .A2(n20328), .B1(n20718), .B2(n10159), .ZN(
        n20319) );
  AOI22_X1 U23220 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20330), .B1(
        n20322), .B2(n20661), .ZN(n20318) );
  OAI211_X1 U23221 ( .C1(n20664), .C2(n20325), .A(n20319), .B(n20318), .ZN(
        P1_U3068) );
  AOI22_X1 U23222 ( .A1(n20328), .A2(n20725), .B1(n20724), .B2(n10159), .ZN(
        n20321) );
  AOI22_X1 U23223 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20330), .B1(
        n20329), .B2(n20726), .ZN(n20320) );
  OAI211_X1 U23224 ( .C1(n20729), .C2(n20358), .A(n20321), .B(n20320), .ZN(
        P1_U3069) );
  AOI22_X1 U23225 ( .A1(n20328), .A2(n20731), .B1(n20730), .B2(n10159), .ZN(
        n20324) );
  AOI22_X1 U23226 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20330), .B1(
        n20322), .B2(n20669), .ZN(n20323) );
  OAI211_X1 U23227 ( .C1(n20672), .C2(n20325), .A(n20324), .B(n20323), .ZN(
        P1_U3070) );
  AOI22_X1 U23228 ( .A1(n20328), .A2(n20737), .B1(n20736), .B2(n10159), .ZN(
        n20327) );
  AOI22_X1 U23229 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20330), .B1(
        n20329), .B2(n20738), .ZN(n20326) );
  OAI211_X1 U23230 ( .C1(n20741), .C2(n20358), .A(n20327), .B(n20326), .ZN(
        P1_U3071) );
  AOI22_X1 U23231 ( .A1(n20328), .A2(n20744), .B1(n20743), .B2(n10159), .ZN(
        n20332) );
  AOI22_X1 U23232 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20330), .B1(
        n20329), .B2(n20746), .ZN(n20331) );
  OAI211_X1 U23233 ( .C1(n20752), .C2(n20358), .A(n20332), .B(n20331), .ZN(
        P1_U3072) );
  NOR2_X1 U23234 ( .A1(n20333), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20338) );
  INV_X1 U23235 ( .A(n20338), .ZN(n20335) );
  NOR2_X1 U23236 ( .A1(n20611), .A2(n20335), .ZN(n20353) );
  AOI21_X1 U23237 ( .B1(n20334), .B2(n20612), .A(n20353), .ZN(n20336) );
  OAI22_X1 U23238 ( .A1(n20336), .A2(n20693), .B1(n20335), .B2(n11268), .ZN(
        n20354) );
  AOI22_X1 U23239 ( .A1(n20692), .A2(n20354), .B1(n20691), .B2(n20353), .ZN(
        n20340) );
  OAI211_X1 U23240 ( .C1(n20403), .C2(n14399), .A(n20701), .B(n20336), .ZN(
        n20337) );
  OAI211_X1 U23241 ( .C1(n20701), .C2(n20338), .A(n20699), .B(n20337), .ZN(
        n20355) );
  AOI22_X1 U23242 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20355), .B1(
        n20393), .B2(n20649), .ZN(n20339) );
  OAI211_X1 U23243 ( .C1(n20652), .C2(n20358), .A(n20340), .B(n20339), .ZN(
        P1_U3073) );
  AOI22_X1 U23244 ( .A1(n20354), .A2(n20707), .B1(n20706), .B2(n20353), .ZN(
        n20342) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20355), .B1(
        n20393), .B2(n20653), .ZN(n20341) );
  OAI211_X1 U23246 ( .C1(n20656), .C2(n20358), .A(n20342), .B(n20341), .ZN(
        P1_U3074) );
  AOI22_X1 U23247 ( .A1(n20354), .A2(n20713), .B1(n20712), .B2(n20353), .ZN(
        n20344) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20355), .B1(
        n20393), .B2(n20657), .ZN(n20343) );
  OAI211_X1 U23249 ( .C1(n20660), .C2(n20358), .A(n20344), .B(n20343), .ZN(
        P1_U3075) );
  AOI22_X1 U23250 ( .A1(n20719), .A2(n20354), .B1(n20718), .B2(n20353), .ZN(
        n20346) );
  AOI22_X1 U23251 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20355), .B1(
        n20393), .B2(n20661), .ZN(n20345) );
  OAI211_X1 U23252 ( .C1(n20664), .C2(n20358), .A(n20346), .B(n20345), .ZN(
        P1_U3076) );
  AOI22_X1 U23253 ( .A1(n20354), .A2(n20725), .B1(n20724), .B2(n20353), .ZN(
        n20348) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20355), .B1(
        n20393), .B2(n20665), .ZN(n20347) );
  OAI211_X1 U23255 ( .C1(n20668), .C2(n20358), .A(n20348), .B(n20347), .ZN(
        P1_U3077) );
  AOI22_X1 U23256 ( .A1(n20354), .A2(n20731), .B1(n20730), .B2(n20353), .ZN(
        n20350) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20355), .B1(
        n20393), .B2(n20669), .ZN(n20349) );
  OAI211_X1 U23258 ( .C1(n20672), .C2(n20358), .A(n20350), .B(n20349), .ZN(
        P1_U3078) );
  AOI22_X1 U23259 ( .A1(n20354), .A2(n20737), .B1(n20736), .B2(n20353), .ZN(
        n20352) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20355), .B1(
        n20393), .B2(n20673), .ZN(n20351) );
  OAI211_X1 U23261 ( .C1(n20676), .C2(n20358), .A(n20352), .B(n20351), .ZN(
        P1_U3079) );
  AOI22_X1 U23262 ( .A1(n20354), .A2(n20744), .B1(n20743), .B2(n20353), .ZN(
        n20357) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20355), .B1(
        n20393), .B2(n20679), .ZN(n20356) );
  OAI211_X1 U23264 ( .C1(n20684), .C2(n20358), .A(n20357), .B(n20356), .ZN(
        P1_U3080) );
  NAND3_X1 U23265 ( .A1(n20391), .A2(n20380), .A3(n20617), .ZN(n20359) );
  NAND2_X1 U23266 ( .A1(n20359), .A2(n20566), .ZN(n20366) );
  NOR2_X1 U23267 ( .A1(n20401), .A2(n14385), .ZN(n20364) );
  INV_X1 U23268 ( .A(n20360), .ZN(n20362) );
  INV_X1 U23269 ( .A(n20639), .ZN(n20361) );
  NAND2_X1 U23270 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20363), .ZN(
        n20404) );
  NOR2_X1 U23271 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20404), .ZN(
        n20377) );
  AOI22_X1 U23272 ( .A1(n20377), .A2(n20691), .B1(n20393), .B2(n20702), .ZN(
        n20370) );
  INV_X1 U23273 ( .A(n20364), .ZN(n20365) );
  INV_X1 U23274 ( .A(n20377), .ZN(n20390) );
  AOI22_X1 U23275 ( .A1(n20366), .A2(n20365), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20390), .ZN(n20368) );
  NAND3_X1 U23276 ( .A1(n20647), .A2(n20368), .A3(n20367), .ZN(n20394) );
  AOI22_X1 U23277 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20394), .B1(
        n20424), .B2(n20649), .ZN(n20369) );
  OAI211_X1 U23278 ( .C1(n20397), .C2(n20493), .A(n20370), .B(n20369), .ZN(
        P1_U3081) );
  OAI22_X1 U23279 ( .A1(n20380), .A2(n20656), .B1(n20577), .B2(n20390), .ZN(
        n20371) );
  INV_X1 U23280 ( .A(n20371), .ZN(n20373) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20394), .B1(
        n20424), .B2(n20653), .ZN(n20372) );
  OAI211_X1 U23282 ( .C1(n20397), .C2(n20497), .A(n20373), .B(n20372), .ZN(
        P1_U3082) );
  OAI22_X1 U23283 ( .A1(n20380), .A2(n20660), .B1(n20581), .B2(n20390), .ZN(
        n20374) );
  INV_X1 U23284 ( .A(n20374), .ZN(n20376) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20394), .B1(
        n20424), .B2(n20657), .ZN(n20375) );
  OAI211_X1 U23286 ( .C1(n20397), .C2(n20501), .A(n20376), .B(n20375), .ZN(
        P1_U3083) );
  AOI22_X1 U23287 ( .A1(n20377), .A2(n20718), .B1(n20424), .B2(n20661), .ZN(
        n20379) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20394), .B1(
        n20393), .B2(n20720), .ZN(n20378) );
  OAI211_X1 U23289 ( .C1(n20397), .C2(n20505), .A(n20379), .B(n20378), .ZN(
        P1_U3084) );
  OAI22_X1 U23290 ( .A1(n20380), .A2(n20668), .B1(n20588), .B2(n20390), .ZN(
        n20381) );
  INV_X1 U23291 ( .A(n20381), .ZN(n20383) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20394), .B1(
        n20424), .B2(n20665), .ZN(n20382) );
  OAI211_X1 U23293 ( .C1(n20397), .C2(n20509), .A(n20383), .B(n20382), .ZN(
        P1_U3085) );
  OAI22_X1 U23294 ( .A1(n20391), .A2(n20735), .B1(n20592), .B2(n20390), .ZN(
        n20384) );
  INV_X1 U23295 ( .A(n20384), .ZN(n20386) );
  INV_X1 U23296 ( .A(n20672), .ZN(n20732) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20394), .B1(
        n20393), .B2(n20732), .ZN(n20385) );
  OAI211_X1 U23298 ( .C1(n20397), .C2(n20514), .A(n20386), .B(n20385), .ZN(
        P1_U3086) );
  OAI22_X1 U23299 ( .A1(n20391), .A2(n20741), .B1(n20596), .B2(n20390), .ZN(
        n20387) );
  INV_X1 U23300 ( .A(n20387), .ZN(n20389) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20394), .B1(
        n20393), .B2(n20738), .ZN(n20388) );
  OAI211_X1 U23302 ( .C1(n20397), .C2(n20518), .A(n20389), .B(n20388), .ZN(
        P1_U3087) );
  OAI22_X1 U23303 ( .A1(n20391), .A2(n20752), .B1(n20601), .B2(n20390), .ZN(
        n20392) );
  INV_X1 U23304 ( .A(n20392), .ZN(n20396) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20394), .B1(
        n20393), .B2(n20746), .ZN(n20395) );
  OAI211_X1 U23306 ( .C1(n20397), .C2(n20525), .A(n20396), .B(n20395), .ZN(
        P1_U3088) );
  INV_X1 U23307 ( .A(n20403), .ZN(n20399) );
  INV_X1 U23308 ( .A(n20540), .ZN(n20398) );
  INV_X1 U23309 ( .A(n20686), .ZN(n20531) );
  OAI21_X1 U23310 ( .B1(n20401), .B2(n20531), .A(n20400), .ZN(n20407) );
  INV_X1 U23311 ( .A(n20407), .ZN(n20402) );
  OAI22_X1 U23312 ( .A1(n20402), .A2(n20693), .B1(n20404), .B2(n11268), .ZN(
        n20423) );
  AOI22_X1 U23313 ( .A1(n20422), .A2(n20691), .B1(n20692), .B2(n20423), .ZN(
        n20409) );
  NAND2_X1 U23314 ( .A1(n20403), .A2(n20617), .ZN(n20406) );
  INV_X1 U23315 ( .A(n20699), .ZN(n20534) );
  AOI21_X1 U23316 ( .B1(n20693), .B2(n20404), .A(n20534), .ZN(n20405) );
  OAI221_X1 U23317 ( .B1(n20407), .B2(n20538), .C1(n20407), .C2(n20406), .A(
        n20405), .ZN(n20425) );
  AOI22_X1 U23318 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20702), .ZN(n20408) );
  OAI211_X1 U23319 ( .C1(n20705), .C2(n20456), .A(n20409), .B(n20408), .ZN(
        P1_U3089) );
  AOI22_X1 U23320 ( .A1(n20423), .A2(n20707), .B1(n20422), .B2(n20706), .ZN(
        n20411) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20708), .ZN(n20410) );
  OAI211_X1 U23322 ( .C1(n20711), .C2(n20456), .A(n20411), .B(n20410), .ZN(
        P1_U3090) );
  AOI22_X1 U23323 ( .A1(n20423), .A2(n20713), .B1(n20422), .B2(n20712), .ZN(
        n20413) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20714), .ZN(n20412) );
  OAI211_X1 U23325 ( .C1(n20717), .C2(n20456), .A(n20413), .B(n20412), .ZN(
        P1_U3091) );
  AOI22_X1 U23326 ( .A1(n20422), .A2(n20718), .B1(n20719), .B2(n20423), .ZN(
        n20415) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20720), .ZN(n20414) );
  OAI211_X1 U23328 ( .C1(n20723), .C2(n20456), .A(n20415), .B(n20414), .ZN(
        P1_U3092) );
  AOI22_X1 U23329 ( .A1(n20423), .A2(n20725), .B1(n20422), .B2(n20724), .ZN(
        n20417) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20726), .ZN(n20416) );
  OAI211_X1 U23331 ( .C1(n20729), .C2(n20456), .A(n20417), .B(n20416), .ZN(
        P1_U3093) );
  AOI22_X1 U23332 ( .A1(n20423), .A2(n20731), .B1(n20422), .B2(n20730), .ZN(
        n20419) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20732), .ZN(n20418) );
  OAI211_X1 U23334 ( .C1(n20735), .C2(n20456), .A(n20419), .B(n20418), .ZN(
        P1_U3094) );
  AOI22_X1 U23335 ( .A1(n20423), .A2(n20737), .B1(n20422), .B2(n20736), .ZN(
        n20421) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20738), .ZN(n20420) );
  OAI211_X1 U23337 ( .C1(n20741), .C2(n20456), .A(n20421), .B(n20420), .ZN(
        P1_U3095) );
  AOI22_X1 U23338 ( .A1(n20423), .A2(n20744), .B1(n20422), .B2(n20743), .ZN(
        n20427) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20746), .ZN(n20426) );
  OAI211_X1 U23340 ( .C1(n20752), .C2(n20456), .A(n20427), .B(n20426), .ZN(
        P1_U3096) );
  AND2_X1 U23341 ( .A1(n20428), .A2(n12991), .ZN(n20527) );
  NAND2_X1 U23342 ( .A1(n20429), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20485) );
  AOI21_X1 U23343 ( .B1(n20527), .B2(n14385), .A(n10161), .ZN(n20434) );
  INV_X1 U23344 ( .A(n20482), .ZN(n20430) );
  NAND2_X1 U23345 ( .A1(n20431), .A2(n20430), .ZN(n20572) );
  OAI22_X1 U23346 ( .A1(n20434), .A2(n20693), .B1(n20432), .B2(n20572), .ZN(
        n20451) );
  AOI22_X1 U23347 ( .A1(n20692), .A2(n20451), .B1(n20691), .B2(n10161), .ZN(
        n20438) );
  INV_X1 U23348 ( .A(n20456), .ZN(n20433) );
  OAI21_X1 U23349 ( .B1(n20452), .B2(n20433), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20435) );
  NAND2_X1 U23350 ( .A1(n20435), .A2(n20434), .ZN(n20436) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20453), .B1(
        n20452), .B2(n20649), .ZN(n20437) );
  OAI211_X1 U23352 ( .C1(n20652), .C2(n20456), .A(n20438), .B(n20437), .ZN(
        P1_U3097) );
  AOI22_X1 U23353 ( .A1(n20451), .A2(n20707), .B1(n10161), .B2(n20706), .ZN(
        n20440) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20453), .B1(
        n20452), .B2(n20653), .ZN(n20439) );
  OAI211_X1 U23355 ( .C1(n20656), .C2(n20456), .A(n20440), .B(n20439), .ZN(
        P1_U3098) );
  AOI22_X1 U23356 ( .A1(n20451), .A2(n20713), .B1(n10161), .B2(n20712), .ZN(
        n20442) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20453), .B1(
        n20452), .B2(n20657), .ZN(n20441) );
  OAI211_X1 U23358 ( .C1(n20660), .C2(n20456), .A(n20442), .B(n20441), .ZN(
        P1_U3099) );
  AOI22_X1 U23359 ( .A1(n20719), .A2(n20451), .B1(n20718), .B2(n10161), .ZN(
        n20444) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20453), .B1(
        n20452), .B2(n20661), .ZN(n20443) );
  OAI211_X1 U23361 ( .C1(n20664), .C2(n20456), .A(n20444), .B(n20443), .ZN(
        P1_U3100) );
  AOI22_X1 U23362 ( .A1(n20451), .A2(n20725), .B1(n10161), .B2(n20724), .ZN(
        n20446) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20453), .B1(
        n20452), .B2(n20665), .ZN(n20445) );
  OAI211_X1 U23364 ( .C1(n20668), .C2(n20456), .A(n20446), .B(n20445), .ZN(
        P1_U3101) );
  AOI22_X1 U23365 ( .A1(n20451), .A2(n20731), .B1(n10161), .B2(n20730), .ZN(
        n20448) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20453), .B1(
        n20452), .B2(n20669), .ZN(n20447) );
  OAI211_X1 U23367 ( .C1(n20672), .C2(n20456), .A(n20448), .B(n20447), .ZN(
        P1_U3102) );
  AOI22_X1 U23368 ( .A1(n20451), .A2(n20737), .B1(n10161), .B2(n20736), .ZN(
        n20450) );
  AOI22_X1 U23369 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20453), .B1(
        n20452), .B2(n20673), .ZN(n20449) );
  OAI211_X1 U23370 ( .C1(n20676), .C2(n20456), .A(n20450), .B(n20449), .ZN(
        P1_U3103) );
  AOI22_X1 U23371 ( .A1(n20451), .A2(n20744), .B1(n10161), .B2(n20743), .ZN(
        n20455) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20453), .B1(
        n20452), .B2(n20679), .ZN(n20454) );
  OAI211_X1 U23373 ( .C1(n20684), .C2(n20456), .A(n20455), .B(n20454), .ZN(
        P1_U3104) );
  NOR2_X1 U23374 ( .A1(n20485), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20460) );
  INV_X1 U23375 ( .A(n20460), .ZN(n20457) );
  NOR2_X1 U23376 ( .A1(n20611), .A2(n20457), .ZN(n20475) );
  AOI21_X1 U23377 ( .B1(n20527), .B2(n20612), .A(n20475), .ZN(n20458) );
  OAI22_X1 U23378 ( .A1(n20458), .A2(n20693), .B1(n20457), .B2(n11268), .ZN(
        n20476) );
  AOI22_X1 U23379 ( .A1(n20692), .A2(n20476), .B1(n20691), .B2(n20475), .ZN(
        n20462) );
  OAI211_X1 U23380 ( .C1(n20541), .C2(n14399), .A(n20701), .B(n20458), .ZN(
        n20459) );
  OAI211_X1 U23381 ( .C1(n20701), .C2(n20460), .A(n20699), .B(n20459), .ZN(
        n20477) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20477), .B1(
        n20511), .B2(n20649), .ZN(n20461) );
  OAI211_X1 U23383 ( .C1(n20652), .C2(n20480), .A(n20462), .B(n20461), .ZN(
        P1_U3105) );
  AOI22_X1 U23384 ( .A1(n20476), .A2(n20707), .B1(n20706), .B2(n20475), .ZN(
        n20464) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20477), .B1(
        n20511), .B2(n20653), .ZN(n20463) );
  OAI211_X1 U23386 ( .C1(n20656), .C2(n20480), .A(n20464), .B(n20463), .ZN(
        P1_U3106) );
  AOI22_X1 U23387 ( .A1(n20476), .A2(n20713), .B1(n20712), .B2(n20475), .ZN(
        n20466) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20477), .B1(
        n20511), .B2(n20657), .ZN(n20465) );
  OAI211_X1 U23389 ( .C1(n20660), .C2(n20480), .A(n20466), .B(n20465), .ZN(
        P1_U3107) );
  AOI22_X1 U23390 ( .A1(n20719), .A2(n20476), .B1(n20718), .B2(n20475), .ZN(
        n20468) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20477), .B1(
        n20511), .B2(n20661), .ZN(n20467) );
  OAI211_X1 U23392 ( .C1(n20664), .C2(n20480), .A(n20468), .B(n20467), .ZN(
        P1_U3108) );
  AOI22_X1 U23393 ( .A1(n20476), .A2(n20725), .B1(n20724), .B2(n20475), .ZN(
        n20470) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20477), .B1(
        n20511), .B2(n20665), .ZN(n20469) );
  OAI211_X1 U23395 ( .C1(n20668), .C2(n20480), .A(n20470), .B(n20469), .ZN(
        P1_U3109) );
  AOI22_X1 U23396 ( .A1(n20476), .A2(n20731), .B1(n20730), .B2(n20475), .ZN(
        n20472) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20477), .B1(
        n20511), .B2(n20669), .ZN(n20471) );
  OAI211_X1 U23398 ( .C1(n20672), .C2(n20480), .A(n20472), .B(n20471), .ZN(
        P1_U3110) );
  AOI22_X1 U23399 ( .A1(n20476), .A2(n20737), .B1(n20736), .B2(n20475), .ZN(
        n20474) );
  AOI22_X1 U23400 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20477), .B1(
        n20511), .B2(n20673), .ZN(n20473) );
  OAI211_X1 U23401 ( .C1(n20676), .C2(n20480), .A(n20474), .B(n20473), .ZN(
        P1_U3111) );
  AOI22_X1 U23402 ( .A1(n20476), .A2(n20744), .B1(n20743), .B2(n20475), .ZN(
        n20479) );
  AOI22_X1 U23403 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20477), .B1(
        n20511), .B2(n20679), .ZN(n20478) );
  OAI211_X1 U23404 ( .C1(n20684), .C2(n20480), .A(n20479), .B(n20478), .ZN(
        P1_U3112) );
  NAND3_X1 U23405 ( .A1(n20563), .A2(n20520), .A3(n20617), .ZN(n20481) );
  NAND2_X1 U23406 ( .A1(n20481), .A2(n20566), .ZN(n20488) );
  AND2_X1 U23407 ( .A1(n20527), .A2(n20638), .ZN(n20486) );
  NAND2_X1 U23408 ( .A1(n20482), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20640) );
  INV_X1 U23409 ( .A(n20640), .ZN(n20484) );
  INV_X1 U23410 ( .A(n20485), .ZN(n20528) );
  NAND2_X1 U23411 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20528), .ZN(
        n20535) );
  NOR2_X1 U23412 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20535), .ZN(
        n20502) );
  AOI22_X1 U23413 ( .A1(n20502), .A2(n20691), .B1(n20511), .B2(n20702), .ZN(
        n20492) );
  INV_X1 U23414 ( .A(n20486), .ZN(n20487) );
  INV_X1 U23415 ( .A(n20502), .ZN(n20519) );
  AOI22_X1 U23416 ( .A1(n20488), .A2(n20487), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20519), .ZN(n20489) );
  NAND2_X1 U23417 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20640), .ZN(n20646) );
  NAND3_X1 U23418 ( .A1(n20490), .A2(n20489), .A3(n20646), .ZN(n20522) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20522), .B1(
        n20546), .B2(n20649), .ZN(n20491) );
  OAI211_X1 U23420 ( .C1(n20526), .C2(n20493), .A(n20492), .B(n20491), .ZN(
        P1_U3113) );
  OAI22_X1 U23421 ( .A1(n20520), .A2(n20656), .B1(n20577), .B2(n20519), .ZN(
        n20494) );
  INV_X1 U23422 ( .A(n20494), .ZN(n20496) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20522), .B1(
        n20546), .B2(n20653), .ZN(n20495) );
  OAI211_X1 U23424 ( .C1(n20526), .C2(n20497), .A(n20496), .B(n20495), .ZN(
        P1_U3114) );
  OAI22_X1 U23425 ( .A1(n20563), .A2(n20717), .B1(n20519), .B2(n20581), .ZN(
        n20498) );
  INV_X1 U23426 ( .A(n20498), .ZN(n20500) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20522), .B1(
        n20511), .B2(n20714), .ZN(n20499) );
  OAI211_X1 U23428 ( .C1(n20526), .C2(n20501), .A(n20500), .B(n20499), .ZN(
        P1_U3115) );
  AOI22_X1 U23429 ( .A1(n20502), .A2(n20718), .B1(n20511), .B2(n20720), .ZN(
        n20504) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20522), .B1(
        n20546), .B2(n20661), .ZN(n20503) );
  OAI211_X1 U23431 ( .C1(n20526), .C2(n20505), .A(n20504), .B(n20503), .ZN(
        P1_U3116) );
  OAI22_X1 U23432 ( .A1(n20563), .A2(n20729), .B1(n20519), .B2(n20588), .ZN(
        n20506) );
  INV_X1 U23433 ( .A(n20506), .ZN(n20508) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20522), .B1(
        n20511), .B2(n20726), .ZN(n20507) );
  OAI211_X1 U23435 ( .C1(n20526), .C2(n20509), .A(n20508), .B(n20507), .ZN(
        P1_U3117) );
  OAI22_X1 U23436 ( .A1(n20563), .A2(n20735), .B1(n20519), .B2(n20592), .ZN(
        n20510) );
  INV_X1 U23437 ( .A(n20510), .ZN(n20513) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20522), .B1(
        n20511), .B2(n20732), .ZN(n20512) );
  OAI211_X1 U23439 ( .C1(n20526), .C2(n20514), .A(n20513), .B(n20512), .ZN(
        P1_U3118) );
  OAI22_X1 U23440 ( .A1(n20520), .A2(n20676), .B1(n20519), .B2(n20596), .ZN(
        n20515) );
  INV_X1 U23441 ( .A(n20515), .ZN(n20517) );
  AOI22_X1 U23442 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20522), .B1(
        n20546), .B2(n20673), .ZN(n20516) );
  OAI211_X1 U23443 ( .C1(n20526), .C2(n20518), .A(n20517), .B(n20516), .ZN(
        P1_U3119) );
  OAI22_X1 U23444 ( .A1(n20520), .A2(n20684), .B1(n20519), .B2(n20601), .ZN(
        n20521) );
  INV_X1 U23445 ( .A(n20521), .ZN(n20524) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20522), .B1(
        n20546), .B2(n20679), .ZN(n20523) );
  OAI211_X1 U23447 ( .C1(n20526), .C2(n20525), .A(n20524), .B(n20523), .ZN(
        P1_U3120) );
  INV_X1 U23448 ( .A(n20527), .ZN(n20532) );
  AND2_X1 U23449 ( .A1(n20529), .A2(n20528), .ZN(n20557) );
  INV_X1 U23450 ( .A(n20557), .ZN(n20530) );
  OAI21_X1 U23451 ( .B1(n20532), .B2(n20531), .A(n20530), .ZN(n20539) );
  INV_X1 U23452 ( .A(n20539), .ZN(n20533) );
  OAI22_X1 U23453 ( .A1(n20533), .A2(n20693), .B1(n20535), .B2(n11268), .ZN(
        n20558) );
  AOI22_X1 U23454 ( .A1(n20692), .A2(n20558), .B1(n20691), .B2(n20557), .ZN(
        n20543) );
  NAND2_X1 U23455 ( .A1(n20541), .A2(n20701), .ZN(n20537) );
  AOI21_X1 U23456 ( .B1(n20693), .B2(n20535), .A(n20534), .ZN(n20536) );
  OAI221_X1 U23457 ( .B1(n20539), .B2(n20538), .C1(n20539), .C2(n20537), .A(
        n20536), .ZN(n20560) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20649), .ZN(n20542) );
  OAI211_X1 U23459 ( .C1(n20652), .C2(n20563), .A(n20543), .B(n20542), .ZN(
        P1_U3121) );
  AOI22_X1 U23460 ( .A1(n20558), .A2(n20707), .B1(n20706), .B2(n20557), .ZN(
        n20545) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20653), .ZN(n20544) );
  OAI211_X1 U23462 ( .C1(n20656), .C2(n20563), .A(n20545), .B(n20544), .ZN(
        P1_U3122) );
  AOI22_X1 U23463 ( .A1(n20558), .A2(n20713), .B1(n20712), .B2(n20557), .ZN(
        n20548) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20560), .B1(
        n20546), .B2(n20714), .ZN(n20547) );
  OAI211_X1 U23465 ( .C1(n20717), .C2(n20608), .A(n20548), .B(n20547), .ZN(
        P1_U3123) );
  AOI22_X1 U23466 ( .A1(n20719), .A2(n20558), .B1(n20718), .B2(n20557), .ZN(
        n20550) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20661), .ZN(n20549) );
  OAI211_X1 U23468 ( .C1(n20664), .C2(n20563), .A(n20550), .B(n20549), .ZN(
        P1_U3124) );
  AOI22_X1 U23469 ( .A1(n20558), .A2(n20725), .B1(n20724), .B2(n20557), .ZN(
        n20552) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20665), .ZN(n20551) );
  OAI211_X1 U23471 ( .C1(n20668), .C2(n20563), .A(n20552), .B(n20551), .ZN(
        P1_U3125) );
  AOI22_X1 U23472 ( .A1(n20558), .A2(n20731), .B1(n20730), .B2(n20557), .ZN(
        n20554) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20669), .ZN(n20553) );
  OAI211_X1 U23474 ( .C1(n20672), .C2(n20563), .A(n20554), .B(n20553), .ZN(
        P1_U3126) );
  AOI22_X1 U23475 ( .A1(n20558), .A2(n20737), .B1(n20736), .B2(n20557), .ZN(
        n20556) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20673), .ZN(n20555) );
  OAI211_X1 U23477 ( .C1(n20676), .C2(n20563), .A(n20556), .B(n20555), .ZN(
        P1_U3127) );
  AOI22_X1 U23478 ( .A1(n20558), .A2(n20744), .B1(n20743), .B2(n20557), .ZN(
        n20562) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20560), .B1(
        n20559), .B2(n20679), .ZN(n20561) );
  OAI211_X1 U23480 ( .C1(n20684), .C2(n20563), .A(n20562), .B(n20561), .ZN(
        P1_U3128) );
  NAND2_X1 U23481 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20688) );
  OR2_X1 U23482 ( .A1(n20564), .A2(n20688), .ZN(n20600) );
  INV_X1 U23483 ( .A(n20600), .ZN(n20585) );
  AOI22_X1 U23484 ( .A1(n20585), .A2(n20691), .B1(n20634), .B2(n20649), .ZN(
        n20576) );
  NAND3_X1 U23485 ( .A1(n20608), .A2(n20617), .A3(n20602), .ZN(n20567) );
  NAND2_X1 U23486 ( .A1(n20567), .A2(n20566), .ZN(n20571) );
  NOR2_X1 U23487 ( .A1(n12991), .A2(n20568), .ZN(n20687) );
  NAND2_X1 U23488 ( .A1(n20687), .A2(n14385), .ZN(n20573) );
  AOI22_X1 U23489 ( .A1(n20571), .A2(n20573), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20572), .ZN(n20569) );
  OAI211_X1 U23490 ( .C1(n20585), .C2(n20570), .A(n20647), .B(n20569), .ZN(
        n20605) );
  INV_X1 U23491 ( .A(n20571), .ZN(n20574) );
  OAI22_X1 U23492 ( .A1(n20574), .A2(n20573), .B1(n20572), .B2(n20639), .ZN(
        n20604) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20605), .B1(
        n20692), .B2(n20604), .ZN(n20575) );
  OAI211_X1 U23494 ( .C1(n20652), .C2(n20608), .A(n20576), .B(n20575), .ZN(
        P1_U3129) );
  OAI22_X1 U23495 ( .A1(n20602), .A2(n20711), .B1(n20577), .B2(n20600), .ZN(
        n20578) );
  INV_X1 U23496 ( .A(n20578), .ZN(n20580) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20605), .B1(
        n20707), .B2(n20604), .ZN(n20579) );
  OAI211_X1 U23498 ( .C1(n20656), .C2(n20608), .A(n20580), .B(n20579), .ZN(
        P1_U3130) );
  OAI22_X1 U23499 ( .A1(n20602), .A2(n20717), .B1(n20581), .B2(n20600), .ZN(
        n20582) );
  INV_X1 U23500 ( .A(n20582), .ZN(n20584) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20605), .B1(
        n20713), .B2(n20604), .ZN(n20583) );
  OAI211_X1 U23502 ( .C1(n20660), .C2(n20608), .A(n20584), .B(n20583), .ZN(
        P1_U3131) );
  AOI22_X1 U23503 ( .A1(n20585), .A2(n20718), .B1(n20634), .B2(n20661), .ZN(
        n20587) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20605), .B1(
        n20719), .B2(n20604), .ZN(n20586) );
  OAI211_X1 U23505 ( .C1(n20664), .C2(n20608), .A(n20587), .B(n20586), .ZN(
        P1_U3132) );
  OAI22_X1 U23506 ( .A1(n20602), .A2(n20729), .B1(n20588), .B2(n20600), .ZN(
        n20589) );
  INV_X1 U23507 ( .A(n20589), .ZN(n20591) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20605), .B1(
        n20725), .B2(n20604), .ZN(n20590) );
  OAI211_X1 U23509 ( .C1(n20668), .C2(n20608), .A(n20591), .B(n20590), .ZN(
        P1_U3133) );
  OAI22_X1 U23510 ( .A1(n20602), .A2(n20735), .B1(n20592), .B2(n20600), .ZN(
        n20593) );
  INV_X1 U23511 ( .A(n20593), .ZN(n20595) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20605), .B1(
        n20731), .B2(n20604), .ZN(n20594) );
  OAI211_X1 U23513 ( .C1(n20672), .C2(n20608), .A(n20595), .B(n20594), .ZN(
        P1_U3134) );
  OAI22_X1 U23514 ( .A1(n20602), .A2(n20741), .B1(n20596), .B2(n20600), .ZN(
        n20597) );
  INV_X1 U23515 ( .A(n20597), .ZN(n20599) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20605), .B1(
        n20737), .B2(n20604), .ZN(n20598) );
  OAI211_X1 U23517 ( .C1(n20676), .C2(n20608), .A(n20599), .B(n20598), .ZN(
        P1_U3135) );
  OAI22_X1 U23518 ( .A1(n20602), .A2(n20752), .B1(n20601), .B2(n20600), .ZN(
        n20603) );
  INV_X1 U23519 ( .A(n20603), .ZN(n20607) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20605), .B1(
        n20744), .B2(n20604), .ZN(n20606) );
  OAI211_X1 U23521 ( .C1(n20684), .C2(n20608), .A(n20607), .B(n20606), .ZN(
        P1_U3136) );
  INV_X1 U23522 ( .A(n20642), .ZN(n20694) );
  INV_X1 U23523 ( .A(n20609), .ZN(n20610) );
  NOR3_X2 U23524 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20611), .A3(
        n20688), .ZN(n20632) );
  AOI21_X1 U23525 ( .B1(n20687), .B2(n20612), .A(n20632), .ZN(n20614) );
  NOR2_X1 U23526 ( .A1(n20688), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20616) );
  INV_X1 U23527 ( .A(n20616), .ZN(n20613) );
  OAI22_X1 U23528 ( .A1(n20614), .A2(n20693), .B1(n20613), .B2(n11268), .ZN(
        n20633) );
  AOI22_X1 U23529 ( .A1(n20692), .A2(n20633), .B1(n20691), .B2(n20632), .ZN(
        n20619) );
  OAI211_X1 U23530 ( .C1(n20642), .C2(n14399), .A(n20617), .B(n20614), .ZN(
        n20615) );
  OAI211_X1 U23531 ( .C1(n20617), .C2(n20616), .A(n20699), .B(n20615), .ZN(
        n20635) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20702), .ZN(n20618) );
  OAI211_X1 U23533 ( .C1(n20705), .C2(n20683), .A(n20619), .B(n20618), .ZN(
        P1_U3137) );
  AOI22_X1 U23534 ( .A1(n20633), .A2(n20707), .B1(n20706), .B2(n20632), .ZN(
        n20621) );
  AOI22_X1 U23535 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20708), .ZN(n20620) );
  OAI211_X1 U23536 ( .C1(n20711), .C2(n20683), .A(n20621), .B(n20620), .ZN(
        P1_U3138) );
  AOI22_X1 U23537 ( .A1(n20633), .A2(n20713), .B1(n20712), .B2(n20632), .ZN(
        n20623) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20714), .ZN(n20622) );
  OAI211_X1 U23539 ( .C1(n20717), .C2(n20683), .A(n20623), .B(n20622), .ZN(
        P1_U3139) );
  AOI22_X1 U23540 ( .A1(n20719), .A2(n20633), .B1(n20718), .B2(n20632), .ZN(
        n20625) );
  AOI22_X1 U23541 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20720), .ZN(n20624) );
  OAI211_X1 U23542 ( .C1(n20723), .C2(n20683), .A(n20625), .B(n20624), .ZN(
        P1_U3140) );
  AOI22_X1 U23543 ( .A1(n20633), .A2(n20725), .B1(n20724), .B2(n20632), .ZN(
        n20627) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20726), .ZN(n20626) );
  OAI211_X1 U23545 ( .C1(n20729), .C2(n20683), .A(n20627), .B(n20626), .ZN(
        P1_U3141) );
  AOI22_X1 U23546 ( .A1(n20633), .A2(n20731), .B1(n20730), .B2(n20632), .ZN(
        n20629) );
  AOI22_X1 U23547 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20732), .ZN(n20628) );
  OAI211_X1 U23548 ( .C1(n20735), .C2(n20683), .A(n20629), .B(n20628), .ZN(
        P1_U3142) );
  AOI22_X1 U23549 ( .A1(n20633), .A2(n20737), .B1(n20736), .B2(n20632), .ZN(
        n20631) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20738), .ZN(n20630) );
  OAI211_X1 U23551 ( .C1(n20741), .C2(n20683), .A(n20631), .B(n20630), .ZN(
        P1_U3143) );
  AOI22_X1 U23552 ( .A1(n20633), .A2(n20744), .B1(n20743), .B2(n20632), .ZN(
        n20637) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20746), .ZN(n20636) );
  OAI211_X1 U23554 ( .C1(n20752), .C2(n20683), .A(n20637), .B(n20636), .ZN(
        P1_U3144) );
  NAND2_X1 U23555 ( .A1(n20687), .A2(n20638), .ZN(n20644) );
  OAI22_X1 U23556 ( .A1(n20644), .A2(n20693), .B1(n20640), .B2(n20639), .ZN(
        n20678) );
  NOR3_X2 U23557 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20689), .A3(
        n20688), .ZN(n20677) );
  AOI22_X1 U23558 ( .A1(n20692), .A2(n20678), .B1(n20691), .B2(n20677), .ZN(
        n20651) );
  INV_X1 U23559 ( .A(n20683), .ZN(n20643) );
  NOR2_X2 U23560 ( .A1(n20642), .A2(n20641), .ZN(n20747) );
  OAI21_X1 U23561 ( .B1(n20643), .B2(n20747), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20645) );
  AOI21_X1 U23562 ( .B1(n20645), .B2(n20644), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20648) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20680), .B1(
        n20747), .B2(n20649), .ZN(n20650) );
  OAI211_X1 U23564 ( .C1(n20652), .C2(n20683), .A(n20651), .B(n20650), .ZN(
        P1_U3145) );
  AOI22_X1 U23565 ( .A1(n20678), .A2(n20707), .B1(n20706), .B2(n20677), .ZN(
        n20655) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20680), .B1(
        n20747), .B2(n20653), .ZN(n20654) );
  OAI211_X1 U23567 ( .C1(n20656), .C2(n20683), .A(n20655), .B(n20654), .ZN(
        P1_U3146) );
  AOI22_X1 U23568 ( .A1(n20678), .A2(n20713), .B1(n20712), .B2(n20677), .ZN(
        n20659) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20680), .B1(
        n20747), .B2(n20657), .ZN(n20658) );
  OAI211_X1 U23570 ( .C1(n20660), .C2(n20683), .A(n20659), .B(n20658), .ZN(
        P1_U3147) );
  AOI22_X1 U23571 ( .A1(n20719), .A2(n20678), .B1(n20718), .B2(n20677), .ZN(
        n20663) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20680), .B1(
        n20747), .B2(n20661), .ZN(n20662) );
  OAI211_X1 U23573 ( .C1(n20664), .C2(n20683), .A(n20663), .B(n20662), .ZN(
        P1_U3148) );
  AOI22_X1 U23574 ( .A1(n20678), .A2(n20725), .B1(n20724), .B2(n20677), .ZN(
        n20667) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20680), .B1(
        n20747), .B2(n20665), .ZN(n20666) );
  OAI211_X1 U23576 ( .C1(n20668), .C2(n20683), .A(n20667), .B(n20666), .ZN(
        P1_U3149) );
  AOI22_X1 U23577 ( .A1(n20678), .A2(n20731), .B1(n20730), .B2(n20677), .ZN(
        n20671) );
  AOI22_X1 U23578 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20680), .B1(
        n20747), .B2(n20669), .ZN(n20670) );
  OAI211_X1 U23579 ( .C1(n20672), .C2(n20683), .A(n20671), .B(n20670), .ZN(
        P1_U3150) );
  AOI22_X1 U23580 ( .A1(n20678), .A2(n20737), .B1(n20736), .B2(n20677), .ZN(
        n20675) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20680), .B1(
        n20747), .B2(n20673), .ZN(n20674) );
  OAI211_X1 U23582 ( .C1(n20676), .C2(n20683), .A(n20675), .B(n20674), .ZN(
        P1_U3151) );
  AOI22_X1 U23583 ( .A1(n20678), .A2(n20744), .B1(n20743), .B2(n20677), .ZN(
        n20682) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20680), .B1(
        n20747), .B2(n20679), .ZN(n20681) );
  OAI211_X1 U23585 ( .C1(n20684), .C2(n20683), .A(n20682), .B(n20681), .ZN(
        P1_U3152) );
  NOR2_X1 U23586 ( .A1(n20685), .A2(n20688), .ZN(n20742) );
  AOI21_X1 U23587 ( .B1(n20687), .B2(n20686), .A(n20742), .ZN(n20695) );
  NOR2_X1 U23588 ( .A1(n20689), .A2(n20688), .ZN(n20700) );
  INV_X1 U23589 ( .A(n20700), .ZN(n20690) );
  OAI22_X1 U23590 ( .A1(n20695), .A2(n20693), .B1(n20690), .B2(n11268), .ZN(
        n20745) );
  AOI22_X1 U23591 ( .A1(n20692), .A2(n20745), .B1(n20691), .B2(n20742), .ZN(
        n20704) );
  NOR2_X1 U23592 ( .A1(n20694), .A2(n20693), .ZN(n20697) );
  OAI21_X1 U23593 ( .B1(n20697), .B2(n20696), .A(n20695), .ZN(n20698) );
  OAI211_X1 U23594 ( .C1(n20701), .C2(n20700), .A(n20699), .B(n20698), .ZN(
        n20748) );
  AOI22_X1 U23595 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20702), .ZN(n20703) );
  OAI211_X1 U23596 ( .C1(n20705), .C2(n20751), .A(n20704), .B(n20703), .ZN(
        P1_U3153) );
  AOI22_X1 U23597 ( .A1(n20745), .A2(n20707), .B1(n20706), .B2(n20742), .ZN(
        n20710) );
  AOI22_X1 U23598 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20708), .ZN(n20709) );
  OAI211_X1 U23599 ( .C1(n20711), .C2(n20751), .A(n20710), .B(n20709), .ZN(
        P1_U3154) );
  AOI22_X1 U23600 ( .A1(n20745), .A2(n20713), .B1(n20712), .B2(n20742), .ZN(
        n20716) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20714), .ZN(n20715) );
  OAI211_X1 U23602 ( .C1(n20717), .C2(n20751), .A(n20716), .B(n20715), .ZN(
        P1_U3155) );
  AOI22_X1 U23603 ( .A1(n20719), .A2(n20745), .B1(n20718), .B2(n20742), .ZN(
        n20722) );
  AOI22_X1 U23604 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20720), .ZN(n20721) );
  OAI211_X1 U23605 ( .C1(n20723), .C2(n20751), .A(n20722), .B(n20721), .ZN(
        P1_U3156) );
  AOI22_X1 U23606 ( .A1(n20745), .A2(n20725), .B1(n20724), .B2(n20742), .ZN(
        n20728) );
  AOI22_X1 U23607 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20726), .ZN(n20727) );
  OAI211_X1 U23608 ( .C1(n20729), .C2(n20751), .A(n20728), .B(n20727), .ZN(
        P1_U3157) );
  AOI22_X1 U23609 ( .A1(n20745), .A2(n20731), .B1(n20730), .B2(n20742), .ZN(
        n20734) );
  AOI22_X1 U23610 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20732), .ZN(n20733) );
  OAI211_X1 U23611 ( .C1(n20735), .C2(n20751), .A(n20734), .B(n20733), .ZN(
        P1_U3158) );
  AOI22_X1 U23612 ( .A1(n20745), .A2(n20737), .B1(n20736), .B2(n20742), .ZN(
        n20740) );
  AOI22_X1 U23613 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20738), .ZN(n20739) );
  OAI211_X1 U23614 ( .C1(n20741), .C2(n20751), .A(n20740), .B(n20739), .ZN(
        P1_U3159) );
  AOI22_X1 U23615 ( .A1(n20745), .A2(n20744), .B1(n20743), .B2(n20742), .ZN(
        n20750) );
  AOI22_X1 U23616 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20748), .B1(
        n20747), .B2(n20746), .ZN(n20749) );
  OAI211_X1 U23617 ( .C1(n20752), .C2(n20751), .A(n20750), .B(n20749), .ZN(
        P1_U3160) );
  NOR2_X1 U23618 ( .A1(n20754), .A2(n20753), .ZN(n20757) );
  INV_X1 U23619 ( .A(n20755), .ZN(n20756) );
  OAI21_X1 U23620 ( .B1(n20757), .B2(n11268), .A(n20756), .ZN(P1_U3163) );
  NOR2_X1 U23621 ( .A1(n20830), .A2(n20758), .ZN(P1_U3164) );
  AND2_X1 U23622 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20759), .ZN(
        P1_U3165) );
  AND2_X1 U23623 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20759), .ZN(
        P1_U3166) );
  AND2_X1 U23624 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20759), .ZN(
        P1_U3167) );
  AND2_X1 U23625 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20759), .ZN(
        P1_U3168) );
  AND2_X1 U23626 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20759), .ZN(
        P1_U3169) );
  AND2_X1 U23627 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20759), .ZN(
        P1_U3170) );
  AND2_X1 U23628 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20759), .ZN(
        P1_U3171) );
  AND2_X1 U23629 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20759), .ZN(
        P1_U3172) );
  AND2_X1 U23630 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20759), .ZN(
        P1_U3173) );
  AND2_X1 U23631 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20759), .ZN(
        P1_U3174) );
  AND2_X1 U23632 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20759), .ZN(
        P1_U3175) );
  AND2_X1 U23633 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20759), .ZN(
        P1_U3176) );
  AND2_X1 U23634 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20759), .ZN(
        P1_U3177) );
  AND2_X1 U23635 ( .A1(n20759), .A2(P1_DATAWIDTH_REG_17__SCAN_IN), .ZN(
        P1_U3178) );
  AND2_X1 U23636 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20759), .ZN(
        P1_U3179) );
  AND2_X1 U23637 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20759), .ZN(
        P1_U3180) );
  AND2_X1 U23638 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20759), .ZN(
        P1_U3181) );
  AND2_X1 U23639 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20759), .ZN(
        P1_U3182) );
  AND2_X1 U23640 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20759), .ZN(
        P1_U3183) );
  AND2_X1 U23641 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20759), .ZN(
        P1_U3184) );
  AND2_X1 U23642 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20759), .ZN(
        P1_U3185) );
  AND2_X1 U23643 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20759), .ZN(P1_U3186) );
  AND2_X1 U23644 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20759), .ZN(P1_U3187) );
  AND2_X1 U23645 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20759), .ZN(P1_U3188) );
  AND2_X1 U23646 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20759), .ZN(P1_U3189) );
  AND2_X1 U23647 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20759), .ZN(P1_U3190) );
  AND2_X1 U23648 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20759), .ZN(P1_U3191) );
  AND2_X1 U23649 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20759), .ZN(P1_U3192) );
  AND2_X1 U23650 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20759), .ZN(P1_U3193) );
  AND2_X1 U23651 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20760), .ZN(n20774) );
  INV_X1 U23652 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20856) );
  NOR2_X1 U23653 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20762) );
  OAI22_X1 U23654 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20767), .B1(n20762), 
        .B2(n20761), .ZN(n20763) );
  NOR2_X1 U23655 ( .A1(n20856), .A2(n20763), .ZN(n20764) );
  OAI22_X1 U23656 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20774), .B1(n20861), 
        .B2(n20764), .ZN(P1_U3194) );
  INV_X1 U23657 ( .A(n20765), .ZN(n20768) );
  NOR2_X1 U23658 ( .A1(n20772), .A2(n20856), .ZN(n20766) );
  OAI22_X1 U23659 ( .A1(n20768), .A2(n20767), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20766), .ZN(n20773) );
  OAI211_X1 U23660 ( .C1(NA), .C2(n20769), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20775), .ZN(n20770) );
  OAI211_X1 U23661 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20856), .A(HOLD), .B(
        n20770), .ZN(n20771) );
  OAI22_X1 U23662 ( .A1(n20774), .A2(n20773), .B1(n20772), .B2(n20771), .ZN(
        P1_U3196) );
  OR2_X1 U23663 ( .A1(n20858), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20818) );
  AOI222_X1 U23664 ( .A1(n20819), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n9595), .ZN(n20776) );
  INV_X1 U23665 ( .A(n20776), .ZN(P1_U3197) );
  INV_X1 U23666 ( .A(n9595), .ZN(n20814) );
  AOI22_X1 U23667 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n20819), .ZN(n20777) );
  OAI21_X1 U23668 ( .B1(n20778), .B2(n20814), .A(n20777), .ZN(P1_U3198) );
  AOI222_X1 U23669 ( .A1(n9595), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20819), .ZN(n20779) );
  INV_X1 U23670 ( .A(n20779), .ZN(P1_U3199) );
  AOI22_X1 U23671 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20819), .ZN(n20780) );
  OAI21_X1 U23672 ( .B1(n20781), .B2(n20814), .A(n20780), .ZN(P1_U3200) );
  AOI22_X1 U23673 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n9595), .ZN(n20782) );
  OAI21_X1 U23674 ( .B1(n20784), .B2(n20818), .A(n20782), .ZN(P1_U3201) );
  AOI22_X1 U23675 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20819), .ZN(n20783) );
  OAI21_X1 U23676 ( .B1(n20784), .B2(n20814), .A(n20783), .ZN(P1_U3202) );
  AOI22_X1 U23677 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n9595), .ZN(n20785) );
  OAI21_X1 U23678 ( .B1(n20787), .B2(n20818), .A(n20785), .ZN(P1_U3203) );
  AOI22_X1 U23679 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20819), .ZN(n20786) );
  OAI21_X1 U23680 ( .B1(n20787), .B2(n20814), .A(n20786), .ZN(P1_U3204) );
  AOI222_X1 U23681 ( .A1(n9595), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20819), .ZN(n20788) );
  INV_X1 U23682 ( .A(n20788), .ZN(P1_U3205) );
  AOI222_X1 U23683 ( .A1(n20819), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n9595), .ZN(n20789) );
  INV_X1 U23684 ( .A(n20789), .ZN(P1_U3206) );
  AOI222_X1 U23685 ( .A1(n9595), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20819), .ZN(n20790) );
  INV_X1 U23686 ( .A(n20790), .ZN(P1_U3207) );
  AOI22_X1 U23687 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n20819), .ZN(n20791) );
  OAI21_X1 U23688 ( .B1(n20792), .B2(n20814), .A(n20791), .ZN(P1_U3208) );
  AOI22_X1 U23689 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n9595), .ZN(n20793) );
  OAI21_X1 U23690 ( .B1(n20794), .B2(n20818), .A(n20793), .ZN(P1_U3209) );
  AOI222_X1 U23691 ( .A1(n20819), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n9595), .ZN(n20795) );
  INV_X1 U23692 ( .A(n20795), .ZN(P1_U3210) );
  AOI222_X1 U23693 ( .A1(n9595), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20819), .ZN(n20796) );
  INV_X1 U23694 ( .A(n20796), .ZN(P1_U3211) );
  AOI222_X1 U23695 ( .A1(n9595), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20819), .ZN(n20797) );
  INV_X1 U23696 ( .A(n20797), .ZN(P1_U3212) );
  AOI22_X1 U23697 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20819), .ZN(n20798) );
  OAI21_X1 U23698 ( .B1(n20799), .B2(n20814), .A(n20798), .ZN(P1_U3213) );
  AOI22_X1 U23699 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n9595), .ZN(n20800) );
  OAI21_X1 U23700 ( .B1(n20802), .B2(n20818), .A(n20800), .ZN(P1_U3214) );
  AOI22_X1 U23701 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20819), .ZN(n20801) );
  OAI21_X1 U23702 ( .B1(n20802), .B2(n20814), .A(n20801), .ZN(P1_U3215) );
  AOI22_X1 U23703 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n9595), .ZN(n20803) );
  OAI21_X1 U23704 ( .B1(n20804), .B2(n20818), .A(n20803), .ZN(P1_U3216) );
  AOI222_X1 U23705 ( .A1(n9595), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20819), .ZN(n20805) );
  INV_X1 U23706 ( .A(n20805), .ZN(P1_U3217) );
  AOI222_X1 U23707 ( .A1(n9595), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20819), .ZN(n20806) );
  INV_X1 U23708 ( .A(n20806), .ZN(P1_U3218) );
  AOI22_X1 U23709 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(n20819), .ZN(n20807) );
  OAI21_X1 U23710 ( .B1(n14192), .B2(n20814), .A(n20807), .ZN(P1_U3219) );
  AOI22_X1 U23711 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(n20858), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(n9595), .ZN(n20808) );
  OAI21_X1 U23712 ( .B1(n20809), .B2(n20818), .A(n20808), .ZN(P1_U3220) );
  AOI222_X1 U23713 ( .A1(n9595), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20819), .ZN(n20810) );
  INV_X1 U23714 ( .A(n20810), .ZN(P1_U3221) );
  AOI222_X1 U23715 ( .A1(n9595), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20819), .ZN(n20811) );
  INV_X1 U23716 ( .A(n20811), .ZN(P1_U3222) );
  AOI222_X1 U23717 ( .A1(n9595), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20819), .ZN(n20812) );
  INV_X1 U23718 ( .A(n20812), .ZN(P1_U3223) );
  AOI222_X1 U23719 ( .A1(n9595), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20819), .ZN(n20813) );
  INV_X1 U23720 ( .A(n20813), .ZN(P1_U3224) );
  OAI222_X1 U23721 ( .A1(n20818), .A2(n20817), .B1(n20816), .B2(n20861), .C1(
        n20815), .C2(n20814), .ZN(P1_U3225) );
  AOI222_X1 U23722 ( .A1(n9595), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20858), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20819), .ZN(n20821) );
  INV_X1 U23723 ( .A(n20821), .ZN(P1_U3226) );
  OAI22_X1 U23724 ( .A1(n20858), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20861), .ZN(n20822) );
  INV_X1 U23725 ( .A(n20822), .ZN(P1_U3458) );
  OAI22_X1 U23726 ( .A1(n20858), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20861), .ZN(n20823) );
  INV_X1 U23727 ( .A(n20823), .ZN(P1_U3459) );
  AOI22_X1 U23728 ( .A1(n20861), .A2(n20825), .B1(n20824), .B2(n20858), .ZN(
        P1_U3460) );
  OAI22_X1 U23729 ( .A1(n20858), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20861), .ZN(n20826) );
  INV_X1 U23730 ( .A(n20826), .ZN(P1_U3461) );
  OAI21_X1 U23731 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20830), .A(n20828), 
        .ZN(n20827) );
  INV_X1 U23732 ( .A(n20827), .ZN(P1_U3464) );
  OAI21_X1 U23733 ( .B1(n20830), .B2(n20829), .A(n20828), .ZN(P1_U3465) );
  INV_X1 U23734 ( .A(n20831), .ZN(n20835) );
  OAI22_X1 U23735 ( .A1(n20835), .A2(n20834), .B1(n20833), .B2(n20832), .ZN(
        n20837) );
  MUX2_X1 U23736 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20837), .S(
        n20836), .Z(P1_U3469) );
  AOI21_X1 U23737 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20839) );
  AOI22_X1 U23738 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20839), .B2(n20838), .ZN(n20841) );
  INV_X1 U23739 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20840) );
  AOI22_X1 U23740 ( .A1(n20842), .A2(n20841), .B1(n20840), .B2(n20845), .ZN(
        P1_U3481) );
  INV_X1 U23741 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20846) );
  NOR2_X1 U23742 ( .A1(n20845), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20843) );
  AOI22_X1 U23743 ( .A1(n20846), .A2(n20845), .B1(n20844), .B2(n20843), .ZN(
        P1_U3482) );
  INV_X1 U23744 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20847) );
  AOI22_X1 U23745 ( .A1(n20861), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20847), 
        .B2(n20858), .ZN(P1_U3483) );
  OAI211_X1 U23746 ( .C1(n20851), .C2(n20850), .A(n20849), .B(n20848), .ZN(
        n20857) );
  OAI211_X1 U23747 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n11172), .A(n20852), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20854) );
  NAND3_X1 U23748 ( .A1(n20857), .A2(n20854), .A3(n20853), .ZN(n20855) );
  OAI21_X1 U23749 ( .B1(n20857), .B2(n20856), .A(n20855), .ZN(P1_U3485) );
  AOI22_X1 U23750 ( .A1(n20861), .A2(n20860), .B1(n20859), .B2(n20858), .ZN(
        P1_U3486) );
  BUF_X1 U11119 ( .A(n10491), .Z(n9602) );
  CLKBUF_X1 U11048 ( .A(n11128), .Z(n13785) );
  CLKBUF_X2 U11058 ( .A(n11138), .Z(n13771) );
  CLKBUF_X1 U11059 ( .A(n11153), .Z(n13054) );
  INV_X2 U11086 ( .A(n12445), .ZN(n16972) );
  INV_X2 U11108 ( .A(n12454), .ZN(n17074) );
  NOR3_X2 U11121 ( .A1(n16381), .A2(n18764), .A3(n13657), .ZN(n15603) );
  CLKBUF_X1 U11168 ( .A(n16362), .Z(n16370) );
  CLKBUF_X1 U11334 ( .A(n11329), .Z(n13773) );
endmodule

