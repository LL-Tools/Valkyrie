

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput63, keyinput62, keyinput61, 
        keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, 
        keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, 
        keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, 
        keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, 
        keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, 
        keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, 
        keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, 
        keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, 
        keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, 
        keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, 
        keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687;

  INV_X1 U3399 ( .A(n5907), .ZN(n5944) );
  CLKBUF_X1 U3400 ( .A(n3469), .Z(n3328) );
  CLKBUF_X1 U3401 ( .A(n3395), .Z(n3308) );
  BUF_X1 U3402 ( .A(n3394), .Z(n3315) );
  CLKBUF_X2 U3403 ( .A(n3239), .Z(n2952) );
  CLKBUF_X1 U3404 ( .A(n3530), .Z(n3945) );
  NOR2_X2 U3405 ( .A1(n4592), .A2(n4474), .ZN(n3348) );
  OR2_X2 U3406 ( .A1(n2982), .A2(n2981), .ZN(n4485) );
  AND2_X1 U3407 ( .A1(n2975), .A2(n4288), .ZN(n3698) );
  AND2_X1 U3408 ( .A1(n2976), .A2(n2975), .ZN(n3314) );
  AND2_X1 U3409 ( .A1(n4067), .A2(n4285), .ZN(n3367) );
  AND2_X1 U3410 ( .A1(n5255), .A2(n4285), .ZN(n3400) );
  AND2_X1 U3411 ( .A1(n2976), .A2(n2974), .ZN(n3723) );
  AND2_X2 U3412 ( .A1(n2973), .A2(n5255), .ZN(n3969) );
  AND2_X2 U3413 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5255) );
  AND4_X1 U3414 ( .A1(n3168), .A2(n3167), .A3(n3166), .A4(n3165), .ZN(n3174)
         );
  AND4_X1 U3415 ( .A1(n3228), .A2(n3227), .A3(n3226), .A4(n3225), .ZN(n2963)
         );
  NOR2_X1 U3416 ( .A1(n3551), .A2(n3550), .ZN(n3552) );
  AND2_X1 U3417 ( .A1(n5799), .A2(n5341), .ZN(n3077) );
  NAND4_X1 U3418 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(n3249)
         );
  AOI21_X1 U3419 ( .B1(n4991), .B2(n5799), .A(n3032), .ZN(n4191) );
  AND2_X1 U3421 ( .A1(n4384), .A2(n4366), .ZN(n4365) );
  NAND2_X1 U3422 ( .A1(n3562), .A2(n2959), .ZN(n4516) );
  NAND2_X1 U3423 ( .A1(n5511), .A2(n5479), .ZN(n5503) );
  AOI211_X1 U3424 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5633), .A(n5387), .B(n5386), .ZN(n5388) );
  INV_X1 U3425 ( .A(n5870), .ZN(n5893) );
  INV_X2 U3427 ( .A(n3423), .ZN(n4507) );
  INV_X2 U3428 ( .A(n5455), .ZN(n5456) );
  NOR2_X2 U3429 ( .A1(n5422), .A2(n5423), .ZN(n5421) );
  AND2_X2 U3430 ( .A1(n3481), .A2(n3510), .ZN(n4216) );
  NAND2_X2 U3431 ( .A1(n5445), .A2(n5275), .ZN(n5455) );
  NAND2_X2 U3432 ( .A1(n4152), .A2(n4151), .ZN(n6041) );
  OR3_X2 U3433 ( .A1(n5448), .A2(n5333), .A3(n5352), .ZN(n2957) );
  NAND2_X1 U3435 ( .A1(n3507), .A2(n3506), .ZN(n4329) );
  INV_X1 U3436 ( .A(n5737), .ZN(n4944) );
  BUF_X2 U3437 ( .A(n3249), .Z(n4491) );
  AND4_X1 U3438 ( .A1(n3010), .A2(n3009), .A3(n3008), .A4(n3007), .ZN(n3021)
         );
  BUF_X2 U3441 ( .A(n3464), .Z(n2951) );
  CLKBUF_X2 U3442 ( .A(n3698), .Z(n3984) );
  BUF_X2 U3443 ( .A(n3400), .Z(n2953) );
  NOR2_X4 U3444 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n2975) );
  INV_X2 U34450 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3444) );
  OAI22_X1 U34460 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n5487), .B1(
        n5497), .B2(n5481), .ZN(n5482) );
  NOR2_X1 U34470 ( .A1(n5201), .A2(n5202), .ZN(n5203) );
  CLKBUF_X1 U34480 ( .A(n5201), .Z(n5207) );
  CLKBUF_X1 U3449 ( .A(n5133), .Z(n5161) );
  INV_X1 U3450 ( .A(n5303), .ZN(n5300) );
  XNOR2_X1 U34510 ( .A(n3649), .B(n3663), .ZN(n4709) );
  NAND2_X1 U34520 ( .A1(n4399), .A2(n4398), .ZN(n4577) );
  NAND2_X1 U34530 ( .A1(n4365), .A2(n3662), .ZN(n4389) );
  CLKBUF_X1 U3454 ( .A(n4365), .Z(n4517) );
  NOR2_X2 U34550 ( .A1(n4329), .A2(n4382), .ZN(n4384) );
  AND2_X2 U34560 ( .A1(n4413), .A2(n4412), .ZN(n5737) );
  XNOR2_X1 U3457 ( .A(n4223), .B(n4222), .ZN(n4561) );
  NAND2_X1 U3458 ( .A1(n4221), .A2(n4220), .ZN(n4223) );
  CLKBUF_X1 U34590 ( .A(n4298), .Z(n4670) );
  AND2_X1 U34610 ( .A1(n3382), .A2(n3418), .ZN(n3415) );
  CLKBUF_X1 U34620 ( .A(n4054), .Z(n5618) );
  CLKBUF_X1 U34630 ( .A(n3387), .Z(n3457) );
  NAND2_X1 U34640 ( .A1(n3289), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U34650 ( .A1(n3028), .A2(n3027), .ZN(n3031) );
  NAND2_X1 U3466 ( .A1(n3351), .A2(n3350), .ZN(n5786) );
  INV_X1 U3467 ( .A(n4503), .ZN(n5437) );
  OR2_X1 U34680 ( .A1(n3334), .A2(n3333), .ZN(n4197) );
  NAND2_X1 U34690 ( .A1(n3423), .A2(n3249), .ZN(n4324) );
  OR2_X1 U34700 ( .A1(n3322), .A2(n3321), .ZN(n4414) );
  AND4_X1 U34710 ( .A1(n3158), .A2(n3157), .A3(n3156), .A4(n3155), .ZN(n3176)
         );
  AND4_X1 U34720 ( .A1(n3018), .A2(n3017), .A3(n3016), .A4(n3015), .ZN(n3019)
         );
  AND4_X1 U34730 ( .A1(n2986), .A2(n2985), .A3(n2984), .A4(n2983), .ZN(n3002)
         );
  AND4_X1 U34740 ( .A1(n2994), .A2(n2993), .A3(n2992), .A4(n2991), .ZN(n3000)
         );
  AND4_X1 U3475 ( .A1(n3006), .A2(n3005), .A3(n3004), .A4(n3003), .ZN(n3022)
         );
  AND4_X1 U3476 ( .A1(n3146), .A2(n3145), .A3(n3144), .A4(n3143), .ZN(n3152)
         );
  AND4_X1 U3477 ( .A1(n3163), .A2(n3162), .A3(n3161), .A4(n3160), .ZN(n3175)
         );
  AND4_X1 U3478 ( .A1(n2990), .A2(n2989), .A3(n2988), .A4(n2987), .ZN(n3001)
         );
  AND4_X1 U3479 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(n3153)
         );
  AND4_X1 U3480 ( .A1(n3138), .A2(n3137), .A3(n3136), .A4(n3135), .ZN(n3154)
         );
  AND4_X1 U3481 ( .A1(n3014), .A2(n3013), .A3(n3012), .A4(n3011), .ZN(n3020)
         );
  BUF_X2 U3482 ( .A(n3367), .Z(n3982) );
  BUF_X2 U3483 ( .A(n3159), .Z(n3983) );
  BUF_X2 U3484 ( .A(n3314), .Z(n3790) );
  AND2_X2 U3485 ( .A1(n6402), .A2(n4307), .ZN(n4378) );
  INV_X2 U3486 ( .A(n6481), .ZN(n6531) );
  AOI22_X1 U3487 ( .A1(n6626), .A2(keyinput34), .B1(n6625), .B2(keyinput12), 
        .ZN(n6624) );
  AND2_X1 U3488 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4285) );
  BUF_X2 U3489 ( .A(n3323), .Z(n2954) );
  AND2_X1 U3490 ( .A1(n2974), .A2(n5255), .ZN(n3239) );
  XNOR2_X1 U3491 ( .A(n4413), .B(n3557), .ZN(n4401) );
  NAND2_X2 U3492 ( .A1(n5457), .A2(n5722), .ZN(n5445) );
  AND2_X2 U3493 ( .A1(n3342), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4067)
         );
  INV_X1 U3494 ( .A(n3024), .ZN(n2956) );
  NAND2_X4 U3495 ( .A1(n4485), .A2(n4474), .ZN(n3024) );
  AOI21_X2 U3496 ( .B1(n5119), .B2(n5118), .A(n5117), .ZN(n5519) );
  NAND2_X2 U3497 ( .A1(n6041), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4202)
         );
  NOR2_X2 U3498 ( .A1(n4351), .A2(n4350), .ZN(n4519) );
  OR2_X2 U3499 ( .A1(n4334), .A2(n4252), .ZN(n4351) );
  NOR3_X4 U3500 ( .A1(n5221), .A2(n5220), .A3(n5219), .ZN(n3103) );
  NAND2_X1 U3501 ( .A1(n5301), .A2(n5342), .ZN(n5303) );
  OAI21_X2 U3502 ( .B1(n5306), .B2(n5305), .A(n5304), .ZN(n5377) );
  NAND2_X1 U3503 ( .A1(n6394), .A2(n6399), .ZN(n4437) );
  NAND2_X1 U3504 ( .A1(n3273), .A2(n3272), .ZN(n4041) );
  INV_X1 U3505 ( .A(n4024), .ZN(n3273) );
  NAND2_X1 U3506 ( .A1(n5133), .A2(n3810), .ZN(n5201) );
  NOR2_X2 U3507 ( .A1(n5145), .A2(n5144), .ZN(n5133) );
  NAND2_X1 U3508 ( .A1(n3643), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3676)
         );
  NAND2_X1 U3509 ( .A1(n4315), .A2(n4188), .ZN(n4187) );
  AND2_X1 U3510 ( .A1(n5115), .A2(n5114), .ZN(n5118) );
  INV_X1 U3511 ( .A(n5116), .ZN(n5117) );
  INV_X1 U3512 ( .A(n3077), .ZN(n3112) );
  INV_X1 U3513 ( .A(n4592), .ZN(n4149) );
  NAND2_X1 U3514 ( .A1(n3360), .A2(n3359), .ZN(n3384) );
  NOR2_X1 U3515 ( .A1(n3357), .A2(n3356), .ZN(n3358) );
  AND2_X2 U3516 ( .A1(n2963), .A2(n2965), .ZN(n3423) );
  OAI21_X1 U3517 ( .B1(n6526), .B2(n4307), .A(n6492), .ZN(n4464) );
  NAND2_X1 U3518 ( .A1(n4149), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3410) );
  NOR2_X1 U3519 ( .A1(n4023), .A2(n4491), .ZN(n3246) );
  NAND2_X1 U3520 ( .A1(n6523), .A2(n3260), .ZN(n5321) );
  INV_X1 U3521 ( .A(n6523), .ZN(n4984) );
  NAND2_X1 U3522 ( .A1(n4365), .A2(n3642), .ZN(n3649) );
  NAND2_X1 U3523 ( .A1(n3525), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3559)
         );
  AND2_X1 U3524 ( .A1(n4138), .A2(n4137), .ZN(n4153) );
  AND2_X1 U3525 ( .A1(n3362), .A2(n3410), .ZN(n3556) );
  XNOR2_X1 U3526 ( .A(n3126), .B(n3125), .ZN(n5534) );
  INV_X1 U3527 ( .A(n5306), .ZN(n3122) );
  OR2_X1 U3528 ( .A1(n4078), .A2(n4077), .ZN(n5963) );
  INV_X1 U3529 ( .A(n5695), .ZN(n5975) );
  OR2_X1 U3530 ( .A1(n4437), .A2(n6359), .ZN(n6042) );
  NOR2_X1 U3531 ( .A1(n6490), .A2(n4066), .ZN(n5254) );
  INV_X1 U3532 ( .A(n6394), .ZN(n4066) );
  INV_X1 U3533 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6402) );
  OR2_X1 U3534 ( .A1(n3406), .A2(n3405), .ZN(n3409) );
  NAND2_X1 U3535 ( .A1(n4740), .A2(n4744), .ZN(n4746) );
  NAND2_X1 U3536 ( .A1(n4739), .A2(n4738), .ZN(n4740) );
  OR2_X1 U3537 ( .A1(n3373), .A2(n3372), .ZN(n4196) );
  NAND2_X1 U3538 ( .A1(n3294), .A2(n3293), .ZN(n4034) );
  AND2_X1 U3539 ( .A1(n4071), .A2(n4503), .ZN(n3271) );
  AND2_X1 U3540 ( .A1(n4592), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3184) );
  AND2_X1 U3541 ( .A1(n5203), .A2(n5216), .ZN(n5215) );
  AND2_X1 U3542 ( .A1(n3808), .A2(n5157), .ZN(n5160) );
  NOR2_X1 U3543 ( .A1(n3714), .A2(n3713), .ZN(n3789) );
  AOI21_X1 U3544 ( .B1(n3426), .B2(n3425), .A(n3424), .ZN(n3449) );
  INV_X1 U3545 ( .A(n3300), .ZN(n4036) );
  AND2_X1 U3546 ( .A1(n5077), .A2(n5082), .ZN(n5115) );
  INV_X1 U3547 ( .A(n4041), .ZN(n4043) );
  OAI221_X1 U3548 ( .B1(n6626), .B2(keyinput34), .C1(n6625), .C2(keyinput12), 
        .A(n6624), .ZN(n6627) );
  INV_X1 U3549 ( .A(n4439), .ZN(n6520) );
  INV_X1 U3550 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3558) );
  INV_X1 U3551 ( .A(n4118), .ZN(n3124) );
  AND2_X1 U3552 ( .A1(n3058), .A2(n3057), .ZN(n4518) );
  INV_X1 U3553 ( .A(n3249), .ZN(n4327) );
  AND2_X1 U3554 ( .A1(n4166), .A2(n5797), .ZN(n5979) );
  OR2_X1 U3555 ( .A1(n3961), .A2(n3960), .ZN(n4011) );
  NOR2_X2 U3556 ( .A1(n5407), .A2(n5337), .ZN(n5357) );
  AND2_X1 U3557 ( .A1(n5421), .A2(n5414), .ZN(n5416) );
  AND2_X1 U3558 ( .A1(n3933), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3934)
         );
  NOR2_X1 U3559 ( .A1(n3892), .A2(n3891), .ZN(n3933) );
  OR2_X1 U3560 ( .A1(n5390), .A2(n5391), .ZN(n5422) );
  NAND2_X1 U3561 ( .A1(n5215), .A2(n5232), .ZN(n5390) );
  CLKBUF_X1 U3562 ( .A(n5215), .Z(n5233) );
  NAND2_X1 U3563 ( .A1(n3853), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3890)
         );
  AND2_X1 U3565 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3715), .ZN(n3716)
         );
  INV_X1 U3566 ( .A(n3750), .ZN(n3715) );
  NAND2_X1 U3567 ( .A1(n3716), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3852)
         );
  AND2_X1 U3568 ( .A1(n5159), .A2(n5158), .ZN(n5236) );
  NOR2_X1 U3569 ( .A1(n3783), .A2(n5819), .ZN(n3751) );
  AND2_X1 U3570 ( .A1(n3789), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3784)
         );
  NAND2_X1 U3571 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n3784), .ZN(n3783)
         );
  NAND2_X1 U3572 ( .A1(n3681), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3714)
         );
  NOR2_X1 U3573 ( .A1(n3676), .A2(n5085), .ZN(n3681) );
  NAND2_X1 U3574 ( .A1(n3665), .A2(n3664), .ZN(n4803) );
  NOR2_X1 U3575 ( .A1(n3625), .A2(n3624), .ZN(n3643) );
  NAND2_X1 U3576 ( .A1(n3594), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3578)
         );
  NAND2_X1 U3577 ( .A1(n4401), .A2(n3425), .ZN(n3562) );
  AOI21_X1 U3578 ( .B1(n4234), .B2(n3425), .A(n3529), .ZN(n4382) );
  INV_X1 U3579 ( .A(n4331), .ZN(n3506) );
  INV_X1 U3580 ( .A(n3482), .ZN(n3483) );
  NAND2_X1 U3581 ( .A1(n3483), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3502)
         );
  CLKBUF_X1 U3582 ( .A(n5457), .Z(n5723) );
  AND2_X1 U3583 ( .A1(n5053), .A2(n4949), .ZN(n5116) );
  NOR2_X2 U3584 ( .A1(n4936), .A2(n4937), .ZN(n4964) );
  AND2_X1 U3585 ( .A1(n5089), .A2(n5093), .ZN(n5079) );
  NAND2_X1 U3586 ( .A1(n4947), .A2(n6059), .ZN(n5089) );
  CLKBUF_X1 U3587 ( .A(n4940), .Z(n4995) );
  AND2_X1 U3588 ( .A1(n3055), .A2(n3054), .ZN(n4350) );
  NAND2_X1 U3589 ( .A1(n4190), .A2(n4332), .ZN(n4334) );
  INV_X1 U3590 ( .A(n4153), .ZN(n4159) );
  AND2_X1 U3591 ( .A1(n5058), .A2(n5062), .ZN(n5284) );
  XNOR2_X1 U3592 ( .A(n3361), .B(n3384), .ZN(n4054) );
  INV_X1 U3593 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3342) );
  CLKBUF_X1 U3594 ( .A(n3342), .Z(n4258) );
  AND2_X1 U3595 ( .A1(n6244), .A2(n4766), .ZN(n4625) );
  NOR2_X1 U3596 ( .A1(n4301), .A2(n3426), .ZN(n6244) );
  AND2_X1 U3597 ( .A1(n4465), .A2(n4464), .ZN(n4508) );
  CLKBUF_X1 U3598 ( .A(n3914), .Z(n4005) );
  OR2_X1 U3599 ( .A1(n4437), .A2(n6346), .ZN(n5628) );
  AND2_X1 U3600 ( .A1(n5321), .A2(n4588), .ZN(n5907) );
  INV_X1 U3601 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5914) );
  NAND2_X1 U3602 ( .A1(n4984), .A2(n3262), .ZN(n5918) );
  INV_X1 U3603 ( .A(n5886), .ZN(n5946) );
  AND2_X1 U3604 ( .A1(n3261), .A2(n3258), .ZN(n5943) );
  CLKBUF_X1 U3605 ( .A(n3440), .Z(n6365) );
  AND2_X1 U3606 ( .A1(n5978), .A2(n4326), .ZN(n5968) );
  OR2_X1 U3607 ( .A1(n5968), .A2(n5971), .ZN(n5974) );
  INV_X1 U3608 ( .A(n5974), .ZN(n4760) );
  NAND2_X1 U3609 ( .A1(n5978), .A2(n4325), .ZN(n5695) );
  NOR2_X1 U3610 ( .A1(n4378), .A2(n5979), .ZN(n5626) );
  INV_X1 U3611 ( .A(n4323), .ZN(n6025) );
  XNOR2_X1 U3612 ( .A(n5357), .B(n5356), .ZN(n5379) );
  INV_X1 U3613 ( .A(n5960), .ZN(n5976) );
  CLKBUF_X1 U3614 ( .A(n4709), .Z(n4711) );
  CLKBUF_X1 U3615 ( .A(n6051), .Z(n6287) );
  INV_X1 U3616 ( .A(n6048), .ZN(n5523) );
  INV_X1 U3617 ( .A(n6040), .ZN(n5525) );
  NAND2_X1 U3618 ( .A1(n5523), .A2(n6047), .ZN(n6040) );
  AND2_X1 U3619 ( .A1(n6042), .A2(n4441), .ZN(n6048) );
  OR2_X1 U3620 ( .A1(n5310), .A2(n5309), .ZN(n5764) );
  NAND2_X1 U3621 ( .A1(n4159), .A2(n6352), .ZN(n5595) );
  CLKBUF_X1 U3622 ( .A(n4299), .Z(n4300) );
  CLKBUF_X1 U3623 ( .A(n4255), .Z(n5621) );
  INV_X1 U3625 ( .A(n5254), .ZN(n6492) );
  AND2_X1 U3626 ( .A1(n4625), .A2(n5009), .ZN(n4648) );
  INV_X1 U3627 ( .A(n6279), .ZN(n6261) );
  INV_X1 U3628 ( .A(n4916), .ZN(n6285) );
  INV_X1 U3629 ( .A(n4930), .ZN(n6299) );
  INV_X1 U3630 ( .A(n4912), .ZN(n6311) );
  INV_X1 U3631 ( .A(n4908), .ZN(n6317) );
  INV_X1 U3632 ( .A(n4900), .ZN(n6329) );
  NOR2_X1 U3633 ( .A1(n6117), .A2(n4815), .ZN(n6339) );
  INV_X1 U3634 ( .A(n4924), .ZN(n6335) );
  NAND2_X1 U3635 ( .A1(n3213), .A2(n3212), .ZN(n6394) );
  OR2_X1 U3636 ( .A1(n3211), .A2(n3255), .ZN(n3212) );
  OAI21_X1 U3637 ( .B1(n3255), .B2(n3556), .A(n3210), .ZN(n3213) );
  AND2_X1 U3638 ( .A1(n6392), .A2(n6391), .ZN(n6486) );
  AOI21_X1 U3639 ( .B1(n5453), .B2(n5870), .A(n4018), .ZN(n4019) );
  BUF_X2 U3641 ( .A(n3316), .Z(n3970) );
  INV_X1 U3642 ( .A(n3103), .ZN(n5394) );
  OR2_X1 U3643 ( .A1(n5379), .A2(n6051), .ZN(n2958) );
  NAND2_X1 U3644 ( .A1(n4341), .A2(n4340), .ZN(n4396) );
  AND2_X1 U3645 ( .A1(n4964), .A2(n4963), .ZN(n4962) );
  AND2_X1 U3646 ( .A1(n2973), .A2(n4288), .ZN(n3464) );
  AND2_X1 U3647 ( .A1(n4191), .A2(n3041), .ZN(n4190) );
  NOR2_X2 U3648 ( .A1(n6287), .A2(n4493), .ZN(n6325) );
  NOR2_X2 U3649 ( .A1(n6287), .A2(n4511), .ZN(n6331) );
  NOR4_X2 U3650 ( .A1(n5811), .A2(n5810), .A3(n5809), .A4(n5808), .ZN(n6510)
         );
  NOR2_X2 U3651 ( .A1(n6287), .A2(n4499), .ZN(n6319) );
  NOR2_X2 U3652 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6521) );
  AND2_X1 U3653 ( .A1(n3561), .A2(n2961), .ZN(n2959) );
  INV_X1 U3654 ( .A(n3680), .ZN(n3425) );
  NAND2_X1 U3655 ( .A1(n6402), .A2(n4464), .ZN(n4770) );
  AND2_X1 U3656 ( .A1(n5434), .A2(n5235), .ZN(n2960) );
  INV_X2 U3657 ( .A(n4474), .ZN(n3276) );
  OR2_X1 U3658 ( .A1(n4581), .A2(n4003), .ZN(n2961) );
  NAND2_X1 U3659 ( .A1(n4947), .A2(n5756), .ZN(n2962) );
  NOR2_X1 U3660 ( .A1(n4994), .A2(n4941), .ZN(n2964) );
  AND2_X1 U3661 ( .A1(n4491), .A2(n4474), .ZN(n4400) );
  AOI21_X1 U3662 ( .B1(n5167), .B2(n6402), .A(n3477), .ZN(n4303) );
  OAI21_X1 U3663 ( .B1(n3457), .B2(n5263), .A(n3393), .ZN(n3455) );
  INV_X1 U3664 ( .A(n4216), .ZN(n4301) );
  AND4_X1 U3665 ( .A1(n3232), .A2(n3231), .A3(n3230), .A4(n3229), .ZN(n2965)
         );
  AND2_X1 U3666 ( .A1(n4214), .A2(n4213), .ZN(n2966) );
  INV_X1 U3667 ( .A(n3234), .ZN(n3836) );
  OAI21_X1 U3668 ( .B1(n3556), .B2(n3276), .A(n4491), .ZN(n3188) );
  OR2_X1 U3669 ( .A1(n4139), .A2(n3024), .ZN(n3298) );
  OR2_X1 U3670 ( .A1(n4324), .A2(n4497), .ZN(n3270) );
  INV_X1 U3671 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n2968) );
  NAND2_X1 U3672 ( .A1(n3271), .A2(n3270), .ZN(n4024) );
  OAI211_X1 U3673 ( .C1(n6346), .C2(n3352), .A(n4155), .B(n5786), .ZN(n3353)
         );
  AOI21_X1 U3674 ( .B1(n3341), .B2(n3438), .A(n4409), .ZN(n3417) );
  INV_X1 U3675 ( .A(n4023), .ZN(n3272) );
  AND2_X1 U3676 ( .A1(n5091), .A2(n4996), .ZN(n4945) );
  AND2_X1 U3677 ( .A1(n3347), .A2(n3346), .ZN(n4056) );
  AND3_X1 U3678 ( .A1(n3305), .A2(n3304), .A3(n3303), .ZN(n3306) );
  AND2_X1 U3679 ( .A1(n3184), .A2(n4497), .ZN(n3337) );
  AND2_X1 U3680 ( .A1(n3809), .A2(n5160), .ZN(n3810) );
  OR2_X1 U3681 ( .A1(n4497), .A2(n6402), .ZN(n3362) );
  INV_X1 U3682 ( .A(n3645), .ZN(n3424) );
  AND4_X1 U3683 ( .A1(n3172), .A2(n3171), .A3(n3170), .A4(n3169), .ZN(n3173)
         );
  OR2_X1 U3684 ( .A1(n3959), .A2(n3958), .ZN(n3961) );
  INV_X1 U3685 ( .A(n4400), .ZN(n4410) );
  AND2_X1 U3686 ( .A1(n4946), .A2(n4945), .ZN(n5077) );
  AND2_X1 U3687 ( .A1(n5318), .A2(n4192), .ZN(n3041) );
  NAND2_X1 U3688 ( .A1(n2956), .A2(n3033), .ZN(n3042) );
  NAND2_X1 U3689 ( .A1(n4034), .A2(n3306), .ZN(n3359) );
  NAND2_X1 U3690 ( .A1(n3423), .A2(n4503), .ZN(n3300) );
  INV_X1 U3691 ( .A(n3337), .ZN(n3553) );
  AOI21_X1 U3692 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6402), .A(n3209), 
        .ZN(n3210) );
  OR2_X1 U3693 ( .A1(n6504), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4439) );
  OR2_X1 U3694 ( .A1(n3042), .A2(EBX_REG_1__SCAN_IN), .ZN(n3028) );
  OR2_X1 U3696 ( .A1(n6366), .A2(n6402), .ZN(n3979) );
  INV_X1 U3697 ( .A(n3033), .ZN(n3064) );
  AND4_X1 U3698 ( .A1(n2998), .A2(n2997), .A3(n2996), .A4(n2995), .ZN(n2999)
         );
  NOR2_X1 U3699 ( .A1(n3852), .A2(n5498), .ZN(n3853) );
  OR2_X1 U3700 ( .A1(n5746), .A2(n5436), .ZN(n5434) );
  NOR2_X1 U3701 ( .A1(n3559), .A2(n3558), .ZN(n3560) );
  NOR2_X1 U3702 ( .A1(n5737), .A2(n5470), .ZN(n5276) );
  INV_X1 U3703 ( .A(n3552), .ZN(n4413) );
  NOR2_X1 U3704 ( .A1(n5009), .A2(n4410), .ZN(n4148) );
  INV_X1 U3705 ( .A(n6170), .ZN(n4767) );
  NAND2_X1 U3706 ( .A1(n3463), .A2(n3462), .ZN(n6207) );
  AND2_X1 U3707 ( .A1(n4592), .A2(n4474), .ZN(n3033) );
  NAND2_X1 U3708 ( .A1(n3934), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3959)
         );
  OR3_X1 U3709 ( .A1(n6451), .A2(n4014), .A3(n5913), .ZN(n4970) );
  INV_X1 U3710 ( .A(n3573), .ZN(n3594) );
  NOR2_X1 U3711 ( .A1(n3502), .A2(n5914), .ZN(n3525) );
  INV_X1 U3712 ( .A(n3024), .ZN(n5237) );
  NAND2_X1 U3713 ( .A1(n5416), .A2(n5405), .ZN(n5407) );
  OR2_X1 U3714 ( .A1(n3890), .A2(n5483), .ZN(n3892) );
  OR2_X1 U3715 ( .A1(n5744), .A2(n5743), .ZN(n5746) );
  NOR2_X1 U3716 ( .A1(n6625), .A2(n3578), .ZN(n3619) );
  AND2_X1 U3717 ( .A1(n4215), .A2(n6031), .ZN(n4560) );
  NAND2_X1 U3718 ( .A1(n5456), .A2(n5276), .ZN(n5465) );
  INV_X1 U3719 ( .A(n5737), .ZN(n5517) );
  NOR2_X1 U3720 ( .A1(n5065), .A2(n5103), .ZN(n5310) );
  NOR2_X2 U3721 ( .A1(n4586), .A2(n4392), .ZN(n4572) );
  NAND2_X1 U3722 ( .A1(n4521), .A2(n4426), .ZN(n4807) );
  NAND2_X1 U3723 ( .A1(n4233), .A2(n4232), .ZN(n4338) );
  OR2_X1 U3724 ( .A1(n5284), .A2(n4245), .ZN(n4958) );
  AND2_X1 U3725 ( .A1(n3109), .A2(n5341), .ZN(n4118) );
  NAND2_X1 U3726 ( .A1(n3478), .A2(n3422), .ZN(n4298) );
  INV_X1 U3727 ( .A(n4300), .ZN(n4766) );
  INV_X1 U3728 ( .A(n6339), .ZN(n4844) );
  AND2_X1 U3730 ( .A1(n5321), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5901) );
  AND2_X1 U3731 ( .A1(n5321), .A2(n4013), .ZN(n5870) );
  NAND2_X1 U3732 ( .A1(n3123), .A2(n3122), .ZN(n3126) );
  NAND2_X1 U3733 ( .A1(n4962), .A2(n5123), .ZN(n5767) );
  AND2_X1 U3734 ( .A1(n4519), .A2(n4518), .ZN(n4521) );
  INV_X1 U3735 ( .A(n5958), .ZN(n5953) );
  AND2_X1 U3736 ( .A1(n5978), .A2(n4328), .ZN(n5971) );
  INV_X1 U3737 ( .A(n5978), .ZN(n5970) );
  AND2_X1 U3738 ( .A1(n5407), .A2(n5406), .ZN(n5696) );
  NAND2_X1 U3739 ( .A1(n3751), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3750)
         );
  AND2_X1 U3740 ( .A1(n5746), .A2(n5745), .ZN(n5969) );
  NAND2_X1 U3741 ( .A1(n4803), .A2(n4802), .ZN(n5145) );
  AND2_X1 U3742 ( .A1(n4433), .A2(n4432), .ZN(n4727) );
  NAND2_X1 U3743 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3482) );
  INV_X1 U3744 ( .A(n5278), .ZN(n5279) );
  OAI211_X1 U3745 ( .C1(n5335), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5334), .B(n2957), .ZN(n5336) );
  OR2_X1 U3746 ( .A1(n5509), .A2(n5508), .ZN(n5511) );
  INV_X1 U3747 ( .A(n6082), .ZN(n6109) );
  INV_X1 U3748 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3388) );
  INV_X1 U3749 ( .A(n5197), .ZN(n4705) );
  INV_X1 U3750 ( .A(n4702), .ZN(n6164) );
  NOR2_X1 U3751 ( .A1(n5010), .A2(n5176), .ZN(n5011) );
  INV_X1 U3752 ( .A(n6177), .ZN(n6200) );
  NOR2_X1 U3753 ( .A1(n4670), .A2(n3479), .ZN(n6172) );
  OR3_X1 U3754 ( .A1(n4528), .A2(n4527), .A3(n4526), .ZN(n4553) );
  INV_X1 U3755 ( .A(n5009), .ZN(n5176) );
  INV_X1 U3756 ( .A(n4890), .ZN(n4932) );
  INV_X1 U3757 ( .A(n6265), .ZN(n6273) );
  AND2_X1 U3758 ( .A1(n4814), .A2(n5009), .ZN(n4884) );
  AND2_X1 U3759 ( .A1(n4814), .A2(n5176), .ZN(n4882) );
  OAI21_X1 U3760 ( .B1(n4821), .B2(n6490), .A(n4820), .ZN(n4843) );
  INV_X1 U3761 ( .A(n4920), .ZN(n6305) );
  INV_X1 U3762 ( .A(n4904), .ZN(n6323) );
  AND2_X1 U3763 ( .A1(n4300), .A2(n5176), .ZN(n6118) );
  INV_X1 U3764 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6403) );
  AND2_X1 U3765 ( .A1(n5628), .A2(n5630), .ZN(n6523) );
  INV_X1 U3766 ( .A(n5901), .ZN(n5945) );
  INV_X1 U3767 ( .A(n5943), .ZN(n5933) );
  AND2_X1 U3768 ( .A1(n4985), .A2(n5893), .ZN(n5951) );
  OR2_X1 U3769 ( .A1(n2960), .A2(n5236), .ZN(n5719) );
  NAND2_X1 U3770 ( .A1(n4323), .A2(n4322), .ZN(n5978) );
  INV_X1 U3771 ( .A(n5979), .ZN(n6007) );
  AND2_X1 U3772 ( .A1(n2958), .A2(n5364), .ZN(n5365) );
  OR2_X1 U3773 ( .A1(n4728), .A2(n4727), .ZN(n5881) );
  XNOR2_X1 U3774 ( .A(n5279), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5366)
         );
  OR2_X1 U3775 ( .A1(n5571), .A2(n5312), .ZN(n5755) );
  INV_X1 U3776 ( .A(n6112), .ZN(n6084) );
  INV_X1 U3777 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5169) );
  INV_X1 U3778 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6382) );
  INV_X1 U3779 ( .A(n4648), .ZN(n4559) );
  NAND2_X1 U3780 ( .A1(n6288), .A2(n6118), .ZN(n6344) );
  INV_X1 U3781 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U3782 ( .A1(n4020), .A2(n4019), .ZN(U2796) );
  AND2_X2 U3783 ( .A1(n3444), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n2976)
         );
  NOR2_X2 U3784 ( .A1(n3388), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n2974)
         );
  AOI22_X1 U3785 ( .A1(n3723), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n2972) );
  AND2_X2 U3786 ( .A1(n2968), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n2973)
         );
  AND2_X2 U3787 ( .A1(n2973), .A2(n2976), .ZN(n3159) );
  AND2_X2 U3788 ( .A1(n2976), .A2(n4285), .ZN(n3323) );
  AOI22_X1 U3789 ( .A1(n3159), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n2954), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n2971) );
  AOI22_X1 U3790 ( .A1(n3969), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3239), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n2970) );
  NOR2_X4 U3792 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4288) );
  AND2_X2 U3793 ( .A1(n4288), .A2(n4285), .ZN(n3224) );
  AOI22_X1 U3794 ( .A1(n3316), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n2969) );
  NAND4_X1 U3795 ( .A1(n2972), .A2(n2971), .A3(n2970), .A4(n2969), .ZN(n2982)
         );
  AND2_X2 U3796 ( .A1(n4067), .A2(n2975), .ZN(n3394) );
  AND2_X2 U3797 ( .A1(n4067), .A2(n2974), .ZN(n3395) );
  AOI22_X1 U3798 ( .A1(n3394), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n2980) );
  AND2_X2 U3799 ( .A1(n2974), .A2(n4288), .ZN(n3530) );
  AOI22_X1 U3800 ( .A1(n3464), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n2979) );
  AND2_X2 U3801 ( .A1(n2975), .A2(n5255), .ZN(n3469) );
  AOI22_X1 U3802 ( .A1(n3698), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n2978) );
  AOI22_X1 U3803 ( .A1(n3314), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n2977) );
  NAND4_X1 U3804 ( .A1(n2980), .A2(n2979), .A3(n2978), .A4(n2977), .ZN(n2981)
         );
  NAND2_X1 U3805 ( .A1(n2954), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n2986)
         );
  NAND2_X1 U3806 ( .A1(n3159), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n2985)
         );
  NAND2_X1 U3807 ( .A1(n3395), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n2984) );
  NAND2_X1 U3808 ( .A1(n3367), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n2983)
         );
  NAND2_X1 U3809 ( .A1(n3464), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n2990) );
  NAND2_X1 U3810 ( .A1(n3969), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n2989)
         );
  NAND2_X1 U3811 ( .A1(n3394), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n2988) );
  NAND2_X1 U3812 ( .A1(n3530), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n2987) );
  NAND2_X1 U3813 ( .A1(n3316), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n2994) );
  NAND2_X1 U3814 ( .A1(n3314), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n2993) );
  NAND2_X1 U3815 ( .A1(n3698), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n2992) );
  NAND2_X1 U3816 ( .A1(n3469), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n2991) );
  NAND2_X1 U3817 ( .A1(n3723), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n2998) );
  NAND2_X1 U3818 ( .A1(n3239), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n2997) );
  NAND2_X1 U3819 ( .A1(n3400), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n2996)
         );
  NAND2_X1 U3820 ( .A1(n3224), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n2995)
         );
  NAND4_X4 U3821 ( .A1(n3002), .A2(n3001), .A3(n3000), .A4(n2999), .ZN(n4474)
         );
  NAND2_X1 U3822 ( .A1(n3394), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3006) );
  NAND2_X1 U3823 ( .A1(n3159), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3005)
         );
  NAND2_X1 U3824 ( .A1(n3395), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3004) );
  NAND2_X1 U3825 ( .A1(n2955), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3003)
         );
  NAND2_X1 U3826 ( .A1(n3464), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3010) );
  NAND2_X1 U3827 ( .A1(n3723), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3009) );
  NAND2_X1 U3828 ( .A1(n3367), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3008)
         );
  NAND2_X1 U3829 ( .A1(n3530), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3007) );
  NAND2_X1 U3830 ( .A1(n3314), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3014) );
  NAND2_X1 U3831 ( .A1(n3969), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3013)
         );
  NAND2_X1 U3832 ( .A1(n3239), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3012) );
  NAND2_X1 U3833 ( .A1(n3400), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3011)
         );
  NAND2_X1 U3834 ( .A1(n3316), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3018) );
  NAND2_X1 U3835 ( .A1(n3698), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3017) );
  NAND2_X1 U3836 ( .A1(n3469), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3016) );
  NAND2_X1 U3837 ( .A1(n3224), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3015)
         );
  NAND4_X4 U3838 ( .A1(n3022), .A2(n3021), .A3(n3020), .A4(n3019), .ZN(n4592)
         );
  INV_X1 U3839 ( .A(n4485), .ZN(n4073) );
  NAND2_X1 U3840 ( .A1(n4073), .A2(n4592), .ZN(n3073) );
  INV_X1 U3841 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3023) );
  NAND2_X1 U3842 ( .A1(n3073), .A2(n3023), .ZN(n3026) );
  NAND2_X1 U3843 ( .A1(n3033), .A2(n4988), .ZN(n3025) );
  NAND3_X1 U3844 ( .A1(n3026), .A2(n5341), .A3(n3025), .ZN(n3027) );
  NAND2_X1 U3845 ( .A1(n3073), .A2(EBX_REG_0__SCAN_IN), .ZN(n3030) );
  INV_X1 U3846 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4123) );
  NAND2_X1 U3847 ( .A1(n5341), .A2(n4123), .ZN(n3029) );
  NAND2_X1 U3848 ( .A1(n3030), .A2(n3029), .ZN(n4116) );
  XNOR2_X1 U3849 ( .A(n3031), .B(n4116), .ZN(n4991) );
  INV_X1 U3850 ( .A(n3031), .ZN(n3032) );
  INV_X1 U3851 ( .A(n3073), .ZN(n3056) );
  NAND2_X1 U3852 ( .A1(n3056), .A2(n3064), .ZN(n3082) );
  NAND2_X1 U3853 ( .A1(n3064), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3034)
         );
  AND2_X1 U3854 ( .A1(n3082), .A2(n3034), .ZN(n3036) );
  MUX2_X1 U3855 ( .A(n3042), .B(n3073), .S(EBX_REG_2__SCAN_IN), .Z(n3035) );
  NAND2_X1 U3856 ( .A1(n3036), .A2(n3035), .ZN(n5318) );
  INV_X1 U3857 ( .A(EBX_REG_3__SCAN_IN), .ZN(n3037) );
  NAND2_X1 U3858 ( .A1(n3077), .A2(n3037), .ZN(n3040) );
  INV_X1 U3859 ( .A(n3056), .ZN(n3109) );
  NAND2_X1 U3860 ( .A1(n5341), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3038)
         );
  OAI211_X1 U3861 ( .C1(n3064), .C2(EBX_REG_3__SCAN_IN), .A(n3109), .B(n3038), 
        .ZN(n3039) );
  AND2_X1 U3862 ( .A1(n3040), .A2(n3039), .ZN(n4192) );
  OR2_X1 U3863 ( .A1(n3120), .A2(EBX_REG_4__SCAN_IN), .ZN(n3047) );
  INV_X1 U3864 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4361) );
  NAND2_X1 U3865 ( .A1(n3073), .A2(n4361), .ZN(n3045) );
  BUF_X2 U3866 ( .A(n3024), .Z(n5341) );
  INV_X1 U3867 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3043) );
  NAND2_X1 U3868 ( .A1(n5799), .A2(n3043), .ZN(n3044) );
  NAND3_X1 U3869 ( .A1(n3045), .A2(n5341), .A3(n3044), .ZN(n3046) );
  NAND2_X1 U3870 ( .A1(n3047), .A2(n3046), .ZN(n4332) );
  BUF_X1 U3871 ( .A(n3064), .Z(n3049) );
  NAND2_X1 U3872 ( .A1(n5341), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3048)
         );
  OAI211_X1 U3873 ( .C1(n3049), .C2(EBX_REG_5__SCAN_IN), .A(n3073), .B(n3048), 
        .ZN(n3050) );
  OAI21_X1 U3874 ( .B1(n3112), .B2(EBX_REG_5__SCAN_IN), .A(n3050), .ZN(n4252)
         );
  OR2_X1 U3875 ( .A1(n3120), .A2(EBX_REG_6__SCAN_IN), .ZN(n3055) );
  INV_X1 U3876 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4346) );
  NAND2_X1 U3877 ( .A1(n3109), .A2(n4346), .ZN(n3053) );
  INV_X1 U3878 ( .A(EBX_REG_6__SCAN_IN), .ZN(n3051) );
  NAND2_X1 U3879 ( .A1(n5799), .A2(n3051), .ZN(n3052) );
  NAND3_X1 U3880 ( .A1(n3053), .A2(n5341), .A3(n3052), .ZN(n3054) );
  MUX2_X1 U3881 ( .A(n3112), .B(n5341), .S(EBX_REG_7__SCAN_IN), .Z(n3058) );
  INV_X1 U3882 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U3883 ( .A1(n6077), .A2(n4118), .ZN(n3057) );
  OR2_X1 U3884 ( .A1(n3120), .A2(EBX_REG_8__SCAN_IN), .ZN(n3062) );
  INV_X1 U3885 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4419) );
  NAND2_X1 U3886 ( .A1(n3109), .A2(n4419), .ZN(n3060) );
  INV_X1 U3887 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4613) );
  NAND2_X1 U3888 ( .A1(n5799), .A2(n4613), .ZN(n3059) );
  NAND3_X1 U3889 ( .A1(n3060), .A2(n5341), .A3(n3059), .ZN(n3061) );
  NAND2_X1 U3890 ( .A1(n3062), .A2(n3061), .ZN(n4426) );
  MUX2_X1 U3891 ( .A(n3112), .B(n3024), .S(EBX_REG_9__SCAN_IN), .Z(n3063) );
  OAI21_X1 U3892 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n3124), .A(n3063), 
        .ZN(n4808) );
  OR2_X2 U3893 ( .A1(n4807), .A2(n4808), .ZN(n4805) );
  MUX2_X1 U3894 ( .A(n3120), .B(n3073), .S(EBX_REG_10__SCAN_IN), .Z(n3066) );
  NAND2_X1 U3895 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n3049), .ZN(n3065) );
  AND3_X1 U3896 ( .A1(n3066), .A2(n3082), .A3(n3065), .ZN(n4584) );
  OR2_X2 U3897 ( .A1(n4805), .A2(n4584), .ZN(n4586) );
  NAND2_X1 U3898 ( .A1(n3024), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3067) );
  OAI211_X1 U3899 ( .C1(n3049), .C2(EBX_REG_11__SCAN_IN), .A(n3073), .B(n3067), 
        .ZN(n3068) );
  OAI21_X1 U3900 ( .B1(n3112), .B2(EBX_REG_11__SCAN_IN), .A(n3068), .ZN(n4392)
         );
  NAND2_X1 U3901 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n3049), .ZN(n3069) );
  AND2_X1 U3902 ( .A1(n3082), .A2(n3069), .ZN(n3071) );
  MUX2_X1 U3903 ( .A(n3120), .B(n3109), .S(EBX_REG_12__SCAN_IN), .Z(n3070) );
  NAND2_X1 U3904 ( .A1(n3071), .A2(n3070), .ZN(n4571) );
  NAND2_X1 U3905 ( .A1(n4572), .A2(n4571), .ZN(n4570) );
  NAND2_X1 U3906 ( .A1(n3024), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3072) );
  OAI211_X1 U3907 ( .C1(n3049), .C2(EBX_REG_13__SCAN_IN), .A(n3073), .B(n3072), 
        .ZN(n3074) );
  OAI21_X1 U3908 ( .B1(n3112), .B2(EBX_REG_13__SCAN_IN), .A(n3074), .ZN(n4712)
         );
  OR2_X2 U3909 ( .A1(n4570), .A2(n4712), .ZN(n4936) );
  MUX2_X1 U3910 ( .A(n3120), .B(n3109), .S(EBX_REG_14__SCAN_IN), .Z(n3076) );
  NAND2_X1 U3911 ( .A1(n3049), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3075) );
  AND3_X1 U3912 ( .A1(n3076), .A2(n3082), .A3(n3075), .ZN(n4937) );
  INV_X1 U3913 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U3914 ( .A1(n3077), .A2(n5964), .ZN(n3080) );
  NAND2_X1 U3915 ( .A1(n3024), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3078) );
  OAI211_X1 U3916 ( .C1(n3049), .C2(EBX_REG_15__SCAN_IN), .A(n3109), .B(n3078), 
        .ZN(n3079) );
  AND2_X1 U3917 ( .A1(n3080), .A2(n3079), .ZN(n4963) );
  NAND2_X1 U3918 ( .A1(n3049), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3081) );
  AND2_X1 U3919 ( .A1(n3082), .A2(n3081), .ZN(n3084) );
  MUX2_X1 U3920 ( .A(n3120), .B(n3109), .S(EBX_REG_16__SCAN_IN), .Z(n3083) );
  NAND2_X1 U3921 ( .A1(n3084), .A2(n3083), .ZN(n5123) );
  NAND2_X1 U3922 ( .A1(n3024), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3085) );
  OAI211_X1 U3923 ( .C1(n3049), .C2(EBX_REG_17__SCAN_IN), .A(n3109), .B(n3085), 
        .ZN(n3086) );
  OAI21_X1 U3924 ( .B1(n3112), .B2(EBX_REG_17__SCAN_IN), .A(n3086), .ZN(n5766)
         );
  OR2_X2 U3925 ( .A1(n5767), .A2(n5766), .ZN(n5769) );
  OR2_X1 U3926 ( .A1(n3120), .A2(EBX_REG_19__SCAN_IN), .ZN(n3089) );
  INV_X1 U3927 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U3928 ( .A1(n3109), .A2(n5762), .ZN(n3087) );
  OAI211_X1 U3929 ( .C1(EBX_REG_19__SCAN_IN), .C2(n3049), .A(n3087), .B(n3024), 
        .ZN(n3088) );
  AND2_X1 U3930 ( .A1(n3089), .A2(n3088), .ZN(n5240) );
  NOR2_X2 U3931 ( .A1(n5769), .A2(n5240), .ZN(n5163) );
  INV_X1 U3932 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5603) );
  NOR2_X1 U3933 ( .A1(n3049), .A2(EBX_REG_20__SCAN_IN), .ZN(n3090) );
  AOI21_X1 U3934 ( .B1(n4118), .B2(n5603), .A(n3090), .ZN(n5164) );
  OR2_X1 U3935 ( .A1(n3124), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3092)
         );
  INV_X1 U3936 ( .A(EBX_REG_18__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U3937 ( .A1(n5799), .A2(n3091), .ZN(n5238) );
  NAND2_X1 U3938 ( .A1(n3092), .A2(n5238), .ZN(n5239) );
  NAND2_X1 U3939 ( .A1(n5237), .A2(EBX_REG_20__SCAN_IN), .ZN(n3094) );
  NAND2_X1 U3940 ( .A1(n5239), .A2(n3024), .ZN(n3093) );
  OAI211_X1 U3941 ( .C1(n5164), .C2(n5239), .A(n3094), .B(n3093), .ZN(n3095)
         );
  INV_X1 U3942 ( .A(n3095), .ZN(n3096) );
  AND2_X2 U3943 ( .A1(n5163), .A2(n3096), .ZN(n5212) );
  MUX2_X1 U3944 ( .A(n3112), .B(n3024), .S(EBX_REG_21__SCAN_IN), .Z(n3098) );
  OR2_X1 U3945 ( .A1(n3124), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3097)
         );
  AND2_X1 U3946 ( .A1(n3098), .A2(n3097), .ZN(n5211) );
  NAND2_X2 U3947 ( .A1(n5212), .A2(n5211), .ZN(n5221) );
  MUX2_X1 U3948 ( .A(n3120), .B(n3109), .S(EBX_REG_22__SCAN_IN), .Z(n3100) );
  NAND2_X1 U3949 ( .A1(n3049), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3099) );
  AND2_X1 U3950 ( .A1(n3100), .A2(n3099), .ZN(n5220) );
  NAND2_X1 U3951 ( .A1(n3024), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3101) );
  OAI211_X1 U3952 ( .C1(EBX_REG_23__SCAN_IN), .C2(n3049), .A(n3109), .B(n3101), 
        .ZN(n3102) );
  OAI21_X1 U3953 ( .B1(n3112), .B2(EBX_REG_23__SCAN_IN), .A(n3102), .ZN(n5219)
         );
  MUX2_X1 U3954 ( .A(n3112), .B(n3024), .S(EBX_REG_25__SCAN_IN), .Z(n3105) );
  OR2_X1 U3955 ( .A1(n3124), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3104)
         );
  AND2_X1 U3956 ( .A1(n3105), .A2(n3104), .ZN(n5395) );
  MUX2_X1 U3957 ( .A(n3120), .B(n3109), .S(EBX_REG_24__SCAN_IN), .Z(n3107) );
  NAND2_X1 U3958 ( .A1(n3049), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3106) );
  NAND2_X1 U3959 ( .A1(n3107), .A2(n3106), .ZN(n5396) );
  NAND2_X1 U3960 ( .A1(n5395), .A2(n5396), .ZN(n3108) );
  NOR2_X2 U3961 ( .A1(n5394), .A2(n3108), .ZN(n5425) );
  MUX2_X1 U3962 ( .A(n3120), .B(n3109), .S(EBX_REG_26__SCAN_IN), .Z(n3111) );
  NAND2_X1 U3963 ( .A1(n3049), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3110) );
  NAND2_X1 U3964 ( .A1(n3111), .A2(n3110), .ZN(n5424) );
  NAND2_X1 U3965 ( .A1(n5425), .A2(n5424), .ZN(n5427) );
  MUX2_X1 U3966 ( .A(n3112), .B(n3024), .S(EBX_REG_27__SCAN_IN), .Z(n3113) );
  OAI21_X1 U3967 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n3124), .A(n3113), 
        .ZN(n5417) );
  OR2_X2 U3968 ( .A1(n5427), .A2(n5417), .ZN(n5419) );
  OR2_X1 U3969 ( .A1(n3120), .A2(EBX_REG_28__SCAN_IN), .ZN(n3118) );
  INV_X1 U3970 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3114) );
  NAND2_X1 U3971 ( .A1(n3109), .A2(n3114), .ZN(n3116) );
  INV_X1 U3972 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U3973 ( .A1(n5799), .A2(n5413), .ZN(n3115) );
  NAND3_X1 U3974 ( .A1(n3116), .A2(n3024), .A3(n3115), .ZN(n3117) );
  AND2_X1 U3975 ( .A1(n3118), .A2(n3117), .ZN(n5408) );
  NOR2_X4 U3976 ( .A1(n5419), .A2(n5408), .ZN(n5301) );
  INV_X1 U3977 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5352) );
  NOR2_X1 U3978 ( .A1(n3049), .A2(EBX_REG_29__SCAN_IN), .ZN(n3119) );
  AOI21_X1 U3979 ( .B1(n4118), .B2(n5352), .A(n3119), .ZN(n5342) );
  OR2_X1 U3980 ( .A1(n3120), .A2(EBX_REG_29__SCAN_IN), .ZN(n5343) );
  INV_X1 U3981 ( .A(n5301), .ZN(n5299) );
  OAI22_X1 U3982 ( .A1(n5303), .A2(n5237), .B1(n5343), .B2(n5299), .ZN(n5347)
         );
  AND2_X1 U3983 ( .A1(n3049), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3121)
         );
  AOI21_X1 U3984 ( .B1(n3124), .B2(EBX_REG_30__SCAN_IN), .A(n3121), .ZN(n5302)
         );
  NAND2_X1 U3985 ( .A1(n5347), .A2(n5302), .ZN(n3123) );
  NOR2_X1 U3986 ( .A1(n5300), .A2(n5237), .ZN(n5306) );
  OAI22_X1 U3987 ( .A1(n3124), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n3049), .ZN(n3125) );
  NAND2_X1 U3988 ( .A1(n5169), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3179) );
  INV_X1 U3989 ( .A(n3179), .ZN(n3177) );
  XNOR2_X1 U3990 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3178) );
  NAND2_X1 U3991 ( .A1(n3177), .A2(n3178), .ZN(n3128) );
  INV_X1 U3992 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U3993 ( .A1(n6374), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3127) );
  NAND2_X1 U3994 ( .A1(n3128), .A2(n3127), .ZN(n3195) );
  XNOR2_X1 U3995 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3193) );
  NAND2_X1 U3996 ( .A1(n3195), .A2(n3193), .ZN(n3130) );
  INV_X1 U3997 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U3998 ( .A1(n5168), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3129) );
  NAND2_X1 U3999 ( .A1(n3130), .A2(n3129), .ZN(n3199) );
  XNOR2_X1 U4000 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3200) );
  NAND2_X1 U4001 ( .A1(n3199), .A2(n3200), .ZN(n3132) );
  NAND2_X1 U4002 ( .A1(n6382), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U4003 ( .A1(n3132), .A2(n3131), .ZN(n3206) );
  INV_X1 U4004 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6381) );
  AND2_X1 U4005 ( .A1(n6381), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3133)
         );
  OR2_X1 U4006 ( .A1(n3206), .A2(n3133), .ZN(n3134) );
  INV_X1 U4007 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4293) );
  NAND2_X1 U4008 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4293), .ZN(n3205) );
  NAND2_X1 U4009 ( .A1(n3134), .A2(n3205), .ZN(n3255) );
  NAND2_X1 U4010 ( .A1(n3314), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U4011 ( .A1(n3969), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3137)
         );
  NAND2_X1 U4012 ( .A1(n3239), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U4013 ( .A1(n3400), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3135)
         );
  NAND2_X1 U4014 ( .A1(n3464), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U4015 ( .A1(n3723), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U4016 ( .A1(n3367), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3140)
         );
  NAND2_X1 U4017 ( .A1(n3530), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3139) );
  NAND2_X1 U4018 ( .A1(n3394), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3146) );
  NAND2_X1 U4019 ( .A1(n3159), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3145)
         );
  NAND2_X1 U4020 ( .A1(n3395), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3144) );
  NAND2_X1 U4021 ( .A1(n2954), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3143)
         );
  NAND2_X1 U4022 ( .A1(n3316), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U4023 ( .A1(n3698), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4024 ( .A1(n3469), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3148) );
  NAND2_X1 U4025 ( .A1(n3224), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3147)
         );
  NAND2_X1 U4027 ( .A1(n3723), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U4028 ( .A1(n3969), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3157)
         );
  NAND2_X1 U4029 ( .A1(n2955), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3156)
         );
  NAND2_X1 U4030 ( .A1(n3464), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3155) );
  NAND2_X1 U4031 ( .A1(n3394), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U4032 ( .A1(n3159), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3162)
         );
  NAND2_X1 U4033 ( .A1(n3395), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U4034 ( .A1(n3530), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3160) );
  NAND2_X1 U4035 ( .A1(n3316), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3168) );
  NAND2_X1 U4036 ( .A1(n3314), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3167) );
  NAND2_X1 U4037 ( .A1(n3239), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U4038 ( .A1(n3698), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U4039 ( .A1(n3367), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3172)
         );
  NAND2_X1 U4040 ( .A1(n3469), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U4041 ( .A1(n3224), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3170)
         );
  NAND2_X1 U4042 ( .A1(n3400), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3169)
         );
  XOR2_X1 U4043 ( .A(n3178), .B(n3177), .Z(n3251) );
  OAI21_X1 U4044 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5169), .A(n3179), 
        .ZN(n3180) );
  NOR2_X1 U4045 ( .A1(n3556), .A2(n3180), .ZN(n3183) );
  INV_X2 U4046 ( .A(n4497), .ZN(n4143) );
  NAND2_X1 U4047 ( .A1(n4143), .A2(n4491), .ZN(n4139) );
  INV_X1 U4048 ( .A(n4139), .ZN(n3181) );
  OAI21_X1 U4049 ( .B1(n3181), .B2(n3180), .A(n3184), .ZN(n3182) );
  OAI21_X1 U4050 ( .B1(n4149), .B2(n4491), .A(n3276), .ZN(n3196) );
  NAND2_X1 U4051 ( .A1(n3182), .A2(n3196), .ZN(n3187) );
  OAI211_X1 U4052 ( .C1(n3188), .C2(n3251), .A(n3183), .B(n3187), .ZN(n3186)
         );
  NAND2_X1 U4053 ( .A1(n3337), .A2(n4400), .ZN(n3211) );
  NAND3_X1 U4054 ( .A1(n3188), .A2(STATE2_REG_0__SCAN_IN), .A3(n3251), .ZN(
        n3185) );
  NAND3_X1 U4055 ( .A1(n3186), .A2(n3211), .A3(n3185), .ZN(n3192) );
  INV_X1 U4056 ( .A(n3187), .ZN(n3190) );
  INV_X1 U4057 ( .A(n3188), .ZN(n3189) );
  NAND3_X1 U4058 ( .A1(n3190), .A2(n3251), .A3(n3189), .ZN(n3191) );
  NAND2_X1 U4059 ( .A1(n3192), .A2(n3191), .ZN(n3202) );
  INV_X1 U4060 ( .A(n3193), .ZN(n3194) );
  XNOR2_X1 U4061 ( .A(n3195), .B(n3194), .ZN(n3252) );
  INV_X1 U4062 ( .A(n3252), .ZN(n3198) );
  AOI211_X1 U4063 ( .C1(n3202), .C2(n3196), .A(n3556), .B(n3198), .ZN(n3204)
         );
  INV_X1 U4064 ( .A(n3196), .ZN(n3197) );
  AOI21_X1 U4065 ( .B1(n3337), .B2(n3198), .A(n3197), .ZN(n3201) );
  XOR2_X1 U4066 ( .A(n3200), .B(n3199), .Z(n3253) );
  OAI22_X1 U4067 ( .A1(n3202), .A2(n3201), .B1(n3253), .B2(n4410), .ZN(n3203)
         );
  OAI22_X1 U4068 ( .A1(n3204), .A2(n3203), .B1(n3337), .B2(n3253), .ZN(n3208)
         );
  OR2_X1 U4069 ( .A1(n3206), .A2(n3205), .ZN(n3256) );
  NOR2_X1 U4070 ( .A1(n3337), .A2(n3256), .ZN(n3207) );
  OAI22_X1 U4071 ( .A1(n3208), .A2(n3207), .B1(n3211), .B2(n3256), .ZN(n3209)
         );
  AND2_X1 U4072 ( .A1(n6403), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4072) );
  AND2_X1 U4073 ( .A1(n4072), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6399) );
  AOI22_X1 U4074 ( .A1(n3723), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3217) );
  AOI22_X1 U4075 ( .A1(n3159), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3216) );
  AOI22_X1 U4076 ( .A1(n3314), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3239), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3215) );
  AOI22_X1 U4077 ( .A1(n3469), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3214) );
  NAND4_X1 U4078 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), .ZN(n3223)
         );
  AOI22_X1 U4079 ( .A1(n3316), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3221) );
  AOI22_X1 U4080 ( .A1(n3464), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U4081 ( .A1(n2955), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3219) );
  AOI22_X1 U4082 ( .A1(n3969), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3218) );
  NAND4_X1 U4083 ( .A1(n3221), .A2(n3220), .A3(n3219), .A4(n3218), .ZN(n3222)
         );
  OR2_X2 U4084 ( .A1(n3223), .A2(n3222), .ZN(n4503) );
  AND2_X2 U4085 ( .A1(n4143), .A2(n4503), .ZN(n3233) );
  AOI22_X1 U4086 ( .A1(n3159), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3314), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4087 ( .A1(n3464), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3723), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3227) );
  AOI22_X1 U4088 ( .A1(n2954), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3226) );
  AOI22_X1 U4089 ( .A1(n3394), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3225) );
  AOI22_X1 U4090 ( .A1(n3367), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3232) );
  AOI22_X1 U4091 ( .A1(n3239), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3231) );
  AOI22_X1 U4092 ( .A1(n3316), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3230) );
  AOI22_X1 U4093 ( .A1(n3969), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3229) );
  NAND2_X2 U4094 ( .A1(n4507), .A2(n4327), .ZN(n4071) );
  NAND2_X2 U4095 ( .A1(n3233), .A2(n4071), .ZN(n3280) );
  INV_X1 U4096 ( .A(n3280), .ZN(n3247) );
  AOI22_X1 U4097 ( .A1(n3316), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3238) );
  INV_X1 U4098 ( .A(n3723), .ZN(n3234) );
  AOI22_X1 U4099 ( .A1(n3723), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4100 ( .A1(n3969), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U4101 ( .A1(n3159), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3235) );
  NAND4_X1 U4102 ( .A1(n3238), .A2(n3237), .A3(n3236), .A4(n3235), .ZN(n3245)
         );
  AOI22_X1 U4103 ( .A1(n3464), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4104 ( .A1(n3314), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3239), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3242) );
  AOI22_X1 U4105 ( .A1(n2954), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4106 ( .A1(n3469), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3400), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3240) );
  NAND4_X1 U4107 ( .A1(n3243), .A2(n3242), .A3(n3241), .A4(n3240), .ZN(n3244)
         );
  OR2_X2 U4108 ( .A1(n3245), .A2(n3244), .ZN(n4466) );
  INV_X2 U4109 ( .A(n4466), .ZN(n4134) );
  NAND2_X1 U4110 ( .A1(n4134), .A2(n4485), .ZN(n4023) );
  AND2_X2 U4111 ( .A1(n3247), .A2(n3246), .ZN(n4141) );
  NAND2_X1 U4112 ( .A1(n4141), .A2(n4592), .ZN(n6346) );
  NAND2_X1 U4113 ( .A1(n4149), .A2(n4466), .ZN(n3248) );
  NOR2_X1 U4114 ( .A1(n3280), .A2(n3248), .ZN(n3250) );
  NAND2_X1 U4115 ( .A1(n4324), .A2(n4485), .ZN(n3302) );
  AND2_X1 U4116 ( .A1(n3302), .A2(n3300), .ZN(n3350) );
  NAND2_X1 U4117 ( .A1(n3250), .A2(n3350), .ZN(n6351) );
  NAND3_X1 U4118 ( .A1(n3253), .A2(n3252), .A3(n3251), .ZN(n3254) );
  NAND2_X1 U4119 ( .A1(n3255), .A2(n3254), .ZN(n3257) );
  AND2_X1 U4120 ( .A1(n3257), .A2(n3256), .ZN(n6349) );
  INV_X1 U4121 ( .A(n6399), .ZN(n6406) );
  OR3_X1 U4122 ( .A1(n6351), .A2(n6349), .A3(n6406), .ZN(n5630) );
  INV_X1 U4123 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5265) );
  NOR2_X1 U4124 ( .A1(n6523), .A2(n5265), .ZN(n3261) );
  NOR2_X1 U4125 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6538) );
  NOR2_X1 U4126 ( .A1(n3049), .A2(n6538), .ZN(n3258) );
  AND2_X2 U4127 ( .A1(n3276), .A2(n4592), .ZN(n4415) );
  NAND2_X1 U4128 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6414) );
  OAI21_X1 U4129 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6414), .ZN(n3275) );
  OR2_X1 U4130 ( .A1(n3275), .A2(STATE_REG_0__SCAN_IN), .ZN(n6420) );
  INV_X1 U4131 ( .A(n6420), .ZN(n5797) );
  NAND2_X1 U4132 ( .A1(n5797), .A2(n6538), .ZN(n6389) );
  AND2_X1 U4133 ( .A1(n4415), .A2(n6389), .ZN(n4594) );
  NOR2_X1 U4134 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6526) );
  INV_X1 U4135 ( .A(n6526), .ZN(n6410) );
  NOR3_X1 U4136 ( .A1(n6402), .A2(n6490), .A3(n6410), .ZN(n6397) );
  NAND2_X1 U4137 ( .A1(n6403), .A2(n6490), .ZN(n6504) );
  NOR2_X1 U4138 ( .A1(n4439), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5516) );
  INV_X1 U4139 ( .A(n5516), .ZN(n4850) );
  INV_X1 U4140 ( .A(n4850), .ZN(n6099) );
  AND2_X1 U4141 ( .A1(n6402), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4438) );
  NOR2_X1 U4142 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3914) );
  AND2_X1 U4143 ( .A1(n4438), .A2(n4005), .ZN(n6409) );
  OR2_X1 U4144 ( .A1(n6099), .A2(n6409), .ZN(n3259) );
  NOR2_X1 U4145 ( .A1(n6397), .A2(n3259), .ZN(n3260) );
  AOI22_X1 U4146 ( .A1(n3261), .A2(n4594), .B1(PHYADDRPOINTER_REG_31__SCAN_IN), 
        .B2(n5901), .ZN(n3268) );
  NAND2_X1 U4147 ( .A1(n3276), .A2(n6420), .ZN(n4131) );
  AND3_X1 U4148 ( .A1(n4131), .A2(n6538), .A3(n4592), .ZN(n3262) );
  INV_X1 U4149 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U4150 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5672) );
  OR2_X1 U4151 ( .A1(n6569), .A2(n5672), .ZN(n4016) );
  NAND3_X1 U4152 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n4015) );
  INV_X1 U4153 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6451) );
  INV_X1 U4154 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6447) );
  INV_X1 U4155 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6445) );
  INV_X1 U4156 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6441) );
  INV_X1 U4157 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6438) );
  INV_X1 U4158 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6434) );
  NAND3_X1 U4159 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5917) );
  NOR2_X1 U4160 ( .A1(n6434), .A2(n5917), .ZN(n5899) );
  NAND2_X1 U4161 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5899), .ZN(n4590) );
  NOR2_X1 U4162 ( .A1(n6438), .A2(n4590), .ZN(n5890) );
  NAND2_X1 U4163 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5890), .ZN(n4609) );
  NOR2_X1 U4164 ( .A1(n6441), .A2(n4609), .ZN(n4611) );
  NAND2_X1 U4165 ( .A1(REIP_REG_9__SCAN_IN), .A2(n4611), .ZN(n5866) );
  NOR2_X1 U4166 ( .A1(n6445), .A2(n5866), .ZN(n4976) );
  NAND2_X1 U4167 ( .A1(REIP_REG_11__SCAN_IN), .A2(n4976), .ZN(n5846) );
  NOR2_X1 U4168 ( .A1(n6447), .A2(n5846), .ZN(n5849) );
  NAND2_X1 U4169 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5849), .ZN(n4014) );
  INV_X1 U4170 ( .A(n5321), .ZN(n5913) );
  NOR2_X1 U4171 ( .A1(n4015), .A2(n4970), .ZN(n5242) );
  NAND4_X1 U4172 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5242), .ZN(n5668) );
  NOR2_X1 U4173 ( .A1(n4016), .A2(n5668), .ZN(n5224) );
  INV_X1 U4174 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6464) );
  INV_X1 U4175 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6468) );
  INV_X1 U4176 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6466) );
  NOR3_X1 U4177 ( .A1(n6464), .A2(n6468), .A3(n6466), .ZN(n4017) );
  NAND2_X1 U4178 ( .A1(n5224), .A2(n4017), .ZN(n3263) );
  NAND2_X1 U4179 ( .A1(n5918), .A2(n5321), .ZN(n5941) );
  AND2_X1 U4180 ( .A1(n3263), .A2(n5941), .ZN(n5655) );
  INV_X1 U4181 ( .A(n5918), .ZN(n5900) );
  NAND2_X1 U4182 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n3264) );
  AND2_X1 U4183 ( .A1(n5900), .A2(n3264), .ZN(n3265) );
  OR2_X1 U4184 ( .A1(n5655), .A2(n3265), .ZN(n5633) );
  INV_X1 U4185 ( .A(n5633), .ZN(n3266) );
  OAI211_X1 U4186 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5918), .A(n3266), .B(
        REIP_REG_30__SCAN_IN), .ZN(n5373) );
  NAND3_X1 U4187 ( .A1(n5373), .A2(REIP_REG_31__SCAN_IN), .A3(n5941), .ZN(
        n3267) );
  OAI211_X1 U4188 ( .C1(n5534), .C2(n5933), .A(n3268), .B(n3267), .ZN(n3269)
         );
  INV_X1 U4189 ( .A(n3269), .ZN(n4020) );
  INV_X2 U4190 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6393) );
  OR2_X1 U4191 ( .A1(n4503), .A2(n6393), .ZN(n3644) );
  INV_X2 U4192 ( .A(n3644), .ZN(n3802) );
  NAND2_X1 U4193 ( .A1(n6393), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4194 ( .A1(n3802), .A2(EAX_REG_31__SCAN_IN), .B1(n3424), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4010) );
  NAND2_X1 U4195 ( .A1(n3280), .A2(n4415), .ZN(n3278) );
  AND2_X1 U4196 ( .A1(n4324), .A2(n4592), .ZN(n3274) );
  NAND2_X1 U4197 ( .A1(n3274), .A2(n3280), .ZN(n4031) );
  NAND2_X1 U4198 ( .A1(n3276), .A2(n3275), .ZN(n3345) );
  NAND2_X1 U4199 ( .A1(n3345), .A2(n4327), .ZN(n3277) );
  NAND4_X1 U4200 ( .A1(n3298), .A2(n3278), .A3(n4031), .A4(n3277), .ZN(n3279)
         );
  NOR2_X1 U4201 ( .A1(n4041), .A2(n3279), .ZN(n3288) );
  NOR2_X1 U4202 ( .A1(n3280), .A2(n4036), .ZN(n3286) );
  NOR2_X1 U4203 ( .A1(n3300), .A2(n4143), .ZN(n3697) );
  INV_X1 U4204 ( .A(n3697), .ZN(n3283) );
  NOR2_X1 U4205 ( .A1(n5437), .A2(n4071), .ZN(n3281) );
  NOR2_X1 U4206 ( .A1(n3281), .A2(n4466), .ZN(n3282) );
  NAND2_X1 U4207 ( .A1(n3283), .A2(n3282), .ZN(n3285) );
  AND2_X1 U4208 ( .A1(n3302), .A2(n3276), .ZN(n3284) );
  OAI211_X1 U4209 ( .C1(n3286), .C2(n4134), .A(n3285), .B(n3284), .ZN(n3287)
         );
  NAND2_X1 U4210 ( .A1(n3287), .A2(n4149), .ZN(n3292) );
  NAND2_X1 U4211 ( .A1(n3288), .A2(n3292), .ZN(n3289) );
  INV_X1 U4212 ( .A(n4072), .ZN(n3392) );
  MUX2_X1 U4213 ( .A(n3392), .B(n6520), .S(n5169), .Z(n3290) );
  INV_X1 U4214 ( .A(n3290), .ZN(n3291) );
  OAI21_X2 U4215 ( .B1(n3387), .B2(n3444), .A(n3291), .ZN(n3360) );
  INV_X1 U4216 ( .A(n3292), .ZN(n3294) );
  OR2_X1 U4217 ( .A1(n4139), .A2(n3276), .ZN(n3293) );
  NAND2_X1 U4218 ( .A1(n4324), .A2(n4497), .ZN(n3295) );
  NAND2_X1 U4219 ( .A1(n3295), .A2(n4485), .ZN(n3296) );
  OAI21_X1 U4220 ( .B1(n4024), .B2(n3296), .A(n4474), .ZN(n3305) );
  NOR2_X1 U4221 ( .A1(n4485), .A2(n4592), .ZN(n3297) );
  NAND2_X1 U4222 ( .A1(n3297), .A2(n4134), .ZN(n4035) );
  OR2_X1 U4223 ( .A1(n6504), .A2(n6402), .ZN(n6405) );
  AOI21_X1 U4224 ( .B1(n4466), .B2(n4592), .A(n6405), .ZN(n3299) );
  OAI211_X1 U4225 ( .C1(n4035), .C2(n3300), .A(n3299), .B(n3298), .ZN(n3301)
         );
  INV_X1 U4226 ( .A(n3301), .ZN(n3304) );
  OAI21_X1 U4227 ( .B1(n3280), .B2(n3302), .A(n4415), .ZN(n3303) );
  INV_X1 U4228 ( .A(n3359), .ZN(n3307) );
  XNOR2_X1 U4229 ( .A(n3360), .B(n3307), .ZN(n3440) );
  NAND2_X1 U4230 ( .A1(n3440), .A2(n6402), .ZN(n3435) );
  AOI22_X1 U4231 ( .A1(n3836), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3982), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4232 ( .A1(n3983), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3312) );
  BUF_X1 U4233 ( .A(n2955), .Z(n3309) );
  AOI22_X1 U4234 ( .A1(n3309), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4235 ( .A1(n2952), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3310) );
  NAND4_X1 U4236 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3322)
         );
  AOI22_X1 U4237 ( .A1(n3790), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3969), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4238 ( .A1(n2951), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4239 ( .A1(n3970), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4240 ( .A1(n3224), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3317) );
  NAND4_X1 U4241 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3321)
         );
  NOR2_X1 U4242 ( .A1(n3362), .A2(n4414), .ZN(n3375) );
  NAND2_X1 U4243 ( .A1(n4143), .A2(n4414), .ZN(n3338) );
  NOR2_X1 U4244 ( .A1(n3338), .A2(n6402), .ZN(n4409) );
  INV_X1 U4245 ( .A(n3234), .ZN(n3901) );
  AOI22_X1 U4246 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n3790), .B1(n3836), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4247 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n3315), .B1(n3308), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4248 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3309), .B1(n3530), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4249 ( .A1(n3970), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3324) );
  NAND4_X1 U4250 ( .A1(n3327), .A2(n3326), .A3(n3325), .A4(n3324), .ZN(n3334)
         );
  AOI22_X1 U4251 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n2951), .B1(n3969), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4252 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3983), .B1(n3982), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4253 ( .A1(n3984), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4254 ( .A1(n2952), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3329) );
  NAND4_X1 U4255 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(n3333)
         );
  INV_X1 U4256 ( .A(n4197), .ZN(n3335) );
  MUX2_X1 U4257 ( .A(n3375), .B(n4409), .S(n3335), .Z(n3336) );
  INV_X1 U4258 ( .A(n3336), .ZN(n3436) );
  NAND2_X1 U4259 ( .A1(n3435), .A2(n3436), .ZN(n3341) );
  INV_X1 U4260 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3340) );
  AOI21_X1 U4261 ( .B1(n4149), .B2(n4197), .A(n6402), .ZN(n3339) );
  OAI211_X1 U4262 ( .C1(n3553), .C2(n3340), .A(n3339), .B(n3338), .ZN(n3438)
         );
  XNOR2_X1 U4263 ( .A(n5169), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6173)
         );
  NAND2_X1 U4264 ( .A1(n6520), .A2(n6173), .ZN(n3344) );
  NAND2_X1 U4265 ( .A1(n3392), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4266 ( .A1(n3344), .A2(n3343), .ZN(n3355) );
  INV_X1 U4267 ( .A(n3355), .ZN(n3354) );
  INV_X1 U4268 ( .A(n3345), .ZN(n3352) );
  INV_X1 U4269 ( .A(n4035), .ZN(n3347) );
  NOR2_X1 U4270 ( .A1(n4491), .A2(n4474), .ZN(n3346) );
  AND2_X1 U4271 ( .A1(n4503), .A2(n4507), .ZN(n4326) );
  NAND2_X1 U4272 ( .A1(n4056), .A2(n4326), .ZN(n4155) );
  NAND2_X1 U4273 ( .A1(n3348), .A2(n4466), .ZN(n3349) );
  NOR2_X1 U4274 ( .A1(n3280), .A2(n3349), .ZN(n3351) );
  NAND2_X1 U4275 ( .A1(n3353), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3357) );
  OAI211_X1 U4276 ( .C1(n3387), .C2(n4258), .A(n3354), .B(n3357), .ZN(n3385)
         );
  NOR2_X1 U4277 ( .A1(n3355), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3356)
         );
  INV_X1 U4278 ( .A(n3358), .ZN(n3383) );
  NAND2_X1 U4279 ( .A1(n3385), .A2(n3383), .ZN(n3361) );
  INV_X1 U4280 ( .A(n3362), .ZN(n4074) );
  BUF_X1 U4281 ( .A(n3969), .Z(n3989) );
  AOI22_X1 U4282 ( .A1(n3989), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n2951), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4283 ( .A1(n3983), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4284 ( .A1(n3315), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4285 ( .A1(n3970), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3363) );
  NAND4_X1 U4286 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3373)
         );
  AOI22_X1 U4287 ( .A1(n3901), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4288 ( .A1(n3982), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4289 ( .A1(n3984), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4290 ( .A1(n3790), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3368) );
  NAND4_X1 U4291 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3372)
         );
  NAND2_X1 U4292 ( .A1(n4074), .A2(n4196), .ZN(n3374) );
  OAI21_X2 U4293 ( .B1(n4054), .B2(STATE2_REG_0__SCAN_IN), .A(n3374), .ZN(
        n3428) );
  INV_X1 U4294 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3379) );
  INV_X1 U4295 ( .A(n3375), .ZN(n3378) );
  INV_X1 U4296 ( .A(n4196), .ZN(n3376) );
  OR2_X1 U4297 ( .A1(n3410), .A2(n3376), .ZN(n3377) );
  OAI211_X1 U4298 ( .C1(n3553), .C2(n3379), .A(n3378), .B(n3377), .ZN(n3427)
         );
  NAND2_X1 U4299 ( .A1(n3428), .A2(n3427), .ZN(n3420) );
  NAND2_X1 U4300 ( .A1(n3417), .A2(n3420), .ZN(n3382) );
  INV_X1 U4301 ( .A(n3428), .ZN(n3381) );
  INV_X1 U4302 ( .A(n3427), .ZN(n3380) );
  NAND2_X1 U4303 ( .A1(n3381), .A2(n3380), .ZN(n3418) );
  NAND2_X1 U4304 ( .A1(n3384), .A2(n3383), .ZN(n3386) );
  NAND2_X1 U4305 ( .A1(n3386), .A2(n3385), .ZN(n3454) );
  AND2_X1 U4306 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3389) );
  NAND2_X1 U4307 ( .A1(n3389), .A2(n5168), .ZN(n6242) );
  INV_X1 U4308 ( .A(n3389), .ZN(n3390) );
  NAND2_X1 U4309 ( .A1(n3390), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3391) );
  NAND2_X1 U4310 ( .A1(n6242), .A2(n3391), .ZN(n4468) );
  AOI22_X1 U4311 ( .A1(n6520), .A2(n4468), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3392), .ZN(n3393) );
  XNOR2_X1 U4312 ( .A(n3454), .B(n3455), .ZN(n4255) );
  NAND2_X1 U4313 ( .A1(n4255), .A2(n6402), .ZN(n3408) );
  AOI22_X1 U4314 ( .A1(n2951), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4315 ( .A1(n3315), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4316 ( .A1(n3983), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4317 ( .A1(n3982), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3396) );
  NAND4_X1 U4318 ( .A1(n3399), .A2(n3398), .A3(n3397), .A4(n3396), .ZN(n3406)
         );
  AOI22_X1 U4319 ( .A1(n3969), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4320 ( .A1(n3970), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4321 ( .A1(n3328), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4322 ( .A1(n3790), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3401) );
  NAND4_X1 U4323 ( .A1(n3404), .A2(n3403), .A3(n3402), .A4(n3401), .ZN(n3405)
         );
  NAND2_X1 U4324 ( .A1(n4074), .A2(n3409), .ZN(n3407) );
  NAND2_X1 U4325 ( .A1(n3408), .A2(n3407), .ZN(n3414) );
  INV_X1 U4326 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3411) );
  INV_X1 U4327 ( .A(n3409), .ZN(n4206) );
  OAI22_X1 U4328 ( .A1(n3553), .A2(n3411), .B1(n3410), .B2(n4206), .ZN(n3412)
         );
  INV_X1 U4329 ( .A(n3412), .ZN(n3413) );
  XNOR2_X1 U4330 ( .A(n3414), .B(n3413), .ZN(n3416) );
  NAND2_X1 U4331 ( .A1(n3415), .A2(n3416), .ZN(n3478) );
  INV_X1 U4332 ( .A(n3416), .ZN(n3421) );
  INV_X1 U4333 ( .A(n3417), .ZN(n3429) );
  NAND2_X1 U4334 ( .A1(n3418), .A2(n3429), .ZN(n3419) );
  NAND3_X1 U4335 ( .A1(n3421), .A2(n3420), .A3(n3419), .ZN(n3422) );
  INV_X1 U4336 ( .A(n4298), .ZN(n3426) );
  NAND2_X1 U4337 ( .A1(n3423), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3680) );
  XNOR2_X1 U4338 ( .A(n3428), .B(n3427), .ZN(n3430) );
  XNOR2_X1 U4339 ( .A(n3430), .B(n3429), .ZN(n4299) );
  NAND2_X1 U4340 ( .A1(n4299), .A2(n3425), .ZN(n3434) );
  AOI22_X1 U4341 ( .A1(n3802), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6393), .ZN(n3432) );
  AND2_X1 U4342 ( .A1(n4326), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3441) );
  NAND2_X1 U4343 ( .A1(n3441), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3431) );
  AND2_X1 U4344 ( .A1(n3432), .A2(n3431), .ZN(n3433) );
  NAND2_X1 U4345 ( .A1(n3434), .A2(n3433), .ZN(n4079) );
  NAND2_X1 U4346 ( .A1(n3435), .A2(n3438), .ZN(n3437) );
  MUX2_X2 U4347 ( .A(n3438), .B(n3437), .S(n3436), .Z(n5009) );
  NAND2_X1 U4348 ( .A1(n5009), .A2(n4036), .ZN(n3439) );
  NAND2_X1 U4349 ( .A1(n3439), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4120) );
  INV_X1 U4350 ( .A(n3441), .ZN(n3501) );
  NAND2_X1 U4351 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n6393), .ZN(n3443)
         );
  NAND2_X1 U4352 ( .A1(n3802), .A2(EAX_REG_0__SCAN_IN), .ZN(n3442) );
  OAI211_X1 U4353 ( .C1(n3501), .C2(n3444), .A(n3443), .B(n3442), .ZN(n3445)
         );
  AOI21_X1 U4354 ( .B1(n6365), .B2(n3425), .A(n3445), .ZN(n4119) );
  OR2_X1 U4355 ( .A1(n4120), .A2(n4119), .ZN(n4122) );
  NAND2_X1 U4356 ( .A1(n4119), .A2(n4005), .ZN(n3446) );
  NAND2_X1 U4357 ( .A1(n4122), .A2(n3446), .ZN(n4080) );
  NAND2_X1 U4358 ( .A1(n4079), .A2(n4080), .ZN(n4082) );
  NAND2_X1 U4359 ( .A1(n3449), .A2(n4082), .ZN(n4313) );
  OAI21_X1 U4360 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3482), .ZN(n6039) );
  AOI22_X1 U4361 ( .A1(n4005), .A2(n6039), .B1(n3424), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3448) );
  NAND2_X1 U4362 ( .A1(n3802), .A2(EAX_REG_2__SCAN_IN), .ZN(n3447) );
  OAI211_X1 U4363 ( .C1(n3501), .C2(n5263), .A(n3448), .B(n3447), .ZN(n4312)
         );
  NAND2_X1 U4364 ( .A1(n4313), .A2(n4312), .ZN(n3453) );
  INV_X1 U4365 ( .A(n4082), .ZN(n3451) );
  INV_X1 U4366 ( .A(n3449), .ZN(n3450) );
  NAND2_X1 U4367 ( .A1(n3451), .A2(n3450), .ZN(n3452) );
  NAND2_X1 U4368 ( .A1(n3453), .A2(n3452), .ZN(n4315) );
  INV_X1 U4369 ( .A(n3454), .ZN(n3456) );
  NAND2_X1 U4370 ( .A1(n3456), .A2(n3455), .ZN(n4290) );
  INV_X1 U4371 ( .A(n3457), .ZN(n3458) );
  NAND2_X1 U4372 ( .A1(n3458), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3463) );
  NAND3_X1 U4373 ( .A1(n6382), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6213) );
  INV_X1 U4374 ( .A(n6213), .ZN(n3459) );
  NAND2_X1 U4375 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3459), .ZN(n6204) );
  NAND2_X1 U4376 ( .A1(n6382), .A2(n6204), .ZN(n3460) );
  NOR3_X1 U4377 ( .A1(n6382), .A2(n5168), .A3(n6374), .ZN(n6294) );
  NAND2_X1 U4378 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6294), .ZN(n6280) );
  NAND2_X1 U4379 ( .A1(n3460), .A2(n6280), .ZN(n4762) );
  OAI22_X1 U4380 ( .A1(n4439), .A2(n4762), .B1(n4072), .B2(n6382), .ZN(n3461)
         );
  INV_X1 U4381 ( .A(n3461), .ZN(n3462) );
  XNOR2_X2 U4382 ( .A(n4290), .B(n6207), .ZN(n5167) );
  AOI22_X1 U4383 ( .A1(n2951), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4384 ( .A1(n3315), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4385 ( .A1(n3983), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4386 ( .A1(n3982), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3465) );
  NAND4_X1 U4387 ( .A1(n3468), .A2(n3467), .A3(n3466), .A4(n3465), .ZN(n3475)
         );
  AOI22_X1 U4388 ( .A1(n3989), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4389 ( .A1(n3970), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4390 ( .A1(n3328), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4391 ( .A1(n3790), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3470) );
  NAND4_X1 U4392 ( .A1(n3473), .A2(n3472), .A3(n3471), .A4(n3470), .ZN(n3474)
         );
  NOR2_X1 U4393 ( .A1(n3475), .A2(n3474), .ZN(n4217) );
  INV_X1 U4394 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3476) );
  OAI22_X1 U4395 ( .A1(n3556), .A2(n4217), .B1(n3476), .B2(n3553), .ZN(n3477)
         );
  NAND2_X1 U4396 ( .A1(n3478), .A2(n4303), .ZN(n3481) );
  INV_X1 U4397 ( .A(n3478), .ZN(n3480) );
  INV_X1 U4398 ( .A(n4303), .ZN(n3479) );
  NAND2_X1 U4399 ( .A1(n3480), .A2(n3479), .ZN(n3510) );
  INV_X1 U4400 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4268) );
  OAI21_X1 U4401 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3483), .A(n3502), 
        .ZN(n5934) );
  AOI22_X1 U4402 ( .A1(n4005), .A2(n5934), .B1(n3424), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3485) );
  NAND2_X1 U4403 ( .A1(n3802), .A2(EAX_REG_3__SCAN_IN), .ZN(n3484) );
  OAI211_X1 U4404 ( .C1(n3501), .C2(n4268), .A(n3485), .B(n3484), .ZN(n3486)
         );
  INV_X1 U4405 ( .A(n3486), .ZN(n3487) );
  OAI21_X1 U4406 ( .B1(n4301), .B2(n3680), .A(n3487), .ZN(n4188) );
  INV_X1 U4407 ( .A(n4187), .ZN(n3507) );
  AOI22_X1 U4408 ( .A1(n3315), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4409 ( .A1(n3983), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U4410 ( .A1(n3989), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4411 ( .A1(n2952), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3488) );
  NAND4_X1 U4412 ( .A1(n3491), .A2(n3490), .A3(n3489), .A4(n3488), .ZN(n3497)
         );
  AOI22_X1 U4413 ( .A1(n3790), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4414 ( .A1(n2951), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3982), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4415 ( .A1(n3970), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4416 ( .A1(n3224), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3492) );
  NAND4_X1 U4417 ( .A1(n3495), .A2(n3494), .A3(n3493), .A4(n3492), .ZN(n3496)
         );
  OR2_X1 U4418 ( .A1(n3497), .A2(n3496), .ZN(n4227) );
  INV_X1 U4419 ( .A(n4227), .ZN(n4235) );
  INV_X1 U4420 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3498) );
  OAI22_X1 U4421 ( .A1(n3556), .A2(n4235), .B1(n3498), .B2(n3553), .ZN(n3508)
         );
  XNOR2_X1 U4422 ( .A(n3510), .B(n3508), .ZN(n4226) );
  INV_X1 U4423 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6621) );
  OAI21_X1 U4424 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6621), .A(n6393), 
        .ZN(n3500) );
  NAND2_X1 U4425 ( .A1(n3802), .A2(EAX_REG_4__SCAN_IN), .ZN(n3499) );
  OAI211_X1 U4426 ( .C1(n3501), .C2(n4293), .A(n3500), .B(n3499), .ZN(n3504)
         );
  AOI21_X1 U4427 ( .B1(n3502), .B2(n5914), .A(n3525), .ZN(n4444) );
  NAND2_X1 U4428 ( .A1(n4444), .A2(n3914), .ZN(n3503) );
  AND2_X1 U4429 ( .A1(n3504), .A2(n3503), .ZN(n3505) );
  AOI21_X1 U4430 ( .B1(n4226), .B2(n3425), .A(n3505), .ZN(n4331) );
  INV_X1 U4431 ( .A(n3508), .ZN(n3509) );
  NOR2_X1 U4432 ( .A1(n3510), .A2(n3509), .ZN(n3523) );
  AOI22_X1 U4433 ( .A1(n2951), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4434 ( .A1(n3315), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4435 ( .A1(n3983), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4436 ( .A1(n3982), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3511) );
  NAND4_X1 U4437 ( .A1(n3514), .A2(n3513), .A3(n3512), .A4(n3511), .ZN(n3520)
         );
  AOI22_X1 U4438 ( .A1(n3989), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4439 ( .A1(n3970), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3517) );
  INV_X1 U4440 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6571) );
  AOI22_X1 U4441 ( .A1(n3328), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4442 ( .A1(n3790), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3515) );
  NAND4_X1 U4443 ( .A1(n3518), .A2(n3517), .A3(n3516), .A4(n3515), .ZN(n3519)
         );
  NOR2_X1 U4444 ( .A1(n3520), .A2(n3519), .ZN(n4239) );
  INV_X1 U4445 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3521) );
  OAI22_X1 U4446 ( .A1(n3556), .A2(n4239), .B1(n3521), .B2(n3553), .ZN(n3522)
         );
  NAND2_X1 U4447 ( .A1(n3523), .A2(n3522), .ZN(n3551) );
  OR2_X1 U4448 ( .A1(n3523), .A2(n3522), .ZN(n3524) );
  AND2_X1 U4449 ( .A1(n3551), .A2(n3524), .ZN(n4234) );
  INV_X1 U4450 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3528) );
  OAI21_X1 U4451 ( .B1(n3525), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3559), 
        .ZN(n5905) );
  NAND2_X1 U4452 ( .A1(n5905), .A2(n4005), .ZN(n3527) );
  NAND2_X1 U4453 ( .A1(n3424), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3526)
         );
  OAI211_X1 U4454 ( .C1(n3644), .C2(n3528), .A(n3527), .B(n3526), .ZN(n3529)
         );
  AOI22_X1 U4455 ( .A1(n3989), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n2951), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4456 ( .A1(n3983), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4457 ( .A1(n3982), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4458 ( .A1(n3984), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3531) );
  NAND4_X1 U4459 ( .A1(n3534), .A2(n3533), .A3(n3532), .A4(n3531), .ZN(n3540)
         );
  AOI22_X1 U4460 ( .A1(n3309), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4461 ( .A1(n3901), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4462 ( .A1(n3970), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4463 ( .A1(n3790), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3535) );
  NAND4_X1 U4464 ( .A1(n3538), .A2(n3537), .A3(n3536), .A4(n3535), .ZN(n3539)
         );
  OR2_X1 U4465 ( .A1(n3540), .A2(n3539), .ZN(n4403) );
  INV_X1 U4466 ( .A(n4403), .ZN(n3542) );
  INV_X1 U4467 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3541) );
  OAI22_X1 U4468 ( .A1(n3556), .A2(n3542), .B1(n3553), .B2(n3541), .ZN(n3543)
         );
  INV_X1 U4469 ( .A(n3543), .ZN(n3550) );
  NAND2_X1 U4470 ( .A1(n3551), .A2(n3550), .ZN(n4342) );
  NAND2_X1 U4471 ( .A1(n4342), .A2(n3425), .ZN(n3549) );
  INV_X1 U4472 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3545) );
  OAI21_X1 U4473 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6621), .A(n6393), 
        .ZN(n3544) );
  OAI21_X1 U4474 ( .B1(n3644), .B2(n3545), .A(n3544), .ZN(n3547) );
  XOR2_X1 U4475 ( .A(n3558), .B(n3559), .Z(n4599) );
  NAND2_X1 U4476 ( .A1(n4599), .A2(n3914), .ZN(n3546) );
  NAND2_X1 U4477 ( .A1(n3547), .A2(n3546), .ZN(n3548) );
  NAND2_X1 U4478 ( .A1(n3549), .A2(n3548), .ZN(n4366) );
  INV_X1 U4479 ( .A(n4414), .ZN(n3555) );
  INV_X1 U4480 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3554) );
  OAI22_X1 U4481 ( .A1(n3556), .A2(n3555), .B1(n3554), .B2(n3553), .ZN(n3557)
         );
  AOI22_X1 U4482 ( .A1(n3802), .A2(EAX_REG_7__SCAN_IN), .B1(n3424), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3561) );
  NAND2_X1 U4483 ( .A1(n3560), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3573)
         );
  OAI21_X1 U4484 ( .B1(n3560), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3573), 
        .ZN(n5892) );
  INV_X1 U4485 ( .A(n5892), .ZN(n4581) );
  INV_X1 U4486 ( .A(n3914), .ZN(n4003) );
  AOI22_X1 U4487 ( .A1(n3989), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4488 ( .A1(n3901), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3982), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4489 ( .A1(n3983), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3564) );
  BUF_X1 U4490 ( .A(n3224), .Z(n3795) );
  AOI22_X1 U4491 ( .A1(n3328), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4492 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3572)
         );
  AOI22_X1 U4493 ( .A1(n2951), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4494 ( .A1(n3315), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4495 ( .A1(n3970), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4496 ( .A1(n3790), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3567) );
  NAND4_X1 U4497 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3571)
         );
  NOR2_X1 U4498 ( .A1(n3572), .A2(n3571), .ZN(n3577) );
  INV_X1 U4499 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6625) );
  XOR2_X1 U4500 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3619), .Z(n5869) );
  INV_X1 U4501 ( .A(n5869), .ZN(n3574) );
  AOI22_X1 U4502 ( .A1(n3424), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n3914), 
        .B2(n3574), .ZN(n3576) );
  NAND2_X1 U4503 ( .A1(n3802), .A2(EAX_REG_10__SCAN_IN), .ZN(n3575) );
  OAI211_X1 U4504 ( .C1(n3680), .C2(n3577), .A(n3576), .B(n3575), .ZN(n4435)
         );
  AOI21_X1 U4505 ( .B1(n3578), .B2(n6625), .A(n3619), .ZN(n5883) );
  OR2_X1 U4506 ( .A1(n5883), .A2(n4003), .ZN(n3593) );
  AOI22_X1 U4507 ( .A1(n2951), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3982), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4508 ( .A1(n3901), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4509 ( .A1(n3984), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4510 ( .A1(n3790), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3579) );
  NAND4_X1 U4511 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n3588)
         );
  AOI22_X1 U4512 ( .A1(n3315), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4513 ( .A1(n3983), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4514 ( .A1(n3989), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4515 ( .A1(n3970), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3583) );
  NAND4_X1 U4516 ( .A1(n3586), .A2(n3585), .A3(n3584), .A4(n3583), .ZN(n3587)
         );
  OAI21_X1 U4517 ( .B1(n3588), .B2(n3587), .A(n3425), .ZN(n3591) );
  NAND2_X1 U4518 ( .A1(n3802), .A2(EAX_REG_9__SCAN_IN), .ZN(n3590) );
  NAND2_X1 U4519 ( .A1(n3424), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3589)
         );
  AND3_X1 U4520 ( .A1(n3591), .A2(n3590), .A3(n3589), .ZN(n3592) );
  AND2_X1 U4521 ( .A1(n3593), .A2(n3592), .ZN(n4725) );
  XOR2_X1 U4522 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3594), .Z(n4616) );
  INV_X1 U4523 ( .A(n4616), .ZN(n4620) );
  AOI22_X1 U4524 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3983), .B1(n3315), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4525 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n3309), .B1(n3945), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4526 ( .A1(n3970), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4527 ( .A1(n3901), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3595) );
  NAND4_X1 U4528 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3604)
         );
  AOI22_X1 U4529 ( .A1(n3989), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n2951), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4530 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3982), .B1(n3308), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4531 ( .A1(n3790), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4532 ( .A1(n3984), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3599) );
  NAND4_X1 U4533 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3603)
         );
  OAI21_X1 U4534 ( .B1(n3604), .B2(n3603), .A(n3425), .ZN(n3607) );
  NAND2_X1 U4535 ( .A1(n3802), .A2(EAX_REG_8__SCAN_IN), .ZN(n3606) );
  NAND2_X1 U4536 ( .A1(n3424), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3605)
         );
  NAND3_X1 U4537 ( .A1(n3607), .A2(n3606), .A3(n3605), .ZN(n3608) );
  AOI21_X1 U4538 ( .B1(n4620), .B2(n3914), .A(n3608), .ZN(n4604) );
  NOR2_X1 U4539 ( .A1(n4725), .A2(n4604), .ZN(n4432) );
  AND2_X1 U4540 ( .A1(n4435), .A2(n4432), .ZN(n4387) );
  AOI22_X1 U4541 ( .A1(n3989), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n2951), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4542 ( .A1(n3982), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4543 ( .A1(n3328), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4544 ( .A1(n2952), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3609) );
  NAND4_X1 U4545 ( .A1(n3612), .A2(n3611), .A3(n3610), .A4(n3609), .ZN(n3618)
         );
  AOI22_X1 U4546 ( .A1(n3790), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4547 ( .A1(n3983), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4548 ( .A1(n3309), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4549 ( .A1(n3970), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3613) );
  NAND4_X1 U4550 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(n3617)
         );
  OAI21_X1 U4551 ( .B1(n3618), .B2(n3617), .A(n3425), .ZN(n3623) );
  NAND2_X1 U4552 ( .A1(n3802), .A2(EAX_REG_11__SCAN_IN), .ZN(n3622) );
  NAND2_X1 U4553 ( .A1(n3619), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3625)
         );
  INV_X1 U4554 ( .A(n3625), .ZN(n3620) );
  XNOR2_X1 U4555 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3620), .ZN(n4999)
         );
  AOI22_X1 U4556 ( .A1(n4005), .A2(n4999), .B1(n3424), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3621) );
  NAND3_X1 U4557 ( .A1(n3623), .A2(n3622), .A3(n3621), .ZN(n4390) );
  AND2_X1 U4558 ( .A1(n4387), .A2(n4390), .ZN(n3661) );
  INV_X1 U4559 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3624) );
  XOR2_X1 U4560 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3643), .Z(n5101) );
  INV_X1 U4561 ( .A(n5101), .ZN(n5857) );
  INV_X1 U4562 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4575) );
  INV_X1 U4563 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5098) );
  OAI22_X1 U4564 ( .A1(n3644), .A2(n4575), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5098), .ZN(n3626) );
  NAND2_X1 U4565 ( .A1(n3626), .A2(n4003), .ZN(n3638) );
  AOI22_X1 U4566 ( .A1(n3989), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4567 ( .A1(n2951), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3982), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4568 ( .A1(n3309), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4569 ( .A1(n3790), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3627) );
  NAND4_X1 U4570 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n3636)
         );
  AOI22_X1 U4571 ( .A1(n3983), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4572 ( .A1(n3315), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4573 ( .A1(n3970), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4574 ( .A1(n3328), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3631) );
  NAND4_X1 U4575 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(n3635)
         );
  OAI21_X1 U4576 ( .B1(n3636), .B2(n3635), .A(n3425), .ZN(n3637) );
  NAND2_X1 U4577 ( .A1(n3638), .A2(n3637), .ZN(n3639) );
  AOI21_X1 U4578 ( .B1(n5857), .B2(n3914), .A(n3639), .ZN(n4567) );
  INV_X1 U4579 ( .A(n4567), .ZN(n3640) );
  AND2_X1 U4580 ( .A1(n3661), .A2(n3640), .ZN(n3641) );
  AND2_X1 U4581 ( .A1(n4516), .A2(n3641), .ZN(n3642) );
  INV_X1 U4582 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5085) );
  XNOR2_X1 U4583 ( .A(n3676), .B(n5085), .ZN(n5084) );
  NAND2_X1 U4584 ( .A1(n5084), .A2(n3914), .ZN(n3648) );
  NOR2_X1 U4585 ( .A1(n3645), .A2(n5085), .ZN(n3646) );
  AOI21_X1 U4586 ( .B1(n3802), .B2(EAX_REG_13__SCAN_IN), .A(n3646), .ZN(n3647)
         );
  NAND2_X1 U4587 ( .A1(n3648), .A2(n3647), .ZN(n3663) );
  AOI22_X1 U4588 ( .A1(n2951), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4589 ( .A1(n3315), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4590 ( .A1(n3983), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4591 ( .A1(n3982), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3650) );
  NAND4_X1 U4592 ( .A1(n3653), .A2(n3652), .A3(n3651), .A4(n3650), .ZN(n3659)
         );
  AOI22_X1 U4593 ( .A1(n3989), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4594 ( .A1(n3970), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4595 ( .A1(n3328), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4596 ( .A1(n3790), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3654) );
  NAND4_X1 U4597 ( .A1(n3657), .A2(n3656), .A3(n3655), .A4(n3654), .ZN(n3658)
         );
  OR2_X1 U4598 ( .A1(n3659), .A2(n3658), .ZN(n3660) );
  AND2_X1 U4599 ( .A1(n3425), .A2(n3660), .ZN(n4710) );
  NAND2_X1 U4600 ( .A1(n4709), .A2(n4710), .ZN(n3665) );
  AND2_X1 U4601 ( .A1(n3661), .A2(n4516), .ZN(n3662) );
  NOR2_X2 U4602 ( .A1(n4389), .A2(n4567), .ZN(n4566) );
  NAND2_X1 U4603 ( .A1(n4566), .A2(n3663), .ZN(n3664) );
  AOI22_X1 U4604 ( .A1(n3989), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4605 ( .A1(n3983), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4606 ( .A1(n3982), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4607 ( .A1(n3970), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3666) );
  NAND4_X1 U4608 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3675)
         );
  AOI22_X1 U4609 ( .A1(n2951), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4610 ( .A1(n3309), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4611 ( .A1(n3984), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4612 ( .A1(n3790), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3670) );
  NAND4_X1 U4613 ( .A1(n3673), .A2(n3672), .A3(n3671), .A4(n3670), .ZN(n3674)
         );
  NOR2_X1 U4614 ( .A1(n3675), .A2(n3674), .ZN(n3679) );
  XNOR2_X1 U4615 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3681), .ZN(n5071)
         );
  AOI22_X1 U4616 ( .A1(n4005), .A2(n5071), .B1(n3424), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3678) );
  NAND2_X1 U4617 ( .A1(n3802), .A2(EAX_REG_14__SCAN_IN), .ZN(n3677) );
  OAI211_X1 U4618 ( .C1(n3680), .C2(n3679), .A(n3678), .B(n3677), .ZN(n4802)
         );
  INV_X1 U4619 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3713) );
  XOR2_X1 U4620 ( .A(n3713), .B(n3714), .Z(n5837) );
  INV_X1 U4621 ( .A(n5837), .ZN(n3696) );
  AOI22_X1 U4622 ( .A1(n2951), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4623 ( .A1(n3983), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4624 ( .A1(n3836), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4625 ( .A1(n3224), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3682) );
  NAND4_X1 U4626 ( .A1(n3685), .A2(n3684), .A3(n3683), .A4(n3682), .ZN(n3691)
         );
  AOI22_X1 U4627 ( .A1(n3989), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3982), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4628 ( .A1(n3395), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4629 ( .A1(n3970), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4630 ( .A1(n3790), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3686) );
  NAND4_X1 U4631 ( .A1(n3689), .A2(n3688), .A3(n3687), .A4(n3686), .ZN(n3690)
         );
  OAI21_X1 U4632 ( .B1(n3691), .B2(n3690), .A(n3425), .ZN(n3694) );
  NAND2_X1 U4633 ( .A1(n3802), .A2(EAX_REG_15__SCAN_IN), .ZN(n3693) );
  NAND2_X1 U4634 ( .A1(n3424), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3692)
         );
  NAND3_X1 U4635 ( .A1(n3694), .A2(n3693), .A3(n3692), .ZN(n3695) );
  AOI21_X1 U4636 ( .B1(n3696), .B2(n3914), .A(n3695), .ZN(n5144) );
  NAND2_X1 U4637 ( .A1(n3697), .A2(n4491), .ZN(n6366) );
  AOI22_X1 U4638 ( .A1(n3790), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n2951), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4639 ( .A1(n3983), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4640 ( .A1(n3394), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4641 ( .A1(n3970), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3699) );
  NAND4_X1 U4642 ( .A1(n3702), .A2(n3701), .A3(n3700), .A4(n3699), .ZN(n3708)
         );
  AOI22_X1 U4643 ( .A1(n3989), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4644 ( .A1(n3982), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4645 ( .A1(n3328), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4646 ( .A1(n2952), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3703) );
  NAND4_X1 U4647 ( .A1(n3706), .A2(n3705), .A3(n3704), .A4(n3703), .ZN(n3707)
         );
  NOR2_X1 U4648 ( .A1(n3708), .A2(n3707), .ZN(n3712) );
  NAND2_X1 U4649 ( .A1(n6393), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3709)
         );
  NAND2_X1 U4650 ( .A1(n4003), .A2(n3709), .ZN(n3710) );
  AOI21_X1 U4651 ( .B1(n3802), .B2(EAX_REG_21__SCAN_IN), .A(n3710), .ZN(n3711)
         );
  OAI21_X1 U4652 ( .B1(n3979), .B2(n3712), .A(n3711), .ZN(n3718) );
  INV_X1 U4653 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5819) );
  OAI21_X1 U4654 ( .B1(n3716), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3852), 
        .ZN(n5679) );
  OR2_X1 U4655 ( .A1(n5679), .A2(n4003), .ZN(n3717) );
  NAND2_X1 U4656 ( .A1(n3718), .A2(n3717), .ZN(n5210) );
  INV_X1 U4657 ( .A(n5210), .ZN(n3809) );
  AOI22_X1 U4658 ( .A1(n3989), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n2951), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4659 ( .A1(n3983), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4660 ( .A1(n3315), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4661 ( .A1(n3469), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4662 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3729)
         );
  AOI22_X1 U4663 ( .A1(n3901), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4664 ( .A1(n3982), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4665 ( .A1(n3970), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4666 ( .A1(n3790), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3724) );
  NAND4_X1 U4667 ( .A1(n3727), .A2(n3726), .A3(n3725), .A4(n3724), .ZN(n3728)
         );
  NOR2_X1 U4668 ( .A1(n3729), .A2(n3728), .ZN(n3733) );
  NAND2_X1 U4669 ( .A1(n6393), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3730)
         );
  NAND2_X1 U4670 ( .A1(n4003), .A2(n3730), .ZN(n3731) );
  AOI21_X1 U4671 ( .B1(n3802), .B2(EAX_REG_20__SCAN_IN), .A(n3731), .ZN(n3732)
         );
  OAI21_X1 U4672 ( .B1(n3979), .B2(n3733), .A(n3732), .ZN(n3735) );
  XNOR2_X1 U4673 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3750), .ZN(n5690)
         );
  NAND2_X1 U4674 ( .A1(n5690), .A2(n4005), .ZN(n3734) );
  AND2_X1 U4675 ( .A1(n3735), .A2(n3734), .ZN(n5162) );
  AOI22_X1 U4676 ( .A1(n2951), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4677 ( .A1(n3983), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4678 ( .A1(n3309), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4679 ( .A1(n3328), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3736) );
  NAND4_X1 U4680 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3745)
         );
  AOI22_X1 U4681 ( .A1(n3982), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4682 ( .A1(n3989), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4683 ( .A1(n3970), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4684 ( .A1(n3790), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3740) );
  NAND4_X1 U4685 ( .A1(n3743), .A2(n3742), .A3(n3741), .A4(n3740), .ZN(n3744)
         );
  NOR2_X1 U4686 ( .A1(n3745), .A2(n3744), .ZN(n3749) );
  NAND2_X1 U4687 ( .A1(n6393), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3746)
         );
  NAND2_X1 U4688 ( .A1(n4003), .A2(n3746), .ZN(n3747) );
  AOI21_X1 U4689 ( .B1(n3802), .B2(EAX_REG_19__SCAN_IN), .A(n3747), .ZN(n3748)
         );
  OAI21_X1 U4690 ( .B1(n3979), .B2(n3749), .A(n3748), .ZN(n3753) );
  OAI21_X1 U4691 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n3751), .A(n3750), 
        .ZN(n5734) );
  OR2_X1 U4692 ( .A1(n4003), .A2(n5734), .ZN(n3752) );
  NAND2_X1 U4693 ( .A1(n3753), .A2(n3752), .ZN(n5235) );
  AOI22_X1 U4694 ( .A1(n3989), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4695 ( .A1(n3309), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4696 ( .A1(n3901), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4697 ( .A1(n3970), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4698 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3763)
         );
  AOI22_X1 U4699 ( .A1(n2951), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3982), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4700 ( .A1(n3983), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4701 ( .A1(n3984), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4702 ( .A1(n3790), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3758) );
  NAND4_X1 U4703 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3762)
         );
  NOR2_X1 U4704 ( .A1(n3763), .A2(n3762), .ZN(n3766) );
  OAI21_X1 U4705 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5819), .A(n4003), .ZN(
        n3764) );
  AOI21_X1 U4706 ( .B1(n3802), .B2(EAX_REG_18__SCAN_IN), .A(n3764), .ZN(n3765)
         );
  OAI21_X1 U4707 ( .B1(n3979), .B2(n3766), .A(n3765), .ZN(n3768) );
  XNOR2_X1 U4708 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3783), .ZN(n5817)
         );
  NAND2_X1 U4709 ( .A1(n5817), .A2(n3914), .ZN(n3767) );
  NAND2_X1 U4710 ( .A1(n3768), .A2(n3767), .ZN(n5436) );
  OR2_X1 U4711 ( .A1(n5235), .A2(n5436), .ZN(n3787) );
  AOI22_X1 U4712 ( .A1(n3790), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3969), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4713 ( .A1(n3901), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3982), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4714 ( .A1(n3315), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4715 ( .A1(n3970), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3769) );
  NAND4_X1 U4716 ( .A1(n3772), .A2(n3771), .A3(n3770), .A4(n3769), .ZN(n3778)
         );
  AOI22_X1 U4717 ( .A1(n3983), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4718 ( .A1(n2951), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4719 ( .A1(n3984), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4720 ( .A1(n2952), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3773) );
  NAND4_X1 U4721 ( .A1(n3776), .A2(n3775), .A3(n3774), .A4(n3773), .ZN(n3777)
         );
  NOR2_X1 U4722 ( .A1(n3778), .A2(n3777), .ZN(n3782) );
  INV_X1 U4723 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3779) );
  OAI21_X1 U4724 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3779), .A(n4003), .ZN(
        n3780) );
  AOI21_X1 U4725 ( .B1(n3802), .B2(EAX_REG_17__SCAN_IN), .A(n3780), .ZN(n3781)
         );
  OAI21_X1 U4726 ( .B1(n3979), .B2(n3782), .A(n3781), .ZN(n3786) );
  OAI21_X1 U4727 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3784), .A(n3783), 
        .ZN(n5826) );
  OR2_X1 U4728 ( .A1(n4003), .A2(n5826), .ZN(n3785) );
  NAND2_X1 U4729 ( .A1(n3786), .A2(n3785), .ZN(n5743) );
  NOR2_X1 U4730 ( .A1(n3787), .A2(n5743), .ZN(n5158) );
  AND2_X1 U4731 ( .A1(n5162), .A2(n5158), .ZN(n3808) );
  INV_X1 U4732 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3788) );
  XNOR2_X1 U4733 ( .A(n3789), .B(n3788), .ZN(n5151) );
  OR2_X1 U4734 ( .A1(n5151), .A2(n4003), .ZN(n3807) );
  AOI22_X1 U4735 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n3982), .B1(n3969), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4736 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3983), .B1(n3315), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4737 ( .A1(n3790), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4738 ( .A1(n3984), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3791) );
  NAND4_X1 U4739 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3801)
         );
  AOI22_X1 U4740 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3395), .B1(n3309), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4741 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n2951), .B1(n3945), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4742 ( .A1(n3970), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4743 ( .A1(n3836), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3796) );
  NAND4_X1 U4744 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n3800)
         );
  NOR2_X1 U4745 ( .A1(n3801), .A2(n3800), .ZN(n3804) );
  AOI22_X1 U4746 ( .A1(n3802), .A2(EAX_REG_16__SCAN_IN), .B1(n3424), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3803) );
  OAI21_X1 U4747 ( .B1(n3979), .B2(n3804), .A(n3803), .ZN(n3805) );
  INV_X1 U4748 ( .A(n3805), .ZN(n3806) );
  NAND2_X1 U4749 ( .A1(n3807), .A2(n3806), .ZN(n5157) );
  AOI22_X1 U4750 ( .A1(n2951), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4751 ( .A1(n3394), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n2955), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4752 ( .A1(n3983), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4753 ( .A1(n3982), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3811) );
  NAND4_X1 U4754 ( .A1(n3814), .A2(n3813), .A3(n3812), .A4(n3811), .ZN(n3820)
         );
  AOI22_X1 U4755 ( .A1(n3989), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4756 ( .A1(n3970), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4757 ( .A1(n3469), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4758 ( .A1(n3790), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3815) );
  NAND4_X1 U4759 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(n3819)
         );
  NOR2_X1 U4760 ( .A1(n3820), .A2(n3819), .ZN(n3823) );
  INV_X1 U4761 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5498) );
  AOI21_X1 U4762 ( .B1(n5498), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3821) );
  AOI21_X1 U4763 ( .B1(n3802), .B2(EAX_REG_22__SCAN_IN), .A(n3821), .ZN(n3822)
         );
  OAI21_X1 U4764 ( .B1(n3979), .B2(n3823), .A(n3822), .ZN(n3825) );
  XNOR2_X1 U4765 ( .A(n3852), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5669)
         );
  NAND2_X1 U4766 ( .A1(n5669), .A2(n4005), .ZN(n3824) );
  NAND2_X1 U4767 ( .A1(n3825), .A2(n3824), .ZN(n5202) );
  AOI22_X1 U4768 ( .A1(n2951), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4769 ( .A1(n3315), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4770 ( .A1(n3159), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4771 ( .A1(n3982), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3826) );
  NAND4_X1 U4772 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n3835)
         );
  AOI22_X1 U4773 ( .A1(n3969), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4774 ( .A1(n3970), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4775 ( .A1(n3469), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4776 ( .A1(n3790), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4777 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3834)
         );
  OR2_X1 U4778 ( .A1(n3835), .A2(n3834), .ZN(n3848) );
  AOI22_X1 U4779 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n2951), .B1(n3901), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4780 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n3309), .B1(n3315), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4781 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3983), .B1(n3308), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4782 ( .A1(n3982), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3837) );
  NAND4_X1 U4783 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3846)
         );
  AOI22_X1 U4784 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3989), .B1(n2952), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4785 ( .A1(n3970), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4786 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n3224), .B1(n3328), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4787 ( .A1(n3790), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3841) );
  NAND4_X1 U4788 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3845)
         );
  OR2_X1 U4789 ( .A1(n3846), .A2(n3845), .ZN(n3847) );
  NAND2_X1 U4790 ( .A1(n3847), .A2(n3848), .ZN(n3885) );
  OAI21_X1 U4791 ( .B1(n3848), .B2(n3847), .A(n3885), .ZN(n3849) );
  OR2_X1 U4792 ( .A1(n3979), .A2(n3849), .ZN(n3857) );
  NAND2_X1 U4793 ( .A1(n6393), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3850)
         );
  NAND2_X1 U4794 ( .A1(n4003), .A2(n3850), .ZN(n3851) );
  AOI21_X1 U4795 ( .B1(n3802), .B2(EAX_REG_23__SCAN_IN), .A(n3851), .ZN(n3856)
         );
  OR2_X1 U4796 ( .A1(n3853), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3854)
         );
  NAND2_X1 U4797 ( .A1(n3890), .A2(n3854), .ZN(n5492) );
  NOR2_X1 U4798 ( .A1(n5492), .A2(n4003), .ZN(n3855) );
  AOI21_X1 U4799 ( .B1(n3857), .B2(n3856), .A(n3855), .ZN(n5216) );
  AOI22_X1 U4800 ( .A1(n2951), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4801 ( .A1(n3982), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n2955), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4802 ( .A1(n3159), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4803 ( .A1(n3970), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3859) );
  NAND4_X1 U4804 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n3868)
         );
  AOI22_X1 U4805 ( .A1(n3969), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4806 ( .A1(n3308), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4807 ( .A1(n3984), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4808 ( .A1(n3790), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3863) );
  NAND4_X1 U4809 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(n3867)
         );
  NOR2_X1 U4810 ( .A1(n3868), .A2(n3867), .ZN(n3886) );
  XNOR2_X1 U4811 ( .A(n3885), .B(n3886), .ZN(n3869) );
  OR2_X1 U4812 ( .A1(n3979), .A2(n3869), .ZN(n3874) );
  XNOR2_X1 U4813 ( .A(n3890), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5659)
         );
  NAND2_X1 U4814 ( .A1(n3802), .A2(EAX_REG_24__SCAN_IN), .ZN(n3871) );
  NAND2_X1 U4815 ( .A1(n3424), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3870)
         );
  OAI211_X1 U4816 ( .C1(n5659), .C2(n4003), .A(n3871), .B(n3870), .ZN(n3872)
         );
  INV_X1 U4817 ( .A(n3872), .ZN(n3873) );
  NAND2_X1 U4818 ( .A1(n3874), .A2(n3873), .ZN(n5232) );
  AOI22_X1 U4819 ( .A1(n2951), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4820 ( .A1(n3315), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n2955), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4821 ( .A1(n3159), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4822 ( .A1(n3982), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3875) );
  NAND4_X1 U4823 ( .A1(n3878), .A2(n3877), .A3(n3876), .A4(n3875), .ZN(n3884)
         );
  AOI22_X1 U4824 ( .A1(n3989), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4825 ( .A1(n3970), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4826 ( .A1(n3328), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4827 ( .A1(n3790), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3879) );
  NAND4_X1 U4828 ( .A1(n3882), .A2(n3881), .A3(n3880), .A4(n3879), .ZN(n3883)
         );
  OR2_X1 U4829 ( .A1(n3884), .A2(n3883), .ZN(n3908) );
  NOR2_X1 U4830 ( .A1(n3886), .A2(n3885), .ZN(n3909) );
  XNOR2_X1 U4831 ( .A(n3908), .B(n3909), .ZN(n3889) );
  INV_X1 U4832 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3891) );
  OAI21_X1 U4833 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3891), .A(n4003), .ZN(
        n3887) );
  AOI21_X1 U4834 ( .B1(n3802), .B2(EAX_REG_25__SCAN_IN), .A(n3887), .ZN(n3888)
         );
  OAI21_X1 U4835 ( .B1(n3979), .B2(n3889), .A(n3888), .ZN(n3896) );
  INV_X1 U4836 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5483) );
  AND2_X1 U4837 ( .A1(n3892), .A2(n3891), .ZN(n3893) );
  OR2_X1 U4838 ( .A1(n3893), .A2(n3933), .ZN(n5727) );
  INV_X1 U4839 ( .A(n5727), .ZN(n3894) );
  NAND2_X1 U4840 ( .A1(n3894), .A2(n4005), .ZN(n3895) );
  NAND2_X1 U4841 ( .A1(n3896), .A2(n3895), .ZN(n5391) );
  AOI22_X1 U4842 ( .A1(n3969), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n2951), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4843 ( .A1(n2955), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4844 ( .A1(n3970), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3698), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4845 ( .A1(n3469), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3897) );
  NAND4_X1 U4846 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3907)
         );
  AOI22_X1 U4847 ( .A1(n3982), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4848 ( .A1(n3159), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4849 ( .A1(n3836), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4850 ( .A1(n3790), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3902) );
  NAND4_X1 U4851 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3906)
         );
  NOR2_X1 U4852 ( .A1(n3907), .A2(n3906), .ZN(n3918) );
  NAND2_X1 U4853 ( .A1(n3909), .A2(n3908), .ZN(n3917) );
  XOR2_X1 U4854 ( .A(n3918), .B(n3917), .Z(n3912) );
  INV_X1 U4855 ( .A(n3979), .ZN(n4000) );
  INV_X1 U4856 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U4857 ( .A1(n3802), .A2(EAX_REG_26__SCAN_IN), .ZN(n3910) );
  OAI211_X1 U4858 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n5658), .A(n3910), .B(
        n4003), .ZN(n3911) );
  AOI21_X1 U4859 ( .B1(n3912), .B2(n4000), .A(n3911), .ZN(n3913) );
  INV_X1 U4860 ( .A(n3913), .ZN(n3916) );
  XNOR2_X1 U4861 ( .A(n3933), .B(n5658), .ZN(n5649) );
  NAND2_X1 U4862 ( .A1(n5649), .A2(n3914), .ZN(n3915) );
  NAND2_X1 U4863 ( .A1(n3916), .A2(n3915), .ZN(n5423) );
  NOR2_X1 U4864 ( .A1(n3918), .A2(n3917), .ZN(n3940) );
  AOI22_X1 U4865 ( .A1(n2951), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4866 ( .A1(n3315), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n2955), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4867 ( .A1(n3159), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4868 ( .A1(n3982), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3919) );
  NAND4_X1 U4869 ( .A1(n3922), .A2(n3921), .A3(n3920), .A4(n3919), .ZN(n3928)
         );
  AOI22_X1 U4870 ( .A1(n3969), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4871 ( .A1(n3970), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4872 ( .A1(n3328), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4873 ( .A1(n3790), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3923) );
  NAND4_X1 U4874 ( .A1(n3926), .A2(n3925), .A3(n3924), .A4(n3923), .ZN(n3927)
         );
  OR2_X1 U4875 ( .A1(n3928), .A2(n3927), .ZN(n3939) );
  INV_X1 U4876 ( .A(n3939), .ZN(n3929) );
  XNOR2_X1 U4877 ( .A(n3940), .B(n3929), .ZN(n3930) );
  NAND2_X1 U4878 ( .A1(n3930), .A2(n4000), .ZN(n3938) );
  NAND2_X1 U4879 ( .A1(n6393), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3931)
         );
  NAND2_X1 U4880 ( .A1(n4003), .A2(n3931), .ZN(n3932) );
  AOI21_X1 U4881 ( .B1(n3802), .B2(EAX_REG_27__SCAN_IN), .A(n3932), .ZN(n3937)
         );
  OR2_X1 U4882 ( .A1(n3934), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3935)
         );
  NAND2_X1 U4883 ( .A1(n3959), .A2(n3935), .ZN(n5641) );
  NOR2_X1 U4884 ( .A1(n5641), .A2(n4003), .ZN(n3936) );
  AOI21_X1 U4885 ( .B1(n3938), .B2(n3937), .A(n3936), .ZN(n5414) );
  NAND2_X1 U4886 ( .A1(n3940), .A2(n3939), .ZN(n3963) );
  AOI22_X1 U4887 ( .A1(n3308), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4888 ( .A1(n2951), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4889 ( .A1(n3984), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4890 ( .A1(n3790), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3941) );
  NAND4_X1 U4891 ( .A1(n3944), .A2(n3943), .A3(n3942), .A4(n3941), .ZN(n3951)
         );
  AOI22_X1 U4892 ( .A1(n3836), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3969), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4893 ( .A1(n3159), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n2955), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4894 ( .A1(n3982), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3945), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4895 ( .A1(n3970), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3946) );
  NAND4_X1 U4896 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(n3950)
         );
  NOR2_X1 U4897 ( .A1(n3951), .A2(n3950), .ZN(n3964) );
  XOR2_X1 U4898 ( .A(n3963), .B(n3964), .Z(n3952) );
  NAND2_X1 U4899 ( .A1(n3952), .A2(n4000), .ZN(n3957) );
  NAND2_X1 U4900 ( .A1(n6393), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3953)
         );
  NAND2_X1 U4901 ( .A1(n4003), .A2(n3953), .ZN(n3954) );
  AOI21_X1 U4902 ( .B1(n3802), .B2(EAX_REG_28__SCAN_IN), .A(n3954), .ZN(n3956)
         );
  XNOR2_X1 U4903 ( .A(n3959), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5634)
         );
  AND2_X1 U4904 ( .A1(n5634), .A2(n4005), .ZN(n3955) );
  AOI21_X1 U4905 ( .B1(n3957), .B2(n3956), .A(n3955), .ZN(n5405) );
  INV_X1 U4906 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3958) );
  INV_X1 U4907 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3960) );
  NAND2_X1 U4908 ( .A1(n3961), .A2(n3960), .ZN(n3962) );
  NAND2_X1 U4909 ( .A1(n4011), .A2(n3962), .ZN(n5381) );
  NOR2_X1 U4910 ( .A1(n3964), .A2(n3963), .ZN(n3997) );
  AOI22_X1 U4911 ( .A1(n2951), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4912 ( .A1(n3394), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n2955), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4913 ( .A1(n3983), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4914 ( .A1(n3982), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3965) );
  NAND4_X1 U4915 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3965), .ZN(n3976)
         );
  AOI22_X1 U4916 ( .A1(n3969), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4917 ( .A1(n3970), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3984), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4918 ( .A1(n3328), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4919 ( .A1(n3790), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3971) );
  NAND4_X1 U4920 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(n3975)
         );
  OR2_X1 U4921 ( .A1(n3976), .A2(n3975), .ZN(n3996) );
  XNOR2_X1 U4922 ( .A(n3997), .B(n3996), .ZN(n3980) );
  AOI21_X1 U4923 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6393), .A(n4005), 
        .ZN(n3978) );
  NAND2_X1 U4924 ( .A1(n3802), .A2(EAX_REG_29__SCAN_IN), .ZN(n3977) );
  OAI211_X1 U4925 ( .C1(n3980), .C2(n3979), .A(n3978), .B(n3977), .ZN(n3981)
         );
  OAI21_X1 U4926 ( .B1(n4003), .B2(n5381), .A(n3981), .ZN(n5337) );
  AOI22_X1 U4927 ( .A1(n2951), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3982), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4928 ( .A1(n3983), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4929 ( .A1(n3984), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3224), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4930 ( .A1(n3790), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3985) );
  NAND4_X1 U4931 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(n3995)
         );
  AOI22_X1 U4932 ( .A1(n3901), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n2955), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4933 ( .A1(n3395), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3394), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4934 ( .A1(n3989), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n2952), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4935 ( .A1(n3970), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3990) );
  NAND4_X1 U4936 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(n3994)
         );
  NOR2_X1 U4937 ( .A1(n3995), .A2(n3994), .ZN(n3999) );
  NAND2_X1 U4938 ( .A1(n3997), .A2(n3996), .ZN(n3998) );
  XOR2_X1 U4939 ( .A(n3999), .B(n3998), .Z(n4001) );
  NAND2_X1 U4940 ( .A1(n4001), .A2(n4000), .ZN(n4008) );
  NAND2_X1 U4941 ( .A1(n6393), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4002)
         );
  NAND2_X1 U4942 ( .A1(n4003), .A2(n4002), .ZN(n4004) );
  AOI21_X1 U4943 ( .B1(n3802), .B2(EAX_REG_30__SCAN_IN), .A(n4004), .ZN(n4007)
         );
  XNOR2_X1 U4944 ( .A(n4011), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5368)
         );
  AND2_X1 U4945 ( .A1(n5368), .A2(n4005), .ZN(n4006) );
  AOI21_X1 U4946 ( .B1(n4008), .B2(n4007), .A(n4006), .ZN(n5356) );
  NAND2_X1 U4947 ( .A1(n5357), .A2(n5356), .ZN(n4009) );
  XOR2_X1 U4948 ( .A(n4010), .B(n4009), .Z(n5453) );
  INV_X1 U4949 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5359) );
  NOR2_X1 U4950 ( .A1(n4011), .A2(n5359), .ZN(n4012) );
  XNOR2_X1 U4951 ( .A(n4012), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5451)
         );
  NOR2_X1 U4952 ( .A1(n5451), .A2(n6403), .ZN(n4013) );
  NOR2_X1 U4953 ( .A1(n5918), .A2(n4014), .ZN(n4968) );
  NAND2_X1 U4954 ( .A1(REIP_REG_14__SCAN_IN), .A2(n4968), .ZN(n5138) );
  NOR2_X1 U4955 ( .A1(n5138), .A2(n4015), .ZN(n5816) );
  AND3_X1 U4956 ( .A1(n5816), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U4957 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5689), .ZN(n5685) );
  NOR2_X1 U4958 ( .A1(n5685), .A2(n4016), .ZN(n5393) );
  AND2_X1 U4959 ( .A1(n5393), .A2(n4017), .ZN(n5643) );
  NAND3_X1 U4960 ( .A1(n5643), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5385) );
  INV_X1 U4961 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5367) );
  INV_X1 U4962 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6476) );
  NOR4_X1 U4963 ( .A1(n5385), .A2(REIP_REG_31__SCAN_IN), .A3(n5367), .A4(n6476), .ZN(n4018) );
  NOR2_X1 U4964 ( .A1(n3348), .A2(n5799), .ZN(n4022) );
  AND2_X1 U4965 ( .A1(n6521), .A2(n6403), .ZN(n5627) );
  OAI21_X1 U4966 ( .B1(n5627), .B2(READREQUEST_REG_SCAN_IN), .A(n6523), .ZN(
        n4021) );
  OAI21_X1 U4967 ( .B1(n6523), .B2(n4022), .A(n4021), .ZN(U3474) );
  NAND2_X1 U4968 ( .A1(n4024), .A2(n5237), .ZN(n4028) );
  NAND2_X1 U4969 ( .A1(n4149), .A2(n4474), .ZN(n4987) );
  OR2_X1 U4970 ( .A1(n4987), .A2(n4466), .ZN(n4046) );
  NAND2_X1 U4971 ( .A1(n4326), .A2(n4149), .ZN(n4025) );
  NAND2_X1 U4972 ( .A1(n4025), .A2(n4466), .ZN(n4026) );
  AND2_X1 U4973 ( .A1(n4046), .A2(n4026), .ZN(n4027) );
  OAI211_X1 U4974 ( .C1(n3272), .C2(n4118), .A(n4028), .B(n4027), .ZN(n4032)
         );
  INV_X1 U4975 ( .A(n4324), .ZN(n4029) );
  NAND2_X1 U4976 ( .A1(n4029), .A2(n4415), .ZN(n4030) );
  NAND2_X1 U4977 ( .A1(n4031), .A2(n4030), .ZN(n4044) );
  NOR2_X1 U4978 ( .A1(n4032), .A2(n4044), .ZN(n4033) );
  NAND2_X1 U4979 ( .A1(n4034), .A2(n4033), .ZN(n4055) );
  OR2_X1 U4980 ( .A1(n6366), .A2(n4035), .ZN(n4276) );
  NAND2_X1 U4981 ( .A1(n4056), .A2(n4036), .ZN(n4037) );
  NAND2_X1 U4982 ( .A1(n4276), .A2(n4037), .ZN(n4038) );
  NOR2_X1 U4983 ( .A1(n4055), .A2(n4038), .ZN(n4157) );
  NOR2_X1 U4984 ( .A1(n6366), .A2(n3276), .ZN(n4125) );
  NAND2_X1 U4985 ( .A1(n4157), .A2(n4125), .ZN(n4257) );
  NOR2_X1 U4986 ( .A1(n6351), .A2(n3276), .ZN(n6369) );
  AOI21_X1 U4987 ( .B1(n3049), .B2(n6420), .A(READY_N), .ZN(n4039) );
  OAI21_X1 U4988 ( .B1(n6369), .B2(n4141), .A(n4039), .ZN(n4040) );
  INV_X1 U4989 ( .A(n4040), .ZN(n4049) );
  NOR2_X1 U4990 ( .A1(READY_N), .A2(n6349), .ZN(n4316) );
  INV_X1 U4991 ( .A(n4316), .ZN(n4047) );
  NAND2_X1 U4992 ( .A1(n6366), .A2(n4149), .ZN(n4042) );
  NAND2_X1 U4993 ( .A1(n4043), .A2(n4042), .ZN(n4140) );
  OR2_X1 U4994 ( .A1(n4140), .A2(n4044), .ZN(n4045) );
  NAND2_X1 U4995 ( .A1(n4045), .A2(n6351), .ZN(n4128) );
  OAI211_X1 U4996 ( .C1(n5786), .C2(n4047), .A(n4128), .B(n4046), .ZN(n4048)
         );
  AOI21_X1 U4997 ( .B1(n6394), .B2(n4049), .A(n4048), .ZN(n4051) );
  INV_X1 U4998 ( .A(n3348), .ZN(n4318) );
  NOR2_X1 U4999 ( .A1(n4140), .A2(n4318), .ZN(n6348) );
  NAND2_X1 U5000 ( .A1(n6394), .A2(n6348), .ZN(n4050) );
  OAI211_X1 U5001 ( .C1(n4257), .C2(n6394), .A(n4051), .B(n4050), .ZN(n6376)
         );
  NAND2_X1 U5002 ( .A1(n6376), .A2(n6399), .ZN(n5785) );
  INV_X1 U5003 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5802) );
  NOR2_X1 U5004 ( .A1(n6403), .A2(n6393), .ZN(n4307) );
  NAND2_X1 U5005 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4307), .ZN(n6487) );
  OR2_X1 U5006 ( .A1(n5802), .A2(n6487), .ZN(n4052) );
  NAND2_X1 U5007 ( .A1(n6402), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6488) );
  AND2_X1 U5008 ( .A1(n4052), .A2(n6488), .ZN(n4053) );
  NAND2_X1 U5009 ( .A1(n5785), .A2(n4053), .ZN(n6502) );
  INV_X1 U5010 ( .A(n6502), .ZN(n5262) );
  INV_X1 U5011 ( .A(n4055), .ZN(n4060) );
  INV_X1 U5012 ( .A(n4141), .ZN(n4058) );
  INV_X1 U5013 ( .A(n4056), .ZN(n4057) );
  AND3_X1 U5014 ( .A1(n4058), .A2(n5786), .A3(n4057), .ZN(n4059) );
  NAND2_X1 U5015 ( .A1(n4060), .A2(n4059), .ZN(n6364) );
  INV_X1 U5016 ( .A(n6364), .ZN(n4061) );
  OR2_X1 U5017 ( .A1(n5618), .A2(n4061), .ZN(n4065) );
  NOR2_X1 U5018 ( .A1(n4288), .A2(n5255), .ZN(n4063) );
  INV_X1 U5019 ( .A(n6366), .ZN(n4062) );
  AOI22_X1 U5020 ( .A1(n6369), .A2(n4258), .B1(n4063), .B2(n4062), .ZN(n4064)
         );
  NAND2_X1 U5021 ( .A1(n4065), .A2(n4064), .ZN(n6371) );
  INV_X1 U5022 ( .A(n6504), .ZN(n5787) );
  INV_X1 U5023 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5528) );
  AOI22_X1 U5024 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5528), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3023), .ZN(n5258) );
  INV_X1 U5025 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6498) );
  NOR2_X1 U5026 ( .A1(n6403), .A2(n6498), .ZN(n5253) );
  AOI222_X1 U5027 ( .A1(n6371), .A2(n5787), .B1(n5258), .B2(n5253), .C1(n4067), 
        .C2(n5254), .ZN(n4069) );
  NOR2_X1 U5028 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6492), .ZN(n6497)
         );
  OAI21_X1 U5029 ( .B1(n5262), .B2(n6497), .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .ZN(n4068) );
  OAI21_X1 U5030 ( .B1(n5262), .B2(n4069), .A(n4068), .ZN(U3460) );
  OR2_X1 U5031 ( .A1(n4257), .A2(n6406), .ZN(n4070) );
  NOR2_X1 U5032 ( .A1(n6394), .A2(n4070), .ZN(n4078) );
  INV_X1 U5033 ( .A(n4071), .ZN(n4076) );
  AND4_X1 U5034 ( .A1(n5437), .A2(n4134), .A3(n4073), .A4(n4072), .ZN(n4075)
         );
  NAND3_X1 U5035 ( .A1(n4076), .A2(n4075), .A3(n4074), .ZN(n4317) );
  NOR2_X1 U5036 ( .A1(n4317), .A2(n3049), .ZN(n4077) );
  AND2_X1 U5037 ( .A1(n5963), .A2(n4503), .ZN(n5954) );
  INV_X2 U5038 ( .A(n5954), .ZN(n5959) );
  OR2_X1 U5039 ( .A1(n4080), .A2(n4079), .ZN(n4081) );
  NAND2_X1 U5040 ( .A1(n4082), .A2(n4081), .ZN(n4993) );
  NAND2_X1 U5041 ( .A1(n5963), .A2(n5437), .ZN(n5958) );
  XNOR2_X1 U5042 ( .A(n4991), .B(n5799), .ZN(n6108) );
  INV_X1 U5043 ( .A(n5963), .ZN(n5319) );
  AOI22_X1 U5044 ( .A1(n5953), .A2(n6108), .B1(n5319), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4083) );
  OAI21_X1 U5045 ( .B1(n5959), .B2(n4993), .A(n4083), .ZN(U2858) );
  NAND2_X1 U5046 ( .A1(n4141), .A2(n4415), .ZN(n6390) );
  OR2_X1 U5047 ( .A1(n4437), .A2(n6390), .ZN(n6028) );
  INV_X2 U5048 ( .A(n6028), .ZN(n6022) );
  NOR2_X1 U5049 ( .A1(n5628), .A2(READY_N), .ZN(n4085) );
  OR2_X1 U5050 ( .A1(n6022), .A2(n4085), .ZN(n4084) );
  INV_X2 U5051 ( .A(n4084), .ZN(n6026) );
  AOI22_X1 U5052 ( .A1(n6026), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6022), .ZN(n4086) );
  NAND2_X1 U5053 ( .A1(n4085), .A2(n4474), .ZN(n4323) );
  NAND2_X1 U5054 ( .A1(n6025), .A2(DATAI_4_), .ZN(n4100) );
  NAND2_X1 U5055 ( .A1(n4086), .A2(n4100), .ZN(U2943) );
  AOI22_X1 U5056 ( .A1(n6026), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6022), .ZN(n4087) );
  NAND2_X1 U5057 ( .A1(n6025), .A2(DATAI_0_), .ZN(n4089) );
  NAND2_X1 U5058 ( .A1(n4087), .A2(n4089), .ZN(U2924) );
  AOI22_X1 U5059 ( .A1(n6026), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6022), .ZN(n4088) );
  INV_X1 U5060 ( .A(DATAI_13_), .ZN(n4761) );
  OR2_X1 U5061 ( .A1(n4323), .A2(n4761), .ZN(n4103) );
  NAND2_X1 U5062 ( .A1(n4088), .A2(n4103), .ZN(U2952) );
  AOI22_X1 U5063 ( .A1(n6026), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6022), .ZN(n4090) );
  NAND2_X1 U5064 ( .A1(n4090), .A2(n4089), .ZN(U2939) );
  AOI22_X1 U5065 ( .A1(n6026), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6022), .ZN(n4091) );
  NAND2_X1 U5066 ( .A1(n6025), .A2(DATAI_3_), .ZN(n4098) );
  NAND2_X1 U5067 ( .A1(n4091), .A2(n4098), .ZN(U2927) );
  AOI22_X1 U5068 ( .A1(n6026), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6022), .ZN(n4092) );
  NAND2_X1 U5069 ( .A1(n6025), .A2(DATAI_2_), .ZN(n4096) );
  NAND2_X1 U5070 ( .A1(n4092), .A2(n4096), .ZN(U2926) );
  AOI22_X1 U5071 ( .A1(n6026), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6022), .ZN(n4093) );
  NAND2_X1 U5072 ( .A1(n6025), .A2(DATAI_7_), .ZN(n4114) );
  NAND2_X1 U5073 ( .A1(n4093), .A2(n4114), .ZN(U2946) );
  AOI22_X1 U5074 ( .A1(n6026), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6022), .ZN(n4094) );
  NAND2_X1 U5075 ( .A1(n6025), .A2(DATAI_5_), .ZN(n4112) );
  NAND2_X1 U5076 ( .A1(n4094), .A2(n4112), .ZN(U2929) );
  AOI22_X1 U5077 ( .A1(n6026), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n6022), .ZN(n4095) );
  NAND2_X1 U5078 ( .A1(n6025), .A2(DATAI_12_), .ZN(n4105) );
  NAND2_X1 U5079 ( .A1(n4095), .A2(n4105), .ZN(U2951) );
  AOI22_X1 U5080 ( .A1(n6026), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6022), .ZN(n4097) );
  NAND2_X1 U5081 ( .A1(n4097), .A2(n4096), .ZN(U2941) );
  AOI22_X1 U5082 ( .A1(n6026), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6022), .ZN(n4099) );
  NAND2_X1 U5083 ( .A1(n4099), .A2(n4098), .ZN(U2942) );
  AOI22_X1 U5084 ( .A1(n6026), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6022), .ZN(n4101) );
  NAND2_X1 U5085 ( .A1(n4101), .A2(n4100), .ZN(U2928) );
  AOI22_X1 U5086 ( .A1(n6026), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6022), .ZN(n4102) );
  NAND2_X1 U5087 ( .A1(n6025), .A2(DATAI_6_), .ZN(n4108) );
  NAND2_X1 U5088 ( .A1(n4102), .A2(n4108), .ZN(U2945) );
  AOI22_X1 U5089 ( .A1(n6026), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6022), .ZN(n4104) );
  NAND2_X1 U5090 ( .A1(n4104), .A2(n4103), .ZN(U2937) );
  AOI22_X1 U5091 ( .A1(n6026), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n6022), .ZN(n4106) );
  NAND2_X1 U5092 ( .A1(n4106), .A2(n4105), .ZN(U2936) );
  AOI22_X1 U5093 ( .A1(n6026), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6022), .ZN(n4107) );
  NAND2_X1 U5094 ( .A1(n6025), .A2(DATAI_1_), .ZN(n4110) );
  NAND2_X1 U5095 ( .A1(n4107), .A2(n4110), .ZN(U2940) );
  AOI22_X1 U5096 ( .A1(n6026), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6022), .ZN(n4109) );
  NAND2_X1 U5097 ( .A1(n4109), .A2(n4108), .ZN(U2930) );
  AOI22_X1 U5098 ( .A1(n6026), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6022), .ZN(n4111) );
  NAND2_X1 U5099 ( .A1(n4111), .A2(n4110), .ZN(U2925) );
  AOI22_X1 U5100 ( .A1(n6026), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6022), .ZN(n4113) );
  NAND2_X1 U5101 ( .A1(n4113), .A2(n4112), .ZN(U2944) );
  AOI22_X1 U5102 ( .A1(n6026), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6022), .ZN(n4115) );
  NAND2_X1 U5103 ( .A1(n4115), .A2(n4114), .ZN(U2931) );
  INV_X1 U5104 ( .A(n4116), .ZN(n4117) );
  AOI21_X1 U5105 ( .B1(n4118), .B2(n6498), .A(n4117), .ZN(n5942) );
  INV_X1 U5106 ( .A(n5942), .ZN(n4124) );
  NAND2_X1 U5107 ( .A1(n4120), .A2(n4119), .ZN(n4121) );
  NAND2_X1 U5108 ( .A1(n4122), .A2(n4121), .ZN(n6052) );
  OAI222_X1 U5109 ( .A1(n4124), .A2(n5958), .B1(n5963), .B2(n4123), .C1(n6052), 
        .C2(n5959), .ZN(U2859) );
  INV_X1 U5110 ( .A(n4125), .ZN(n4129) );
  NAND2_X1 U5111 ( .A1(n4474), .A2(n6420), .ZN(n4126) );
  NAND3_X1 U5112 ( .A1(n4126), .A2(n4316), .A3(n4466), .ZN(n4127) );
  OAI211_X1 U5113 ( .C1(n6394), .C2(n4129), .A(n4128), .B(n4127), .ZN(n4130)
         );
  NAND2_X1 U5114 ( .A1(n4130), .A2(n6399), .ZN(n4138) );
  INV_X1 U5115 ( .A(READY_N), .ZN(n6572) );
  NAND3_X1 U5116 ( .A1(n4141), .A2(n4131), .A3(n6572), .ZN(n4133) );
  INV_X1 U5117 ( .A(n4326), .ZN(n4132) );
  NAND3_X1 U5118 ( .A1(n4133), .A2(n4592), .A3(n4132), .ZN(n4135) );
  NAND2_X1 U5119 ( .A1(n4135), .A2(n4134), .ZN(n4136) );
  OR2_X1 U5120 ( .A1(n4437), .A2(n4136), .ZN(n4137) );
  OR2_X1 U5121 ( .A1(n4140), .A2(n4139), .ZN(n6359) );
  NAND2_X1 U5122 ( .A1(n4141), .A2(n5799), .ZN(n4142) );
  OAI211_X1 U5123 ( .C1(n4155), .C2(n4143), .A(n4142), .B(n5786), .ZN(n4144)
         );
  INV_X1 U5124 ( .A(n4144), .ZN(n4145) );
  NAND2_X1 U5125 ( .A1(n6359), .A2(n4145), .ZN(n4146) );
  NOR2_X1 U5126 ( .A1(n6348), .A2(n4146), .ZN(n4147) );
  NOR2_X2 U5127 ( .A1(n4153), .A2(n4147), .ZN(n6112) );
  INV_X1 U5128 ( .A(n4148), .ZN(n4152) );
  INV_X1 U5129 ( .A(n4415), .ZN(n6525) );
  NAND2_X1 U5130 ( .A1(n4149), .A2(n4485), .ZN(n4207) );
  OAI21_X1 U5131 ( .B1(n6525), .B2(n4197), .A(n4207), .ZN(n4150) );
  INV_X1 U5132 ( .A(n4150), .ZN(n4151) );
  NAND2_X1 U5133 ( .A1(n4153), .A2(n4850), .ZN(n4247) );
  INV_X1 U5134 ( .A(n4247), .ZN(n4154) );
  NAND2_X1 U5135 ( .A1(n4159), .A2(n6369), .ZN(n5058) );
  INV_X1 U5136 ( .A(n5058), .ZN(n5776) );
  AOI211_X1 U5137 ( .C1(n6112), .C2(n4202), .A(n4154), .B(n5776), .ZN(n4163)
         );
  OAI21_X1 U5138 ( .B1(n4155), .B2(n4497), .A(n6390), .ZN(n4156) );
  NAND2_X1 U5139 ( .A1(n4159), .A2(n4156), .ZN(n6082) );
  INV_X1 U5140 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6512) );
  NOR2_X1 U5141 ( .A1(n4850), .A2(n6512), .ZN(n6045) );
  INV_X1 U5142 ( .A(n4257), .ZN(n6352) );
  INV_X1 U5143 ( .A(n4157), .ZN(n4158) );
  NAND2_X1 U5144 ( .A1(n4159), .A2(n4158), .ZN(n5062) );
  NAND2_X1 U5145 ( .A1(n5595), .A2(n5062), .ZN(n5061) );
  NAND2_X1 U5146 ( .A1(n6498), .A2(n5061), .ZN(n4248) );
  INV_X1 U5147 ( .A(n4248), .ZN(n4160) );
  AOI211_X1 U5148 ( .C1(n6109), .C2(n5942), .A(n6045), .B(n4160), .ZN(n4162)
         );
  NAND3_X1 U5149 ( .A1(n6112), .A2(n6041), .A3(n4202), .ZN(n4161) );
  OAI211_X1 U5150 ( .C1(n4163), .C2(n6498), .A(n4162), .B(n4161), .ZN(U3018)
         );
  INV_X1 U5151 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4168) );
  INV_X1 U5152 ( .A(n6369), .ZN(n4164) );
  OR2_X1 U5153 ( .A1(n4437), .A2(n4164), .ZN(n4165) );
  NAND2_X1 U5154 ( .A1(n6028), .A2(n4165), .ZN(n4166) );
  NAND2_X1 U5155 ( .A1(n5979), .A2(n4592), .ZN(n4380) );
  AOI22_X1 U5156 ( .A1(n4378), .A2(UWORD_REG_7__SCAN_IN), .B1(n5626), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4167) );
  OAI21_X1 U5157 ( .B1(n4168), .B2(n4380), .A(n4167), .ZN(U2900) );
  INV_X1 U5158 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5159 ( .A1(n4378), .A2(UWORD_REG_12__SCAN_IN), .B1(n5626), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4169) );
  OAI21_X1 U5160 ( .B1(n4170), .B2(n4380), .A(n4169), .ZN(U2895) );
  INV_X1 U5161 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5162 ( .A1(n4378), .A2(UWORD_REG_3__SCAN_IN), .B1(n5626), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4171) );
  OAI21_X1 U5163 ( .B1(n4172), .B2(n4380), .A(n4171), .ZN(U2904) );
  INV_X1 U5164 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5165 ( .A1(n4378), .A2(UWORD_REG_5__SCAN_IN), .B1(n5626), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4173) );
  OAI21_X1 U5166 ( .B1(n4174), .B2(n4380), .A(n4173), .ZN(U2902) );
  INV_X1 U5167 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5168 ( .A1(n4378), .A2(UWORD_REG_11__SCAN_IN), .B1(n5626), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4175) );
  OAI21_X1 U5169 ( .B1(n4176), .B2(n4380), .A(n4175), .ZN(U2896) );
  INV_X1 U5170 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U5171 ( .A1(n4378), .A2(UWORD_REG_4__SCAN_IN), .B1(n5626), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4177) );
  OAI21_X1 U5172 ( .B1(n4178), .B2(n4380), .A(n4177), .ZN(U2903) );
  INV_X1 U5173 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U5174 ( .A1(n4378), .A2(UWORD_REG_6__SCAN_IN), .B1(n5626), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4179) );
  OAI21_X1 U5175 ( .B1(n4180), .B2(n4380), .A(n4179), .ZN(U2901) );
  INV_X1 U5176 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4182) );
  AOI22_X1 U5177 ( .A1(n4378), .A2(UWORD_REG_2__SCAN_IN), .B1(n5626), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4181) );
  OAI21_X1 U5178 ( .B1(n4182), .B2(n4380), .A(n4181), .ZN(U2905) );
  INV_X1 U5179 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4184) );
  AOI22_X1 U5180 ( .A1(n4378), .A2(UWORD_REG_9__SCAN_IN), .B1(n5626), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4183) );
  OAI21_X1 U5181 ( .B1(n4184), .B2(n4380), .A(n4183), .ZN(U2898) );
  INV_X1 U5182 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U5183 ( .A1(n4378), .A2(UWORD_REG_8__SCAN_IN), .B1(n5626), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4185) );
  OAI21_X1 U5184 ( .B1(n4186), .B2(n4380), .A(n4185), .ZN(U2899) );
  OR2_X1 U5185 ( .A1(n4315), .A2(n4188), .ZN(n4189) );
  NAND2_X1 U5186 ( .A1(n4187), .A2(n4189), .ZN(n5935) );
  CLKBUF_X1 U5187 ( .A(n4191), .Z(n5317) );
  AOI21_X1 U5188 ( .B1(n5317), .B2(n5318), .A(n4192), .ZN(n4193) );
  OR2_X1 U5189 ( .A1(n4190), .A2(n4193), .ZN(n6081) );
  INV_X1 U5190 ( .A(n6081), .ZN(n4194) );
  AOI22_X1 U5191 ( .A1(n5953), .A2(n4194), .B1(n5319), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4195) );
  OAI21_X1 U5192 ( .B1(n5935), .B2(n5959), .A(n4195), .ZN(U2856) );
  XNOR2_X2 U5193 ( .A(n4202), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4718)
         );
  NAND2_X1 U5194 ( .A1(n4299), .A2(n4400), .ZN(n4201) );
  NAND2_X1 U5195 ( .A1(n4196), .A2(n4197), .ZN(n4205) );
  OAI21_X1 U5196 ( .B1(n4197), .B2(n4196), .A(n4205), .ZN(n4198) );
  OAI211_X1 U5197 ( .C1(n4198), .C2(n6525), .A(n3272), .B(n4491), .ZN(n4199)
         );
  INV_X1 U5198 ( .A(n4199), .ZN(n4200) );
  NAND2_X1 U5199 ( .A1(n4201), .A2(n4200), .ZN(n4717) );
  NAND2_X1 U5200 ( .A1(n4718), .A2(n4717), .ZN(n4716) );
  INV_X1 U5201 ( .A(n4202), .ZN(n6043) );
  NAND2_X1 U5202 ( .A1(n6043), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4203)
         );
  AND2_X1 U5203 ( .A1(n4716), .A2(n4203), .ZN(n6032) );
  INV_X1 U5204 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4210) );
  OR2_X1 U5205 ( .A1(n4410), .A2(n4210), .ZN(n4204) );
  OR2_X1 U5206 ( .A1(n4298), .A2(n4204), .ZN(n4212) );
  NAND2_X1 U5207 ( .A1(n4205), .A2(n4206), .ZN(n4218) );
  OAI21_X1 U5208 ( .B1(n4206), .B2(n4205), .A(n4218), .ZN(n4209) );
  INV_X1 U5209 ( .A(n4207), .ZN(n4208) );
  AOI21_X1 U5210 ( .B1(n4209), .B2(n4415), .A(n4208), .ZN(n4213) );
  OR2_X1 U5211 ( .A1(n4210), .A2(n4213), .ZN(n4211) );
  AND2_X1 U5212 ( .A1(n4212), .A2(n4211), .ZN(n6030) );
  NAND2_X1 U5213 ( .A1(n6032), .A2(n6030), .ZN(n4215) );
  OR2_X1 U5214 ( .A1(n4298), .A2(n4410), .ZN(n4214) );
  NAND2_X1 U5215 ( .A1(n2966), .A2(n4210), .ZN(n6031) );
  NAND2_X1 U5216 ( .A1(n4216), .A2(n4400), .ZN(n4221) );
  INV_X1 U5217 ( .A(n4217), .ZN(n4219) );
  NAND2_X1 U5218 ( .A1(n4218), .A2(n4219), .ZN(n4236) );
  OAI211_X1 U5219 ( .C1(n4219), .C2(n4218), .A(n4236), .B(n4415), .ZN(n4220)
         );
  INV_X1 U5220 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4222) );
  NAND2_X1 U5221 ( .A1(n4560), .A2(n4561), .ZN(n4225) );
  NAND2_X1 U5222 ( .A1(n4223), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4224)
         );
  NAND2_X1 U5223 ( .A1(n4225), .A2(n4224), .ZN(n4357) );
  NAND2_X1 U5224 ( .A1(n4226), .A2(n4400), .ZN(n4230) );
  XNOR2_X1 U5225 ( .A(n4236), .B(n4227), .ZN(n4228) );
  NAND2_X1 U5226 ( .A1(n4228), .A2(n4415), .ZN(n4229) );
  NAND2_X1 U5227 ( .A1(n4230), .A2(n4229), .ZN(n4231) );
  XNOR2_X1 U5228 ( .A(n4231), .B(n4361), .ZN(n4358) );
  NAND2_X1 U5229 ( .A1(n4357), .A2(n4358), .ZN(n4233) );
  NAND2_X1 U5230 ( .A1(n4231), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4232)
         );
  NAND2_X1 U5231 ( .A1(n4234), .A2(n4400), .ZN(n4243) );
  NOR2_X1 U5232 ( .A1(n4236), .A2(n4235), .ZN(n4238) );
  INV_X1 U5233 ( .A(n4239), .ZN(n4237) );
  NAND2_X1 U5234 ( .A1(n4238), .A2(n4237), .ZN(n4402) );
  INV_X1 U5235 ( .A(n4238), .ZN(n4240) );
  AOI21_X1 U5236 ( .B1(n4240), .B2(n4239), .A(n6525), .ZN(n4241) );
  NAND2_X1 U5237 ( .A1(n4402), .A2(n4241), .ZN(n4242) );
  NAND2_X1 U5238 ( .A1(n4243), .A2(n4242), .ZN(n4339) );
  INV_X1 U5239 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4244) );
  XNOR2_X1 U5240 ( .A(n4339), .B(n4244), .ZN(n4337) );
  XNOR2_X1 U5241 ( .A(n4338), .B(n4337), .ZN(n4459) );
  NAND2_X1 U5242 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4420) );
  INV_X1 U5243 ( .A(n4420), .ZN(n4360) );
  NAND2_X1 U5244 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U5245 ( .A1(n4210), .A2(n6093), .ZN(n6092) );
  NAND2_X1 U5246 ( .A1(n4360), .A2(n6092), .ZN(n4422) );
  NOR2_X1 U5247 ( .A1(n4210), .A2(n3023), .ZN(n4347) );
  NAND2_X1 U5248 ( .A1(n5058), .A2(n6498), .ZN(n6105) );
  INV_X1 U5249 ( .A(n6105), .ZN(n4245) );
  INV_X1 U5250 ( .A(n4958), .ZN(n6100) );
  NAND2_X1 U5251 ( .A1(n4347), .A2(n6100), .ZN(n4246) );
  OAI22_X1 U5252 ( .A1(n5595), .A2(n4422), .B1(n4420), .B2(n4246), .ZN(n4250)
         );
  NAND2_X1 U5253 ( .A1(n5284), .A2(n5595), .ZN(n6106) );
  INV_X1 U5254 ( .A(n6106), .ZN(n5297) );
  NOR2_X1 U5255 ( .A1(n4244), .A2(n4422), .ZN(n4249) );
  NAND2_X1 U5256 ( .A1(n4248), .A2(n4247), .ZN(n6110) );
  NAND2_X1 U5257 ( .A1(n5595), .A2(n6110), .ZN(n5285) );
  OAI21_X1 U5258 ( .B1(n5284), .B2(n4347), .A(n5285), .ZN(n6098) );
  INV_X1 U5259 ( .A(n6098), .ZN(n4359) );
  OAI21_X1 U5260 ( .B1(n5297), .B2(n4249), .A(n4359), .ZN(n4349) );
  OAI21_X1 U5261 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4250), .A(n4349), 
        .ZN(n4254) );
  INV_X1 U5262 ( .A(n4351), .ZN(n4251) );
  AOI21_X1 U5263 ( .B1(n4252), .B2(n4334), .A(n4251), .ZN(n5904) );
  INV_X1 U5264 ( .A(n4850), .ZN(n6107) );
  AND2_X1 U5265 ( .A1(n6107), .A2(REIP_REG_5__SCAN_IN), .ZN(n4455) );
  AOI21_X1 U5266 ( .B1(n6109), .B2(n5904), .A(n4455), .ZN(n4253) );
  OAI211_X1 U5267 ( .C1(n6084), .C2(n4459), .A(n4254), .B(n4253), .ZN(U3013)
         );
  OR2_X1 U5268 ( .A1(n6376), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4267)
         );
  INV_X1 U5269 ( .A(n6348), .ZN(n4256) );
  NAND2_X1 U5270 ( .A1(n4257), .A2(n4256), .ZN(n4279) );
  INV_X1 U5271 ( .A(n5255), .ZN(n5251) );
  NAND2_X1 U5272 ( .A1(n5251), .A2(n5263), .ZN(n4269) );
  NAND2_X1 U5273 ( .A1(n5255), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4270) );
  NAND2_X1 U5274 ( .A1(n4269), .A2(n4270), .ZN(n4259) );
  NAND2_X1 U5275 ( .A1(n4279), .A2(n4259), .ZN(n4264) );
  XNOR2_X1 U5276 ( .A(n4258), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4262)
         );
  INV_X1 U5277 ( .A(n4276), .ZN(n4261) );
  INV_X1 U5278 ( .A(n4259), .ZN(n4260) );
  AOI22_X1 U5279 ( .A1(n6369), .A2(n4262), .B1(n4261), .B2(n4260), .ZN(n4263)
         );
  NAND2_X1 U5280 ( .A1(n4264), .A2(n4263), .ZN(n4265) );
  AOI21_X1 U5281 ( .B1(n5621), .B2(n6364), .A(n4265), .ZN(n5252) );
  NAND2_X1 U5282 ( .A1(n6376), .A2(n5252), .ZN(n4266) );
  AND2_X1 U5283 ( .A1(n4267), .A2(n4266), .ZN(n6363) );
  OR2_X1 U5284 ( .A1(n6376), .A2(n4268), .ZN(n4283) );
  NAND2_X1 U5285 ( .A1(n5167), .A2(n6364), .ZN(n4281) );
  XNOR2_X1 U5286 ( .A(n4269), .B(n4268), .ZN(n4278) );
  AND2_X1 U5287 ( .A1(n4270), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4271)
         );
  NOR2_X1 U5288 ( .A1(n2952), .A2(n4271), .ZN(n6493) );
  NAND2_X1 U5289 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4272) );
  INV_X1 U5290 ( .A(n4272), .ZN(n4273) );
  MUX2_X1 U5291 ( .A(n4273), .B(n4272), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4274) );
  NAND2_X1 U5292 ( .A1(n6369), .A2(n4274), .ZN(n4275) );
  OAI21_X1 U5293 ( .B1(n6493), .B2(n4276), .A(n4275), .ZN(n4277) );
  AOI21_X1 U5294 ( .B1(n4279), .B2(n4278), .A(n4277), .ZN(n4280) );
  NAND2_X1 U5295 ( .A1(n4281), .A2(n4280), .ZN(n6491) );
  NAND2_X1 U5296 ( .A1(n6376), .A2(n6491), .ZN(n4282) );
  NAND2_X1 U5297 ( .A1(n4283), .A2(n4282), .ZN(n6383) );
  NAND3_X1 U5298 ( .A1(n6363), .A2(n6403), .A3(n6383), .ZN(n4287) );
  NAND2_X1 U5299 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5802), .ZN(n4294) );
  INV_X1 U5300 ( .A(n4294), .ZN(n4284) );
  NAND2_X1 U5301 ( .A1(n4285), .A2(n4284), .ZN(n4286) );
  NAND2_X1 U5302 ( .A1(n4287), .A2(n4286), .ZN(n6361) );
  INV_X1 U5303 ( .A(n4288), .ZN(n4289) );
  NAND2_X1 U5304 ( .A1(n6361), .A2(n4289), .ZN(n4308) );
  INV_X1 U5305 ( .A(n6207), .ZN(n4768) );
  NOR2_X1 U5306 ( .A1(n4290), .A2(n4768), .ZN(n4291) );
  XNOR2_X1 U5307 ( .A(n4291), .B(n4293), .ZN(n5916) );
  INV_X1 U5308 ( .A(n5916), .ZN(n4292) );
  OAI22_X1 U5309 ( .A1(n6376), .A2(n4293), .B1(n4292), .B2(n5786), .ZN(n4296)
         );
  NOR2_X1 U5310 ( .A1(n4294), .A2(n4293), .ZN(n4295) );
  AOI21_X1 U5311 ( .B1(n4296), .B2(n6403), .A(n4295), .ZN(n6360) );
  AND3_X1 U5312 ( .A1(n4308), .A2(n6360), .A3(n5802), .ZN(n4297) );
  INV_X1 U5313 ( .A(n4770), .ZN(n4677) );
  OAI21_X1 U5314 ( .B1(n4297), .B2(n6487), .A(n4770), .ZN(n6116) );
  OR2_X1 U5315 ( .A1(n4670), .A2(n4303), .ZN(n6117) );
  NOR2_X1 U5316 ( .A1(n6117), .A2(n4300), .ZN(n4814) );
  NAND2_X1 U5317 ( .A1(n4814), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4857) );
  INV_X1 U5318 ( .A(n4857), .ZN(n4302) );
  NOR2_X1 U5319 ( .A1(n4302), .A2(n6244), .ZN(n4652) );
  AND2_X1 U5320 ( .A1(n4300), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6243) );
  NAND2_X1 U5321 ( .A1(n6172), .A2(n6243), .ZN(n6210) );
  INV_X1 U5322 ( .A(n6521), .ZN(n6284) );
  AOI21_X1 U5323 ( .B1(n4652), .B2(n6210), .A(n6284), .ZN(n4305) );
  AND2_X1 U5324 ( .A1(n6521), .A2(n6621), .ZN(n6290) );
  INV_X1 U5325 ( .A(n6290), .ZN(n4672) );
  INV_X1 U5326 ( .A(n5167), .ZN(n5931) );
  AND2_X1 U5327 ( .A1(n6490), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5622) );
  OAI22_X1 U5328 ( .A1(n4301), .A2(n4672), .B1(n5931), .B2(n5622), .ZN(n4304)
         );
  OAI21_X1 U5329 ( .B1(n4305), .B2(n4304), .A(n6116), .ZN(n4306) );
  OAI21_X1 U5330 ( .B1(n6116), .B2(n6382), .A(n4306), .ZN(U3462) );
  NAND3_X1 U5331 ( .A1(n4308), .A2(n6360), .A3(n4307), .ZN(n6401) );
  INV_X1 U5332 ( .A(n6401), .ZN(n4310) );
  INV_X1 U5333 ( .A(n6365), .ZN(n6206) );
  OAI22_X1 U5334 ( .A1(n5009), .A2(n6284), .B1(n6206), .B2(n5622), .ZN(n4309)
         );
  OAI21_X1 U5335 ( .B1(n4310), .B2(n4309), .A(n6116), .ZN(n4311) );
  OAI21_X1 U5336 ( .B1(n6116), .B2(n5169), .A(n4311), .ZN(U3465) );
  NOR2_X1 U5337 ( .A1(n4313), .A2(n4312), .ZN(n4314) );
  OR2_X1 U5338 ( .A1(n4315), .A2(n4314), .ZN(n6029) );
  INV_X1 U5339 ( .A(n4437), .ZN(n4321) );
  NAND2_X1 U5340 ( .A1(n6399), .A2(n4316), .ZN(n4319) );
  OAI22_X1 U5341 ( .A1(n5786), .A2(n4319), .B1(n4318), .B2(n4317), .ZN(n4320)
         );
  AOI21_X1 U5342 ( .B1(n4321), .B2(n6348), .A(n4320), .ZN(n4322) );
  NAND2_X1 U5343 ( .A1(n4324), .A2(n4503), .ZN(n4325) );
  AND2_X1 U5344 ( .A1(n4327), .A2(n4503), .ZN(n4328) );
  INV_X1 U5345 ( .A(DATAI_2_), .ZN(n4467) );
  INV_X1 U5346 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6563) );
  OAI222_X1 U5347 ( .A1(n6029), .A2(n5695), .B1(n4760), .B2(n4467), .C1(n5978), 
        .C2(n6563), .ZN(U2889) );
  INV_X1 U5348 ( .A(DATAI_0_), .ZN(n4480) );
  INV_X1 U5349 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6008) );
  OAI222_X1 U5350 ( .A1(n6052), .A2(n5695), .B1(n4760), .B2(n4480), .C1(n5978), 
        .C2(n6008), .ZN(U2891) );
  INV_X1 U5351 ( .A(DATAI_1_), .ZN(n4475) );
  INV_X1 U5352 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6004) );
  OAI222_X1 U5353 ( .A1(n4993), .A2(n5695), .B1(n4760), .B2(n4475), .C1(n5978), 
        .C2(n6004), .ZN(U2890) );
  INV_X1 U5354 ( .A(DATAI_3_), .ZN(n4486) );
  INV_X1 U5355 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6001) );
  OAI222_X1 U5356 ( .A1(n5935), .A2(n5695), .B1(n4760), .B2(n4486), .C1(n5978), 
        .C2(n6001), .ZN(U2888) );
  INV_X1 U5357 ( .A(n4329), .ZN(n4330) );
  AOI21_X1 U5358 ( .B1(n4331), .B2(n4187), .A(n4330), .ZN(n5924) );
  INV_X1 U5359 ( .A(n5924), .ZN(n4356) );
  OR2_X1 U5360 ( .A1(n4190), .A2(n4332), .ZN(n4333) );
  NAND2_X1 U5361 ( .A1(n4334), .A2(n4333), .ZN(n5921) );
  INV_X1 U5362 ( .A(n5921), .ZN(n4335) );
  AOI22_X1 U5363 ( .A1(n5953), .A2(n4335), .B1(n5319), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4336) );
  OAI21_X1 U5364 ( .B1(n4356), .B2(n5959), .A(n4336), .ZN(U2855) );
  NAND2_X1 U5365 ( .A1(n4338), .A2(n4337), .ZN(n4341) );
  NAND2_X1 U5366 ( .A1(n4339), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4340)
         );
  NAND3_X1 U5367 ( .A1(n4413), .A2(n4342), .A3(n4400), .ZN(n4345) );
  XNOR2_X1 U5368 ( .A(n4402), .B(n4403), .ZN(n4343) );
  NAND2_X1 U5369 ( .A1(n4343), .A2(n4415), .ZN(n4344) );
  NAND2_X1 U5370 ( .A1(n4345), .A2(n4344), .ZN(n4397) );
  XNOR2_X1 U5371 ( .A(n4397), .B(n4346), .ZN(n4395) );
  XNOR2_X1 U5372 ( .A(n4396), .B(n4395), .ZN(n4454) );
  NOR3_X1 U5373 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4244), .A3(n4422), 
        .ZN(n4348) );
  INV_X1 U5374 ( .A(n4347), .ZN(n4421) );
  OAI21_X1 U5375 ( .B1(n4421), .B2(n4958), .A(n5595), .ZN(n4428) );
  AOI22_X1 U5376 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4349), .B1(n4348), 
        .B2(n4428), .ZN(n4355) );
  AND2_X1 U5377 ( .A1(n4351), .A2(n4350), .ZN(n4352) );
  OR2_X1 U5378 ( .A1(n4352), .A2(n4519), .ZN(n4589) );
  OAI22_X1 U5379 ( .A1(n6082), .A2(n4589), .B1(n6438), .B2(n4850), .ZN(n4353)
         );
  INV_X1 U5380 ( .A(n4353), .ZN(n4354) );
  OAI211_X1 U5381 ( .C1(n6084), .C2(n4454), .A(n4355), .B(n4354), .ZN(U3012)
         );
  INV_X1 U5382 ( .A(DATAI_4_), .ZN(n4498) );
  INV_X1 U5383 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5999) );
  OAI222_X1 U5384 ( .A1(n4356), .A2(n5695), .B1(n4760), .B2(n4498), .C1(n5978), 
        .C2(n5999), .ZN(U2887) );
  XNOR2_X1 U5385 ( .A(n4357), .B(n4358), .ZN(n4448) );
  OAI21_X1 U5386 ( .B1(n5595), .B2(n6092), .A(n4359), .ZN(n6079) );
  OAI22_X1 U5387 ( .A1(n6082), .A2(n5921), .B1(n6434), .B2(n4850), .ZN(n4363)
         );
  NAND2_X1 U5388 ( .A1(n6092), .A2(n4428), .ZN(n6088) );
  AOI211_X1 U5389 ( .C1(n4222), .C2(n4361), .A(n4360), .B(n6088), .ZN(n4362)
         );
  AOI211_X1 U5390 ( .C1(n6079), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4363), 
        .B(n4362), .ZN(n4364) );
  OAI21_X1 U5391 ( .B1(n6084), .B2(n4448), .A(n4364), .ZN(U3014) );
  NOR2_X1 U5392 ( .A1(n4384), .A2(n4366), .ZN(n4367) );
  OR2_X1 U5393 ( .A1(n4517), .A2(n4367), .ZN(n4601) );
  INV_X1 U5394 ( .A(n4589), .ZN(n4368) );
  AOI22_X1 U5395 ( .A1(n5953), .A2(n4368), .B1(n5319), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4369) );
  OAI21_X1 U5396 ( .B1(n4601), .B2(n5959), .A(n4369), .ZN(U2853) );
  INV_X1 U5397 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4371) );
  AOI22_X1 U5398 ( .A1(n4378), .A2(UWORD_REG_1__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4370) );
  OAI21_X1 U5399 ( .B1(n4371), .B2(n4380), .A(n4370), .ZN(U2906) );
  INV_X1 U5400 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4373) );
  AOI22_X1 U5401 ( .A1(n4378), .A2(UWORD_REG_13__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4372) );
  OAI21_X1 U5402 ( .B1(n4373), .B2(n4380), .A(n4372), .ZN(U2894) );
  INV_X1 U5403 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4375) );
  AOI22_X1 U5404 ( .A1(n4378), .A2(UWORD_REG_10__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4374) );
  OAI21_X1 U5405 ( .B1(n4375), .B2(n4380), .A(n4374), .ZN(U2897) );
  INV_X1 U5406 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U5407 ( .A1(n4378), .A2(UWORD_REG_0__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4376) );
  OAI21_X1 U5408 ( .B1(n4377), .B2(n4380), .A(n4376), .ZN(U2907) );
  INV_X1 U5409 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4381) );
  AOI22_X1 U5410 ( .A1(n4378), .A2(UWORD_REG_14__SCAN_IN), .B1(
        DATAO_REG_30__SCAN_IN), .B2(n6005), .ZN(n4379) );
  OAI21_X1 U5411 ( .B1(n4381), .B2(n4380), .A(n4379), .ZN(U2893) );
  AND2_X1 U5412 ( .A1(n4329), .A2(n4382), .ZN(n4383) );
  NOR2_X1 U5413 ( .A1(n4384), .A2(n4383), .ZN(n5908) );
  INV_X1 U5414 ( .A(n5908), .ZN(n4386) );
  AOI22_X1 U5415 ( .A1(n5953), .A2(n5904), .B1(n5319), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4385) );
  OAI21_X1 U5416 ( .B1(n4386), .B2(n5959), .A(n4385), .ZN(U2854) );
  INV_X1 U5417 ( .A(DATAI_6_), .ZN(n4510) );
  OAI222_X1 U5418 ( .A1(n4601), .A2(n5695), .B1(n4760), .B2(n4510), .C1(n5978), 
        .C2(n3545), .ZN(U2885) );
  INV_X1 U5419 ( .A(DATAI_5_), .ZN(n4492) );
  OAI222_X1 U5420 ( .A1(n4386), .A2(n5695), .B1(n4760), .B2(n4492), .C1(n5978), 
        .C2(n3528), .ZN(U2886) );
  AND2_X1 U5421 ( .A1(n4387), .A2(n4516), .ZN(n4388) );
  NAND2_X1 U5422 ( .A1(n4517), .A2(n4388), .ZN(n4434) );
  INV_X1 U5423 ( .A(n4434), .ZN(n4391) );
  OAI21_X1 U5424 ( .B1(n4391), .B2(n4390), .A(n4389), .ZN(n5003) );
  AOI21_X1 U5425 ( .B1(n4392), .B2(n4586), .A(n4572), .ZN(n6054) );
  AOI22_X1 U5426 ( .A1(n5953), .A2(n6054), .B1(n5319), .B2(EBX_REG_11__SCAN_IN), .ZN(n4393) );
  OAI21_X1 U5427 ( .B1(n5003), .B2(n5959), .A(n4393), .ZN(U2848) );
  AOI22_X1 U5428 ( .A1(n5974), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n5970), .ZN(n4394) );
  OAI21_X1 U5429 ( .B1(n5003), .B2(n5695), .A(n4394), .ZN(U2880) );
  NAND2_X1 U5430 ( .A1(n4396), .A2(n4395), .ZN(n4399) );
  NAND2_X1 U5431 ( .A1(n4397), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4398)
         );
  NAND2_X1 U5432 ( .A1(n4401), .A2(n4400), .ZN(n4407) );
  INV_X1 U5433 ( .A(n4402), .ZN(n4404) );
  NAND2_X1 U5434 ( .A1(n4404), .A2(n4403), .ZN(n4417) );
  XNOR2_X1 U5435 ( .A(n4417), .B(n4414), .ZN(n4405) );
  NAND2_X1 U5436 ( .A1(n4405), .A2(n4415), .ZN(n4406) );
  NAND2_X1 U5437 ( .A1(n4407), .A2(n4406), .ZN(n4408) );
  XNOR2_X1 U5438 ( .A(n4408), .B(n6077), .ZN(n4578) );
  NAND2_X1 U5439 ( .A1(n4577), .A2(n4578), .ZN(n4743) );
  NAND2_X1 U5440 ( .A1(n4408), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4741)
         );
  NAND2_X1 U5441 ( .A1(n4743), .A2(n4741), .ZN(n4730) );
  INV_X1 U5442 ( .A(n4409), .ZN(n4411) );
  NOR2_X1 U5443 ( .A1(n4411), .A2(n4410), .ZN(n4412) );
  NAND2_X1 U5444 ( .A1(n4415), .A2(n4414), .ZN(n4416) );
  OR2_X1 U5445 ( .A1(n4417), .A2(n4416), .ZN(n4418) );
  NAND2_X1 U5446 ( .A1(n4944), .A2(n4418), .ZN(n4731) );
  XNOR2_X1 U5447 ( .A(n4731), .B(n4419), .ZN(n4745) );
  XNOR2_X1 U5448 ( .A(n4730), .B(n4745), .ZN(n4624) );
  INV_X1 U5449 ( .A(n5285), .ZN(n4425) );
  NAND2_X1 U5450 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4423) );
  NOR3_X1 U5451 ( .A1(n4421), .A2(n4420), .A3(n4423), .ZN(n4957) );
  NOR2_X1 U5452 ( .A1(n4423), .A2(n4422), .ZN(n4955) );
  OAI22_X1 U5453 ( .A1(n5284), .A2(n4957), .B1(n4955), .B2(n5595), .ZN(n4424)
         );
  NOR2_X1 U5454 ( .A1(n4425), .A2(n4424), .ZN(n6078) );
  INV_X1 U5455 ( .A(n6078), .ZN(n4753) );
  OR2_X1 U5456 ( .A1(n4521), .A2(n4426), .ZN(n4427) );
  NAND2_X1 U5457 ( .A1(n4807), .A2(n4427), .ZN(n4610) );
  OAI22_X1 U5458 ( .A1(n6082), .A2(n4610), .B1(n6441), .B2(n4850), .ZN(n4430)
         );
  NOR2_X1 U5459 ( .A1(n6077), .A2(n4419), .ZN(n4752) );
  NAND2_X1 U5460 ( .A1(n4955), .A2(n4428), .ZN(n6073) );
  AOI211_X1 U5461 ( .C1(n6077), .C2(n4419), .A(n4752), .B(n6073), .ZN(n4429)
         );
  AOI211_X1 U5462 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n4753), .A(n4430), 
        .B(n4429), .ZN(n4431) );
  OAI21_X1 U5463 ( .B1(n6084), .B2(n4624), .A(n4431), .ZN(U3010) );
  AND2_X1 U5464 ( .A1(n4517), .A2(n4516), .ZN(n4433) );
  OAI21_X1 U5465 ( .B1(n4727), .B2(n4435), .A(n4434), .ZN(n5868) );
  AOI22_X1 U5466 ( .A1(n5974), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5970), .ZN(n4436) );
  OAI21_X1 U5467 ( .B1(n5868), .B2(n5695), .A(n4436), .ZN(U2881) );
  NAND2_X1 U5468 ( .A1(n4438), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6411) );
  OR2_X1 U5469 ( .A1(n6411), .A2(n6284), .ZN(n6051) );
  INV_X1 U5470 ( .A(n6051), .ZN(n6036) );
  NAND2_X1 U5471 ( .A1(n6284), .A2(n4439), .ZN(n4440) );
  NAND2_X1 U5472 ( .A1(n4440), .A2(n6402), .ZN(n4441) );
  NAND2_X1 U5473 ( .A1(n6402), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4443) );
  NAND2_X1 U5474 ( .A1(n6621), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4442) );
  NAND2_X1 U5475 ( .A1(n4443), .A2(n4442), .ZN(n6047) );
  INV_X1 U5476 ( .A(n4444), .ZN(n5927) );
  AOI22_X1 U5477 ( .A1(n6048), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6107), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4445) );
  OAI21_X1 U5478 ( .B1(n6040), .B2(n5927), .A(n4445), .ZN(n4446) );
  AOI21_X1 U5479 ( .B1(n5924), .B2(n6036), .A(n4446), .ZN(n4447) );
  OAI21_X1 U5480 ( .B1(n6042), .B2(n4448), .A(n4447), .ZN(U2982) );
  INV_X1 U5481 ( .A(n4601), .ZN(n4452) );
  INV_X1 U5482 ( .A(n4599), .ZN(n4450) );
  AOI22_X1 U5483 ( .A1(n6048), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6107), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n4449) );
  OAI21_X1 U5484 ( .B1(n6040), .B2(n4450), .A(n4449), .ZN(n4451) );
  AOI21_X1 U5485 ( .B1(n4452), .B2(n6036), .A(n4451), .ZN(n4453) );
  OAI21_X1 U5486 ( .B1(n6042), .B2(n4454), .A(n4453), .ZN(U2980) );
  AOI21_X1 U5487 ( .B1(n6048), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4455), 
        .ZN(n4456) );
  OAI21_X1 U5488 ( .B1(n6040), .B2(n5905), .A(n4456), .ZN(n4457) );
  AOI21_X1 U5489 ( .B1(n5908), .B2(n6036), .A(n4457), .ZN(n4458) );
  OAI21_X1 U5490 ( .B1(n6042), .B2(n4459), .A(n4458), .ZN(U2981) );
  AND2_X1 U5491 ( .A1(n5621), .A2(n5618), .ZN(n4856) );
  INV_X1 U5492 ( .A(n4884), .ZN(n4460) );
  NAND2_X1 U5493 ( .A1(n6244), .A2(n6118), .ZN(n6279) );
  AOI21_X1 U5494 ( .B1(n4460), .B2(n6279), .A(n6621), .ZN(n4461) );
  AOI211_X1 U5495 ( .C1(n4856), .C2(n5167), .A(n6284), .B(n4461), .ZN(n4463)
         );
  OR3_X1 U5496 ( .A1(n5168), .A2(n6382), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4860) );
  NOR2_X1 U5497 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4860), .ZN(n4509)
         );
  NOR2_X1 U5498 ( .A1(n4468), .A2(n6393), .ZN(n6180) );
  INV_X1 U5499 ( .A(n6180), .ZN(n6119) );
  OR2_X1 U5500 ( .A1(n6173), .A2(n4762), .ZN(n4529) );
  AOI21_X1 U5501 ( .B1(n4529), .B2(STATE2_REG_2__SCAN_IN), .A(n4770), .ZN(
        n4525) );
  OAI211_X1 U5502 ( .C1(n6490), .C2(n4509), .A(n6119), .B(n4525), .ZN(n4462)
         );
  NOR2_X1 U5503 ( .A1(n4463), .A2(n4462), .ZN(n4515) );
  INV_X1 U5504 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4473) );
  INV_X1 U5505 ( .A(n6488), .ZN(n4465) );
  NAND2_X1 U5506 ( .A1(n4508), .A2(n4466), .ZN(n4920) );
  NAND2_X1 U5507 ( .A1(n6036), .A2(DATAI_18_), .ZN(n6310) );
  INV_X1 U5508 ( .A(n6310), .ZN(n6257) );
  AOI22_X1 U5509 ( .A1(n6305), .A2(n4509), .B1(n6257), .B2(n4884), .ZN(n4472)
         );
  NOR2_X1 U5510 ( .A1(n4467), .A2(n4770), .ZN(n6306) );
  NOR2_X1 U5511 ( .A1(n5931), .A2(n6284), .ZN(n4813) );
  INV_X1 U5512 ( .A(n4813), .ZN(n4530) );
  INV_X1 U5513 ( .A(n4856), .ZN(n4469) );
  AND2_X1 U5514 ( .A1(n4468), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6174) );
  INV_X1 U5515 ( .A(n6174), .ZN(n4811) );
  OAI22_X1 U5516 ( .A1(n4530), .A2(n4469), .B1(n4811), .B2(n4529), .ZN(n4512)
         );
  INV_X1 U5517 ( .A(DATAI_26_), .ZN(n4470) );
  NOR2_X1 U5518 ( .A1(n6287), .A2(n4470), .ZN(n6307) );
  AOI22_X1 U5519 ( .A1(n6306), .A2(n4512), .B1(n6307), .B2(n6261), .ZN(n4471)
         );
  OAI211_X1 U5520 ( .C1(n4515), .C2(n4473), .A(n4472), .B(n4471), .ZN(U3118)
         );
  INV_X1 U5521 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4479) );
  NAND2_X1 U5522 ( .A1(n4508), .A2(n4474), .ZN(n4930) );
  NAND2_X1 U5523 ( .A1(n6036), .A2(DATAI_17_), .ZN(n6304) );
  INV_X1 U5524 ( .A(n6304), .ZN(n6253) );
  AOI22_X1 U5525 ( .A1(n6299), .A2(n4509), .B1(n6253), .B2(n4884), .ZN(n4478)
         );
  NOR2_X1 U5526 ( .A1(n4475), .A2(n4770), .ZN(n6300) );
  INV_X1 U5527 ( .A(DATAI_25_), .ZN(n4476) );
  NOR2_X1 U5528 ( .A1(n6287), .A2(n4476), .ZN(n6301) );
  AOI22_X1 U5529 ( .A1(n6300), .A2(n4512), .B1(n6301), .B2(n6261), .ZN(n4477)
         );
  OAI211_X1 U5530 ( .C1(n4515), .C2(n4479), .A(n4478), .B(n4477), .ZN(U3117)
         );
  INV_X1 U5531 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4484) );
  NAND2_X1 U5532 ( .A1(n4508), .A2(n4592), .ZN(n4916) );
  NAND2_X1 U5533 ( .A1(n6036), .A2(DATAI_16_), .ZN(n6298) );
  INV_X1 U5534 ( .A(n6298), .ZN(n6205) );
  AOI22_X1 U5535 ( .A1(n6285), .A2(n4509), .B1(n6205), .B2(n4884), .ZN(n4483)
         );
  NOR2_X1 U5536 ( .A1(n4480), .A2(n4770), .ZN(n6286) );
  INV_X1 U5537 ( .A(DATAI_24_), .ZN(n4481) );
  NOR2_X1 U5538 ( .A1(n6287), .A2(n4481), .ZN(n6295) );
  AOI22_X1 U5539 ( .A1(n6286), .A2(n4512), .B1(n6295), .B2(n6261), .ZN(n4482)
         );
  OAI211_X1 U5540 ( .C1(n4515), .C2(n4484), .A(n4483), .B(n4482), .ZN(U3116)
         );
  INV_X1 U5541 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4490) );
  NAND2_X1 U5542 ( .A1(n4508), .A2(n4485), .ZN(n4912) );
  NAND2_X1 U5543 ( .A1(n6036), .A2(DATAI_19_), .ZN(n6316) );
  INV_X1 U5544 ( .A(n6316), .ZN(n6262) );
  AOI22_X1 U5545 ( .A1(n6311), .A2(n4509), .B1(n6262), .B2(n4884), .ZN(n4489)
         );
  NOR2_X1 U5546 ( .A1(n4486), .A2(n4770), .ZN(n6312) );
  INV_X1 U5547 ( .A(DATAI_27_), .ZN(n4487) );
  NOR2_X1 U5548 ( .A1(n6287), .A2(n4487), .ZN(n6313) );
  AOI22_X1 U5549 ( .A1(n6312), .A2(n4512), .B1(n6313), .B2(n6261), .ZN(n4488)
         );
  OAI211_X1 U5550 ( .C1(n4515), .C2(n4490), .A(n4489), .B(n4488), .ZN(U3119)
         );
  INV_X1 U5551 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U5552 ( .A1(n4508), .A2(n4491), .ZN(n4904) );
  NAND2_X1 U5553 ( .A1(n6036), .A2(DATAI_21_), .ZN(n6328) );
  INV_X1 U5554 ( .A(n6328), .ZN(n6142) );
  AOI22_X1 U5555 ( .A1(n6323), .A2(n4509), .B1(n6142), .B2(n4884), .ZN(n4495)
         );
  NOR2_X1 U5556 ( .A1(n4492), .A2(n4770), .ZN(n6324) );
  INV_X1 U5557 ( .A(DATAI_29_), .ZN(n4493) );
  AOI22_X1 U5558 ( .A1(n6324), .A2(n4512), .B1(n6325), .B2(n6261), .ZN(n4494)
         );
  OAI211_X1 U5559 ( .C1(n4515), .C2(n4496), .A(n4495), .B(n4494), .ZN(U3121)
         );
  INV_X1 U5560 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4502) );
  NAND2_X1 U5561 ( .A1(n4508), .A2(n4497), .ZN(n4908) );
  NAND2_X1 U5562 ( .A1(n6036), .A2(DATAI_20_), .ZN(n6322) );
  INV_X1 U5563 ( .A(n6322), .ZN(n6138) );
  AOI22_X1 U5564 ( .A1(n6317), .A2(n4509), .B1(n6138), .B2(n4884), .ZN(n4501)
         );
  NOR2_X1 U5565 ( .A1(n4498), .A2(n4770), .ZN(n6318) );
  INV_X1 U5566 ( .A(DATAI_28_), .ZN(n4499) );
  AOI22_X1 U5567 ( .A1(n6318), .A2(n4512), .B1(n6319), .B2(n6261), .ZN(n4500)
         );
  OAI211_X1 U5568 ( .C1(n4515), .C2(n4502), .A(n4501), .B(n4500), .ZN(U3120)
         );
  INV_X1 U5569 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U5570 ( .A1(n4508), .A2(n4503), .ZN(n4924) );
  NAND2_X1 U5571 ( .A1(n6036), .A2(DATAI_23_), .ZN(n6345) );
  INV_X1 U5572 ( .A(n6345), .ZN(n6234) );
  AOI22_X1 U5573 ( .A1(n6335), .A2(n4509), .B1(n6234), .B2(n4884), .ZN(n4505)
         );
  INV_X1 U5574 ( .A(DATAI_7_), .ZN(n4523) );
  NOR2_X1 U5575 ( .A1(n4523), .A2(n4770), .ZN(n6338) );
  INV_X1 U5576 ( .A(DATAI_31_), .ZN(n6589) );
  NOR2_X1 U5577 ( .A1(n6287), .A2(n6589), .ZN(n6340) );
  AOI22_X1 U5578 ( .A1(n6338), .A2(n4512), .B1(n6340), .B2(n6261), .ZN(n4504)
         );
  OAI211_X1 U5579 ( .C1(n4515), .C2(n4506), .A(n4505), .B(n4504), .ZN(U3123)
         );
  INV_X1 U5580 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U5581 ( .A1(n4508), .A2(n4507), .ZN(n4900) );
  NAND2_X1 U5582 ( .A1(n6036), .A2(DATAI_22_), .ZN(n6334) );
  INV_X1 U5583 ( .A(n6334), .ZN(n6146) );
  AOI22_X1 U5584 ( .A1(n6329), .A2(n4509), .B1(n6146), .B2(n4884), .ZN(n4514)
         );
  NOR2_X1 U5585 ( .A1(n4510), .A2(n4770), .ZN(n6330) );
  INV_X1 U5586 ( .A(DATAI_30_), .ZN(n4511) );
  AOI22_X1 U5587 ( .A1(n6330), .A2(n4512), .B1(n6331), .B2(n6261), .ZN(n4513)
         );
  OAI211_X1 U5588 ( .C1(n4515), .C2(n6640), .A(n4514), .B(n4513), .ZN(U3122)
         );
  NAND2_X1 U5589 ( .A1(n4517), .A2(n4516), .ZN(n4603) );
  OAI21_X1 U5590 ( .B1(n4517), .B2(n4516), .A(n4603), .ZN(n5894) );
  INV_X1 U5591 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4522) );
  NOR2_X1 U5592 ( .A1(n4519), .A2(n4518), .ZN(n4520) );
  OR2_X1 U5593 ( .A1(n4521), .A2(n4520), .ZN(n5888) );
  OAI222_X1 U5594 ( .A1(n5894), .A2(n5959), .B1(n5963), .B2(n4522), .C1(n5888), 
        .C2(n5958), .ZN(U2852) );
  INV_X1 U5595 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5995) );
  OAI222_X1 U5596 ( .A1(n5894), .A2(n5695), .B1(n4760), .B2(n4523), .C1(n5978), 
        .C2(n5995), .ZN(U2884) );
  NAND2_X1 U5597 ( .A1(n6172), .A2(n6118), .ZN(n6232) );
  INV_X1 U5598 ( .A(n6232), .ZN(n6233) );
  INV_X1 U5599 ( .A(n5618), .ZN(n4810) );
  OR2_X1 U5600 ( .A1(n5621), .A2(n4810), .ZN(n6121) );
  OR2_X1 U5601 ( .A1(n5167), .A2(n6284), .ZN(n6176) );
  INV_X1 U5602 ( .A(n6176), .ZN(n4765) );
  AOI21_X1 U5603 ( .B1(n6521), .B2(n6121), .A(n4765), .ZN(n4524) );
  NOR3_X1 U5604 ( .A1(n4648), .A2(n6233), .A3(n4524), .ZN(n4528) );
  NAND3_X1 U5605 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5168), .A3(n6374), .ZN(n4629) );
  NOR2_X1 U5606 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4629), .ZN(n4531)
         );
  OAI211_X1 U5607 ( .C1(n6490), .C2(n4531), .A(n4811), .B(n4525), .ZN(n4527)
         );
  INV_X1 U5608 ( .A(n6121), .ZN(n4626) );
  NOR2_X1 U5609 ( .A1(n4626), .A2(n4672), .ZN(n4526) );
  NAND2_X1 U5610 ( .A1(n4553), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4534) );
  OAI22_X1 U5611 ( .A1(n4530), .A2(n6121), .B1(n6119), .B2(n4529), .ZN(n4556)
         );
  INV_X1 U5612 ( .A(n4531), .ZN(n4554) );
  INV_X1 U5613 ( .A(n6307), .ZN(n6260) );
  OAI22_X1 U5614 ( .A1(n4920), .A2(n4554), .B1(n6260), .B2(n6232), .ZN(n4532)
         );
  AOI21_X1 U5615 ( .B1(n6306), .B2(n4556), .A(n4532), .ZN(n4533) );
  OAI211_X1 U5616 ( .C1(n4559), .C2(n6310), .A(n4534), .B(n4533), .ZN(U3086)
         );
  NAND2_X1 U5617 ( .A1(n4553), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4537) );
  INV_X1 U5618 ( .A(n6301), .ZN(n6256) );
  OAI22_X1 U5619 ( .A1(n4930), .A2(n4554), .B1(n6256), .B2(n6232), .ZN(n4535)
         );
  AOI21_X1 U5620 ( .B1(n6300), .B2(n4556), .A(n4535), .ZN(n4536) );
  OAI211_X1 U5621 ( .C1(n4559), .C2(n6304), .A(n4537), .B(n4536), .ZN(U3085)
         );
  NAND2_X1 U5622 ( .A1(n4553), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4540) );
  INV_X1 U5623 ( .A(n6295), .ZN(n6218) );
  OAI22_X1 U5624 ( .A1(n4916), .A2(n4554), .B1(n6218), .B2(n6232), .ZN(n4538)
         );
  AOI21_X1 U5625 ( .B1(n6286), .B2(n4556), .A(n4538), .ZN(n4539) );
  OAI211_X1 U5626 ( .C1(n4559), .C2(n6298), .A(n4540), .B(n4539), .ZN(U3084)
         );
  NAND2_X1 U5627 ( .A1(n4553), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4543) );
  INV_X1 U5628 ( .A(n6313), .ZN(n6266) );
  OAI22_X1 U5629 ( .A1(n4912), .A2(n4554), .B1(n6266), .B2(n6232), .ZN(n4541)
         );
  AOI21_X1 U5630 ( .B1(n6312), .B2(n4556), .A(n4541), .ZN(n4542) );
  OAI211_X1 U5631 ( .C1(n4559), .C2(n6316), .A(n4543), .B(n4542), .ZN(U3087)
         );
  NAND2_X1 U5632 ( .A1(n4553), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4546) );
  INV_X1 U5633 ( .A(n6340), .ZN(n6241) );
  OAI22_X1 U5634 ( .A1(n4924), .A2(n4554), .B1(n6241), .B2(n6232), .ZN(n4544)
         );
  AOI21_X1 U5635 ( .B1(n6338), .B2(n4556), .A(n4544), .ZN(n4545) );
  OAI211_X1 U5636 ( .C1(n4559), .C2(n6345), .A(n4546), .B(n4545), .ZN(U3091)
         );
  NAND2_X1 U5637 ( .A1(n4553), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4549) );
  INV_X1 U5638 ( .A(n6331), .ZN(n6149) );
  OAI22_X1 U5639 ( .A1(n4900), .A2(n4554), .B1(n6149), .B2(n6232), .ZN(n4547)
         );
  AOI21_X1 U5640 ( .B1(n6330), .B2(n4556), .A(n4547), .ZN(n4548) );
  OAI211_X1 U5641 ( .C1(n4559), .C2(n6334), .A(n4549), .B(n4548), .ZN(U3090)
         );
  NAND2_X1 U5642 ( .A1(n4553), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4552) );
  INV_X1 U5643 ( .A(n6325), .ZN(n6145) );
  OAI22_X1 U5644 ( .A1(n4904), .A2(n4554), .B1(n6145), .B2(n6232), .ZN(n4550)
         );
  AOI21_X1 U5645 ( .B1(n6324), .B2(n4556), .A(n4550), .ZN(n4551) );
  OAI211_X1 U5646 ( .C1(n4559), .C2(n6328), .A(n4552), .B(n4551), .ZN(U3089)
         );
  NAND2_X1 U5647 ( .A1(n4553), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4558) );
  INV_X1 U5648 ( .A(n6319), .ZN(n6141) );
  OAI22_X1 U5649 ( .A1(n4908), .A2(n4554), .B1(n6141), .B2(n6232), .ZN(n4555)
         );
  AOI21_X1 U5650 ( .B1(n6318), .B2(n4556), .A(n4555), .ZN(n4557) );
  OAI211_X1 U5651 ( .C1(n4559), .C2(n6322), .A(n4558), .B(n4557), .ZN(U3088)
         );
  XNOR2_X1 U5652 ( .A(n4560), .B(n4561), .ZN(n6085) );
  INV_X1 U5653 ( .A(n5935), .ZN(n4564) );
  NAND2_X1 U5654 ( .A1(n5516), .A2(REIP_REG_3__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U5655 ( .A1(n6048), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4562)
         );
  OAI211_X1 U5656 ( .C1(n6040), .C2(n5934), .A(n6080), .B(n4562), .ZN(n4563)
         );
  AOI21_X1 U5657 ( .B1(n4564), .B2(n6036), .A(n4563), .ZN(n4565) );
  OAI21_X1 U5658 ( .B1(n6085), .B2(n6042), .A(n4565), .ZN(U2983) );
  INV_X1 U5659 ( .A(n4566), .ZN(n4569) );
  NAND2_X1 U5660 ( .A1(n4389), .A2(n4567), .ZN(n4568) );
  NAND2_X1 U5661 ( .A1(n4569), .A2(n4568), .ZN(n5858) );
  INV_X1 U5662 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4574) );
  OR2_X1 U5663 ( .A1(n4572), .A2(n4571), .ZN(n4573) );
  NAND2_X1 U5664 ( .A1(n4570), .A2(n4573), .ZN(n5854) );
  OAI222_X1 U5665 ( .A1(n5858), .A2(n5959), .B1(n5963), .B2(n4574), .C1(n5958), 
        .C2(n5854), .ZN(U2847) );
  INV_X1 U5666 ( .A(DATAI_12_), .ZN(n4576) );
  OAI222_X1 U5667 ( .A1(n5858), .A2(n5695), .B1(n4576), .B2(n4760), .C1(n4575), 
        .C2(n5978), .ZN(U2879) );
  XOR2_X1 U5668 ( .A(n4577), .B(n4578), .Z(n6075) );
  INV_X1 U5669 ( .A(n6042), .ZN(n6034) );
  NAND2_X1 U5670 ( .A1(n6075), .A2(n6034), .ZN(n4583) );
  INV_X1 U5671 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4579) );
  NAND2_X1 U5672 ( .A1(n5516), .A2(REIP_REG_7__SCAN_IN), .ZN(n6071) );
  OAI21_X1 U5673 ( .B1(n5523), .B2(n4579), .A(n6071), .ZN(n4580) );
  AOI21_X1 U5674 ( .B1(n5525), .B2(n4581), .A(n4580), .ZN(n4582) );
  OAI211_X1 U5675 ( .C1(n6051), .C2(n5894), .A(n4583), .B(n4582), .ZN(U2979)
         );
  INV_X1 U5676 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4587) );
  NAND2_X1 U5677 ( .A1(n4805), .A2(n4584), .ZN(n4585) );
  AND2_X1 U5678 ( .A1(n4586), .A2(n4585), .ZN(n5865) );
  INV_X1 U5679 ( .A(n5865), .ZN(n4754) );
  OAI222_X1 U5680 ( .A1(n5868), .A2(n5959), .B1(n5963), .B2(n4587), .C1(n5958), 
        .C2(n4754), .ZN(U2849) );
  AND2_X1 U5681 ( .A1(n5451), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4588) );
  NAND2_X1 U5682 ( .A1(n5900), .A2(n6438), .ZN(n5898) );
  OAI22_X1 U5683 ( .A1(n5933), .A2(n4589), .B1(n4590), .B2(n5898), .ZN(n4598)
         );
  OAI21_X1 U5684 ( .B1(n5913), .B2(n4590), .A(n5941), .ZN(n5911) );
  NOR2_X1 U5685 ( .A1(n6538), .A2(EBX_REG_31__SCAN_IN), .ZN(n4591) );
  AND2_X1 U5686 ( .A1(n4592), .A2(n4591), .ZN(n4593) );
  NOR2_X1 U5687 ( .A1(n4594), .A2(n4593), .ZN(n4595) );
  OR2_X1 U5688 ( .A1(n6523), .A2(n4595), .ZN(n5886) );
  AOI22_X1 U5689 ( .A1(EBX_REG_6__SCAN_IN), .A2(n5946), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n5901), .ZN(n4596) );
  OAI211_X1 U5690 ( .C1(n6438), .C2(n5911), .A(n4596), .B(n4850), .ZN(n4597)
         );
  AOI211_X1 U5691 ( .C1(n5907), .C2(n4599), .A(n4598), .B(n4597), .ZN(n4600)
         );
  OAI21_X1 U5692 ( .B1(n5893), .B2(n4601), .A(n4600), .ZN(U2821) );
  OR2_X1 U5693 ( .A1(n4603), .A2(n4604), .ZN(n4726) );
  INV_X1 U5694 ( .A(n4726), .ZN(n4602) );
  AOI21_X1 U5695 ( .B1(n4604), .B2(n4603), .A(n4602), .ZN(n4622) );
  INV_X1 U5696 ( .A(n4622), .ZN(n4618) );
  AOI22_X1 U5697 ( .A1(n5974), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n5970), .ZN(n4605) );
  OAI21_X1 U5698 ( .B1(n4618), .B2(n5695), .A(n4605), .ZN(U2883) );
  INV_X1 U5699 ( .A(n4610), .ZN(n4606) );
  AOI22_X1 U5700 ( .A1(n5953), .A2(n4606), .B1(n5319), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4607) );
  OAI21_X1 U5701 ( .B1(n4618), .B2(n5959), .A(n4607), .ZN(U2851) );
  INV_X1 U5702 ( .A(n4611), .ZN(n5872) );
  NAND2_X1 U5703 ( .A1(n5900), .A2(n5872), .ZN(n4608) );
  OAI22_X1 U5704 ( .A1(n5933), .A2(n4610), .B1(n4609), .B2(n4608), .ZN(n4615)
         );
  OAI21_X1 U5705 ( .B1(n5918), .B2(n4611), .A(n5321), .ZN(n5878) );
  AOI22_X1 U5706 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n5901), .B1(
        REIP_REG_8__SCAN_IN), .B2(n5878), .ZN(n4612) );
  OAI211_X1 U5707 ( .C1(n5886), .C2(n4613), .A(n4612), .B(n4850), .ZN(n4614)
         );
  AOI211_X1 U5708 ( .C1(n4616), .C2(n5907), .A(n4615), .B(n4614), .ZN(n4617)
         );
  OAI21_X1 U5709 ( .B1(n5893), .B2(n4618), .A(n4617), .ZN(U2819) );
  AOI22_X1 U5710 ( .A1(n6048), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6107), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4619) );
  OAI21_X1 U5711 ( .B1(n6040), .B2(n4620), .A(n4619), .ZN(n4621) );
  AOI21_X1 U5712 ( .B1(n4622), .B2(n6036), .A(n4621), .ZN(n4623) );
  OAI21_X1 U5713 ( .B1(n6042), .B2(n4624), .A(n4623), .ZN(U2978) );
  NAND2_X1 U5714 ( .A1(n4625), .A2(n5176), .ZN(n4890) );
  AOI21_X1 U5715 ( .B1(n5169), .B2(STATE2_REG_3__SCAN_IN), .A(n4770), .ZN(
        n6293) );
  AND2_X1 U5716 ( .A1(n5167), .A2(n6365), .ZN(n6282) );
  NOR2_X1 U5717 ( .A1(n5169), .A2(n4629), .ZN(n4649) );
  AOI21_X1 U5718 ( .B1(n6282), .B2(n4626), .A(n4649), .ZN(n4631) );
  NOR2_X1 U5719 ( .A1(n4300), .A2(n6621), .ZN(n5004) );
  AOI21_X1 U5720 ( .B1(n6244), .B2(n5004), .A(n6284), .ZN(n4628) );
  AOI22_X1 U5721 ( .A1(n4631), .A2(n4628), .B1(n6284), .B2(n4629), .ZN(n4627)
         );
  NAND2_X1 U5722 ( .A1(n6293), .A2(n4627), .ZN(n4647) );
  INV_X1 U5723 ( .A(n4628), .ZN(n4630) );
  OAI22_X1 U5724 ( .A1(n4631), .A2(n4630), .B1(n6393), .B2(n4629), .ZN(n4646)
         );
  AOI22_X1 U5725 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4647), .B1(n6306), 
        .B2(n4646), .ZN(n4633) );
  AOI22_X1 U5726 ( .A1(n6305), .A2(n4649), .B1(n4648), .B2(n6307), .ZN(n4632)
         );
  OAI211_X1 U5727 ( .C1(n6310), .C2(n4890), .A(n4633), .B(n4632), .ZN(U3094)
         );
  AOI22_X1 U5728 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4647), .B1(n6330), 
        .B2(n4646), .ZN(n4635) );
  AOI22_X1 U5729 ( .A1(n6329), .A2(n4649), .B1(n4648), .B2(n6331), .ZN(n4634)
         );
  OAI211_X1 U5730 ( .C1(n6334), .C2(n4890), .A(n4635), .B(n4634), .ZN(U3098)
         );
  AOI22_X1 U5731 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4647), .B1(n6338), 
        .B2(n4646), .ZN(n4637) );
  AOI22_X1 U5732 ( .A1(n6335), .A2(n4649), .B1(n4648), .B2(n6340), .ZN(n4636)
         );
  OAI211_X1 U5733 ( .C1(n6345), .C2(n4890), .A(n4637), .B(n4636), .ZN(U3099)
         );
  AOI22_X1 U5734 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4647), .B1(n6318), 
        .B2(n4646), .ZN(n4639) );
  AOI22_X1 U5735 ( .A1(n6317), .A2(n4649), .B1(n4648), .B2(n6319), .ZN(n4638)
         );
  OAI211_X1 U5736 ( .C1(n6322), .C2(n4890), .A(n4639), .B(n4638), .ZN(U3096)
         );
  AOI22_X1 U5737 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4647), .B1(n6286), 
        .B2(n4646), .ZN(n4641) );
  AOI22_X1 U5738 ( .A1(n6285), .A2(n4649), .B1(n4648), .B2(n6295), .ZN(n4640)
         );
  OAI211_X1 U5739 ( .C1(n6298), .C2(n4890), .A(n4641), .B(n4640), .ZN(U3092)
         );
  AOI22_X1 U5740 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4647), .B1(n6300), 
        .B2(n4646), .ZN(n4643) );
  AOI22_X1 U5741 ( .A1(n6299), .A2(n4649), .B1(n4648), .B2(n6301), .ZN(n4642)
         );
  OAI211_X1 U5742 ( .C1(n6304), .C2(n4890), .A(n4643), .B(n4642), .ZN(U3093)
         );
  AOI22_X1 U5743 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4647), .B1(n6312), 
        .B2(n4646), .ZN(n4645) );
  AOI22_X1 U5744 ( .A1(n6311), .A2(n4649), .B1(n4648), .B2(n6313), .ZN(n4644)
         );
  OAI211_X1 U5745 ( .C1(n6316), .C2(n4890), .A(n4645), .B(n4644), .ZN(U3095)
         );
  AOI22_X1 U5746 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4647), .B1(n6324), 
        .B2(n4646), .ZN(n4651) );
  AOI22_X1 U5747 ( .A1(n6323), .A2(n4649), .B1(n4648), .B2(n6325), .ZN(n4650)
         );
  OAI211_X1 U5748 ( .C1(n6328), .C2(n4890), .A(n4651), .B(n4650), .ZN(U3097)
         );
  NAND3_X1 U5749 ( .A1(n4652), .A2(n6243), .A3(n4670), .ZN(n4653) );
  NAND2_X1 U5750 ( .A1(n4653), .A2(n6521), .ZN(n4658) );
  NOR2_X1 U5751 ( .A1(n5621), .A2(n5618), .ZN(n4892) );
  AND2_X1 U5752 ( .A1(n5931), .A2(n4892), .ZN(n4673) );
  NOR2_X1 U5753 ( .A1(n6242), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6165)
         );
  AOI21_X1 U5754 ( .B1(n4673), .B2(n6365), .A(n6165), .ZN(n4654) );
  NAND3_X1 U5755 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6382), .A3(n5168), .ZN(n4676) );
  OAI22_X1 U5756 ( .A1(n4658), .A2(n4654), .B1(n4676), .B2(n6393), .ZN(n6166)
         );
  INV_X1 U5757 ( .A(n6166), .ZN(n4668) );
  INV_X1 U5758 ( .A(n6300), .ZN(n5044) );
  INV_X1 U5759 ( .A(n4654), .ZN(n4657) );
  INV_X1 U5760 ( .A(n6293), .ZN(n4655) );
  AOI21_X1 U5761 ( .B1(n6284), .B2(n4676), .A(n4655), .ZN(n4656) );
  OAI21_X1 U5762 ( .B1(n4658), .B2(n4657), .A(n4656), .ZN(n6167) );
  NAND2_X1 U5763 ( .A1(n4300), .A2(n5009), .ZN(n4815) );
  INV_X1 U5764 ( .A(n4815), .ZN(n6171) );
  NAND3_X1 U5765 ( .A1(n4301), .A2(n6171), .A3(n4670), .ZN(n4702) );
  NAND3_X1 U5766 ( .A1(n4301), .A2(n6118), .A3(n4670), .ZN(n6170) );
  AOI22_X1 U5767 ( .A1(n6299), .A2(n6165), .B1(n6253), .B2(n4767), .ZN(n4659)
         );
  OAI21_X1 U5768 ( .B1(n6256), .B2(n4702), .A(n4659), .ZN(n4660) );
  AOI21_X1 U5769 ( .B1(n6167), .B2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n4660), 
        .ZN(n4661) );
  OAI21_X1 U5770 ( .B1(n4668), .B2(n5044), .A(n4661), .ZN(U3045) );
  INV_X1 U5771 ( .A(n6286), .ZN(n5020) );
  AOI22_X1 U5772 ( .A1(n6285), .A2(n6165), .B1(n6205), .B2(n4767), .ZN(n4662)
         );
  OAI21_X1 U5773 ( .B1(n6218), .B2(n4702), .A(n4662), .ZN(n4663) );
  AOI21_X1 U5774 ( .B1(n6167), .B2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4663), 
        .ZN(n4664) );
  OAI21_X1 U5775 ( .B1(n4668), .B2(n5020), .A(n4664), .ZN(U3044) );
  INV_X1 U5776 ( .A(n6312), .ZN(n5051) );
  AOI22_X1 U5777 ( .A1(n6311), .A2(n6165), .B1(n6262), .B2(n4767), .ZN(n4665)
         );
  OAI21_X1 U5778 ( .B1(n6266), .B2(n4702), .A(n4665), .ZN(n4666) );
  AOI21_X1 U5779 ( .B1(n6167), .B2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4666), 
        .ZN(n4667) );
  OAI21_X1 U5780 ( .B1(n4668), .B2(n5051), .A(n4667), .ZN(U3047) );
  NOR2_X1 U5781 ( .A1(n6119), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4669)
         );
  AOI22_X1 U5782 ( .A1(n4673), .A2(n6521), .B1(n6173), .B2(n4669), .ZN(n4708)
         );
  INV_X1 U5783 ( .A(n6338), .ZN(n5028) );
  AND2_X1 U5784 ( .A1(n4670), .A2(n4766), .ZN(n4671) );
  NAND2_X1 U5785 ( .A1(n4671), .A2(n4301), .ZN(n5177) );
  INV_X1 U5786 ( .A(n5177), .ZN(n5171) );
  NAND2_X1 U5787 ( .A1(n5171), .A2(n5176), .ZN(n5197) );
  OAI21_X1 U5788 ( .B1(n4705), .B2(n6164), .A(n4672), .ZN(n4675) );
  INV_X1 U5789 ( .A(n4673), .ZN(n4674) );
  AOI21_X1 U5790 ( .B1(n4675), .B2(n4674), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4678) );
  NOR2_X1 U5791 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4676), .ZN(n4679)
         );
  OAI21_X1 U5792 ( .B1(n6173), .B2(n6393), .A(n4677), .ZN(n6179) );
  NOR2_X1 U5793 ( .A1(n6174), .A2(n6179), .ZN(n4897) );
  OAI21_X1 U5794 ( .B1(n4678), .B2(n4679), .A(n4897), .ZN(n4701) );
  NAND2_X1 U5795 ( .A1(n4701), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4682) );
  INV_X1 U5796 ( .A(n4679), .ZN(n4703) );
  OAI22_X1 U5797 ( .A1(n4924), .A2(n4703), .B1(n6345), .B2(n4702), .ZN(n4680)
         );
  AOI21_X1 U5798 ( .B1(n6340), .B2(n4705), .A(n4680), .ZN(n4681) );
  OAI211_X1 U5799 ( .C1(n4708), .C2(n5028), .A(n4682), .B(n4681), .ZN(U3043)
         );
  INV_X1 U5800 ( .A(n6330), .ZN(n5032) );
  NAND2_X1 U5801 ( .A1(n4701), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4685) );
  OAI22_X1 U5802 ( .A1(n4900), .A2(n4703), .B1(n6334), .B2(n4702), .ZN(n4683)
         );
  AOI21_X1 U5803 ( .B1(n6331), .B2(n4705), .A(n4683), .ZN(n4684) );
  OAI211_X1 U5804 ( .C1(n4708), .C2(n5032), .A(n4685), .B(n4684), .ZN(U3042)
         );
  INV_X1 U5805 ( .A(n6324), .ZN(n5040) );
  NAND2_X1 U5806 ( .A1(n4701), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4688) );
  OAI22_X1 U5807 ( .A1(n4904), .A2(n4703), .B1(n6328), .B2(n4702), .ZN(n4686)
         );
  AOI21_X1 U5808 ( .B1(n6325), .B2(n4705), .A(n4686), .ZN(n4687) );
  OAI211_X1 U5809 ( .C1(n4708), .C2(n5040), .A(n4688), .B(n4687), .ZN(U3041)
         );
  INV_X1 U5810 ( .A(n6318), .ZN(n5036) );
  NAND2_X1 U5811 ( .A1(n4701), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4691) );
  OAI22_X1 U5812 ( .A1(n4908), .A2(n4703), .B1(n6322), .B2(n4702), .ZN(n4689)
         );
  AOI21_X1 U5813 ( .B1(n6319), .B2(n4705), .A(n4689), .ZN(n4690) );
  OAI211_X1 U5814 ( .C1(n4708), .C2(n5036), .A(n4691), .B(n4690), .ZN(U3040)
         );
  NAND2_X1 U5815 ( .A1(n4701), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4694) );
  OAI22_X1 U5816 ( .A1(n4912), .A2(n4703), .B1(n6316), .B2(n4702), .ZN(n4692)
         );
  AOI21_X1 U5817 ( .B1(n6313), .B2(n4705), .A(n4692), .ZN(n4693) );
  OAI211_X1 U5818 ( .C1(n4708), .C2(n5051), .A(n4694), .B(n4693), .ZN(U3039)
         );
  NAND2_X1 U5819 ( .A1(n4701), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4697) );
  OAI22_X1 U5820 ( .A1(n4916), .A2(n4703), .B1(n6298), .B2(n4702), .ZN(n4695)
         );
  AOI21_X1 U5821 ( .B1(n6295), .B2(n4705), .A(n4695), .ZN(n4696) );
  OAI211_X1 U5822 ( .C1(n4708), .C2(n5020), .A(n4697), .B(n4696), .ZN(U3036)
         );
  INV_X1 U5823 ( .A(n6306), .ZN(n5024) );
  NAND2_X1 U5824 ( .A1(n4701), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4700) );
  OAI22_X1 U5825 ( .A1(n4920), .A2(n4703), .B1(n6310), .B2(n4702), .ZN(n4698)
         );
  AOI21_X1 U5826 ( .B1(n6307), .B2(n4705), .A(n4698), .ZN(n4699) );
  OAI211_X1 U5827 ( .C1(n4708), .C2(n5024), .A(n4700), .B(n4699), .ZN(U3038)
         );
  NAND2_X1 U5828 ( .A1(n4701), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4707) );
  OAI22_X1 U5829 ( .A1(n4930), .A2(n4703), .B1(n6304), .B2(n4702), .ZN(n4704)
         );
  AOI21_X1 U5830 ( .B1(n6301), .B2(n4705), .A(n4704), .ZN(n4706) );
  OAI211_X1 U5831 ( .C1(n4708), .C2(n5044), .A(n4707), .B(n4706), .ZN(U3037)
         );
  XNOR2_X1 U5832 ( .A(n4711), .B(n4710), .ZN(n5843) );
  NAND2_X1 U5833 ( .A1(n4570), .A2(n4712), .ZN(n4713) );
  NAND2_X1 U5834 ( .A1(n4936), .A2(n4713), .ZN(n5840) );
  INV_X1 U5835 ( .A(n5840), .ZN(n4714) );
  AOI22_X1 U5836 ( .A1(n4714), .A2(n5953), .B1(n5319), .B2(EBX_REG_13__SCAN_IN), .ZN(n4715) );
  OAI21_X1 U5837 ( .B1(n5843), .B2(n5959), .A(n4715), .ZN(U2846) );
  OAI21_X1 U5838 ( .B1(n4718), .B2(n4717), .A(n4716), .ZN(n4719) );
  INV_X1 U5839 ( .A(n4719), .ZN(n6111) );
  INV_X1 U5840 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4720) );
  NAND2_X1 U5841 ( .A1(n5525), .A2(n4720), .ZN(n4722) );
  AOI22_X1 U5842 ( .A1(n6048), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6107), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4721) );
  OAI211_X1 U5843 ( .C1(n4993), .C2(n6051), .A(n4722), .B(n4721), .ZN(n4723)
         );
  AOI21_X1 U5844 ( .B1(n6034), .B2(n6111), .A(n4723), .ZN(n4724) );
  INV_X1 U5845 ( .A(n4724), .ZN(U2985) );
  AND2_X1 U5846 ( .A1(n4726), .A2(n4725), .ZN(n4728) );
  AOI22_X1 U5847 ( .A1(n5974), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n5970), .ZN(n4729) );
  OAI21_X1 U5848 ( .B1(n5881), .B2(n5695), .A(n4729), .ZN(U2882) );
  NAND2_X1 U5849 ( .A1(n4730), .A2(n4745), .ZN(n4732) );
  NAND2_X1 U5850 ( .A1(n4731), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4739)
         );
  NAND2_X1 U5851 ( .A1(n4732), .A2(n4739), .ZN(n4734) );
  INV_X1 U5852 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6068) );
  XNOR2_X1 U5853 ( .A(n5517), .B(n6068), .ZN(n4733) );
  XNOR2_X1 U5854 ( .A(n4734), .B(n4733), .ZN(n6065) );
  NAND2_X1 U5855 ( .A1(n6065), .A2(n6034), .ZN(n4737) );
  NAND2_X1 U5856 ( .A1(n5516), .A2(REIP_REG_9__SCAN_IN), .ZN(n6061) );
  OAI21_X1 U5857 ( .B1(n5523), .B2(n6625), .A(n6061), .ZN(n4735) );
  AOI21_X1 U5858 ( .B1(n5525), .B2(n5883), .A(n4735), .ZN(n4736) );
  OAI211_X1 U5859 ( .C1(n6287), .C2(n5881), .A(n4737), .B(n4736), .ZN(U2977)
         );
  OR2_X1 U5860 ( .A1(n4944), .A2(n6068), .ZN(n4738) );
  NAND2_X1 U5861 ( .A1(n4947), .A2(n6068), .ZN(n4744) );
  AND2_X1 U5862 ( .A1(n4741), .A2(n4746), .ZN(n4742) );
  NAND2_X1 U5863 ( .A1(n4743), .A2(n4742), .ZN(n4749) );
  NAND2_X1 U5864 ( .A1(n4745), .A2(n4744), .ZN(n4747) );
  NAND2_X1 U5865 ( .A1(n4747), .A2(n4746), .ZN(n4748) );
  NAND2_X1 U5866 ( .A1(n4749), .A2(n4748), .ZN(n4940) );
  INV_X1 U5867 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6650) );
  AND2_X1 U5868 ( .A1(n5517), .A2(n6650), .ZN(n4994) );
  INV_X1 U5869 ( .A(n4994), .ZN(n4750) );
  NAND2_X1 U5870 ( .A1(n5737), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4996) );
  NAND2_X1 U5871 ( .A1(n4750), .A2(n4996), .ZN(n4751) );
  XNOR2_X1 U5872 ( .A(n4995), .B(n4751), .ZN(n4855) );
  INV_X1 U5873 ( .A(n4752), .ZN(n4954) );
  AOI21_X1 U5874 ( .B1(n4954), .B2(n6106), .A(n4753), .ZN(n6069) );
  NOR2_X1 U5875 ( .A1(n4954), .A2(n6073), .ZN(n6064) );
  NAND2_X1 U5876 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4953) );
  OAI211_X1 U5877 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6064), .B(n4953), .ZN(n4757) );
  OAI22_X1 U5878 ( .A1(n6082), .A2(n4754), .B1(n6445), .B2(n4850), .ZN(n4755)
         );
  INV_X1 U5879 ( .A(n4755), .ZN(n4756) );
  OAI211_X1 U5880 ( .C1(n6069), .C2(n6650), .A(n4757), .B(n4756), .ZN(n4758)
         );
  INV_X1 U5881 ( .A(n4758), .ZN(n4759) );
  OAI21_X1 U5882 ( .B1(n4855), .B2(n6084), .A(n4759), .ZN(U3008) );
  INV_X1 U5883 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5984) );
  OAI222_X1 U5884 ( .A1(n5695), .A2(n5843), .B1(n5978), .B2(n5984), .C1(n4761), 
        .C2(n4760), .ZN(U2878) );
  INV_X1 U5885 ( .A(n4762), .ZN(n4763) );
  OR2_X1 U5886 ( .A1(n6173), .A2(n4763), .ZN(n6120) );
  INV_X1 U5887 ( .A(n6120), .ZN(n4764) );
  AOI22_X1 U5888 ( .A1(n4765), .A2(n4856), .B1(n6174), .B2(n4764), .ZN(n4801)
         );
  NAND3_X1 U5889 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6382), .A3(n6374), .ZN(n5013) );
  NOR2_X1 U5890 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5013), .ZN(n4774)
         );
  NAND2_X1 U5891 ( .A1(n6172), .A2(n4766), .ZN(n5010) );
  OAI21_X1 U5892 ( .B1(n5011), .B2(n4767), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4769) );
  NAND2_X1 U5893 ( .A1(n4856), .A2(n4768), .ZN(n5005) );
  AND2_X1 U5894 ( .A1(n4769), .A2(n5005), .ZN(n4772) );
  AOI21_X1 U5895 ( .B1(n6120), .B2(STATE2_REG_2__SCAN_IN), .A(n4770), .ZN(
        n4771) );
  INV_X1 U5896 ( .A(n4771), .ZN(n6123) );
  AOI211_X1 U5897 ( .C1(n6521), .C2(n4772), .A(n6180), .B(n6123), .ZN(n4773)
         );
  OAI21_X1 U5898 ( .B1(n4774), .B2(n6490), .A(n4773), .ZN(n4796) );
  NAND2_X1 U5899 ( .A1(n4796), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4777) );
  INV_X1 U5900 ( .A(n4774), .ZN(n4797) );
  OAI22_X1 U5901 ( .A1(n4920), .A2(n4797), .B1(n6260), .B2(n6170), .ZN(n4775)
         );
  AOI21_X1 U5902 ( .B1(n6257), .B2(n5011), .A(n4775), .ZN(n4776) );
  OAI211_X1 U5903 ( .C1(n4801), .C2(n5024), .A(n4777), .B(n4776), .ZN(U3054)
         );
  NAND2_X1 U5904 ( .A1(n4796), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4780) );
  OAI22_X1 U5905 ( .A1(n4900), .A2(n4797), .B1(n6149), .B2(n6170), .ZN(n4778)
         );
  AOI21_X1 U5906 ( .B1(n6146), .B2(n5011), .A(n4778), .ZN(n4779) );
  OAI211_X1 U5907 ( .C1(n4801), .C2(n5032), .A(n4780), .B(n4779), .ZN(U3058)
         );
  NAND2_X1 U5908 ( .A1(n4796), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4783) );
  OAI22_X1 U5909 ( .A1(n4908), .A2(n4797), .B1(n6141), .B2(n6170), .ZN(n4781)
         );
  AOI21_X1 U5910 ( .B1(n6138), .B2(n5011), .A(n4781), .ZN(n4782) );
  OAI211_X1 U5911 ( .C1(n4801), .C2(n5036), .A(n4783), .B(n4782), .ZN(U3056)
         );
  NAND2_X1 U5912 ( .A1(n4796), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4786) );
  OAI22_X1 U5913 ( .A1(n4916), .A2(n4797), .B1(n6218), .B2(n6170), .ZN(n4784)
         );
  AOI21_X1 U5914 ( .B1(n6205), .B2(n5011), .A(n4784), .ZN(n4785) );
  OAI211_X1 U5915 ( .C1(n4801), .C2(n5020), .A(n4786), .B(n4785), .ZN(U3052)
         );
  NAND2_X1 U5916 ( .A1(n4796), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4789) );
  OAI22_X1 U5917 ( .A1(n4912), .A2(n4797), .B1(n6266), .B2(n6170), .ZN(n4787)
         );
  AOI21_X1 U5918 ( .B1(n6262), .B2(n5011), .A(n4787), .ZN(n4788) );
  OAI211_X1 U5919 ( .C1(n4801), .C2(n5051), .A(n4789), .B(n4788), .ZN(U3055)
         );
  NAND2_X1 U5920 ( .A1(n4796), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4792) );
  OAI22_X1 U5921 ( .A1(n4930), .A2(n4797), .B1(n6256), .B2(n6170), .ZN(n4790)
         );
  AOI21_X1 U5922 ( .B1(n6253), .B2(n5011), .A(n4790), .ZN(n4791) );
  OAI211_X1 U5923 ( .C1(n4801), .C2(n5044), .A(n4792), .B(n4791), .ZN(U3053)
         );
  NAND2_X1 U5924 ( .A1(n4796), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4795) );
  OAI22_X1 U5925 ( .A1(n4924), .A2(n4797), .B1(n6241), .B2(n6170), .ZN(n4793)
         );
  AOI21_X1 U5926 ( .B1(n6234), .B2(n5011), .A(n4793), .ZN(n4794) );
  OAI211_X1 U5927 ( .C1(n4801), .C2(n5028), .A(n4795), .B(n4794), .ZN(U3059)
         );
  NAND2_X1 U5928 ( .A1(n4796), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4800) );
  OAI22_X1 U5929 ( .A1(n4904), .A2(n4797), .B1(n6145), .B2(n6170), .ZN(n4798)
         );
  AOI21_X1 U5930 ( .B1(n6142), .B2(n5011), .A(n4798), .ZN(n4799) );
  OAI211_X1 U5931 ( .C1(n4801), .C2(n5040), .A(n4800), .B(n4799), .ZN(U3057)
         );
  OAI21_X1 U5932 ( .B1(n4803), .B2(n4802), .A(n5145), .ZN(n5076) );
  AOI22_X1 U5933 ( .A1(n5974), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n5970), .ZN(n4804) );
  OAI21_X1 U5934 ( .B1(n5076), .B2(n5695), .A(n4804), .ZN(U2877) );
  INV_X1 U5935 ( .A(n4805), .ZN(n4806) );
  AOI21_X1 U5936 ( .B1(n4808), .B2(n4807), .A(n4806), .ZN(n6063) );
  INV_X1 U5937 ( .A(n6063), .ZN(n4809) );
  INV_X1 U5938 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5887) );
  OAI222_X1 U5939 ( .A1(n4809), .A2(n5958), .B1(n5963), .B2(n5887), .C1(n5959), 
        .C2(n5881), .ZN(U2850) );
  AND2_X1 U5940 ( .A1(n5621), .A2(n4810), .ZN(n6281) );
  NOR2_X1 U5941 ( .A1(n4811), .A2(n6382), .ZN(n4812) );
  AOI22_X1 U5942 ( .A1(n4813), .A2(n6281), .B1(n6173), .B2(n4812), .ZN(n4849)
         );
  INV_X1 U5943 ( .A(n6294), .ZN(n6283) );
  NOR2_X1 U5944 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6283), .ZN(n4821)
         );
  INV_X1 U5945 ( .A(n4882), .ZN(n4816) );
  AOI21_X1 U5946 ( .B1(n4816), .B2(n4844), .A(n6621), .ZN(n4818) );
  INV_X1 U5947 ( .A(n6281), .ZN(n6208) );
  NAND2_X1 U5948 ( .A1(n6208), .A2(n6521), .ZN(n4817) );
  NOR2_X1 U5949 ( .A1(n4818), .A2(n4817), .ZN(n4819) );
  NOR4_X1 U5950 ( .A1(n6382), .A2(n6180), .A3(n4819), .A4(n6179), .ZN(n4820)
         );
  NAND2_X1 U5951 ( .A1(n4843), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4824)
         );
  INV_X1 U5952 ( .A(n4821), .ZN(n4845) );
  OAI22_X1 U5953 ( .A1(n4924), .A2(n4845), .B1(n4844), .B2(n6345), .ZN(n4822)
         );
  AOI21_X1 U5954 ( .B1(n4882), .B2(n6340), .A(n4822), .ZN(n4823) );
  OAI211_X1 U5955 ( .C1(n4849), .C2(n5028), .A(n4824), .B(n4823), .ZN(U3139)
         );
  NAND2_X1 U5956 ( .A1(n4843), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4827)
         );
  OAI22_X1 U5957 ( .A1(n4916), .A2(n4845), .B1(n6298), .B2(n4844), .ZN(n4825)
         );
  AOI21_X1 U5958 ( .B1(n6295), .B2(n4882), .A(n4825), .ZN(n4826) );
  OAI211_X1 U5959 ( .C1(n4849), .C2(n5020), .A(n4827), .B(n4826), .ZN(U3132)
         );
  NAND2_X1 U5960 ( .A1(n4843), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4830)
         );
  OAI22_X1 U5961 ( .A1(n4908), .A2(n4845), .B1(n4844), .B2(n6322), .ZN(n4828)
         );
  AOI21_X1 U5962 ( .B1(n4882), .B2(n6319), .A(n4828), .ZN(n4829) );
  OAI211_X1 U5963 ( .C1(n4849), .C2(n5036), .A(n4830), .B(n4829), .ZN(U3136)
         );
  NAND2_X1 U5964 ( .A1(n4843), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4833)
         );
  OAI22_X1 U5965 ( .A1(n4900), .A2(n4845), .B1(n4844), .B2(n6334), .ZN(n4831)
         );
  AOI21_X1 U5966 ( .B1(n4882), .B2(n6331), .A(n4831), .ZN(n4832) );
  OAI211_X1 U5967 ( .C1(n4849), .C2(n5032), .A(n4833), .B(n4832), .ZN(U3138)
         );
  NAND2_X1 U5968 ( .A1(n4843), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4836)
         );
  OAI22_X1 U5969 ( .A1(n4920), .A2(n4845), .B1(n4844), .B2(n6310), .ZN(n4834)
         );
  AOI21_X1 U5970 ( .B1(n4882), .B2(n6307), .A(n4834), .ZN(n4835) );
  OAI211_X1 U5971 ( .C1(n4849), .C2(n5024), .A(n4836), .B(n4835), .ZN(U3134)
         );
  NAND2_X1 U5972 ( .A1(n4843), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4839)
         );
  OAI22_X1 U5973 ( .A1(n4930), .A2(n4845), .B1(n4844), .B2(n6304), .ZN(n4837)
         );
  AOI21_X1 U5974 ( .B1(n4882), .B2(n6301), .A(n4837), .ZN(n4838) );
  OAI211_X1 U5975 ( .C1(n4849), .C2(n5044), .A(n4839), .B(n4838), .ZN(U3133)
         );
  NAND2_X1 U5976 ( .A1(n4843), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4842)
         );
  OAI22_X1 U5977 ( .A1(n4912), .A2(n4845), .B1(n4844), .B2(n6316), .ZN(n4840)
         );
  AOI21_X1 U5978 ( .B1(n4882), .B2(n6313), .A(n4840), .ZN(n4841) );
  OAI211_X1 U5979 ( .C1(n4849), .C2(n5051), .A(n4842), .B(n4841), .ZN(U3135)
         );
  NAND2_X1 U5980 ( .A1(n4843), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4848)
         );
  OAI22_X1 U5981 ( .A1(n4904), .A2(n4845), .B1(n4844), .B2(n6328), .ZN(n4846)
         );
  AOI21_X1 U5982 ( .B1(n4882), .B2(n6325), .A(n4846), .ZN(n4847) );
  OAI211_X1 U5983 ( .C1(n4849), .C2(n5040), .A(n4848), .B(n4847), .ZN(U3137)
         );
  INV_X1 U5984 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4851) );
  OAI22_X1 U5985 ( .A1(n5523), .A2(n4851), .B1(n4850), .B2(n6445), .ZN(n4853)
         );
  NOR2_X1 U5986 ( .A1(n5868), .A2(n6287), .ZN(n4852) );
  AOI211_X1 U5987 ( .C1(n5525), .C2(n5869), .A(n4853), .B(n4852), .ZN(n4854)
         );
  OAI21_X1 U5988 ( .B1(n6042), .B2(n4855), .A(n4854), .ZN(U2976) );
  NOR2_X1 U5989 ( .A1(n5169), .A2(n4860), .ZN(n4883) );
  AOI21_X1 U5990 ( .B1(n6282), .B2(n4856), .A(n4883), .ZN(n4861) );
  NAND2_X1 U5991 ( .A1(n4861), .A2(n4857), .ZN(n4858) );
  NOR2_X1 U5992 ( .A1(n6284), .A2(n4858), .ZN(n4859) );
  AOI211_X2 U5993 ( .C1(n6284), .C2(n4860), .A(n4859), .B(n4655), .ZN(n4889)
         );
  INV_X1 U5994 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4864) );
  AOI22_X1 U5995 ( .A1(n6323), .A2(n4883), .B1(n4882), .B2(n6142), .ZN(n4863)
         );
  OAI22_X1 U5996 ( .A1(n4861), .A2(n6284), .B1(n4860), .B2(n6393), .ZN(n4885)
         );
  AOI22_X1 U5997 ( .A1(n6324), .A2(n4885), .B1(n6325), .B2(n4884), .ZN(n4862)
         );
  OAI211_X1 U5998 ( .C1(n4889), .C2(n4864), .A(n4863), .B(n4862), .ZN(U3129)
         );
  INV_X1 U5999 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4867) );
  AOI22_X1 U6000 ( .A1(n6317), .A2(n4883), .B1(n4882), .B2(n6138), .ZN(n4866)
         );
  AOI22_X1 U6001 ( .A1(n6318), .A2(n4885), .B1(n6319), .B2(n4884), .ZN(n4865)
         );
  OAI211_X1 U6002 ( .C1(n4889), .C2(n4867), .A(n4866), .B(n4865), .ZN(U3128)
         );
  INV_X1 U6003 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6586) );
  AOI22_X1 U6004 ( .A1(n6285), .A2(n4883), .B1(n4882), .B2(n6205), .ZN(n4869)
         );
  AOI22_X1 U6005 ( .A1(n6286), .A2(n4885), .B1(n6295), .B2(n4884), .ZN(n4868)
         );
  OAI211_X1 U6006 ( .C1(n4889), .C2(n6586), .A(n4869), .B(n4868), .ZN(U3124)
         );
  INV_X1 U6007 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4872) );
  AOI22_X1 U6008 ( .A1(n6299), .A2(n4883), .B1(n4882), .B2(n6253), .ZN(n4871)
         );
  AOI22_X1 U6009 ( .A1(n6300), .A2(n4885), .B1(n6301), .B2(n4884), .ZN(n4870)
         );
  OAI211_X1 U6010 ( .C1(n4889), .C2(n4872), .A(n4871), .B(n4870), .ZN(U3125)
         );
  INV_X1 U6011 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4875) );
  AOI22_X1 U6012 ( .A1(n6329), .A2(n4883), .B1(n4882), .B2(n6146), .ZN(n4874)
         );
  AOI22_X1 U6013 ( .A1(n6330), .A2(n4885), .B1(n6331), .B2(n4884), .ZN(n4873)
         );
  OAI211_X1 U6014 ( .C1(n4889), .C2(n4875), .A(n4874), .B(n4873), .ZN(U3130)
         );
  INV_X1 U6015 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4878) );
  AOI22_X1 U6016 ( .A1(n6305), .A2(n4883), .B1(n4882), .B2(n6257), .ZN(n4877)
         );
  AOI22_X1 U6017 ( .A1(n6306), .A2(n4885), .B1(n6307), .B2(n4884), .ZN(n4876)
         );
  OAI211_X1 U6018 ( .C1(n4889), .C2(n4878), .A(n4877), .B(n4876), .ZN(U3126)
         );
  INV_X1 U6019 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4881) );
  AOI22_X1 U6020 ( .A1(n6335), .A2(n4883), .B1(n4882), .B2(n6234), .ZN(n4880)
         );
  AOI22_X1 U6021 ( .A1(n6338), .A2(n4885), .B1(n6340), .B2(n4884), .ZN(n4879)
         );
  OAI211_X1 U6022 ( .C1(n4889), .C2(n4881), .A(n4880), .B(n4879), .ZN(U3131)
         );
  INV_X1 U6023 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4888) );
  AOI22_X1 U6024 ( .A1(n6311), .A2(n4883), .B1(n4882), .B2(n6262), .ZN(n4887)
         );
  AOI22_X1 U6025 ( .A1(n6312), .A2(n4885), .B1(n6313), .B2(n4884), .ZN(n4886)
         );
  OAI211_X1 U6026 ( .C1(n4889), .C2(n4888), .A(n4887), .B(n4886), .ZN(U3127)
         );
  NAND2_X1 U6027 ( .A1(n6244), .A2(n6171), .ZN(n6265) );
  OAI21_X1 U6028 ( .B1(n4932), .B2(n6273), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4891) );
  NAND2_X1 U6029 ( .A1(n4891), .A2(n6521), .ZN(n4898) );
  INV_X1 U6030 ( .A(n4898), .ZN(n4894) );
  AND2_X1 U6031 ( .A1(n4892), .A2(n5167), .ZN(n6245) );
  NOR2_X1 U6032 ( .A1(n6119), .A2(n6382), .ZN(n4893) );
  AOI22_X1 U6033 ( .A1(n4894), .A2(n6245), .B1(n6173), .B2(n4893), .ZN(n4935)
         );
  NAND3_X1 U6034 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n5168), .ZN(n6248) );
  NOR2_X1 U6035 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6248), .ZN(n4899)
         );
  OAI22_X1 U6036 ( .A1(n6393), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n6490), .B2(n4899), .ZN(n4895) );
  INV_X1 U6037 ( .A(n4895), .ZN(n4896) );
  OAI211_X1 U6038 ( .C1(n4898), .C2(n6245), .A(n4897), .B(n4896), .ZN(n4928)
         );
  NAND2_X1 U6039 ( .A1(n4928), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4903)
         );
  INV_X1 U6040 ( .A(n4899), .ZN(n4929) );
  OAI22_X1 U6041 ( .A1(n4900), .A2(n4929), .B1(n6334), .B2(n6265), .ZN(n4901)
         );
  AOI21_X1 U6042 ( .B1(n6331), .B2(n4932), .A(n4901), .ZN(n4902) );
  OAI211_X1 U6043 ( .C1(n4935), .C2(n5032), .A(n4903), .B(n4902), .ZN(U3106)
         );
  NAND2_X1 U6044 ( .A1(n4928), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4907)
         );
  OAI22_X1 U6045 ( .A1(n4904), .A2(n4929), .B1(n6328), .B2(n6265), .ZN(n4905)
         );
  AOI21_X1 U6046 ( .B1(n6325), .B2(n4932), .A(n4905), .ZN(n4906) );
  OAI211_X1 U6047 ( .C1(n4935), .C2(n5040), .A(n4907), .B(n4906), .ZN(U3105)
         );
  NAND2_X1 U6048 ( .A1(n4928), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4911)
         );
  OAI22_X1 U6049 ( .A1(n4908), .A2(n4929), .B1(n6322), .B2(n6265), .ZN(n4909)
         );
  AOI21_X1 U6050 ( .B1(n6319), .B2(n4932), .A(n4909), .ZN(n4910) );
  OAI211_X1 U6051 ( .C1(n4935), .C2(n5036), .A(n4911), .B(n4910), .ZN(U3104)
         );
  NAND2_X1 U6052 ( .A1(n4928), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4915)
         );
  OAI22_X1 U6053 ( .A1(n4912), .A2(n4929), .B1(n6316), .B2(n6265), .ZN(n4913)
         );
  AOI21_X1 U6054 ( .B1(n6313), .B2(n4932), .A(n4913), .ZN(n4914) );
  OAI211_X1 U6055 ( .C1(n4935), .C2(n5051), .A(n4915), .B(n4914), .ZN(U3103)
         );
  NAND2_X1 U6056 ( .A1(n4928), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4919)
         );
  OAI22_X1 U6057 ( .A1(n4916), .A2(n4929), .B1(n6298), .B2(n6265), .ZN(n4917)
         );
  AOI21_X1 U6058 ( .B1(n6295), .B2(n4932), .A(n4917), .ZN(n4918) );
  OAI211_X1 U6059 ( .C1(n4935), .C2(n5020), .A(n4919), .B(n4918), .ZN(U3100)
         );
  NAND2_X1 U6060 ( .A1(n4928), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4923)
         );
  OAI22_X1 U6061 ( .A1(n4920), .A2(n4929), .B1(n6310), .B2(n6265), .ZN(n4921)
         );
  AOI21_X1 U6062 ( .B1(n6307), .B2(n4932), .A(n4921), .ZN(n4922) );
  OAI211_X1 U6063 ( .C1(n4935), .C2(n5024), .A(n4923), .B(n4922), .ZN(U3102)
         );
  NAND2_X1 U6064 ( .A1(n4928), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4927)
         );
  OAI22_X1 U6065 ( .A1(n4924), .A2(n4929), .B1(n6345), .B2(n6265), .ZN(n4925)
         );
  AOI21_X1 U6066 ( .B1(n6340), .B2(n4932), .A(n4925), .ZN(n4926) );
  OAI211_X1 U6067 ( .C1(n4935), .C2(n5028), .A(n4927), .B(n4926), .ZN(U3107)
         );
  NAND2_X1 U6068 ( .A1(n4928), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4934)
         );
  OAI22_X1 U6069 ( .A1(n4930), .A2(n4929), .B1(n6304), .B2(n6265), .ZN(n4931)
         );
  AOI21_X1 U6070 ( .B1(n6301), .B2(n4932), .A(n4931), .ZN(n4933) );
  OAI211_X1 U6071 ( .C1(n4935), .C2(n5044), .A(n4934), .B(n4933), .ZN(U3101)
         );
  AOI21_X1 U6072 ( .B1(n4937), .B2(n4936), .A(n4964), .ZN(n5057) );
  INV_X1 U6073 ( .A(n5057), .ZN(n4939) );
  INV_X1 U6074 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4938) );
  OAI222_X1 U6075 ( .A1(n4939), .A2(n5958), .B1(n5963), .B2(n4938), .C1(n5959), 
        .C2(n5076), .ZN(U2845) );
  INV_X1 U6076 ( .A(n4940), .ZN(n4942) );
  INV_X1 U6077 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6059) );
  INV_X1 U6078 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U6079 ( .A1(n4947), .A2(n4943), .ZN(n5093) );
  INV_X1 U6080 ( .A(n5079), .ZN(n4941) );
  NAND2_X1 U6081 ( .A1(n4942), .A2(n2964), .ZN(n5119) );
  NOR2_X1 U6082 ( .A1(n4944), .A2(n4943), .ZN(n5095) );
  INV_X1 U6083 ( .A(n5095), .ZN(n4946) );
  NAND2_X1 U6084 ( .A1(n5737), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5091) );
  INV_X1 U6085 ( .A(n5737), .ZN(n4947) );
  XNOR2_X1 U6086 ( .A(n4947), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5082)
         );
  NAND2_X1 U6087 ( .A1(n5737), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5113) );
  AND2_X1 U6088 ( .A1(n5115), .A2(n5113), .ZN(n4948) );
  NAND2_X1 U6089 ( .A1(n5119), .A2(n4948), .ZN(n4950) );
  INV_X1 U6090 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U6091 ( .A1(n5517), .A2(n5783), .ZN(n5053) );
  INV_X1 U6092 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6560) );
  NAND2_X1 U6093 ( .A1(n5517), .A2(n6560), .ZN(n4949) );
  NAND2_X1 U6094 ( .A1(n4950), .A2(n5116), .ZN(n4952) );
  INV_X1 U6095 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5120) );
  XNOR2_X1 U6096 ( .A(n5517), .B(n5120), .ZN(n4951) );
  XNOR2_X1 U6097 ( .A(n4952), .B(n4951), .ZN(n5149) );
  NOR2_X1 U6098 ( .A1(n4954), .A2(n4953), .ZN(n4956) );
  NAND2_X1 U6099 ( .A1(n4956), .A2(n4955), .ZN(n5289) );
  NOR2_X1 U6100 ( .A1(n5595), .A2(n5289), .ZN(n5065) );
  NAND2_X1 U6101 ( .A1(n4957), .A2(n4956), .ZN(n5282) );
  NOR2_X1 U6102 ( .A1(n5282), .A2(n4958), .ZN(n5103) );
  NAND2_X1 U6103 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5063) );
  NOR2_X1 U6104 ( .A1(n5783), .A2(n5063), .ZN(n5059) );
  NAND2_X1 U6105 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5059), .ZN(n5125) );
  NOR2_X1 U6106 ( .A1(n5310), .A2(n5125), .ZN(n4961) );
  INV_X1 U6107 ( .A(n5595), .ZN(n6096) );
  INV_X1 U6108 ( .A(n5282), .ZN(n5774) );
  OAI21_X1 U6109 ( .B1(n5284), .B2(n5774), .A(n5285), .ZN(n4959) );
  AOI21_X1 U6110 ( .B1(n6096), .B2(n5289), .A(n4959), .ZN(n6060) );
  AOI22_X1 U6111 ( .A1(n4961), .A2(n5120), .B1(n5125), .B2(n6106), .ZN(n4960)
         );
  NAND2_X1 U6112 ( .A1(n6060), .A2(n4960), .ZN(n5130) );
  OAI21_X1 U6113 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n4961), .A(n5130), 
        .ZN(n4967) );
  NOR2_X1 U6114 ( .A1(n4964), .A2(n4963), .ZN(n4965) );
  OR2_X1 U6115 ( .A1(n4962), .A2(n4965), .ZN(n5957) );
  INV_X1 U6116 ( .A(n5957), .ZN(n5832) );
  AND2_X1 U6117 ( .A1(n6107), .A2(REIP_REG_15__SCAN_IN), .ZN(n5143) );
  AOI21_X1 U6118 ( .B1(n5832), .B2(n6109), .A(n5143), .ZN(n4966) );
  OAI211_X1 U6119 ( .C1(n5149), .C2(n6084), .A(n4967), .B(n4966), .ZN(U3003)
         );
  INV_X1 U6120 ( .A(n4968), .ZN(n4969) );
  OAI22_X1 U6121 ( .A1(n4969), .A2(REIP_REG_14__SCAN_IN), .B1(n5071), .B2(
        n5944), .ZN(n4974) );
  INV_X1 U6122 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4972) );
  AND2_X1 U6123 ( .A1(n5941), .A2(n4970), .ZN(n5836) );
  AOI22_X1 U6124 ( .A1(EBX_REG_14__SCAN_IN), .A2(n5946), .B1(
        REIP_REG_14__SCAN_IN), .B2(n5836), .ZN(n4971) );
  OAI211_X1 U6125 ( .C1(n5945), .C2(n4972), .A(n4971), .B(n4850), .ZN(n4973)
         );
  AOI211_X1 U6126 ( .C1(n5057), .C2(n5943), .A(n4974), .B(n4973), .ZN(n4975)
         );
  OAI21_X1 U6127 ( .B1(n5076), .B2(n5893), .A(n4975), .ZN(U2813) );
  NAND2_X1 U6128 ( .A1(n5900), .A2(n5846), .ZN(n4978) );
  INV_X1 U6129 ( .A(n4976), .ZN(n4977) );
  OAI22_X1 U6130 ( .A1(n4978), .A2(n4977), .B1(n4999), .B2(n5944), .ZN(n4982)
         );
  INV_X1 U6131 ( .A(EBX_REG_11__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U6132 ( .A1(n5321), .A2(n4978), .ZN(n5856) );
  AOI22_X1 U6133 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n5901), .B1(
        REIP_REG_11__SCAN_IN), .B2(n5856), .ZN(n4979) );
  OAI211_X1 U6134 ( .C1(n5886), .C2(n4980), .A(n4979), .B(n4850), .ZN(n4981)
         );
  AOI211_X1 U6135 ( .C1(n6054), .C2(n5943), .A(n4982), .B(n4981), .ZN(n4983)
         );
  OAI21_X1 U6136 ( .B1(n5893), .B2(n5003), .A(n4983), .ZN(U2816) );
  NAND2_X1 U6137 ( .A1(n4984), .A2(n3348), .ZN(n4985) );
  OR2_X1 U6138 ( .A1(n5918), .A2(REIP_REG_1__SCAN_IN), .ZN(n5322) );
  AOI22_X1 U6139 ( .A1(n5901), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5913), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4986) );
  OAI211_X1 U6140 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n5944), .A(n5322), 
        .B(n4986), .ZN(n4990) );
  NOR2_X1 U6141 ( .A1(n6523), .A2(n4987), .ZN(n5947) );
  INV_X1 U6142 ( .A(n5947), .ZN(n5932) );
  INV_X1 U6143 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4988) );
  OAI22_X1 U6144 ( .A1(n5618), .A2(n5932), .B1(n5886), .B2(n4988), .ZN(n4989)
         );
  AOI211_X1 U6145 ( .C1(n5943), .C2(n4991), .A(n4990), .B(n4989), .ZN(n4992)
         );
  OAI21_X1 U6146 ( .B1(n5951), .B2(n4993), .A(n4992), .ZN(U2826) );
  OR2_X1 U6147 ( .A1(n4995), .A2(n4994), .ZN(n5078) );
  NAND2_X1 U6148 ( .A1(n5078), .A2(n4996), .ZN(n5090) );
  NAND2_X1 U6149 ( .A1(n5091), .A2(n5089), .ZN(n4997) );
  XNOR2_X1 U6150 ( .A(n5090), .B(n4997), .ZN(n6056) );
  NAND2_X1 U6151 ( .A1(n6056), .A2(n6034), .ZN(n5002) );
  INV_X1 U6152 ( .A(REIP_REG_11__SCAN_IN), .ZN(n4998) );
  NOR2_X1 U6153 ( .A1(n4850), .A2(n4998), .ZN(n6053) );
  NOR2_X1 U6154 ( .A1(n6040), .A2(n4999), .ZN(n5000) );
  AOI211_X1 U6155 ( .C1(n6048), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6053), 
        .B(n5000), .ZN(n5001) );
  OAI211_X1 U6156 ( .C1(n6051), .C2(n5003), .A(n5002), .B(n5001), .ZN(U2975)
         );
  AOI21_X1 U6157 ( .B1(n6172), .B2(n5004), .A(n6284), .ZN(n5015) );
  OR2_X1 U6158 ( .A1(n5005), .A2(n6206), .ZN(n5007) );
  NOR2_X1 U6159 ( .A1(n5169), .A2(n5013), .ZN(n5046) );
  INV_X1 U6160 ( .A(n5046), .ZN(n5006) );
  NAND2_X1 U6161 ( .A1(n5007), .A2(n5006), .ZN(n5012) );
  INV_X1 U6162 ( .A(n5013), .ZN(n5008) );
  AOI22_X1 U6163 ( .A1(n5015), .A2(n5012), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5008), .ZN(n5052) );
  OR2_X1 U6164 ( .A1(n5010), .A2(n5009), .ZN(n6177) );
  INV_X1 U6165 ( .A(n5011), .ZN(n5048) );
  INV_X1 U6166 ( .A(n5012), .ZN(n5014) );
  AOI22_X1 U6167 ( .A1(n5015), .A2(n5014), .B1(n5013), .B2(n6284), .ZN(n5016)
         );
  NAND2_X1 U6168 ( .A1(n6293), .A2(n5016), .ZN(n5045) );
  AOI22_X1 U6169 ( .A1(n6285), .A2(n5046), .B1(INSTQUEUE_REG_5__0__SCAN_IN), 
        .B2(n5045), .ZN(n5017) );
  OAI21_X1 U6170 ( .B1(n6218), .B2(n5048), .A(n5017), .ZN(n5018) );
  AOI21_X1 U6171 ( .B1(n6205), .B2(n6200), .A(n5018), .ZN(n5019) );
  OAI21_X1 U6172 ( .B1(n5052), .B2(n5020), .A(n5019), .ZN(U3060) );
  AOI22_X1 U6173 ( .A1(n6305), .A2(n5046), .B1(INSTQUEUE_REG_5__2__SCAN_IN), 
        .B2(n5045), .ZN(n5021) );
  OAI21_X1 U6174 ( .B1(n6260), .B2(n5048), .A(n5021), .ZN(n5022) );
  AOI21_X1 U6175 ( .B1(n6257), .B2(n6200), .A(n5022), .ZN(n5023) );
  OAI21_X1 U6176 ( .B1(n5052), .B2(n5024), .A(n5023), .ZN(U3062) );
  AOI22_X1 U6177 ( .A1(n6335), .A2(n5046), .B1(INSTQUEUE_REG_5__7__SCAN_IN), 
        .B2(n5045), .ZN(n5025) );
  OAI21_X1 U6178 ( .B1(n6241), .B2(n5048), .A(n5025), .ZN(n5026) );
  AOI21_X1 U6179 ( .B1(n6234), .B2(n6200), .A(n5026), .ZN(n5027) );
  OAI21_X1 U6180 ( .B1(n5052), .B2(n5028), .A(n5027), .ZN(U3067) );
  AOI22_X1 U6181 ( .A1(n6329), .A2(n5046), .B1(INSTQUEUE_REG_5__6__SCAN_IN), 
        .B2(n5045), .ZN(n5029) );
  OAI21_X1 U6182 ( .B1(n6149), .B2(n5048), .A(n5029), .ZN(n5030) );
  AOI21_X1 U6183 ( .B1(n6146), .B2(n6200), .A(n5030), .ZN(n5031) );
  OAI21_X1 U6184 ( .B1(n5052), .B2(n5032), .A(n5031), .ZN(U3066) );
  AOI22_X1 U6185 ( .A1(n6317), .A2(n5046), .B1(INSTQUEUE_REG_5__4__SCAN_IN), 
        .B2(n5045), .ZN(n5033) );
  OAI21_X1 U6186 ( .B1(n6141), .B2(n5048), .A(n5033), .ZN(n5034) );
  AOI21_X1 U6187 ( .B1(n6138), .B2(n6200), .A(n5034), .ZN(n5035) );
  OAI21_X1 U6188 ( .B1(n5052), .B2(n5036), .A(n5035), .ZN(U3064) );
  AOI22_X1 U6189 ( .A1(n6323), .A2(n5046), .B1(INSTQUEUE_REG_5__5__SCAN_IN), 
        .B2(n5045), .ZN(n5037) );
  OAI21_X1 U6190 ( .B1(n6145), .B2(n5048), .A(n5037), .ZN(n5038) );
  AOI21_X1 U6191 ( .B1(n6142), .B2(n6200), .A(n5038), .ZN(n5039) );
  OAI21_X1 U6192 ( .B1(n5052), .B2(n5040), .A(n5039), .ZN(U3065) );
  AOI22_X1 U6193 ( .A1(n6299), .A2(n5046), .B1(INSTQUEUE_REG_5__1__SCAN_IN), 
        .B2(n5045), .ZN(n5041) );
  OAI21_X1 U6194 ( .B1(n6256), .B2(n5048), .A(n5041), .ZN(n5042) );
  AOI21_X1 U6195 ( .B1(n6253), .B2(n6200), .A(n5042), .ZN(n5043) );
  OAI21_X1 U6196 ( .B1(n5052), .B2(n5044), .A(n5043), .ZN(U3061) );
  AOI22_X1 U6197 ( .A1(n6311), .A2(n5046), .B1(INSTQUEUE_REG_5__3__SCAN_IN), 
        .B2(n5045), .ZN(n5047) );
  OAI21_X1 U6198 ( .B1(n6266), .B2(n5048), .A(n5047), .ZN(n5049) );
  AOI21_X1 U6199 ( .B1(n6262), .B2(n6200), .A(n5049), .ZN(n5050) );
  OAI21_X1 U6200 ( .B1(n5052), .B2(n5051), .A(n5050), .ZN(U3063) );
  NAND2_X1 U6201 ( .A1(n5119), .A2(n5115), .ZN(n5081) );
  NAND2_X1 U6202 ( .A1(n5081), .A2(n5053), .ZN(n5055) );
  XNOR2_X1 U6203 ( .A(n5517), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5054)
         );
  XNOR2_X1 U6204 ( .A(n5055), .B(n5054), .ZN(n5070) );
  INV_X1 U6205 ( .A(n5070), .ZN(n5069) );
  NOR2_X1 U6206 ( .A1(n4850), .A2(n6451), .ZN(n5073) );
  INV_X1 U6207 ( .A(n5310), .ZN(n6055) );
  AND3_X1 U6208 ( .A1(n6560), .A2(n6055), .A3(n5059), .ZN(n5056) );
  AOI211_X1 U6209 ( .C1(n6109), .C2(n5057), .A(n5073), .B(n5056), .ZN(n5068)
         );
  OAI21_X1 U6210 ( .B1(n5059), .B2(n5058), .A(n6060), .ZN(n5060) );
  AOI21_X1 U6211 ( .B1(n5061), .B2(n5063), .A(n5060), .ZN(n5784) );
  NOR3_X1 U6212 ( .A1(n6498), .A2(n5062), .A3(n5282), .ZN(n5064) );
  NOR2_X1 U6213 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5063), .ZN(n5775)
         );
  OAI21_X1 U6214 ( .B1(n5065), .B2(n5064), .A(n5775), .ZN(n5781) );
  AOI21_X1 U6215 ( .B1(n5784), .B2(n5781), .A(n6560), .ZN(n5066) );
  INV_X1 U6216 ( .A(n5066), .ZN(n5067) );
  OAI211_X1 U6217 ( .C1(n5069), .C2(n6084), .A(n5068), .B(n5067), .ZN(U3004)
         );
  NAND2_X1 U6218 ( .A1(n5070), .A2(n6034), .ZN(n5075) );
  NOR2_X1 U6219 ( .A1(n6040), .A2(n5071), .ZN(n5072) );
  AOI211_X1 U6220 ( .C1(n6048), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5073), 
        .B(n5072), .ZN(n5074) );
  OAI211_X1 U6221 ( .C1(n6287), .C2(n5076), .A(n5075), .B(n5074), .ZN(U2972)
         );
  NAND2_X1 U6222 ( .A1(n5078), .A2(n5077), .ZN(n5080) );
  NAND2_X1 U6223 ( .A1(n5080), .A2(n5079), .ZN(n5083) );
  OAI21_X1 U6224 ( .B1(n5083), .B2(n5082), .A(n5081), .ZN(n5780) );
  NAND2_X1 U6225 ( .A1(n5780), .A2(n6034), .ZN(n5088) );
  INV_X1 U6226 ( .A(n5084), .ZN(n5844) );
  NAND2_X1 U6227 ( .A1(n5516), .A2(REIP_REG_13__SCAN_IN), .ZN(n5777) );
  OAI21_X1 U6228 ( .B1(n5523), .B2(n5085), .A(n5777), .ZN(n5086) );
  AOI21_X1 U6229 ( .B1(n5525), .B2(n5844), .A(n5086), .ZN(n5087) );
  OAI211_X1 U6230 ( .C1(n5843), .C2(n6051), .A(n5088), .B(n5087), .ZN(U2973)
         );
  NAND2_X1 U6231 ( .A1(n5090), .A2(n5089), .ZN(n5092) );
  NAND2_X1 U6232 ( .A1(n5092), .A2(n5091), .ZN(n5097) );
  INV_X1 U6233 ( .A(n5093), .ZN(n5094) );
  NOR2_X1 U6234 ( .A1(n5095), .A2(n5094), .ZN(n5096) );
  XNOR2_X1 U6235 ( .A(n5097), .B(n5096), .ZN(n5111) );
  NAND2_X1 U6236 ( .A1(n6099), .A2(REIP_REG_12__SCAN_IN), .ZN(n5105) );
  OAI21_X1 U6237 ( .B1(n5523), .B2(n5098), .A(n5105), .ZN(n5100) );
  NOR2_X1 U6238 ( .A1(n5858), .A2(n6287), .ZN(n5099) );
  AOI211_X1 U6239 ( .C1(n5525), .C2(n5101), .A(n5100), .B(n5099), .ZN(n5102)
         );
  OAI21_X1 U6240 ( .B1(n5111), .B2(n6042), .A(n5102), .ZN(U2974) );
  OAI21_X1 U6241 ( .B1(n6096), .B2(n5103), .A(n6059), .ZN(n5104) );
  AOI21_X1 U6242 ( .B1(n6060), .B2(n5104), .A(n4943), .ZN(n5109) );
  INV_X1 U6243 ( .A(n5105), .ZN(n5108) );
  NOR2_X1 U6244 ( .A1(n6082), .A2(n5854), .ZN(n5107) );
  NOR3_X1 U6245 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5310), .A3(n6059), 
        .ZN(n5106) );
  NOR4_X1 U6246 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n5110)
         );
  OAI21_X1 U6247 ( .B1(n5111), .B2(n6084), .A(n5110), .ZN(U3006) );
  NAND2_X1 U6248 ( .A1(n5737), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5112) );
  AND2_X1 U6249 ( .A1(n5113), .A2(n5112), .ZN(n5114) );
  NAND2_X1 U6250 ( .A1(n4947), .A2(n5120), .ZN(n5121) );
  NAND2_X1 U6251 ( .A1(n5519), .A2(n5121), .ZN(n5267) );
  XNOR2_X1 U6252 ( .A(n5517), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5122)
         );
  XNOR2_X1 U6253 ( .A(n5267), .B(n5122), .ZN(n5150) );
  INV_X1 U6254 ( .A(n5150), .ZN(n5132) );
  OR2_X1 U6255 ( .A1(n4962), .A2(n5123), .ZN(n5124) );
  NAND2_X1 U6256 ( .A1(n5767), .A2(n5124), .ZN(n5200) );
  NOR2_X1 U6257 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5310), .ZN(n5127)
         );
  NOR2_X1 U6258 ( .A1(n5120), .A2(n5125), .ZN(n5281) );
  INV_X1 U6259 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5126) );
  NOR2_X1 U6260 ( .A1(n4850), .A2(n5126), .ZN(n5154) );
  AOI21_X1 U6261 ( .B1(n5127), .B2(n5281), .A(n5154), .ZN(n5128) );
  OAI21_X1 U6262 ( .B1(n5200), .B2(n6082), .A(n5128), .ZN(n5129) );
  AOI21_X1 U6263 ( .B1(n5130), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5129), 
        .ZN(n5131) );
  OAI21_X1 U6264 ( .B1(n5132), .B2(n6084), .A(n5131), .ZN(U3002) );
  NAND2_X1 U6265 ( .A1(n5161), .A2(n5157), .ZN(n5744) );
  OAI21_X1 U6266 ( .B1(n5161), .B2(n5157), .A(n5744), .ZN(n5198) );
  AOI22_X1 U6267 ( .A1(n5968), .A2(DATAI_16_), .B1(n5970), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5135) );
  NAND2_X1 U6268 ( .A1(n5971), .A2(DATAI_0_), .ZN(n5134) );
  OAI211_X1 U6269 ( .C1(n5198), .C2(n5695), .A(n5135), .B(n5134), .ZN(U2875)
         );
  NOR2_X1 U6270 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5138), .ZN(n5835) );
  AOI22_X1 U6271 ( .A1(EBX_REG_16__SCAN_IN), .A2(n5946), .B1(n5151), .B2(n5907), .ZN(n5136) );
  OAI211_X1 U6272 ( .C1(n5945), .C2(n3788), .A(n5136), .B(n4850), .ZN(n5137)
         );
  AOI221_X1 U6273 ( .B1(n5836), .B2(REIP_REG_16__SCAN_IN), .C1(n5835), .C2(
        REIP_REG_16__SCAN_IN), .A(n5137), .ZN(n5141) );
  INV_X1 U6274 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6453) );
  NOR2_X1 U6275 ( .A1(n5138), .A2(n6453), .ZN(n5824) );
  INV_X1 U6276 ( .A(n5200), .ZN(n5139) );
  AOI22_X1 U6277 ( .A1(n5824), .A2(n5126), .B1(n5943), .B2(n5139), .ZN(n5140)
         );
  OAI211_X1 U6278 ( .C1(n5198), .C2(n5893), .A(n5141), .B(n5140), .ZN(U2811)
         );
  AND2_X1 U6279 ( .A1(n6048), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5142)
         );
  AOI211_X1 U6280 ( .C1(n5525), .C2(n5837), .A(n5143), .B(n5142), .ZN(n5148)
         );
  AND2_X1 U6281 ( .A1(n5145), .A2(n5144), .ZN(n5146) );
  OR2_X1 U6282 ( .A1(n5146), .A2(n5161), .ZN(n5960) );
  NAND2_X1 U6283 ( .A1(n5976), .A2(n6036), .ZN(n5147) );
  OAI211_X1 U6284 ( .C1(n5149), .C2(n6042), .A(n5148), .B(n5147), .ZN(U2971)
         );
  NAND2_X1 U6285 ( .A1(n5150), .A2(n6034), .ZN(n5156) );
  INV_X1 U6286 ( .A(n5151), .ZN(n5152) );
  NOR2_X1 U6287 ( .A1(n6040), .A2(n5152), .ZN(n5153) );
  AOI211_X1 U6288 ( .C1(n6048), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5154), 
        .B(n5153), .ZN(n5155) );
  OAI211_X1 U6289 ( .C1(n6051), .C2(n5198), .A(n5156), .B(n5155), .ZN(U2970)
         );
  AND2_X1 U6290 ( .A1(n5161), .A2(n5157), .ZN(n5159) );
  NAND2_X1 U6291 ( .A1(n5161), .A2(n5160), .ZN(n5209) );
  OAI21_X1 U6292 ( .B1(n5236), .B2(n5162), .A(n5209), .ZN(n5686) );
  MUX2_X1 U6293 ( .A(n3024), .B(n5239), .S(n5163), .Z(n5165) );
  XNOR2_X1 U6294 ( .A(n5165), .B(n5164), .ZN(n5687) );
  AOI22_X1 U6295 ( .A1(n5687), .A2(n5953), .B1(EBX_REG_20__SCAN_IN), .B2(n5319), .ZN(n5166) );
  OAI21_X1 U6296 ( .B1(n5686), .B2(n5959), .A(n5166), .ZN(U2839) );
  OR2_X1 U6297 ( .A1(n6121), .A2(n5167), .ZN(n6126) );
  INV_X1 U6298 ( .A(n6126), .ZN(n5170) );
  NAND3_X1 U6299 ( .A1(n6382), .A2(n5168), .A3(n6374), .ZN(n6122) );
  NOR2_X1 U6300 ( .A1(n5169), .A2(n6122), .ZN(n5194) );
  AOI21_X1 U6301 ( .B1(n5170), .B2(n6365), .A(n5194), .ZN(n5175) );
  AOI21_X1 U6302 ( .B1(n5171), .B2(STATEBS16_REG_SCAN_IN), .A(n6284), .ZN(
        n5173) );
  AOI22_X1 U6303 ( .A1(n5175), .A2(n5173), .B1(n6284), .B2(n6122), .ZN(n5172)
         );
  NAND2_X1 U6304 ( .A1(n6293), .A2(n5172), .ZN(n5193) );
  INV_X1 U6305 ( .A(n5173), .ZN(n5174) );
  OAI22_X1 U6306 ( .A1(n5175), .A2(n5174), .B1(n6393), .B2(n6122), .ZN(n5192)
         );
  AOI22_X1 U6307 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5193), .B1(n6338), 
        .B2(n5192), .ZN(n5179) );
  NOR2_X2 U6308 ( .A1(n5177), .A2(n5176), .ZN(n6152) );
  AOI22_X1 U6309 ( .A1(n6335), .A2(n5194), .B1(n6340), .B2(n6152), .ZN(n5178)
         );
  OAI211_X1 U6310 ( .C1(n6345), .C2(n5197), .A(n5179), .B(n5178), .ZN(U3035)
         );
  AOI22_X1 U6311 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5193), .B1(n6324), 
        .B2(n5192), .ZN(n5181) );
  AOI22_X1 U6312 ( .A1(n6323), .A2(n5194), .B1(n6325), .B2(n6152), .ZN(n5180)
         );
  OAI211_X1 U6313 ( .C1(n6328), .C2(n5197), .A(n5181), .B(n5180), .ZN(U3033)
         );
  AOI22_X1 U6314 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5193), .B1(n6318), 
        .B2(n5192), .ZN(n5183) );
  AOI22_X1 U6315 ( .A1(n6317), .A2(n5194), .B1(n6319), .B2(n6152), .ZN(n5182)
         );
  OAI211_X1 U6316 ( .C1(n6322), .C2(n5197), .A(n5183), .B(n5182), .ZN(U3032)
         );
  AOI22_X1 U6317 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5193), .B1(n6330), 
        .B2(n5192), .ZN(n5185) );
  AOI22_X1 U6318 ( .A1(n6329), .A2(n5194), .B1(n6331), .B2(n6152), .ZN(n5184)
         );
  OAI211_X1 U6319 ( .C1(n6334), .C2(n5197), .A(n5185), .B(n5184), .ZN(U3034)
         );
  AOI22_X1 U6320 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5193), .B1(n6306), 
        .B2(n5192), .ZN(n5187) );
  AOI22_X1 U6321 ( .A1(n6305), .A2(n5194), .B1(n6307), .B2(n6152), .ZN(n5186)
         );
  OAI211_X1 U6322 ( .C1(n6310), .C2(n5197), .A(n5187), .B(n5186), .ZN(U3030)
         );
  AOI22_X1 U6323 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5193), .B1(n6300), 
        .B2(n5192), .ZN(n5189) );
  AOI22_X1 U6324 ( .A1(n6299), .A2(n5194), .B1(n6301), .B2(n6152), .ZN(n5188)
         );
  OAI211_X1 U6325 ( .C1(n6304), .C2(n5197), .A(n5189), .B(n5188), .ZN(U3029)
         );
  AOI22_X1 U6326 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5193), .B1(n6312), 
        .B2(n5192), .ZN(n5191) );
  AOI22_X1 U6327 ( .A1(n6311), .A2(n5194), .B1(n6313), .B2(n6152), .ZN(n5190)
         );
  OAI211_X1 U6328 ( .C1(n6316), .C2(n5197), .A(n5191), .B(n5190), .ZN(U3031)
         );
  AOI22_X1 U6329 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5193), .B1(n6286), 
        .B2(n5192), .ZN(n5196) );
  AOI22_X1 U6330 ( .A1(n6285), .A2(n5194), .B1(n6295), .B2(n6152), .ZN(n5195)
         );
  OAI211_X1 U6331 ( .C1(n6298), .C2(n5197), .A(n5196), .B(n5195), .ZN(U3028)
         );
  INV_X1 U6332 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5199) );
  OAI222_X1 U6333 ( .A1(n5200), .A2(n5958), .B1(n5963), .B2(n5199), .C1(n5959), 
        .C2(n5198), .ZN(U2843) );
  AND2_X1 U6334 ( .A1(n5207), .A2(n5202), .ZN(n5204) );
  OR2_X1 U6335 ( .A1(n5204), .A2(n5217), .ZN(n5670) );
  INV_X1 U6336 ( .A(n5220), .ZN(n5205) );
  XNOR2_X1 U6337 ( .A(n5221), .B(n5205), .ZN(n5671) );
  AOI22_X1 U6338 ( .A1(n5671), .A2(n5953), .B1(EBX_REG_22__SCAN_IN), .B2(n5319), .ZN(n5206) );
  OAI21_X1 U6339 ( .B1(n5670), .B2(n5959), .A(n5206), .ZN(U2837) );
  INV_X1 U6340 ( .A(n5207), .ZN(n5208) );
  AOI21_X1 U6341 ( .B1(n5210), .B2(n5209), .A(n5208), .ZN(n5713) );
  INV_X1 U6342 ( .A(n5713), .ZN(n5214) );
  INV_X1 U6343 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5213) );
  OAI21_X1 U6344 ( .B1(n5212), .B2(n5211), .A(n5221), .ZN(n5681) );
  OAI222_X1 U6345 ( .A1(n5214), .A2(n5959), .B1(n5963), .B2(n5213), .C1(n5681), 
        .C2(n5958), .ZN(U2838) );
  NOR2_X1 U6346 ( .A1(n5217), .A2(n5216), .ZN(n5218) );
  OR2_X1 U6347 ( .A1(n5233), .A2(n5218), .ZN(n5490) );
  OAI21_X1 U6348 ( .B1(n5221), .B2(n5220), .A(n5219), .ZN(n5222) );
  AND2_X1 U6349 ( .A1(n5222), .A2(n5394), .ZN(n5574) );
  AOI22_X1 U6350 ( .A1(n5574), .A2(n5953), .B1(n5319), .B2(EBX_REG_23__SCAN_IN), .ZN(n5223) );
  OAI21_X1 U6351 ( .B1(n5490), .B2(n5959), .A(n5223), .ZN(U2836) );
  OAI21_X1 U6352 ( .B1(n5685), .B2(n5672), .A(n6569), .ZN(n5230) );
  INV_X1 U6353 ( .A(n5941), .ZN(n5243) );
  NOR2_X1 U6354 ( .A1(n5243), .A2(n5224), .ZN(n5660) );
  INV_X1 U6355 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5225) );
  OAI22_X1 U6356 ( .A1(n5225), .A2(n5945), .B1(n5492), .B2(n5944), .ZN(n5229)
         );
  INV_X1 U6357 ( .A(n5574), .ZN(n5227) );
  INV_X1 U6358 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5226) );
  OAI22_X1 U6359 ( .A1(n5227), .A2(n5933), .B1(n5886), .B2(n5226), .ZN(n5228)
         );
  AOI211_X1 U6360 ( .C1(n5230), .C2(n5660), .A(n5229), .B(n5228), .ZN(n5231)
         );
  OAI21_X1 U6361 ( .B1(n5490), .B2(n5893), .A(n5231), .ZN(U2804) );
  OAI21_X1 U6362 ( .B1(n5233), .B2(n5232), .A(n5390), .ZN(n5661) );
  XOR2_X1 U6363 ( .A(n5396), .B(n5394), .Z(n5662) );
  INV_X1 U6364 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5234) );
  OAI222_X1 U6365 ( .A1(n5959), .A2(n5661), .B1(n5958), .B2(n5662), .C1(n5234), 
        .C2(n5963), .ZN(U2835) );
  MUX2_X1 U6366 ( .A(n5239), .B(n5238), .S(n5237), .Z(n5431) );
  NOR2_X1 U6367 ( .A1(n5769), .A2(n5431), .ZN(n5432) );
  XNOR2_X1 U6368 ( .A(n5432), .B(n5240), .ZN(n5758) );
  AOI22_X1 U6369 ( .A1(n5758), .A2(n5953), .B1(EBX_REG_19__SCAN_IN), .B2(n5319), .ZN(n5241) );
  OAI21_X1 U6370 ( .B1(n5719), .B2(n5959), .A(n5241), .ZN(U2840) );
  NOR2_X1 U6371 ( .A1(n5243), .A2(n5242), .ZN(n5825) );
  AOI22_X1 U6372 ( .A1(EBX_REG_19__SCAN_IN), .A2(n5946), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n5901), .ZN(n5244) );
  INV_X1 U6373 ( .A(n5244), .ZN(n5245) );
  AOI211_X1 U6374 ( .C1(REIP_REG_19__SCAN_IN), .C2(n5825), .A(n6107), .B(n5245), .ZN(n5248) );
  NAND2_X1 U6375 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5246) );
  OAI211_X1 U6376 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5816), .B(n5246), .ZN(n5247) );
  OAI211_X1 U6377 ( .C1(n5944), .C2(n5734), .A(n5248), .B(n5247), .ZN(n5249)
         );
  AOI21_X1 U6378 ( .B1(n5943), .B2(n5758), .A(n5249), .ZN(n5250) );
  OAI21_X1 U6379 ( .B1(n5719), .B2(n5893), .A(n5250), .ZN(U2808) );
  AOI21_X1 U6380 ( .B1(n5254), .B2(n5251), .A(n5262), .ZN(n5264) );
  INV_X1 U6381 ( .A(n5252), .ZN(n5260) );
  INV_X1 U6382 ( .A(n5253), .ZN(n5257) );
  NAND3_X1 U6383 ( .A1(n5255), .A2(n5254), .A3(n5263), .ZN(n5256) );
  OAI21_X1 U6384 ( .B1(n5258), .B2(n5257), .A(n5256), .ZN(n5259) );
  AOI21_X1 U6385 ( .B1(n5260), .B2(n5787), .A(n5259), .ZN(n5261) );
  OAI22_X1 U6386 ( .A1(n5264), .A2(n5263), .B1(n5262), .B2(n5261), .ZN(U3459)
         );
  OAI22_X1 U6387 ( .A1(n5534), .A2(n5958), .B1(n5265), .B2(n5963), .ZN(U2828)
         );
  INV_X1 U6388 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5735) );
  AND2_X1 U6389 ( .A1(n5517), .A2(n5735), .ZN(n5266) );
  OR2_X2 U6390 ( .A1(n5267), .A2(n5266), .ZN(n5736) );
  INV_X1 U6391 ( .A(n5736), .ZN(n5268) );
  NAND2_X1 U6392 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U6393 ( .A1(n5268), .A2(n2962), .ZN(n5477) );
  INV_X1 U6394 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U6395 ( .A1(n5599), .A2(n5735), .ZN(n5518) );
  OAI21_X1 U6396 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5518), .A(n5737), 
        .ZN(n5269) );
  NAND2_X1 U6397 ( .A1(n5477), .A2(n5269), .ZN(n5271) );
  INV_X1 U6398 ( .A(n5271), .ZN(n5270) );
  NAND2_X1 U6399 ( .A1(n5270), .A2(n5762), .ZN(n5729) );
  NOR2_X1 U6400 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5581) );
  INV_X1 U6401 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5562) );
  INV_X1 U6402 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5569) );
  NAND4_X1 U6403 ( .A1(n5581), .A2(n5562), .A3(n5603), .A4(n5569), .ZN(n5274)
         );
  NAND2_X1 U6404 ( .A1(n5271), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5728) );
  AND2_X1 U6405 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5580) );
  NAND4_X1 U6406 ( .A1(n5580), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_24__SCAN_IN), .A4(INSTADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n5272) );
  OAI21_X2 U6407 ( .B1(n5728), .B2(n5272), .A(n5517), .ZN(n5273) );
  OAI21_X1 U6408 ( .B1(n5729), .B2(n5274), .A(n5273), .ZN(n5457) );
  XNOR2_X1 U6409 ( .A(n5517), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5722)
         );
  INV_X1 U6410 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6411 ( .A1(n4947), .A2(n5280), .ZN(n5275) );
  INV_X1 U6412 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6413 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5542) );
  NOR2_X2 U6414 ( .A1(n5465), .A2(n5542), .ZN(n5448) );
  NOR2_X1 U6415 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5544) );
  NAND3_X1 U6416 ( .A1(n5737), .A2(n5544), .A3(n5470), .ZN(n5446) );
  INV_X1 U6417 ( .A(n5446), .ZN(n5277) );
  NAND2_X1 U6418 ( .A1(n5455), .A2(n5277), .ZN(n5332) );
  NOR2_X1 U6419 ( .A1(n5332), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5331)
         );
  AOI21_X1 U6420 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5448), .A(n5331), 
        .ZN(n5278) );
  AND2_X1 U6421 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5529) );
  NOR2_X1 U6422 ( .A1(n5280), .A2(n5470), .ZN(n5558) );
  INV_X1 U6423 ( .A(n5580), .ZN(n5294) );
  NAND2_X1 U6424 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5281), .ZN(n5309) );
  NOR2_X1 U6425 ( .A1(n5282), .A2(n5309), .ZN(n5283) );
  OR2_X1 U6426 ( .A1(n5284), .A2(n5283), .ZN(n5286) );
  NAND2_X1 U6427 ( .A1(n5286), .A2(n5285), .ZN(n5598) );
  INV_X1 U6428 ( .A(n5598), .ZN(n5293) );
  INV_X1 U6429 ( .A(n5756), .ZN(n5288) );
  AND2_X1 U6430 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6431 ( .A1(n5288), .A2(n5287), .ZN(n5311) );
  INV_X1 U6432 ( .A(n5311), .ZN(n5290) );
  NOR2_X1 U6433 ( .A1(n5309), .A2(n5289), .ZN(n5596) );
  NAND2_X1 U6434 ( .A1(n5290), .A2(n5596), .ZN(n5291) );
  NAND2_X1 U6435 ( .A1(n6106), .A2(n5291), .ZN(n5292) );
  NAND2_X1 U6436 ( .A1(n5293), .A2(n5292), .ZN(n5587) );
  AOI21_X1 U6437 ( .B1(n5294), .B2(n6106), .A(n5587), .ZN(n5570) );
  NAND2_X1 U6438 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5312) );
  OAI21_X1 U6439 ( .B1(n6100), .B2(n6096), .A(n5312), .ZN(n5295) );
  NAND2_X1 U6440 ( .A1(n5570), .A2(n5295), .ZN(n5749) );
  INV_X1 U6441 ( .A(n5749), .ZN(n5296) );
  OAI21_X1 U6442 ( .B1(n5558), .B2(n5297), .A(n5296), .ZN(n5550) );
  AOI21_X1 U6443 ( .B1(n5542), .B2(n6106), .A(n5550), .ZN(n5348) );
  OAI21_X1 U6444 ( .B1(n5529), .B2(n5297), .A(n5348), .ZN(n5533) );
  NAND2_X1 U6445 ( .A1(n5516), .A2(REIP_REG_30__SCAN_IN), .ZN(n5358) );
  INV_X1 U6446 ( .A(n5358), .ZN(n5308) );
  INV_X1 U6447 ( .A(n5302), .ZN(n5298) );
  OAI21_X1 U6448 ( .B1(n5300), .B2(n5299), .A(n5298), .ZN(n5305) );
  OAI211_X1 U6449 ( .C1(n5410), .C2(n3024), .A(n5303), .B(n5302), .ZN(n5304)
         );
  NOR2_X1 U6450 ( .A1(n5377), .A2(n6082), .ZN(n5307) );
  AOI211_X1 U6451 ( .C1(INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n5533), .A(n5308), .B(n5307), .ZN(n5316) );
  NOR2_X1 U6452 ( .A1(n5764), .A2(n5311), .ZN(n5592) );
  NAND2_X1 U6453 ( .A1(n5592), .A2(n5580), .ZN(n5571) );
  INV_X1 U6454 ( .A(n5755), .ZN(n5313) );
  NAND2_X1 U6455 ( .A1(n5313), .A2(n5558), .ZN(n5551) );
  NOR2_X1 U6456 ( .A1(n5551), .A2(n5542), .ZN(n5530) );
  INV_X1 U6457 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5314) );
  NAND3_X1 U6458 ( .A1(n5530), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5314), .ZN(n5315) );
  OAI211_X1 U6459 ( .C1(n5366), .C2(n6084), .A(n5316), .B(n5315), .ZN(U2988)
         );
  XOR2_X1 U6460 ( .A(n5318), .B(n5317), .Z(n6094) );
  AOI22_X1 U6461 ( .A1(n5953), .A2(n6094), .B1(n5319), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5320) );
  OAI21_X1 U6462 ( .B1(n6029), .B2(n5959), .A(n5320), .ZN(U2857) );
  NAND2_X1 U6463 ( .A1(n5322), .A2(n5321), .ZN(n5929) );
  AOI22_X1 U6464 ( .A1(EBX_REG_2__SCAN_IN), .A2(n5946), .B1(n5947), .B2(n5621), 
        .ZN(n5328) );
  INV_X1 U6465 ( .A(n6039), .ZN(n5323) );
  AOI22_X1 U6466 ( .A1(n5323), .A2(n5907), .B1(n5901), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6467 ( .A1(n5943), .A2(n6094), .ZN(n5326) );
  INV_X1 U6468 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U6469 ( .A1(n5928), .A2(REIP_REG_1__SCAN_IN), .ZN(n5324) );
  OR2_X1 U6470 ( .A1(n5918), .A2(n5324), .ZN(n5325) );
  NAND4_X1 U6471 ( .A1(n5328), .A2(n5327), .A3(n5326), .A4(n5325), .ZN(n5329)
         );
  AOI21_X1 U6472 ( .B1(REIP_REG_2__SCAN_IN), .B2(n5929), .A(n5329), .ZN(n5330)
         );
  OAI21_X1 U6473 ( .B1(n5951), .B2(n6029), .A(n5330), .ZN(U2825) );
  INV_X1 U6474 ( .A(n5448), .ZN(n5335) );
  INV_X1 U6475 ( .A(n5331), .ZN(n5334) );
  INV_X1 U6476 ( .A(n5332), .ZN(n5333) );
  INV_X1 U6477 ( .A(n5336), .ZN(n5355) );
  AOI21_X1 U6478 ( .B1(n5337), .B2(n5407), .A(n5357), .ZN(n5380) );
  AND2_X1 U6479 ( .A1(n6107), .A2(REIP_REG_29__SCAN_IN), .ZN(n5350) );
  AOI21_X1 U6480 ( .B1(n6048), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5350), 
        .ZN(n5338) );
  OAI21_X1 U6481 ( .B1(n6040), .B2(n5381), .A(n5338), .ZN(n5339) );
  AOI21_X1 U6482 ( .B1(n5380), .B2(n6036), .A(n5339), .ZN(n5340) );
  OAI21_X1 U6483 ( .B1(n5355), .B2(n6042), .A(n5340), .ZN(U2957) );
  NAND2_X1 U6484 ( .A1(n5342), .A2(n3024), .ZN(n5344) );
  NAND2_X1 U6485 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  NOR2_X1 U6486 ( .A1(n5410), .A2(n5345), .ZN(n5346) );
  OR2_X2 U6487 ( .A1(n5347), .A2(n5346), .ZN(n5403) );
  INV_X1 U6488 ( .A(n5403), .ZN(n5351) );
  NOR2_X1 U6489 ( .A1(n5348), .A2(n5352), .ZN(n5349) );
  AOI211_X1 U6490 ( .C1(n5351), .C2(n6109), .A(n5350), .B(n5349), .ZN(n5354)
         );
  NAND2_X1 U6491 ( .A1(n5530), .A2(n5352), .ZN(n5353) );
  OAI211_X1 U6492 ( .C1(n5355), .C2(n6084), .A(n5354), .B(n5353), .ZN(U2989)
         );
  INV_X1 U6493 ( .A(n5368), .ZN(n5362) );
  OAI21_X1 U6494 ( .B1(n5523), .B2(n5359), .A(n5358), .ZN(n5360) );
  INV_X1 U6495 ( .A(n5360), .ZN(n5361) );
  OAI21_X1 U6496 ( .B1(n5362), .B2(n6040), .A(n5361), .ZN(n5363) );
  INV_X1 U6497 ( .A(n5363), .ZN(n5364) );
  OAI21_X1 U6498 ( .B1(n5366), .B2(n6042), .A(n5365), .ZN(U2956) );
  OAI21_X1 U6499 ( .B1(n5385), .B2(n6476), .A(n5367), .ZN(n5372) );
  AOI22_X1 U6500 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n5901), .B1(n5907), 
        .B2(n5368), .ZN(n5370) );
  NAND2_X1 U6501 ( .A1(n5946), .A2(EBX_REG_30__SCAN_IN), .ZN(n5369) );
  OAI211_X1 U6502 ( .C1(n5377), .C2(n5933), .A(n5370), .B(n5369), .ZN(n5371)
         );
  AOI21_X1 U6503 ( .B1(n5373), .B2(n5372), .A(n5371), .ZN(n5374) );
  OAI21_X1 U6504 ( .B1(n5379), .B2(n5893), .A(n5374), .ZN(U2797) );
  AOI22_X1 U6505 ( .A1(n5968), .A2(DATAI_30_), .B1(n5970), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6506 ( .A1(n5971), .A2(DATAI_14_), .ZN(n5375) );
  OAI211_X1 U6507 ( .C1(n5379), .C2(n5695), .A(n5376), .B(n5375), .ZN(U2861)
         );
  INV_X1 U6508 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5378) );
  OAI222_X1 U6509 ( .A1(n5959), .A2(n5379), .B1(n5963), .B2(n5378), .C1(n5377), 
        .C2(n5958), .ZN(U2829) );
  INV_X1 U6510 ( .A(n5380), .ZN(n5442) );
  INV_X1 U6511 ( .A(n5381), .ZN(n5382) );
  AOI22_X1 U6512 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n5901), .B1(n5907), 
        .B2(n5382), .ZN(n5384) );
  NAND2_X1 U6513 ( .A1(n5946), .A2(EBX_REG_29__SCAN_IN), .ZN(n5383) );
  OAI211_X1 U6514 ( .C1(n5403), .C2(n5933), .A(n5384), .B(n5383), .ZN(n5387)
         );
  NOR2_X1 U6515 ( .A1(n5385), .A2(REIP_REG_29__SCAN_IN), .ZN(n5386) );
  OAI21_X1 U6516 ( .B1(n5442), .B2(n5893), .A(n5388), .ZN(U2798) );
  INV_X1 U6517 ( .A(n5422), .ZN(n5389) );
  AOI21_X1 U6518 ( .B1(n5391), .B2(n5390), .A(n5389), .ZN(n5724) );
  INV_X1 U6519 ( .A(n5724), .ZN(n5430) );
  NAND2_X1 U6520 ( .A1(n6464), .A2(n5393), .ZN(n5664) );
  INV_X1 U6521 ( .A(n5664), .ZN(n5392) );
  OAI21_X1 U6522 ( .B1(n5660), .B2(n5392), .A(REIP_REG_25__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6523 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5393), .ZN(n5650) );
  OAI22_X1 U6524 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5650), .B1(n5727), .B2(
        n5944), .ZN(n5400) );
  AOI21_X1 U6525 ( .B1(n3103), .B2(n5396), .A(n5395), .ZN(n5397) );
  OR2_X1 U6526 ( .A1(n5397), .A2(n5425), .ZN(n5750) );
  AOI22_X1 U6527 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5946), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5901), .ZN(n5398) );
  OAI21_X1 U6528 ( .B1(n5750), .B2(n5933), .A(n5398), .ZN(n5399) );
  NOR2_X1 U6529 ( .A1(n5400), .A2(n5399), .ZN(n5401) );
  OAI211_X1 U6530 ( .C1(n5430), .C2(n5893), .A(n5402), .B(n5401), .ZN(U2802)
         );
  INV_X1 U6531 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5404) );
  OAI222_X1 U6532 ( .A1(n5404), .A2(n5963), .B1(n5958), .B2(n5403), .C1(n5442), 
        .C2(n5959), .ZN(U2830) );
  OR2_X1 U6533 ( .A1(n5416), .A2(n5405), .ZN(n5406) );
  NAND2_X1 U6534 ( .A1(n5696), .A2(n5954), .ZN(n5412) );
  AND2_X1 U6535 ( .A1(n5419), .A2(n5408), .ZN(n5409) );
  NOR2_X1 U6536 ( .A1(n5410), .A2(n5409), .ZN(n5635) );
  NAND2_X1 U6537 ( .A1(n5635), .A2(n5953), .ZN(n5411) );
  OAI211_X1 U6538 ( .C1(n5413), .C2(n5963), .A(n5412), .B(n5411), .ZN(U2831)
         );
  NOR2_X1 U6539 ( .A1(n5421), .A2(n5414), .ZN(n5415) );
  OR2_X1 U6540 ( .A1(n5416), .A2(n5415), .ZN(n5645) );
  INV_X1 U6541 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6542 ( .A1(n5427), .A2(n5417), .ZN(n5418) );
  NAND2_X1 U6543 ( .A1(n5419), .A2(n5418), .ZN(n5644) );
  OAI222_X1 U6544 ( .A1(n5959), .A2(n5645), .B1(n5963), .B2(n5420), .C1(n5644), 
        .C2(n5958), .ZN(U2832) );
  AOI21_X1 U6545 ( .B1(n5423), .B2(n5422), .A(n5421), .ZN(n5475) );
  INV_X1 U6546 ( .A(n5475), .ZN(n5652) );
  INV_X1 U6547 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5428) );
  OR2_X1 U6548 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  NAND2_X1 U6549 ( .A1(n5427), .A2(n5426), .ZN(n5651) );
  OAI222_X1 U6550 ( .A1(n5959), .A2(n5652), .B1(n5963), .B2(n5428), .C1(n5651), 
        .C2(n5958), .ZN(U2833) );
  INV_X1 U6551 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5429) );
  OAI222_X1 U6552 ( .A1(n5430), .A2(n5959), .B1(n5963), .B2(n5429), .C1(n5750), 
        .C2(n5958), .ZN(U2834) );
  AND2_X1 U6553 ( .A1(n5769), .A2(n5431), .ZN(n5433) );
  OR2_X1 U6554 ( .A1(n5433), .A2(n5432), .ZN(n5823) );
  INV_X1 U6555 ( .A(n5434), .ZN(n5435) );
  AOI21_X1 U6556 ( .B1(n5436), .B2(n5746), .A(n5435), .ZN(n5965) );
  INV_X1 U6557 ( .A(n5965), .ZN(n5527) );
  OAI222_X1 U6558 ( .A1(n5823), .A2(n5958), .B1(n5963), .B2(n3091), .C1(n5959), 
        .C2(n5527), .ZN(U2841) );
  NAND3_X1 U6559 ( .A1(n5453), .A2(n5437), .A3(n5978), .ZN(n5439) );
  AOI22_X1 U6560 ( .A1(n5968), .A2(DATAI_31_), .B1(n5970), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U6561 ( .A1(n5439), .A2(n5438), .ZN(U2860) );
  AOI22_X1 U6562 ( .A1(n5968), .A2(DATAI_29_), .B1(n5970), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6563 ( .A1(n5971), .A2(DATAI_13_), .ZN(n5440) );
  OAI211_X1 U6564 ( .C1(n5442), .C2(n5695), .A(n5441), .B(n5440), .ZN(U2862)
         );
  AOI22_X1 U6565 ( .A1(n5971), .A2(DATAI_10_), .B1(n5970), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6566 ( .A1(n5968), .A2(DATAI_26_), .ZN(n5443) );
  OAI211_X1 U6567 ( .C1(n5652), .C2(n5695), .A(n5444), .B(n5443), .ZN(U2865)
         );
  NOR4_X1 U6568 ( .A1(n5445), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n5446), .ZN(n5447) );
  AOI21_X1 U6569 ( .B1(n5448), .B2(n5529), .A(n5447), .ZN(n5449) );
  XNOR2_X1 U6570 ( .A(n5449), .B(n5528), .ZN(n5538) );
  AND2_X1 U6571 ( .A1(n6107), .A2(REIP_REG_31__SCAN_IN), .ZN(n5532) );
  AOI21_X1 U6572 ( .B1(n6048), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5532), 
        .ZN(n5450) );
  OAI21_X1 U6573 ( .B1(n6040), .B2(n5451), .A(n5450), .ZN(n5452) );
  AOI21_X1 U6574 ( .B1(n5453), .B2(n6036), .A(n5452), .ZN(n5454) );
  OAI21_X1 U6575 ( .B1(n5538), .B2(n6042), .A(n5454), .ZN(U2955) );
  NAND3_X1 U6576 ( .A1(n5456), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n4947), .ZN(n5458) );
  NOR2_X1 U6577 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5557) );
  NAND3_X1 U6578 ( .A1(n5723), .A2(n5737), .A3(n5557), .ZN(n5464) );
  AOI22_X1 U6579 ( .A1(n5458), .A2(n5464), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5470), .ZN(n5459) );
  XNOR2_X1 U6580 ( .A(n5459), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5547)
         );
  INV_X1 U6581 ( .A(n5634), .ZN(n5461) );
  AND2_X1 U6582 ( .A1(n6107), .A2(REIP_REG_28__SCAN_IN), .ZN(n5541) );
  AOI21_X1 U6583 ( .B1(n6048), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5541), 
        .ZN(n5460) );
  OAI21_X1 U6584 ( .B1(n6040), .B2(n5461), .A(n5460), .ZN(n5462) );
  AOI21_X1 U6585 ( .B1(n5696), .B2(n6036), .A(n5462), .ZN(n5463) );
  OAI21_X1 U6586 ( .B1(n6042), .B2(n5547), .A(n5463), .ZN(U2958) );
  NAND2_X1 U6587 ( .A1(n5465), .A2(n5464), .ZN(n5466) );
  XNOR2_X1 U6588 ( .A(n5466), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5554)
         );
  INV_X1 U6589 ( .A(n5645), .ZN(n5699) );
  AND2_X1 U6590 ( .A1(n6107), .A2(REIP_REG_27__SCAN_IN), .ZN(n5549) );
  AOI21_X1 U6591 ( .B1(n6048), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5549), 
        .ZN(n5467) );
  OAI21_X1 U6592 ( .B1(n6040), .B2(n5641), .A(n5467), .ZN(n5468) );
  AOI21_X1 U6593 ( .B1(n5699), .B2(n6036), .A(n5468), .ZN(n5469) );
  OAI21_X1 U6594 ( .B1(n5554), .B2(n6042), .A(n5469), .ZN(U2959) );
  XNOR2_X1 U6595 ( .A(n5517), .B(n5470), .ZN(n5471) );
  XNOR2_X1 U6596 ( .A(n5455), .B(n5471), .ZN(n5561) );
  INV_X1 U6597 ( .A(n5649), .ZN(n5473) );
  AND2_X1 U6598 ( .A1(n6107), .A2(REIP_REG_26__SCAN_IN), .ZN(n5556) );
  AOI21_X1 U6599 ( .B1(n6048), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5556), 
        .ZN(n5472) );
  OAI21_X1 U6600 ( .B1(n6040), .B2(n5473), .A(n5472), .ZN(n5474) );
  AOI21_X1 U6601 ( .B1(n5475), .B2(n6036), .A(n5474), .ZN(n5476) );
  OAI21_X1 U6602 ( .B1(n6042), .B2(n5561), .A(n5476), .ZN(U2960) );
  OAI21_X1 U6603 ( .B1(n5477), .B2(n5762), .A(n5517), .ZN(n5478) );
  NAND2_X1 U6604 ( .A1(n5729), .A2(n5478), .ZN(n5509) );
  XNOR2_X1 U6605 ( .A(n5517), .B(n5603), .ZN(n5508) );
  NAND2_X1 U6606 ( .A1(n5737), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5479) );
  INV_X1 U6607 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5591) );
  XNOR2_X1 U6608 ( .A(n5517), .B(n5591), .ZN(n5504) );
  NOR2_X1 U6609 ( .A1(n5503), .A2(n5504), .ZN(n5502) );
  NOR2_X1 U6610 ( .A1(n5517), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5495)
         );
  NAND2_X1 U6611 ( .A1(n5502), .A2(n5495), .ZN(n5487) );
  INV_X1 U6612 ( .A(n5502), .ZN(n5480) );
  OAI21_X1 U6613 ( .B1(n5737), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5480), 
        .ZN(n5497) );
  NAND3_X1 U6614 ( .A1(n4947), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5481) );
  XNOR2_X1 U6615 ( .A(n5482), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5567)
         );
  NAND2_X1 U6616 ( .A1(n5516), .A2(REIP_REG_24__SCAN_IN), .ZN(n5563) );
  OAI21_X1 U6617 ( .B1(n5523), .B2(n5483), .A(n5563), .ZN(n5485) );
  NOR2_X1 U6618 ( .A1(n5661), .A2(n6287), .ZN(n5484) );
  AOI211_X1 U6619 ( .C1(n5525), .C2(n5659), .A(n5485), .B(n5484), .ZN(n5486)
         );
  OAI21_X1 U6620 ( .B1(n5567), .B2(n6042), .A(n5486), .ZN(U2962) );
  NAND2_X1 U6621 ( .A1(n5580), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5488) );
  OAI21_X1 U6622 ( .B1(n5511), .B2(n5488), .A(n5487), .ZN(n5489) );
  XNOR2_X1 U6623 ( .A(n5489), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5576)
         );
  INV_X1 U6624 ( .A(n5490), .ZN(n5707) );
  NAND2_X1 U6625 ( .A1(n6099), .A2(REIP_REG_23__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U6626 ( .A1(n6048), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5491)
         );
  OAI211_X1 U6627 ( .C1(n6040), .C2(n5492), .A(n5568), .B(n5491), .ZN(n5493)
         );
  AOI21_X1 U6628 ( .B1(n5707), .B2(n6036), .A(n5493), .ZN(n5494) );
  OAI21_X1 U6629 ( .B1(n5576), .B2(n6042), .A(n5494), .ZN(U2963) );
  AOI21_X1 U6630 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5517), .A(n5495), 
        .ZN(n5496) );
  XNOR2_X1 U6631 ( .A(n5497), .B(n5496), .ZN(n5586) );
  NAND2_X1 U6632 ( .A1(n5516), .A2(REIP_REG_22__SCAN_IN), .ZN(n5577) );
  OAI21_X1 U6633 ( .B1(n5523), .B2(n5498), .A(n5577), .ZN(n5500) );
  NOR2_X1 U6634 ( .A1(n5670), .A2(n6287), .ZN(n5499) );
  AOI211_X1 U6635 ( .C1(n5525), .C2(n5669), .A(n5500), .B(n5499), .ZN(n5501)
         );
  OAI21_X1 U6636 ( .B1(n5586), .B2(n6042), .A(n5501), .ZN(U2964) );
  AOI21_X1 U6637 ( .B1(n5504), .B2(n5503), .A(n5502), .ZN(n5594) );
  NAND2_X1 U6638 ( .A1(n6099), .A2(REIP_REG_21__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U6639 ( .A1(n6048), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5505)
         );
  OAI211_X1 U6640 ( .C1(n6040), .C2(n5679), .A(n5589), .B(n5505), .ZN(n5506)
         );
  AOI21_X1 U6641 ( .B1(n5713), .B2(n6036), .A(n5506), .ZN(n5507) );
  OAI21_X1 U6642 ( .B1(n5594), .B2(n6042), .A(n5507), .ZN(U2965) );
  NAND2_X1 U6643 ( .A1(n5509), .A2(n5508), .ZN(n5510) );
  NAND2_X1 U6644 ( .A1(n5511), .A2(n5510), .ZN(n5608) );
  INV_X1 U6645 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U6646 ( .A1(n5516), .A2(REIP_REG_20__SCAN_IN), .ZN(n5602) );
  OAI21_X1 U6647 ( .B1(n5523), .B2(n5512), .A(n5602), .ZN(n5514) );
  NOR2_X1 U6648 ( .A1(n5686), .A2(n6287), .ZN(n5513) );
  AOI211_X1 U6649 ( .C1(n5525), .C2(n5690), .A(n5514), .B(n5513), .ZN(n5515)
         );
  OAI21_X1 U6650 ( .B1(n6042), .B2(n5608), .A(n5515), .ZN(U2966) );
  NAND2_X1 U6651 ( .A1(n5516), .A2(REIP_REG_18__SCAN_IN), .ZN(n5609) );
  INV_X1 U6652 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5616) );
  OR3_X1 U6653 ( .A1(n5519), .A2(n5518), .A3(n5517), .ZN(n5740) );
  INV_X1 U6654 ( .A(n5740), .ZN(n5520) );
  NOR3_X1 U6655 ( .A1(n5736), .A2(n5737), .A3(n5599), .ZN(n5741) );
  NOR2_X1 U6656 ( .A1(n5520), .A2(n5741), .ZN(n5521) );
  XOR2_X1 U6657 ( .A(n5616), .B(n5521), .Z(n5612) );
  NAND2_X1 U6658 ( .A1(n6034), .A2(n5612), .ZN(n5522) );
  OAI211_X1 U6659 ( .C1(n5523), .C2(n5819), .A(n5609), .B(n5522), .ZN(n5524)
         );
  AOI21_X1 U6660 ( .B1(n5525), .B2(n5817), .A(n5524), .ZN(n5526) );
  OAI21_X1 U6661 ( .B1(n5527), .B2(n6287), .A(n5526), .ZN(U2968) );
  AND3_X1 U6662 ( .A1(n5530), .A2(n5529), .A3(n5528), .ZN(n5531) );
  AOI211_X1 U6663 ( .C1(INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n5533), .A(n5532), .B(n5531), .ZN(n5537) );
  INV_X1 U6664 ( .A(n5534), .ZN(n5535) );
  NAND2_X1 U6665 ( .A1(n5535), .A2(n6109), .ZN(n5536) );
  OAI211_X1 U6666 ( .C1(n5538), .C2(n6084), .A(n5537), .B(n5536), .ZN(U2987)
         );
  INV_X1 U6667 ( .A(n5635), .ZN(n5539) );
  NOR2_X1 U6668 ( .A1(n5539), .A2(n6082), .ZN(n5540) );
  AOI211_X1 U6669 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5550), .A(n5541), .B(n5540), .ZN(n5546) );
  INV_X1 U6670 ( .A(n5542), .ZN(n5543) );
  OR3_X1 U6671 ( .A1(n5551), .A2(n5544), .A3(n5543), .ZN(n5545) );
  OAI211_X1 U6672 ( .C1(n5547), .C2(n6084), .A(n5546), .B(n5545), .ZN(U2990)
         );
  NOR2_X1 U6673 ( .A1(n5644), .A2(n6082), .ZN(n5548) );
  AOI211_X1 U6674 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5550), .A(n5549), .B(n5548), .ZN(n5553) );
  OR2_X1 U6675 ( .A1(n5551), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5552)
         );
  OAI211_X1 U6676 ( .C1(n5554), .C2(n6084), .A(n5553), .B(n5552), .ZN(U2991)
         );
  NOR2_X1 U6677 ( .A1(n5651), .A2(n6082), .ZN(n5555) );
  AOI211_X1 U6678 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5749), .A(n5556), .B(n5555), .ZN(n5560) );
  OR3_X1 U6679 ( .A1(n5755), .A2(n5558), .A3(n5557), .ZN(n5559) );
  OAI211_X1 U6680 ( .C1(n5561), .C2(n6084), .A(n5560), .B(n5559), .ZN(U2992)
         );
  OAI21_X1 U6681 ( .B1(n5571), .B2(n5569), .A(n5562), .ZN(n5565) );
  OAI21_X1 U6682 ( .B1(n5662), .B2(n6082), .A(n5563), .ZN(n5564) );
  AOI21_X1 U6683 ( .B1(n5565), .B2(n5749), .A(n5564), .ZN(n5566) );
  OAI21_X1 U6684 ( .B1(n5567), .B2(n6084), .A(n5566), .ZN(U2994) );
  OAI21_X1 U6685 ( .B1(n5570), .B2(n5569), .A(n5568), .ZN(n5573) );
  NOR2_X1 U6686 ( .A1(n5571), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5572)
         );
  AOI211_X1 U6687 ( .C1(n6109), .C2(n5574), .A(n5573), .B(n5572), .ZN(n5575)
         );
  OAI21_X1 U6688 ( .B1(n5576), .B2(n6084), .A(n5575), .ZN(U2995) );
  INV_X1 U6689 ( .A(n5587), .ZN(n5579) );
  INV_X1 U6690 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5578) );
  OAI21_X1 U6691 ( .B1(n5579), .B2(n5578), .A(n5577), .ZN(n5584) );
  INV_X1 U6692 ( .A(n5592), .ZN(n5582) );
  NOR3_X1 U6693 ( .A1(n5582), .A2(n5581), .A3(n5580), .ZN(n5583) );
  AOI211_X1 U6694 ( .C1(n6109), .C2(n5671), .A(n5584), .B(n5583), .ZN(n5585)
         );
  OAI21_X1 U6695 ( .B1(n5586), .B2(n6084), .A(n5585), .ZN(U2996) );
  NAND2_X1 U6696 ( .A1(n5587), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5588) );
  OAI211_X1 U6697 ( .C1(n5681), .C2(n6082), .A(n5589), .B(n5588), .ZN(n5590)
         );
  AOI21_X1 U6698 ( .B1(n5592), .B2(n5591), .A(n5590), .ZN(n5593) );
  OAI21_X1 U6699 ( .B1(n5594), .B2(n6084), .A(n5593), .ZN(U2997) );
  AOI21_X1 U6700 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5596), .A(n5595), 
        .ZN(n5597) );
  NOR2_X1 U6701 ( .A1(n5598), .A2(n5597), .ZN(n5773) );
  NAND2_X1 U6702 ( .A1(n6100), .A2(n5599), .ZN(n5600) );
  AND2_X1 U6703 ( .A1(n5773), .A2(n5600), .ZN(n5617) );
  NAND2_X1 U6704 ( .A1(n6106), .A2(n5616), .ZN(n5601) );
  AND2_X1 U6705 ( .A1(n5617), .A2(n5601), .ZN(n5763) );
  OAI21_X1 U6706 ( .B1(n5763), .B2(n5603), .A(n5602), .ZN(n5606) );
  XNOR2_X1 U6707 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .B(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5604) );
  NOR3_X1 U6708 ( .A1(n5764), .A2(n5756), .A3(n5604), .ZN(n5605) );
  AOI211_X1 U6709 ( .C1(n6109), .C2(n5687), .A(n5606), .B(n5605), .ZN(n5607)
         );
  OAI21_X1 U6710 ( .B1(n5608), .B2(n6084), .A(n5607), .ZN(U2998) );
  INV_X1 U6711 ( .A(n5609), .ZN(n5611) );
  NOR3_X1 U6712 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5599), .A3(n5764), 
        .ZN(n5610) );
  AOI211_X1 U6713 ( .C1(n6112), .C2(n5612), .A(n5611), .B(n5610), .ZN(n5615)
         );
  INV_X1 U6714 ( .A(n5823), .ZN(n5613) );
  NAND2_X1 U6715 ( .A1(n5613), .A2(n6109), .ZN(n5614) );
  OAI211_X1 U6716 ( .C1(n5617), .C2(n5616), .A(n5615), .B(n5614), .ZN(U3000)
         );
  OAI21_X1 U6717 ( .B1(n4300), .B2(STATEBS16_REG_SCAN_IN), .A(n6521), .ZN(
        n5619) );
  OAI22_X1 U6718 ( .A1(n5619), .A2(n6243), .B1(n5618), .B2(n5622), .ZN(n5620)
         );
  MUX2_X1 U6719 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5620), .S(n6116), 
        .Z(U3464) );
  XNOR2_X1 U6720 ( .A(n3426), .B(n6243), .ZN(n5624) );
  INV_X1 U6721 ( .A(n5621), .ZN(n5623) );
  OAI22_X1 U6722 ( .A1(n5624), .A2(n6284), .B1(n5623), .B2(n5622), .ZN(n5625)
         );
  MUX2_X1 U6723 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5625), .S(n6116), 
        .Z(U3463) );
  AND2_X1 U6724 ( .A1(n5626), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6725 ( .A(n5627), .ZN(n5632) );
  INV_X1 U6726 ( .A(n5628), .ZN(n5629) );
  AOI21_X1 U6727 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5630), .A(n5629), .ZN(
        n5631) );
  NAND2_X1 U6728 ( .A1(n5632), .A2(n5631), .ZN(U2788) );
  AOI22_X1 U6729 ( .A1(EBX_REG_28__SCAN_IN), .A2(n5946), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n5901), .ZN(n5639) );
  AOI22_X1 U6730 ( .A1(n5634), .A2(n5907), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5633), .ZN(n5638) );
  AOI22_X1 U6731 ( .A1(n5696), .A2(n5870), .B1(n5635), .B2(n5943), .ZN(n5637)
         );
  INV_X1 U6732 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6663) );
  NAND3_X1 U6733 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5643), .A3(n6663), .ZN(
        n5636) );
  NAND4_X1 U6734 ( .A1(n5639), .A2(n5638), .A3(n5637), .A4(n5636), .ZN(U2799)
         );
  INV_X1 U6735 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6471) );
  AOI22_X1 U6736 ( .A1(EBX_REG_27__SCAN_IN), .A2(n5946), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5901), .ZN(n5640) );
  OAI21_X1 U6737 ( .B1(n5641), .B2(n5944), .A(n5640), .ZN(n5642) );
  AOI221_X1 U6738 ( .B1(n5655), .B2(REIP_REG_27__SCAN_IN), .C1(n5643), .C2(
        n6471), .A(n5642), .ZN(n5648) );
  OAI22_X1 U6739 ( .A1(n5645), .A2(n5893), .B1(n5644), .B2(n5933), .ZN(n5646)
         );
  INV_X1 U6740 ( .A(n5646), .ZN(n5647) );
  NAND2_X1 U6741 ( .A1(n5648), .A2(n5647), .ZN(U2800) );
  AOI22_X1 U6742 ( .A1(EBX_REG_26__SCAN_IN), .A2(n5946), .B1(n5649), .B2(n5907), .ZN(n5657) );
  OAI21_X1 U6743 ( .B1(n6466), .B2(n5650), .A(n6468), .ZN(n5654) );
  OAI22_X1 U6744 ( .A1(n5652), .A2(n5893), .B1(n5651), .B2(n5933), .ZN(n5653)
         );
  AOI21_X1 U6745 ( .B1(n5655), .B2(n5654), .A(n5653), .ZN(n5656) );
  OAI211_X1 U6746 ( .C1(n5658), .C2(n5945), .A(n5657), .B(n5656), .ZN(U2801)
         );
  AOI22_X1 U6747 ( .A1(EBX_REG_24__SCAN_IN), .A2(n5946), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5901), .ZN(n5667) );
  AOI22_X1 U6748 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5660), .B1(n5659), .B2(
        n5907), .ZN(n5666) );
  INV_X1 U6749 ( .A(n5661), .ZN(n5704) );
  INV_X1 U6750 ( .A(n5662), .ZN(n5663) );
  AOI22_X1 U6751 ( .A1(n5704), .A2(n5870), .B1(n5943), .B2(n5663), .ZN(n5665)
         );
  NAND4_X1 U6752 ( .A1(n5667), .A2(n5666), .A3(n5665), .A4(n5664), .ZN(U2803)
         );
  AOI22_X1 U6753 ( .A1(EBX_REG_22__SCAN_IN), .A2(n5946), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5901), .ZN(n5677) );
  AND2_X1 U6754 ( .A1(n5941), .A2(n5668), .ZN(n5688) );
  AOI22_X1 U6755 ( .A1(n5669), .A2(n5907), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5688), .ZN(n5676) );
  INV_X1 U6756 ( .A(n5670), .ZN(n5710) );
  AOI22_X1 U6757 ( .A1(n5710), .A2(n5870), .B1(n5943), .B2(n5671), .ZN(n5675)
         );
  INV_X1 U6758 ( .A(n5685), .ZN(n5673) );
  OAI211_X1 U6759 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5673), .B(n5672), .ZN(n5674) );
  NAND4_X1 U6760 ( .A1(n5677), .A2(n5676), .A3(n5675), .A4(n5674), .ZN(U2805)
         );
  AOI22_X1 U6761 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5946), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5901), .ZN(n5678) );
  OAI21_X1 U6762 ( .B1(n5679), .B2(n5944), .A(n5678), .ZN(n5680) );
  AOI21_X1 U6763 ( .B1(REIP_REG_21__SCAN_IN), .B2(n5688), .A(n5680), .ZN(n5684) );
  INV_X1 U6764 ( .A(n5681), .ZN(n5682) );
  AOI22_X1 U6765 ( .A1(n5713), .A2(n5870), .B1(n5943), .B2(n5682), .ZN(n5683)
         );
  OAI211_X1 U6766 ( .C1(REIP_REG_21__SCAN_IN), .C2(n5685), .A(n5684), .B(n5683), .ZN(U2806) );
  AOI22_X1 U6767 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5946), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n5901), .ZN(n5694) );
  INV_X1 U6768 ( .A(n5686), .ZN(n5716) );
  AOI22_X1 U6769 ( .A1(n5716), .A2(n5870), .B1(n5943), .B2(n5687), .ZN(n5693)
         );
  OAI21_X1 U6770 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5689), .A(n5688), .ZN(n5692) );
  NAND2_X1 U6771 ( .A1(n5690), .A2(n5907), .ZN(n5691) );
  NAND4_X1 U6772 ( .A1(n5694), .A2(n5693), .A3(n5692), .A4(n5691), .ZN(U2807)
         );
  AOI22_X1 U6773 ( .A1(n5696), .A2(n5975), .B1(n5968), .B2(DATAI_28_), .ZN(
        n5698) );
  AOI22_X1 U6774 ( .A1(n5971), .A2(DATAI_12_), .B1(n5970), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U6775 ( .A1(n5698), .A2(n5697), .ZN(U2863) );
  AOI22_X1 U6776 ( .A1(n5699), .A2(n5975), .B1(n5968), .B2(DATAI_27_), .ZN(
        n5701) );
  AOI22_X1 U6777 ( .A1(n5971), .A2(DATAI_11_), .B1(n5970), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U6778 ( .A1(n5701), .A2(n5700), .ZN(U2864) );
  AOI22_X1 U6779 ( .A1(n5724), .A2(n5975), .B1(n5968), .B2(DATAI_25_), .ZN(
        n5703) );
  AOI22_X1 U6780 ( .A1(n5971), .A2(DATAI_9_), .B1(n5970), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U6781 ( .A1(n5703), .A2(n5702), .ZN(U2866) );
  AOI22_X1 U6782 ( .A1(n5704), .A2(n5975), .B1(n5968), .B2(DATAI_24_), .ZN(
        n5706) );
  AOI22_X1 U6783 ( .A1(n5971), .A2(DATAI_8_), .B1(n5970), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U6784 ( .A1(n5706), .A2(n5705), .ZN(U2867) );
  AOI22_X1 U6785 ( .A1(n5707), .A2(n5975), .B1(n5968), .B2(DATAI_23_), .ZN(
        n5709) );
  AOI22_X1 U6786 ( .A1(n5971), .A2(DATAI_7_), .B1(n5970), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U6787 ( .A1(n5709), .A2(n5708), .ZN(U2868) );
  AOI22_X1 U6788 ( .A1(n5710), .A2(n5975), .B1(n5968), .B2(DATAI_22_), .ZN(
        n5712) );
  AOI22_X1 U6789 ( .A1(n5971), .A2(DATAI_6_), .B1(n5970), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U6790 ( .A1(n5712), .A2(n5711), .ZN(U2869) );
  AOI22_X1 U6791 ( .A1(n5713), .A2(n5975), .B1(n5968), .B2(DATAI_21_), .ZN(
        n5715) );
  AOI22_X1 U6792 ( .A1(n5971), .A2(DATAI_5_), .B1(n5970), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U6793 ( .A1(n5715), .A2(n5714), .ZN(U2870) );
  AOI22_X1 U6794 ( .A1(n5716), .A2(n5975), .B1(n5968), .B2(DATAI_20_), .ZN(
        n5718) );
  AOI22_X1 U6795 ( .A1(n5971), .A2(DATAI_4_), .B1(n5970), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5717) );
  NAND2_X1 U6796 ( .A1(n5718), .A2(n5717), .ZN(U2871) );
  INV_X1 U6797 ( .A(n5719), .ZN(n5731) );
  AOI22_X1 U6798 ( .A1(n5731), .A2(n5975), .B1(n5968), .B2(DATAI_19_), .ZN(
        n5721) );
  AOI22_X1 U6799 ( .A1(n5971), .A2(DATAI_3_), .B1(n5970), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U6800 ( .A1(n5721), .A2(n5720), .ZN(U2872) );
  AOI22_X1 U6801 ( .A1(n6107), .A2(REIP_REG_25__SCAN_IN), .B1(n6048), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5726) );
  OAI21_X1 U6802 ( .B1(n5723), .B2(n5722), .A(n5445), .ZN(n5752) );
  AOI22_X1 U6803 ( .A1(n5724), .A2(n6036), .B1(n6034), .B2(n5752), .ZN(n5725)
         );
  OAI211_X1 U6804 ( .C1(n6040), .C2(n5727), .A(n5726), .B(n5725), .ZN(U2961)
         );
  AOI22_X1 U6805 ( .A1(n6107), .A2(REIP_REG_19__SCAN_IN), .B1(n6048), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U6806 ( .A1(n5729), .A2(n5728), .ZN(n5730) );
  XNOR2_X1 U6807 ( .A(n5730), .B(n5737), .ZN(n5759) );
  AOI22_X1 U6808 ( .A1(n5759), .A2(n6034), .B1(n6036), .B2(n5731), .ZN(n5732)
         );
  OAI211_X1 U6809 ( .C1(n6040), .C2(n5734), .A(n5733), .B(n5732), .ZN(U2967)
         );
  AOI22_X1 U6810 ( .A1(n6107), .A2(REIP_REG_17__SCAN_IN), .B1(n6048), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U6811 ( .A1(n5737), .A2(n5735), .ZN(n5739) );
  AOI21_X1 U6812 ( .B1(n5737), .B2(n5599), .A(n5736), .ZN(n5738) );
  AOI21_X1 U6813 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5739), .A(n5738), 
        .ZN(n5742) );
  OAI21_X1 U6814 ( .B1(n5742), .B2(n5741), .A(n5740), .ZN(n5770) );
  NAND2_X1 U6815 ( .A1(n5744), .A2(n5743), .ZN(n5745) );
  AOI22_X1 U6816 ( .A1(n5770), .A2(n6034), .B1(n6036), .B2(n5969), .ZN(n5747)
         );
  OAI211_X1 U6817 ( .C1(n6040), .C2(n5826), .A(n5748), .B(n5747), .ZN(U2969)
         );
  AOI22_X1 U6818 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n5749), .B1(n6099), .B2(REIP_REG_25__SCAN_IN), .ZN(n5754) );
  INV_X1 U6819 ( .A(n5750), .ZN(n5751) );
  AOI22_X1 U6820 ( .A1(n5752), .A2(n6112), .B1(n6109), .B2(n5751), .ZN(n5753)
         );
  OAI211_X1 U6821 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5755), .A(n5754), .B(n5753), .ZN(U2993) );
  NOR2_X1 U6822 ( .A1(n5756), .A2(n5764), .ZN(n5757) );
  AOI22_X1 U6823 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6099), .B1(n5757), .B2(
        n5762), .ZN(n5761) );
  AOI22_X1 U6824 ( .A1(n5759), .A2(n6112), .B1(n6109), .B2(n5758), .ZN(n5760)
         );
  OAI211_X1 U6825 ( .C1(n5763), .C2(n5762), .A(n5761), .B(n5760), .ZN(U2999)
         );
  INV_X1 U6826 ( .A(n5764), .ZN(n5765) );
  AOI22_X1 U6827 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6099), .B1(n5765), .B2(
        n5599), .ZN(n5772) );
  NAND2_X1 U6828 ( .A1(n5767), .A2(n5766), .ZN(n5768) );
  AND2_X1 U6829 ( .A1(n5769), .A2(n5768), .ZN(n5952) );
  AOI22_X1 U6830 ( .A1(n5770), .A2(n6112), .B1(n6109), .B2(n5952), .ZN(n5771)
         );
  OAI211_X1 U6831 ( .C1(n5773), .C2(n5599), .A(n5772), .B(n5771), .ZN(U3001)
         );
  NAND3_X1 U6832 ( .A1(n5776), .A2(n5775), .A3(n5774), .ZN(n5778) );
  OAI211_X1 U6833 ( .C1(n6082), .C2(n5840), .A(n5778), .B(n5777), .ZN(n5779)
         );
  AOI21_X1 U6834 ( .B1(n5780), .B2(n6112), .A(n5779), .ZN(n5782) );
  OAI211_X1 U6835 ( .C1(n5784), .C2(n5783), .A(n5782), .B(n5781), .ZN(U3005)
         );
  INV_X1 U6836 ( .A(n5785), .ZN(n5789) );
  INV_X1 U6837 ( .A(n5786), .ZN(n5788) );
  NAND4_X1 U6838 ( .A1(n5789), .A2(n5788), .A3(n5787), .A4(n5916), .ZN(n5790)
         );
  OAI21_X1 U6839 ( .B1(n6502), .B2(n4293), .A(n5790), .ZN(U3455) );
  INV_X1 U6840 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6421) );
  NOR2_X1 U6841 ( .A1(n6421), .A2(STATE_REG_0__SCAN_IN), .ZN(n6481) );
  OAI21_X1 U6842 ( .B1(STATE_REG_2__SCAN_IN), .B2(n6421), .A(
        STATE_REG_0__SCAN_IN), .ZN(n5795) );
  NOR2_X1 U6843 ( .A1(ADS_N_REG_SCAN_IN), .A2(n5795), .ZN(n5791) );
  NOR2_X1 U6844 ( .A1(n6481), .A2(n5791), .ZN(U2789) );
  OAI21_X1 U6845 ( .B1(n6351), .B2(n6349), .A(n6346), .ZN(n5792) );
  OAI21_X1 U6846 ( .B1(n6394), .B2(n3348), .A(n5792), .ZN(n5801) );
  OAI21_X1 U6847 ( .B1(n5801), .B2(n6406), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5793) );
  OAI21_X1 U6848 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6405), .A(n5793), .ZN(
        U2790) );
  INV_X1 U6849 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6583) );
  NOR2_X1 U6850 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5796) );
  NOR2_X1 U6851 ( .A1(n6481), .A2(n5796), .ZN(n5794) );
  AOI22_X1 U6852 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6481), .B1(n6583), .B2(
        n5794), .ZN(U2791) );
  NAND2_X1 U6853 ( .A1(n6531), .A2(n5795), .ZN(n6683) );
  INV_X1 U6854 ( .A(n6683), .ZN(n6485) );
  OAI21_X1 U6855 ( .B1(BS16_N), .B2(n5796), .A(n6485), .ZN(n6483) );
  OAI21_X1 U6856 ( .B1(n6485), .B2(n6621), .A(n6483), .ZN(U2792) );
  OR3_X1 U6857 ( .A1(n5799), .A2(n3348), .A3(n5797), .ZN(n5800) );
  AND2_X1 U6858 ( .A1(n5800), .A2(n6572), .ZN(n6524) );
  NOR2_X1 U6859 ( .A1(n5801), .A2(n6524), .ZN(n6357) );
  NOR2_X1 U6860 ( .A1(n6357), .A2(n6406), .ZN(n6519) );
  OAI21_X1 U6861 ( .B1(n6519), .B2(n5802), .A(n6042), .ZN(U2793) );
  NOR2_X1 U6862 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6537) );
  AOI211_X1 U6863 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_6__SCAN_IN), .B(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n5803) );
  INV_X1 U6864 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6626) );
  INV_X1 U6865 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6623) );
  NAND4_X1 U6866 ( .A1(n6537), .A2(n5803), .A3(n6626), .A4(n6623), .ZN(n5811)
         );
  OR4_X1 U6867 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_11__SCAN_IN), 
        .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(
        n5810) );
  OR4_X1 U6868 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n5809) );
  NOR4_X1 U6869 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5807) );
  NOR4_X1 U6870 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n5806) );
  NOR4_X1 U6871 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n5805) );
  NOR4_X1 U6872 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5804) );
  NAND4_X1 U6873 ( .A1(n5807), .A2(n5806), .A3(n5805), .A4(n5804), .ZN(n5808)
         );
  INV_X1 U6874 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5813) );
  NOR3_X1 U6875 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5814) );
  OAI21_X1 U6876 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5814), .A(n6510), .ZN(n5812)
         );
  OAI21_X1 U6877 ( .B1(n6510), .B2(n5813), .A(n5812), .ZN(U2794) );
  INV_X1 U6878 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6506) );
  INV_X1 U6879 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6484) );
  AOI21_X1 U6880 ( .B1(n6506), .B2(n6484), .A(n5814), .ZN(n5815) );
  INV_X1 U6881 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6647) );
  INV_X1 U6882 ( .A(n6510), .ZN(n6513) );
  AOI22_X1 U6883 ( .A1(n6510), .A2(n5815), .B1(n6647), .B2(n6513), .ZN(U2795)
         );
  INV_X1 U6884 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6457) );
  AOI22_X1 U6885 ( .A1(n5817), .A2(n5907), .B1(n5816), .B2(n6457), .ZN(n5822)
         );
  AOI22_X1 U6886 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5946), .B1(
        REIP_REG_18__SCAN_IN), .B2(n5825), .ZN(n5818) );
  OAI211_X1 U6887 ( .C1(n5945), .C2(n5819), .A(n5818), .B(n4850), .ZN(n5820)
         );
  AOI21_X1 U6888 ( .B1(n5965), .B2(n5870), .A(n5820), .ZN(n5821) );
  OAI211_X1 U6889 ( .C1(n5933), .C2(n5823), .A(n5822), .B(n5821), .ZN(U2809)
         );
  AOI21_X1 U6890 ( .B1(REIP_REG_16__SCAN_IN), .B2(n5824), .A(
        REIP_REG_17__SCAN_IN), .ZN(n5831) );
  INV_X1 U6891 ( .A(n5825), .ZN(n5830) );
  OAI22_X1 U6892 ( .A1(n3779), .A2(n5945), .B1(n5826), .B2(n5944), .ZN(n5827)
         );
  AOI211_X1 U6893 ( .C1(n5946), .C2(EBX_REG_17__SCAN_IN), .A(n6107), .B(n5827), 
        .ZN(n5829) );
  AOI22_X1 U6894 ( .A1(n5969), .A2(n5870), .B1(n5943), .B2(n5952), .ZN(n5828)
         );
  OAI211_X1 U6895 ( .C1(n5831), .C2(n5830), .A(n5829), .B(n5828), .ZN(U2810)
         );
  AOI22_X1 U6896 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n5901), .B1(n5943), 
        .B2(n5832), .ZN(n5833) );
  OAI211_X1 U6897 ( .C1(n5886), .C2(n5964), .A(n5833), .B(n4850), .ZN(n5834)
         );
  AOI211_X1 U6898 ( .C1(n5836), .C2(REIP_REG_15__SCAN_IN), .A(n5835), .B(n5834), .ZN(n5839) );
  AOI22_X1 U6899 ( .A1(n5976), .A2(n5870), .B1(n5907), .B2(n5837), .ZN(n5838)
         );
  NAND2_X1 U6900 ( .A1(n5839), .A2(n5838), .ZN(U2812) );
  INV_X1 U6901 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5841) );
  OAI22_X1 U6902 ( .A1(n5841), .A2(n5886), .B1(n5933), .B2(n5840), .ZN(n5842)
         );
  AOI211_X1 U6903 ( .C1(n5901), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6107), 
        .B(n5842), .ZN(n5853) );
  INV_X1 U6904 ( .A(n5843), .ZN(n5845) );
  AOI22_X1 U6905 ( .A1(n5845), .A2(n5870), .B1(n5907), .B2(n5844), .ZN(n5852)
         );
  INV_X1 U6906 ( .A(n5846), .ZN(n5847) );
  NAND2_X1 U6907 ( .A1(n6447), .A2(n5847), .ZN(n5848) );
  NOR2_X1 U6908 ( .A1(n5918), .A2(n5848), .ZN(n5860) );
  OAI21_X1 U6909 ( .B1(n5860), .B2(n5856), .A(REIP_REG_13__SCAN_IN), .ZN(n5851) );
  INV_X1 U6910 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6449) );
  NAND3_X1 U6911 ( .A1(n5900), .A2(n6449), .A3(n5849), .ZN(n5850) );
  NAND4_X1 U6912 ( .A1(n5853), .A2(n5852), .A3(n5851), .A4(n5850), .ZN(U2814)
         );
  OAI21_X1 U6913 ( .B1(n5933), .B2(n5854), .A(n4850), .ZN(n5855) );
  AOI21_X1 U6914 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n5901), .A(n5855), 
        .ZN(n5864) );
  AOI22_X1 U6915 ( .A1(EBX_REG_12__SCAN_IN), .A2(n5946), .B1(
        REIP_REG_12__SCAN_IN), .B2(n5856), .ZN(n5863) );
  OAI22_X1 U6916 ( .A1(n5858), .A2(n5893), .B1(n5857), .B2(n5944), .ZN(n5859)
         );
  INV_X1 U6917 ( .A(n5859), .ZN(n5862) );
  INV_X1 U6918 ( .A(n5860), .ZN(n5861) );
  NAND4_X1 U6919 ( .A1(n5864), .A2(n5863), .A3(n5862), .A4(n5861), .ZN(U2815)
         );
  AOI22_X1 U6920 ( .A1(EBX_REG_10__SCAN_IN), .A2(n5946), .B1(n5943), .B2(n5865), .ZN(n5876) );
  NOR3_X1 U6921 ( .A1(n5918), .A2(REIP_REG_10__SCAN_IN), .A3(n5866), .ZN(n5867) );
  AOI211_X1 U6922 ( .C1(n5901), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6107), 
        .B(n5867), .ZN(n5875) );
  INV_X1 U6923 ( .A(n5868), .ZN(n5871) );
  AOI22_X1 U6924 ( .A1(n5871), .A2(n5870), .B1(n5907), .B2(n5869), .ZN(n5874)
         );
  NOR3_X1 U6925 ( .A1(n5918), .A2(REIP_REG_9__SCAN_IN), .A3(n5872), .ZN(n5877)
         );
  OAI21_X1 U6926 ( .B1(n5877), .B2(n5878), .A(REIP_REG_10__SCAN_IN), .ZN(n5873) );
  NAND4_X1 U6927 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(U2817)
         );
  AOI21_X1 U6928 ( .B1(REIP_REG_9__SCAN_IN), .B2(n5878), .A(n5877), .ZN(n5885)
         );
  OAI21_X1 U6929 ( .B1(n5945), .B2(n6625), .A(n4850), .ZN(n5879) );
  AOI21_X1 U6930 ( .B1(n5943), .B2(n6063), .A(n5879), .ZN(n5880) );
  OAI21_X1 U6931 ( .B1(n5881), .B2(n5893), .A(n5880), .ZN(n5882) );
  AOI21_X1 U6932 ( .B1(n5883), .B2(n5907), .A(n5882), .ZN(n5884) );
  OAI211_X1 U6933 ( .C1(n5887), .C2(n5886), .A(n5885), .B(n5884), .ZN(U2818)
         );
  INV_X1 U6934 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6440) );
  INV_X1 U6935 ( .A(n5888), .ZN(n6070) );
  NOR2_X1 U6936 ( .A1(n5918), .A2(REIP_REG_7__SCAN_IN), .ZN(n5889) );
  AOI22_X1 U6937 ( .A1(n5943), .A2(n6070), .B1(n5890), .B2(n5889), .ZN(n5891)
         );
  OAI211_X1 U6938 ( .C1(n5945), .C2(n4579), .A(n5891), .B(n4850), .ZN(n5896)
         );
  OAI22_X1 U6939 ( .A1(n5894), .A2(n5893), .B1(n5892), .B2(n5944), .ZN(n5895)
         );
  AOI211_X1 U6940 ( .C1(EBX_REG_7__SCAN_IN), .C2(n5946), .A(n5896), .B(n5895), 
        .ZN(n5897) );
  OAI221_X1 U6941 ( .B1(n6440), .B2(n5911), .C1(n6440), .C2(n5898), .A(n5897), 
        .ZN(U2820) );
  AOI21_X1 U6942 ( .B1(n5900), .B2(n5899), .A(REIP_REG_5__SCAN_IN), .ZN(n5912)
         );
  AOI22_X1 U6943 ( .A1(EBX_REG_5__SCAN_IN), .A2(n5946), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n5901), .ZN(n5902) );
  INV_X1 U6944 ( .A(n5902), .ZN(n5903) );
  AOI211_X1 U6945 ( .C1(n5943), .C2(n5904), .A(n6107), .B(n5903), .ZN(n5910)
         );
  INV_X1 U6946 ( .A(n5951), .ZN(n5923) );
  INV_X1 U6947 ( .A(n5905), .ZN(n5906) );
  AOI22_X1 U6948 ( .A1(n5908), .A2(n5923), .B1(n5907), .B2(n5906), .ZN(n5909)
         );
  OAI211_X1 U6949 ( .C1(n5912), .C2(n5911), .A(n5910), .B(n5909), .ZN(U2822)
         );
  OAI21_X1 U6950 ( .B1(n5913), .B2(n5917), .A(n5941), .ZN(n5940) );
  OAI22_X1 U6951 ( .A1(n5914), .A2(n5945), .B1(n6434), .B2(n5940), .ZN(n5915)
         );
  AOI211_X1 U6952 ( .C1(n5916), .C2(n5947), .A(n6107), .B(n5915), .ZN(n5926)
         );
  NOR3_X1 U6953 ( .A1(n5918), .A2(REIP_REG_4__SCAN_IN), .A3(n5917), .ZN(n5919)
         );
  AOI21_X1 U6954 ( .B1(n5946), .B2(EBX_REG_4__SCAN_IN), .A(n5919), .ZN(n5920)
         );
  OAI21_X1 U6955 ( .B1(n5933), .B2(n5921), .A(n5920), .ZN(n5922) );
  AOI21_X1 U6956 ( .B1(n5924), .B2(n5923), .A(n5922), .ZN(n5925) );
  OAI211_X1 U6957 ( .C1(n5927), .C2(n5944), .A(n5926), .B(n5925), .ZN(U2823)
         );
  INV_X1 U6958 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6433) );
  OR2_X1 U6959 ( .A1(n5929), .A2(n5928), .ZN(n5939) );
  INV_X1 U6960 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5930) );
  OAI222_X1 U6961 ( .A1(n5933), .A2(n6081), .B1(n5932), .B2(n5931), .C1(n5945), 
        .C2(n5930), .ZN(n5937) );
  OAI22_X1 U6962 ( .A1(n5951), .A2(n5935), .B1(n5934), .B2(n5944), .ZN(n5936)
         );
  AOI211_X1 U6963 ( .C1(EBX_REG_3__SCAN_IN), .C2(n5946), .A(n5937), .B(n5936), 
        .ZN(n5938) );
  OAI221_X1 U6964 ( .B1(n5940), .B2(n6433), .C1(n5940), .C2(n5939), .A(n5938), 
        .ZN(U2824) );
  AOI22_X1 U6965 ( .A1(n5943), .A2(n5942), .B1(REIP_REG_0__SCAN_IN), .B2(n5941), .ZN(n5950) );
  NAND2_X1 U6966 ( .A1(n5945), .A2(n5944), .ZN(n5948) );
  AOI222_X1 U6967 ( .A1(n5948), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n6365), 
        .B2(n5947), .C1(EBX_REG_0__SCAN_IN), .C2(n5946), .ZN(n5949) );
  OAI211_X1 U6968 ( .C1(n5951), .C2(n6052), .A(n5950), .B(n5949), .ZN(U2827)
         );
  INV_X1 U6969 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5956) );
  AOI22_X1 U6970 ( .A1(n5969), .A2(n5954), .B1(n5953), .B2(n5952), .ZN(n5955)
         );
  OAI21_X1 U6971 ( .B1(n5956), .B2(n5963), .A(n5955), .ZN(U2842) );
  OAI22_X1 U6972 ( .A1(n5960), .A2(n5959), .B1(n5958), .B2(n5957), .ZN(n5961)
         );
  INV_X1 U6973 ( .A(n5961), .ZN(n5962) );
  OAI21_X1 U6974 ( .B1(n5964), .B2(n5963), .A(n5962), .ZN(U2844) );
  AOI22_X1 U6975 ( .A1(n5965), .A2(n5975), .B1(n5968), .B2(DATAI_18_), .ZN(
        n5967) );
  AOI22_X1 U6976 ( .A1(n5971), .A2(DATAI_2_), .B1(n5970), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U6977 ( .A1(n5967), .A2(n5966), .ZN(U2873) );
  AOI22_X1 U6978 ( .A1(n5969), .A2(n5975), .B1(n5968), .B2(DATAI_17_), .ZN(
        n5973) );
  AOI22_X1 U6979 ( .A1(n5971), .A2(DATAI_1_), .B1(n5970), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U6980 ( .A1(n5973), .A2(n5972), .ZN(U2874) );
  INV_X1 U6981 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U6982 ( .A1(n5976), .A2(n5975), .B1(DATAI_15_), .B2(n5974), .ZN(
        n5977) );
  OAI21_X1 U6983 ( .B1(n6671), .B2(n5978), .A(n5977), .ZN(U2876) );
  AOI22_X1 U6984 ( .A1(n4378), .A2(LWORD_REG_15__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5980) );
  OAI21_X1 U6985 ( .B1(n6671), .B2(n6007), .A(n5980), .ZN(U2908) );
  INV_X1 U6986 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5982) );
  AOI22_X1 U6987 ( .A1(n4378), .A2(LWORD_REG_14__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5981) );
  OAI21_X1 U6988 ( .B1(n5982), .B2(n6007), .A(n5981), .ZN(U2909) );
  AOI22_X1 U6989 ( .A1(n4378), .A2(LWORD_REG_13__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5983) );
  OAI21_X1 U6990 ( .B1(n5984), .B2(n6007), .A(n5983), .ZN(U2910) );
  AOI22_X1 U6991 ( .A1(n4378), .A2(LWORD_REG_12__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5985) );
  OAI21_X1 U6992 ( .B1(n4575), .B2(n6007), .A(n5985), .ZN(U2911) );
  INV_X1 U6993 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5987) );
  AOI22_X1 U6994 ( .A1(n4378), .A2(LWORD_REG_11__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5986) );
  OAI21_X1 U6995 ( .B1(n5987), .B2(n6007), .A(n5986), .ZN(U2912) );
  INV_X1 U6996 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5989) );
  AOI22_X1 U6997 ( .A1(n4378), .A2(LWORD_REG_10__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5988) );
  OAI21_X1 U6998 ( .B1(n5989), .B2(n6007), .A(n5988), .ZN(U2913) );
  INV_X1 U6999 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5991) );
  AOI22_X1 U7000 ( .A1(n4378), .A2(LWORD_REG_9__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5990) );
  OAI21_X1 U7001 ( .B1(n5991), .B2(n6007), .A(n5990), .ZN(U2914) );
  INV_X1 U7002 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5993) );
  AOI22_X1 U7003 ( .A1(n4378), .A2(LWORD_REG_8__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5992) );
  OAI21_X1 U7004 ( .B1(n5993), .B2(n6007), .A(n5992), .ZN(U2915) );
  AOI22_X1 U7005 ( .A1(n4378), .A2(LWORD_REG_7__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5994) );
  OAI21_X1 U7006 ( .B1(n5995), .B2(n6007), .A(n5994), .ZN(U2916) );
  AOI22_X1 U7007 ( .A1(n4378), .A2(LWORD_REG_6__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5996) );
  OAI21_X1 U7008 ( .B1(n3545), .B2(n6007), .A(n5996), .ZN(U2917) );
  AOI22_X1 U7009 ( .A1(n4378), .A2(LWORD_REG_5__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5997) );
  OAI21_X1 U7010 ( .B1(n3528), .B2(n6007), .A(n5997), .ZN(U2918) );
  AOI22_X1 U7011 ( .A1(n4378), .A2(LWORD_REG_4__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5998) );
  OAI21_X1 U7012 ( .B1(n5999), .B2(n6007), .A(n5998), .ZN(U2919) );
  AOI22_X1 U7013 ( .A1(n4378), .A2(LWORD_REG_3__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6000) );
  OAI21_X1 U7014 ( .B1(n6001), .B2(n6007), .A(n6000), .ZN(U2920) );
  AOI22_X1 U7015 ( .A1(n4378), .A2(LWORD_REG_2__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6002) );
  OAI21_X1 U7016 ( .B1(n6563), .B2(n6007), .A(n6002), .ZN(U2921) );
  AOI22_X1 U7017 ( .A1(n4378), .A2(LWORD_REG_1__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6003) );
  OAI21_X1 U7018 ( .B1(n6004), .B2(n6007), .A(n6003), .ZN(U2922) );
  AOI22_X1 U7019 ( .A1(n4378), .A2(LWORD_REG_0__SCAN_IN), .B1(n6005), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6006) );
  OAI21_X1 U7020 ( .B1(n6008), .B2(n6007), .A(n6006), .ZN(U2923) );
  AOI22_X1 U7021 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6022), .B1(n6026), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7022 ( .A1(n6025), .A2(DATAI_8_), .ZN(n6014) );
  NAND2_X1 U7023 ( .A1(n6009), .A2(n6014), .ZN(U2932) );
  AOI22_X1 U7024 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6022), .B1(n6026), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7025 ( .A1(n6025), .A2(DATAI_9_), .ZN(n6016) );
  NAND2_X1 U7026 ( .A1(n6010), .A2(n6016), .ZN(U2933) );
  AOI22_X1 U7027 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6022), .B1(n6026), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7028 ( .A1(n6025), .A2(DATAI_10_), .ZN(n6018) );
  NAND2_X1 U7029 ( .A1(n6011), .A2(n6018), .ZN(U2934) );
  AOI22_X1 U7030 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6022), .B1(n6026), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7031 ( .A1(n6025), .A2(DATAI_11_), .ZN(n6020) );
  NAND2_X1 U7032 ( .A1(n6012), .A2(n6020), .ZN(U2935) );
  AOI22_X1 U7033 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6022), .B1(n6026), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7034 ( .A1(n6025), .A2(DATAI_14_), .ZN(n6023) );
  NAND2_X1 U7035 ( .A1(n6013), .A2(n6023), .ZN(U2938) );
  AOI22_X1 U7036 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6022), .B1(n6026), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7037 ( .A1(n6015), .A2(n6014), .ZN(U2947) );
  AOI22_X1 U7038 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6022), .B1(n6026), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7039 ( .A1(n6017), .A2(n6016), .ZN(U2948) );
  AOI22_X1 U7040 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6022), .B1(n6026), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7041 ( .A1(n6019), .A2(n6018), .ZN(U2949) );
  AOI22_X1 U7042 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6022), .B1(n6026), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7043 ( .A1(n6021), .A2(n6020), .ZN(U2950) );
  AOI22_X1 U7044 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6022), .B1(n6026), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7045 ( .A1(n6024), .A2(n6023), .ZN(U2953) );
  AOI22_X1 U7046 ( .A1(n6026), .A2(LWORD_REG_15__SCAN_IN), .B1(n6025), .B2(
        DATAI_15_), .ZN(n6027) );
  OAI21_X1 U7047 ( .B1(n6671), .B2(n6028), .A(n6027), .ZN(U2954) );
  AOI22_X1 U7048 ( .A1(n6107), .A2(REIP_REG_2__SCAN_IN), .B1(n6048), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6038) );
  INV_X1 U7049 ( .A(n6029), .ZN(n6035) );
  AND2_X1 U7050 ( .A1(n6031), .A2(n6030), .ZN(n6033) );
  XNOR2_X1 U7051 ( .A(n6033), .B(n6032), .ZN(n6097) );
  AOI22_X1 U7052 ( .A1(n6036), .A2(n6035), .B1(n6097), .B2(n6034), .ZN(n6037)
         );
  OAI211_X1 U7053 ( .C1(n6040), .C2(n6039), .A(n6038), .B(n6037), .ZN(U2984)
         );
  INV_X1 U7054 ( .A(n6041), .ZN(n6044) );
  AOI211_X1 U7055 ( .C1(n6044), .C2(n6498), .A(n6043), .B(n6042), .ZN(n6046)
         );
  NOR2_X1 U7056 ( .A1(n6046), .A2(n6045), .ZN(n6050) );
  OAI21_X1 U7057 ( .B1(n6048), .B2(n6047), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6049) );
  OAI211_X1 U7058 ( .C1(n6052), .C2(n6051), .A(n6050), .B(n6049), .ZN(U2986)
         );
  AOI21_X1 U7059 ( .B1(n6109), .B2(n6054), .A(n6053), .ZN(n6058) );
  AOI22_X1 U7060 ( .A1(n6112), .A2(n6056), .B1(n6059), .B2(n6055), .ZN(n6057)
         );
  OAI211_X1 U7061 ( .C1(n6060), .C2(n6059), .A(n6058), .B(n6057), .ZN(U3007)
         );
  INV_X1 U7062 ( .A(n6061), .ZN(n6062) );
  AOI21_X1 U7063 ( .B1(n6109), .B2(n6063), .A(n6062), .ZN(n6067) );
  AOI22_X1 U7064 ( .A1(n6065), .A2(n6112), .B1(n6064), .B2(n6068), .ZN(n6066)
         );
  OAI211_X1 U7065 ( .C1(n6069), .C2(n6068), .A(n6067), .B(n6066), .ZN(U3009)
         );
  NAND2_X1 U7066 ( .A1(n6109), .A2(n6070), .ZN(n6072) );
  OAI211_X1 U7067 ( .C1(n6073), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6072), 
        .B(n6071), .ZN(n6074) );
  AOI21_X1 U7068 ( .B1(n6075), .B2(n6112), .A(n6074), .ZN(n6076) );
  OAI21_X1 U7069 ( .B1(n6078), .B2(n6077), .A(n6076), .ZN(U3011) );
  INV_X1 U7070 ( .A(n6079), .ZN(n6091) );
  OAI21_X1 U7071 ( .B1(n6082), .B2(n6081), .A(n6080), .ZN(n6083) );
  INV_X1 U7072 ( .A(n6083), .ZN(n6087) );
  OR2_X1 U7073 ( .A1(n6085), .A2(n6084), .ZN(n6086) );
  OAI211_X1 U7074 ( .C1(n6088), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6087), 
        .B(n6086), .ZN(n6089) );
  INV_X1 U7075 ( .A(n6089), .ZN(n6090) );
  OAI21_X1 U7076 ( .B1(n6091), .B2(n4222), .A(n6090), .ZN(U3015) );
  OAI21_X1 U7077 ( .B1(n6093), .B2(n4210), .A(n6092), .ZN(n6095) );
  AOI22_X1 U7078 ( .A1(n6096), .A2(n6095), .B1(n6109), .B2(n6094), .ZN(n6104)
         );
  AOI22_X1 U7079 ( .A1(n6098), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6112), 
        .B2(n6097), .ZN(n6103) );
  NAND2_X1 U7080 ( .A1(n6099), .A2(REIP_REG_2__SCAN_IN), .ZN(n6102) );
  NAND3_X1 U7081 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6100), .A3(n4210), 
        .ZN(n6101) );
  NAND4_X1 U7082 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(U3016)
         );
  NAND2_X1 U7083 ( .A1(n6106), .A2(n6105), .ZN(n6115) );
  AOI22_X1 U7084 ( .A1(n6109), .A2(n6108), .B1(n6107), .B2(REIP_REG_1__SCAN_IN), .ZN(n6114) );
  AOI22_X1 U7085 ( .A1(n6112), .A2(n6111), .B1(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .B2(n6110), .ZN(n6113) );
  OAI211_X1 U7086 ( .C1(INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n6115), .A(n6114), 
        .B(n6113), .ZN(U3017) );
  NOR2_X1 U7087 ( .A1(n6381), .A2(n6116), .ZN(U3019) );
  INV_X1 U7088 ( .A(n6117), .ZN(n6288) );
  OAI22_X1 U7089 ( .A1(n6176), .A2(n6121), .B1(n6120), .B2(n6119), .ZN(n6151)
         );
  NOR2_X1 U7090 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6122), .ZN(n6150)
         );
  AOI22_X1 U7091 ( .A1(n6286), .A2(n6151), .B1(n6285), .B2(n6150), .ZN(n6131)
         );
  INV_X1 U7092 ( .A(n6150), .ZN(n6124) );
  AOI211_X1 U7093 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6124), .A(n6174), .B(
        n6123), .ZN(n6129) );
  INV_X1 U7094 ( .A(n6344), .ZN(n6125) );
  OAI21_X1 U7095 ( .B1(n6152), .B2(n6125), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6127) );
  NAND3_X1 U7096 ( .A1(n6127), .A2(n6521), .A3(n6126), .ZN(n6128) );
  NAND2_X1 U7097 ( .A1(n6129), .A2(n6128), .ZN(n6153) );
  AOI22_X1 U7098 ( .A1(n6153), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n6205), 
        .B2(n6152), .ZN(n6130) );
  OAI211_X1 U7099 ( .C1(n6218), .C2(n6344), .A(n6131), .B(n6130), .ZN(U3020)
         );
  AOI22_X1 U7100 ( .A1(n6300), .A2(n6151), .B1(n6299), .B2(n6150), .ZN(n6133)
         );
  AOI22_X1 U7101 ( .A1(n6153), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n6253), 
        .B2(n6152), .ZN(n6132) );
  OAI211_X1 U7102 ( .C1(n6256), .C2(n6344), .A(n6133), .B(n6132), .ZN(U3021)
         );
  AOI22_X1 U7103 ( .A1(n6306), .A2(n6151), .B1(n6305), .B2(n6150), .ZN(n6135)
         );
  AOI22_X1 U7104 ( .A1(n6153), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n6257), 
        .B2(n6152), .ZN(n6134) );
  OAI211_X1 U7105 ( .C1(n6260), .C2(n6344), .A(n6135), .B(n6134), .ZN(U3022)
         );
  AOI22_X1 U7106 ( .A1(n6312), .A2(n6151), .B1(n6311), .B2(n6150), .ZN(n6137)
         );
  AOI22_X1 U7107 ( .A1(n6153), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n6262), 
        .B2(n6152), .ZN(n6136) );
  OAI211_X1 U7108 ( .C1(n6266), .C2(n6344), .A(n6137), .B(n6136), .ZN(U3023)
         );
  AOI22_X1 U7109 ( .A1(n6318), .A2(n6151), .B1(n6317), .B2(n6150), .ZN(n6140)
         );
  AOI22_X1 U7110 ( .A1(n6153), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n6138), 
        .B2(n6152), .ZN(n6139) );
  OAI211_X1 U7111 ( .C1(n6141), .C2(n6344), .A(n6140), .B(n6139), .ZN(U3024)
         );
  AOI22_X1 U7112 ( .A1(n6324), .A2(n6151), .B1(n6323), .B2(n6150), .ZN(n6144)
         );
  AOI22_X1 U7113 ( .A1(n6153), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n6142), 
        .B2(n6152), .ZN(n6143) );
  OAI211_X1 U7114 ( .C1(n6145), .C2(n6344), .A(n6144), .B(n6143), .ZN(U3025)
         );
  AOI22_X1 U7115 ( .A1(n6330), .A2(n6151), .B1(n6329), .B2(n6150), .ZN(n6148)
         );
  AOI22_X1 U7116 ( .A1(n6153), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n6146), 
        .B2(n6152), .ZN(n6147) );
  OAI211_X1 U7117 ( .C1(n6149), .C2(n6344), .A(n6148), .B(n6147), .ZN(U3026)
         );
  AOI22_X1 U7118 ( .A1(n6338), .A2(n6151), .B1(n6335), .B2(n6150), .ZN(n6155)
         );
  AOI22_X1 U7119 ( .A1(n6153), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n6234), 
        .B2(n6152), .ZN(n6154) );
  OAI211_X1 U7120 ( .C1(n6241), .C2(n6344), .A(n6155), .B(n6154), .ZN(U3027)
         );
  AOI22_X1 U7121 ( .A1(n6305), .A2(n6165), .B1(n6307), .B2(n6164), .ZN(n6157)
         );
  AOI22_X1 U7122 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6167), .B1(n6306), 
        .B2(n6166), .ZN(n6156) );
  OAI211_X1 U7123 ( .C1(n6310), .C2(n6170), .A(n6157), .B(n6156), .ZN(U3046)
         );
  AOI22_X1 U7124 ( .A1(n6317), .A2(n6165), .B1(n6319), .B2(n6164), .ZN(n6159)
         );
  AOI22_X1 U7125 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6167), .B1(n6318), 
        .B2(n6166), .ZN(n6158) );
  OAI211_X1 U7126 ( .C1(n6322), .C2(n6170), .A(n6159), .B(n6158), .ZN(U3048)
         );
  AOI22_X1 U7127 ( .A1(n6323), .A2(n6165), .B1(n6325), .B2(n6164), .ZN(n6161)
         );
  AOI22_X1 U7128 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6167), .B1(n6324), 
        .B2(n6166), .ZN(n6160) );
  OAI211_X1 U7129 ( .C1(n6328), .C2(n6170), .A(n6161), .B(n6160), .ZN(U3049)
         );
  AOI22_X1 U7130 ( .A1(n6329), .A2(n6165), .B1(n6331), .B2(n6164), .ZN(n6163)
         );
  AOI22_X1 U7131 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6167), .B1(n6330), 
        .B2(n6166), .ZN(n6162) );
  OAI211_X1 U7132 ( .C1(n6334), .C2(n6170), .A(n6163), .B(n6162), .ZN(U3050)
         );
  AOI22_X1 U7133 ( .A1(n6335), .A2(n6165), .B1(n6340), .B2(n6164), .ZN(n6169)
         );
  AOI22_X1 U7134 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6167), .B1(n6338), 
        .B2(n6166), .ZN(n6168) );
  OAI211_X1 U7135 ( .C1(n6345), .C2(n6170), .A(n6169), .B(n6168), .ZN(U3051)
         );
  NAND2_X1 U7136 ( .A1(n6172), .A2(n6171), .ZN(n6240) );
  NAND3_X1 U7137 ( .A1(n6174), .A2(n6173), .A3(n6382), .ZN(n6175) );
  OAI21_X1 U7138 ( .B1(n6208), .B2(n6176), .A(n6175), .ZN(n6199) );
  NOR2_X1 U7139 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6213), .ZN(n6198)
         );
  AOI22_X1 U7140 ( .A1(n6286), .A2(n6199), .B1(n6285), .B2(n6198), .ZN(n6185)
         );
  INV_X1 U7141 ( .A(n6240), .ZN(n6229) );
  NOR2_X1 U7142 ( .A1(n6229), .A2(n6284), .ZN(n6178) );
  AOI21_X1 U7143 ( .B1(n6178), .B2(n6177), .A(n6290), .ZN(n6183) );
  INV_X1 U7144 ( .A(n6198), .ZN(n6181) );
  AOI211_X1 U7145 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6181), .A(n6180), .B(
        n6179), .ZN(n6182) );
  OAI211_X1 U7146 ( .C1(n6281), .C2(n6183), .A(n6182), .B(n6382), .ZN(n6201)
         );
  AOI22_X1 U7147 ( .A1(n6201), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6295), 
        .B2(n6200), .ZN(n6184) );
  OAI211_X1 U7148 ( .C1(n6298), .C2(n6240), .A(n6185), .B(n6184), .ZN(U3068)
         );
  AOI22_X1 U7149 ( .A1(n6300), .A2(n6199), .B1(n6299), .B2(n6198), .ZN(n6187)
         );
  AOI22_X1 U7150 ( .A1(n6201), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6301), 
        .B2(n6200), .ZN(n6186) );
  OAI211_X1 U7151 ( .C1(n6304), .C2(n6240), .A(n6187), .B(n6186), .ZN(U3069)
         );
  AOI22_X1 U7152 ( .A1(n6306), .A2(n6199), .B1(n6305), .B2(n6198), .ZN(n6189)
         );
  AOI22_X1 U7153 ( .A1(n6201), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6307), 
        .B2(n6200), .ZN(n6188) );
  OAI211_X1 U7154 ( .C1(n6310), .C2(n6240), .A(n6189), .B(n6188), .ZN(U3070)
         );
  AOI22_X1 U7155 ( .A1(n6312), .A2(n6199), .B1(n6311), .B2(n6198), .ZN(n6191)
         );
  AOI22_X1 U7156 ( .A1(n6201), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6313), 
        .B2(n6200), .ZN(n6190) );
  OAI211_X1 U7157 ( .C1(n6316), .C2(n6240), .A(n6191), .B(n6190), .ZN(U3071)
         );
  AOI22_X1 U7158 ( .A1(n6318), .A2(n6199), .B1(n6317), .B2(n6198), .ZN(n6193)
         );
  AOI22_X1 U7159 ( .A1(n6201), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6319), 
        .B2(n6200), .ZN(n6192) );
  OAI211_X1 U7160 ( .C1(n6322), .C2(n6240), .A(n6193), .B(n6192), .ZN(U3072)
         );
  AOI22_X1 U7161 ( .A1(n6324), .A2(n6199), .B1(n6323), .B2(n6198), .ZN(n6195)
         );
  AOI22_X1 U7162 ( .A1(n6201), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6325), 
        .B2(n6200), .ZN(n6194) );
  OAI211_X1 U7163 ( .C1(n6328), .C2(n6240), .A(n6195), .B(n6194), .ZN(U3073)
         );
  AOI22_X1 U7164 ( .A1(n6330), .A2(n6199), .B1(n6329), .B2(n6198), .ZN(n6197)
         );
  AOI22_X1 U7165 ( .A1(n6201), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6331), 
        .B2(n6200), .ZN(n6196) );
  OAI211_X1 U7166 ( .C1(n6334), .C2(n6240), .A(n6197), .B(n6196), .ZN(U3074)
         );
  AOI22_X1 U7167 ( .A1(n6338), .A2(n6199), .B1(n6335), .B2(n6198), .ZN(n6203)
         );
  AOI22_X1 U7168 ( .A1(n6201), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6340), 
        .B2(n6200), .ZN(n6202) );
  OAI211_X1 U7169 ( .C1(n6345), .C2(n6240), .A(n6203), .B(n6202), .ZN(U3075)
         );
  INV_X1 U7170 ( .A(n6204), .ZN(n6235) );
  AOI22_X1 U7171 ( .A1(n6285), .A2(n6235), .B1(n6205), .B2(n6233), .ZN(n6217)
         );
  NOR3_X1 U7172 ( .A1(n6208), .A2(n6207), .A3(n6206), .ZN(n6209) );
  NOR2_X1 U7173 ( .A1(n6209), .A2(n6235), .ZN(n6215) );
  AND2_X1 U7174 ( .A1(n6210), .A2(n6521), .ZN(n6212) );
  AOI22_X1 U7175 ( .A1(n6215), .A2(n6212), .B1(n6213), .B2(n6284), .ZN(n6211)
         );
  NAND2_X1 U7176 ( .A1(n6293), .A2(n6211), .ZN(n6237) );
  INV_X1 U7177 ( .A(n6212), .ZN(n6214) );
  OAI22_X1 U7178 ( .A1(n6215), .A2(n6214), .B1(n6393), .B2(n6213), .ZN(n6236)
         );
  AOI22_X1 U7179 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6237), .B1(n6286), 
        .B2(n6236), .ZN(n6216) );
  OAI211_X1 U7180 ( .C1(n6218), .C2(n6240), .A(n6217), .B(n6216), .ZN(U3076)
         );
  AOI22_X1 U7181 ( .A1(n6299), .A2(n6235), .B1(n6253), .B2(n6233), .ZN(n6220)
         );
  AOI22_X1 U7182 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6237), .B1(n6300), 
        .B2(n6236), .ZN(n6219) );
  OAI211_X1 U7183 ( .C1(n6256), .C2(n6240), .A(n6220), .B(n6219), .ZN(U3077)
         );
  AOI22_X1 U7184 ( .A1(n6305), .A2(n6235), .B1(n6307), .B2(n6229), .ZN(n6222)
         );
  AOI22_X1 U7185 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6237), .B1(n6306), 
        .B2(n6236), .ZN(n6221) );
  OAI211_X1 U7186 ( .C1(n6310), .C2(n6232), .A(n6222), .B(n6221), .ZN(U3078)
         );
  AOI22_X1 U7187 ( .A1(n6311), .A2(n6235), .B1(n6262), .B2(n6233), .ZN(n6224)
         );
  AOI22_X1 U7188 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6237), .B1(n6312), 
        .B2(n6236), .ZN(n6223) );
  OAI211_X1 U7189 ( .C1(n6266), .C2(n6240), .A(n6224), .B(n6223), .ZN(U3079)
         );
  AOI22_X1 U7190 ( .A1(n6317), .A2(n6235), .B1(n6319), .B2(n6229), .ZN(n6226)
         );
  AOI22_X1 U7191 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6237), .B1(n6318), 
        .B2(n6236), .ZN(n6225) );
  OAI211_X1 U7192 ( .C1(n6322), .C2(n6232), .A(n6226), .B(n6225), .ZN(U3080)
         );
  AOI22_X1 U7193 ( .A1(n6323), .A2(n6235), .B1(n6325), .B2(n6229), .ZN(n6228)
         );
  AOI22_X1 U7194 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6237), .B1(n6324), 
        .B2(n6236), .ZN(n6227) );
  OAI211_X1 U7195 ( .C1(n6328), .C2(n6232), .A(n6228), .B(n6227), .ZN(U3081)
         );
  AOI22_X1 U7196 ( .A1(n6329), .A2(n6235), .B1(n6331), .B2(n6229), .ZN(n6231)
         );
  AOI22_X1 U7197 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6237), .B1(n6330), 
        .B2(n6236), .ZN(n6230) );
  OAI211_X1 U7198 ( .C1(n6334), .C2(n6232), .A(n6231), .B(n6230), .ZN(U3082)
         );
  AOI22_X1 U7199 ( .A1(n6335), .A2(n6235), .B1(n6234), .B2(n6233), .ZN(n6239)
         );
  AOI22_X1 U7200 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6237), .B1(n6338), 
        .B2(n6236), .ZN(n6238) );
  OAI211_X1 U7201 ( .C1(n6241), .C2(n6240), .A(n6239), .B(n6238), .ZN(U3083)
         );
  NOR2_X1 U7202 ( .A1(n6242), .A2(n6382), .ZN(n6274) );
  AOI22_X1 U7203 ( .A1(n6285), .A2(n6274), .B1(n6295), .B2(n6273), .ZN(n6252)
         );
  AOI21_X1 U7204 ( .B1(n6244), .B2(n6243), .A(n6284), .ZN(n6247) );
  AOI21_X1 U7205 ( .B1(n6245), .B2(n6365), .A(n6274), .ZN(n6249) );
  AOI22_X1 U7206 ( .A1(n6247), .A2(n6249), .B1(n6248), .B2(n6284), .ZN(n6246)
         );
  NAND2_X1 U7207 ( .A1(n6293), .A2(n6246), .ZN(n6276) );
  INV_X1 U7208 ( .A(n6247), .ZN(n6250) );
  OAI22_X1 U7209 ( .A1(n6250), .A2(n6249), .B1(n6248), .B2(n6393), .ZN(n6275)
         );
  AOI22_X1 U7210 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6276), .B1(n6286), 
        .B2(n6275), .ZN(n6251) );
  OAI211_X1 U7211 ( .C1(n6298), .C2(n6279), .A(n6252), .B(n6251), .ZN(U3108)
         );
  AOI22_X1 U7212 ( .A1(n6299), .A2(n6274), .B1(n6253), .B2(n6261), .ZN(n6255)
         );
  AOI22_X1 U7213 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6276), .B1(n6300), 
        .B2(n6275), .ZN(n6254) );
  OAI211_X1 U7214 ( .C1(n6256), .C2(n6265), .A(n6255), .B(n6254), .ZN(U3109)
         );
  AOI22_X1 U7215 ( .A1(n6305), .A2(n6274), .B1(n6257), .B2(n6261), .ZN(n6259)
         );
  AOI22_X1 U7216 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6276), .B1(n6306), 
        .B2(n6275), .ZN(n6258) );
  OAI211_X1 U7217 ( .C1(n6260), .C2(n6265), .A(n6259), .B(n6258), .ZN(U3110)
         );
  AOI22_X1 U7218 ( .A1(n6311), .A2(n6274), .B1(n6262), .B2(n6261), .ZN(n6264)
         );
  AOI22_X1 U7219 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6276), .B1(n6312), 
        .B2(n6275), .ZN(n6263) );
  OAI211_X1 U7220 ( .C1(n6266), .C2(n6265), .A(n6264), .B(n6263), .ZN(U3111)
         );
  AOI22_X1 U7221 ( .A1(n6317), .A2(n6274), .B1(n6319), .B2(n6273), .ZN(n6268)
         );
  AOI22_X1 U7222 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6276), .B1(n6318), 
        .B2(n6275), .ZN(n6267) );
  OAI211_X1 U7223 ( .C1(n6322), .C2(n6279), .A(n6268), .B(n6267), .ZN(U3112)
         );
  AOI22_X1 U7224 ( .A1(n6323), .A2(n6274), .B1(n6325), .B2(n6273), .ZN(n6270)
         );
  AOI22_X1 U7225 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6276), .B1(n6324), 
        .B2(n6275), .ZN(n6269) );
  OAI211_X1 U7226 ( .C1(n6328), .C2(n6279), .A(n6270), .B(n6269), .ZN(U3113)
         );
  AOI22_X1 U7227 ( .A1(n6329), .A2(n6274), .B1(n6331), .B2(n6273), .ZN(n6272)
         );
  AOI22_X1 U7228 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6276), .B1(n6330), 
        .B2(n6275), .ZN(n6271) );
  OAI211_X1 U7229 ( .C1(n6334), .C2(n6279), .A(n6272), .B(n6271), .ZN(U3114)
         );
  AOI22_X1 U7230 ( .A1(n6335), .A2(n6274), .B1(n6340), .B2(n6273), .ZN(n6278)
         );
  AOI22_X1 U7231 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6276), .B1(n6338), 
        .B2(n6275), .ZN(n6277) );
  OAI211_X1 U7232 ( .C1(n6345), .C2(n6279), .A(n6278), .B(n6277), .ZN(U3115)
         );
  INV_X1 U7233 ( .A(n6280), .ZN(n6336) );
  AOI21_X1 U7234 ( .B1(n6282), .B2(n6281), .A(n6336), .ZN(n6289) );
  OAI22_X1 U7235 ( .A1(n6289), .A2(n6284), .B1(n6393), .B2(n6283), .ZN(n6337)
         );
  AOI22_X1 U7236 ( .A1(n6286), .A2(n6337), .B1(n6336), .B2(n6285), .ZN(n6297)
         );
  AOI21_X1 U7237 ( .B1(n6288), .B2(n4300), .A(n6287), .ZN(n6291) );
  OAI21_X1 U7238 ( .B1(n6291), .B2(n6290), .A(n6289), .ZN(n6292) );
  OAI211_X1 U7239 ( .C1(n6294), .C2(n6521), .A(n6293), .B(n6292), .ZN(n6341)
         );
  AOI22_X1 U7240 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6341), .B1(n6295), 
        .B2(n6339), .ZN(n6296) );
  OAI211_X1 U7241 ( .C1(n6298), .C2(n6344), .A(n6297), .B(n6296), .ZN(U3140)
         );
  AOI22_X1 U7242 ( .A1(n6300), .A2(n6337), .B1(n6336), .B2(n6299), .ZN(n6303)
         );
  AOI22_X1 U7243 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6341), .B1(n6301), 
        .B2(n6339), .ZN(n6302) );
  OAI211_X1 U7244 ( .C1(n6304), .C2(n6344), .A(n6303), .B(n6302), .ZN(U3141)
         );
  AOI22_X1 U7245 ( .A1(n6306), .A2(n6337), .B1(n6336), .B2(n6305), .ZN(n6309)
         );
  AOI22_X1 U7246 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6341), .B1(n6307), 
        .B2(n6339), .ZN(n6308) );
  OAI211_X1 U7247 ( .C1(n6310), .C2(n6344), .A(n6309), .B(n6308), .ZN(U3142)
         );
  AOI22_X1 U7248 ( .A1(n6312), .A2(n6337), .B1(n6336), .B2(n6311), .ZN(n6315)
         );
  AOI22_X1 U7249 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6341), .B1(n6313), 
        .B2(n6339), .ZN(n6314) );
  OAI211_X1 U7250 ( .C1(n6316), .C2(n6344), .A(n6315), .B(n6314), .ZN(U3143)
         );
  AOI22_X1 U7251 ( .A1(n6318), .A2(n6337), .B1(n6336), .B2(n6317), .ZN(n6321)
         );
  AOI22_X1 U7252 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6341), .B1(n6319), 
        .B2(n6339), .ZN(n6320) );
  OAI211_X1 U7253 ( .C1(n6322), .C2(n6344), .A(n6321), .B(n6320), .ZN(U3144)
         );
  AOI22_X1 U7254 ( .A1(n6324), .A2(n6337), .B1(n6336), .B2(n6323), .ZN(n6327)
         );
  AOI22_X1 U7255 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6341), .B1(n6325), 
        .B2(n6339), .ZN(n6326) );
  OAI211_X1 U7256 ( .C1(n6328), .C2(n6344), .A(n6327), .B(n6326), .ZN(U3145)
         );
  AOI22_X1 U7257 ( .A1(n6330), .A2(n6337), .B1(n6336), .B2(n6329), .ZN(n6333)
         );
  AOI22_X1 U7258 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6341), .B1(n6331), 
        .B2(n6339), .ZN(n6332) );
  OAI211_X1 U7259 ( .C1(n6334), .C2(n6344), .A(n6333), .B(n6332), .ZN(U3146)
         );
  AOI22_X1 U7260 ( .A1(n6338), .A2(n6337), .B1(n6336), .B2(n6335), .ZN(n6343)
         );
  AOI22_X1 U7261 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6341), .B1(n6340), 
        .B2(n6339), .ZN(n6342) );
  OAI211_X1 U7262 ( .C1(n6345), .C2(n6344), .A(n6343), .B(n6342), .ZN(U3147)
         );
  NAND2_X1 U7263 ( .A1(n6359), .A2(n6346), .ZN(n6347) );
  NOR2_X1 U7264 ( .A1(n6348), .A2(n6347), .ZN(n6355) );
  INV_X1 U7265 ( .A(n6349), .ZN(n6350) );
  OR2_X1 U7266 ( .A1(n6351), .A2(n6350), .ZN(n6354) );
  NAND2_X1 U7267 ( .A1(n6394), .A2(n6352), .ZN(n6353) );
  OAI211_X1 U7268 ( .C1(n6394), .C2(n6355), .A(n6354), .B(n6353), .ZN(n6356)
         );
  INV_X1 U7269 ( .A(n6356), .ZN(n6518) );
  OAI21_X1 U7270 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6357), 
        .ZN(n6358) );
  NAND4_X1 U7271 ( .A1(n6360), .A2(n6518), .A3(n6359), .A4(n6358), .ZN(n6362)
         );
  NOR2_X1 U7272 ( .A1(n6362), .A2(n6361), .ZN(n6387) );
  INV_X1 U7273 ( .A(n6363), .ZN(n6378) );
  NAND2_X1 U7274 ( .A1(n6365), .A2(n6364), .ZN(n6368) );
  OR2_X1 U7275 ( .A1(n6366), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6367)
         );
  NAND2_X1 U7276 ( .A1(n6368), .A2(n6367), .ZN(n6496) );
  NAND2_X1 U7277 ( .A1(n6369), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U7278 ( .A1(n6505), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6370) );
  OR2_X1 U7279 ( .A1(n6496), .A2(n6370), .ZN(n6373) );
  OAI21_X1 U7280 ( .B1(n6373), .B2(n6374), .A(n6371), .ZN(n6372) );
  INV_X1 U7281 ( .A(n6372), .ZN(n6375) );
  AOI22_X1 U7282 ( .A1(n6376), .A2(n6375), .B1(n6374), .B2(n6373), .ZN(n6377)
         );
  OAI21_X1 U7283 ( .B1(n6378), .B2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n6377), 
        .ZN(n6380) );
  NAND2_X1 U7284 ( .A1(n6378), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6379) );
  AOI22_X1 U7285 ( .A1(n6380), .A2(n6379), .B1(n6382), .B2(n6383), .ZN(n6385)
         );
  OAI21_X1 U7286 ( .B1(n6383), .B2(n6382), .A(n6381), .ZN(n6384) );
  OR2_X1 U7287 ( .A1(n6385), .A2(n6384), .ZN(n6386) );
  NAND2_X1 U7288 ( .A1(n6387), .A2(n6386), .ZN(n6398) );
  NAND2_X1 U7289 ( .A1(READY_N), .A2(n4378), .ZN(n6388) );
  OAI21_X1 U7290 ( .B1(n6398), .B2(n6406), .A(n6388), .ZN(n6392) );
  OR2_X1 U7291 ( .A1(n6390), .A2(n6389), .ZN(n6391) );
  AOI21_X1 U7292 ( .B1(READY_N), .B2(n6393), .A(n6486), .ZN(n6404) );
  NOR2_X1 U7293 ( .A1(n6490), .A2(n6410), .ZN(n6395) );
  AOI211_X1 U7294 ( .C1(n6395), .C2(n6394), .A(STATE2_REG_0__SCAN_IN), .B(
        n6486), .ZN(n6396) );
  AOI211_X1 U7295 ( .C1(n6399), .C2(n6398), .A(n6397), .B(n6396), .ZN(n6400)
         );
  OAI221_X1 U7296 ( .B1(n6402), .B2(n6404), .C1(n6402), .C2(n6401), .A(n6400), 
        .ZN(U3148) );
  NOR2_X1 U7297 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6413) );
  NOR3_X1 U7298 ( .A1(n6413), .A2(n6404), .A3(n6403), .ZN(n6408) );
  AOI221_X1 U7299 ( .B1(READY_N), .B2(n6406), .C1(n6405), .C2(n6406), .A(n6486), .ZN(n6407) );
  OR3_X1 U7300 ( .A1(n6409), .A2(n6408), .A3(n6407), .ZN(U3149) );
  OAI211_X1 U7301 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6572), .A(n6487), .B(
        n6410), .ZN(n6412) );
  OAI21_X1 U7302 ( .B1(n6413), .B2(n6412), .A(n6411), .ZN(U3150) );
  AND2_X1 U7303 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6683), .ZN(U3151) );
  AND2_X1 U7304 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6683), .ZN(U3152) );
  AND2_X1 U7305 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6683), .ZN(U3153) );
  AND2_X1 U7306 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6683), .ZN(U3154) );
  AND2_X1 U7307 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6683), .ZN(U3155) );
  AND2_X1 U7308 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6683), .ZN(U3156) );
  AND2_X1 U7309 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6683), .ZN(U3157) );
  AND2_X1 U7310 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6683), .ZN(U3158) );
  AND2_X1 U7311 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6683), .ZN(U3159) );
  AND2_X1 U7312 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6683), .ZN(U3160) );
  INV_X1 U7313 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6574) );
  NOR2_X1 U7314 ( .A1(n6485), .A2(n6574), .ZN(U3161) );
  AND2_X1 U7315 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6683), .ZN(U3162) );
  AND2_X1 U7316 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6683), .ZN(U3163) );
  AND2_X1 U7317 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6683), .ZN(U3164) );
  AND2_X1 U7318 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6683), .ZN(U3165) );
  AND2_X1 U7319 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6683), .ZN(U3166) );
  INV_X1 U7320 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6590) );
  NOR2_X1 U7321 ( .A1(n6485), .A2(n6590), .ZN(U3167) );
  AND2_X1 U7322 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6683), .ZN(U3168) );
  AND2_X1 U7323 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6683), .ZN(U3169) );
  AND2_X1 U7324 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6683), .ZN(U3170) );
  AND2_X1 U7325 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6683), .ZN(U3171) );
  NOR2_X1 U7326 ( .A1(n6485), .A2(n6626), .ZN(U3172) );
  AND2_X1 U7327 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6683), .ZN(U3173) );
  AND2_X1 U7328 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6683), .ZN(U3174) );
  AND2_X1 U7329 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6683), .ZN(U3175) );
  AND2_X1 U7330 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6683), .ZN(U3177) );
  AND2_X1 U7331 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6683), .ZN(U3178) );
  AND2_X1 U7332 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6683), .ZN(U3179) );
  NOR2_X1 U7333 ( .A1(n6485), .A2(n6623), .ZN(U3180) );
  INV_X1 U7334 ( .A(n6414), .ZN(n6423) );
  AOI22_X1 U7335 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6427) );
  AND2_X1 U7336 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6418) );
  INV_X1 U7337 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6416) );
  INV_X1 U7338 ( .A(NA_N), .ZN(n6424) );
  AOI211_X1 U7339 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6424), .A(
        STATE_REG_0__SCAN_IN), .B(n6423), .ZN(n6429) );
  AOI221_X1 U7340 ( .B1(n6418), .B2(n6531), .C1(n6416), .C2(n6531), .A(n6429), 
        .ZN(n6415) );
  OAI21_X1 U7341 ( .B1(n6423), .B2(n6427), .A(n6415), .ZN(U3181) );
  INV_X1 U7342 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6620) );
  NOR2_X1 U7343 ( .A1(n6620), .A2(n6416), .ZN(n6425) );
  NAND2_X1 U7344 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6417) );
  OAI21_X1 U7345 ( .B1(n6425), .B2(n6418), .A(n6417), .ZN(n6419) );
  OAI211_X1 U7346 ( .C1(n6421), .C2(n6572), .A(n6420), .B(n6419), .ZN(U3182)
         );
  AOI221_X1 U7347 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6572), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6422) );
  AOI221_X1 U7348 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6422), .C2(HOLD), .A(n6620), .ZN(n6428) );
  AOI21_X1 U7349 ( .B1(n6425), .B2(n6424), .A(n6423), .ZN(n6426) );
  OAI22_X1 U7350 ( .A1(n6429), .A2(n6428), .B1(n6427), .B2(n6426), .ZN(U3183)
         );
  AND2_X1 U7351 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6481), .ZN(n6477) );
  INV_X1 U7352 ( .A(n6477), .ZN(n6475) );
  NOR2_X1 U7353 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6531), .ZN(n6473) );
  AOI22_X1 U7354 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6473), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6531), .ZN(n6430) );
  OAI21_X1 U7355 ( .B1(n6506), .B2(n6475), .A(n6430), .ZN(U3184) );
  CLKBUF_X1 U7356 ( .A(n6473), .Z(n6469) );
  AOI222_X1 U7357 ( .A1(n6477), .A2(REIP_REG_2__SCAN_IN), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6531), .C1(REIP_REG_3__SCAN_IN), .C2(
        n6469), .ZN(n6431) );
  INV_X1 U7358 ( .A(n6431), .ZN(U3185) );
  AOI22_X1 U7359 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6469), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6531), .ZN(n6432) );
  OAI21_X1 U7360 ( .B1(n6433), .B2(n6475), .A(n6432), .ZN(U3186) );
  INV_X1 U7361 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6656) );
  INV_X1 U7362 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6436) );
  INV_X1 U7363 ( .A(n6473), .ZN(n6479) );
  OAI222_X1 U7364 ( .A1(n6475), .A2(n6434), .B1(n6656), .B2(n6481), .C1(n6436), 
        .C2(n6479), .ZN(U3187) );
  AOI22_X1 U7365 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6469), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6531), .ZN(n6435) );
  OAI21_X1 U7366 ( .B1(n6436), .B2(n6475), .A(n6435), .ZN(U3188) );
  AOI22_X1 U7367 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6469), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6531), .ZN(n6437) );
  OAI21_X1 U7368 ( .B1(n6438), .B2(n6475), .A(n6437), .ZN(U3189) );
  AOI22_X1 U7369 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6473), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6531), .ZN(n6439) );
  OAI21_X1 U7370 ( .B1(n6440), .B2(n6475), .A(n6439), .ZN(U3190) );
  INV_X1 U7371 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6584) );
  INV_X1 U7372 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6443) );
  OAI222_X1 U7373 ( .A1(n6475), .A2(n6441), .B1(n6584), .B2(n6481), .C1(n6443), 
        .C2(n6479), .ZN(U3191) );
  AOI22_X1 U7374 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6473), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6531), .ZN(n6442) );
  OAI21_X1 U7375 ( .B1(n6443), .B2(n6475), .A(n6442), .ZN(U3192) );
  AOI22_X1 U7376 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6473), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6531), .ZN(n6444) );
  OAI21_X1 U7377 ( .B1(n6445), .B2(n6475), .A(n6444), .ZN(U3193) );
  AOI22_X1 U7378 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6469), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6531), .ZN(n6446) );
  OAI21_X1 U7379 ( .B1(n4998), .B2(n6475), .A(n6446), .ZN(U3194) );
  INV_X1 U7380 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6618) );
  OAI222_X1 U7381 ( .A1(n6475), .A2(n6447), .B1(n6618), .B2(n6481), .C1(n6449), 
        .C2(n6479), .ZN(U3195) );
  AOI22_X1 U7382 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6469), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6531), .ZN(n6448) );
  OAI21_X1 U7383 ( .B1(n6449), .B2(n6475), .A(n6448), .ZN(U3196) );
  AOI22_X1 U7384 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6469), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6531), .ZN(n6450) );
  OAI21_X1 U7385 ( .B1(n6451), .B2(n6475), .A(n6450), .ZN(U3197) );
  AOI22_X1 U7386 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6473), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6531), .ZN(n6452) );
  OAI21_X1 U7387 ( .B1(n6453), .B2(n6475), .A(n6452), .ZN(U3198) );
  AOI22_X1 U7388 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6469), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6531), .ZN(n6454) );
  OAI21_X1 U7389 ( .B1(n5126), .B2(n6475), .A(n6454), .ZN(U3199) );
  AOI22_X1 U7390 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6477), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6531), .ZN(n6455) );
  OAI21_X1 U7391 ( .B1(n6457), .B2(n6479), .A(n6455), .ZN(U3200) );
  AOI22_X1 U7392 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6469), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6531), .ZN(n6456) );
  OAI21_X1 U7393 ( .B1(n6457), .B2(n6475), .A(n6456), .ZN(U3201) );
  INV_X1 U7394 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6577) );
  AOI22_X1 U7395 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6477), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6531), .ZN(n6458) );
  OAI21_X1 U7396 ( .B1(n6577), .B2(n6479), .A(n6458), .ZN(U3202) );
  AOI22_X1 U7397 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6473), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6531), .ZN(n6459) );
  OAI21_X1 U7398 ( .B1(n6577), .B2(n6475), .A(n6459), .ZN(U3203) );
  INV_X1 U7399 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6461) );
  AOI22_X1 U7400 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6473), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6531), .ZN(n6460) );
  OAI21_X1 U7401 ( .B1(n6461), .B2(n6475), .A(n6460), .ZN(U3204) );
  AOI22_X1 U7402 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6477), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6531), .ZN(n6462) );
  OAI21_X1 U7403 ( .B1(n6569), .B2(n6479), .A(n6462), .ZN(U3205) );
  AOI22_X1 U7404 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6473), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6531), .ZN(n6463) );
  OAI21_X1 U7405 ( .B1(n6569), .B2(n6475), .A(n6463), .ZN(U3206) );
  INV_X1 U7406 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6555) );
  OAI222_X1 U7407 ( .A1(n6479), .A2(n6466), .B1(n6555), .B2(n6481), .C1(n6464), 
        .C2(n6475), .ZN(U3207) );
  AOI22_X1 U7408 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6469), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6531), .ZN(n6465) );
  OAI21_X1 U7409 ( .B1(n6466), .B2(n6475), .A(n6465), .ZN(U3208) );
  AOI22_X1 U7410 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6469), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6531), .ZN(n6467) );
  OAI21_X1 U7411 ( .B1(n6468), .B2(n6475), .A(n6467), .ZN(U3209) );
  AOI22_X1 U7412 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6469), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6531), .ZN(n6470) );
  OAI21_X1 U7413 ( .B1(n6471), .B2(n6475), .A(n6470), .ZN(U3210) );
  AOI22_X1 U7414 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6477), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6531), .ZN(n6472) );
  OAI21_X1 U7415 ( .B1(n6476), .B2(n6479), .A(n6472), .ZN(U3211) );
  AOI22_X1 U7416 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6473), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6531), .ZN(n6474) );
  OAI21_X1 U7417 ( .B1(n6476), .B2(n6475), .A(n6474), .ZN(U3212) );
  INV_X1 U7418 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6480) );
  AOI22_X1 U7419 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6477), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6531), .ZN(n6478) );
  OAI21_X1 U7420 ( .B1(n6480), .B2(n6479), .A(n6478), .ZN(U3213) );
  MUX2_X1 U7421 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6531), .Z(U3445) );
  INV_X1 U7422 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6508) );
  INV_X1 U7423 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n6651) );
  AOI22_X1 U7424 ( .A1(n6481), .A2(n6508), .B1(n6651), .B2(n6531), .ZN(U3446)
         );
  MUX2_X1 U7425 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6531), .Z(U3447) );
  INV_X1 U7426 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6514) );
  INV_X1 U7427 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6653) );
  AOI22_X1 U7428 ( .A1(n6481), .A2(n6514), .B1(n6653), .B2(n6531), .ZN(U3448)
         );
  OAI21_X1 U7429 ( .B1(n6485), .B2(DATAWIDTH_REG_0__SCAN_IN), .A(n6483), .ZN(
        n6482) );
  INV_X1 U7430 ( .A(n6482), .ZN(U3451) );
  OAI21_X1 U7431 ( .B1(n6485), .B2(n6484), .A(n6483), .ZN(U3452) );
  INV_X1 U7432 ( .A(n6486), .ZN(n6489) );
  OAI211_X1 U7433 ( .C1(n6490), .C2(n6489), .A(n6488), .B(n6487), .ZN(U3453)
         );
  INV_X1 U7434 ( .A(n6491), .ZN(n6494) );
  OAI22_X1 U7435 ( .A1(n6494), .A2(n6504), .B1(n6493), .B2(n6492), .ZN(n6495)
         );
  MUX2_X1 U7436 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6495), .S(n6502), 
        .Z(U3456) );
  INV_X1 U7437 ( .A(n6496), .ZN(n6500) );
  AOI21_X1 U7438 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6498), .A(n6497), .ZN(
        n6499) );
  OAI211_X1 U7439 ( .C1(n6500), .C2(n6504), .A(n6502), .B(n6499), .ZN(n6501)
         );
  OAI21_X1 U7440 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6502), .A(n6501), 
        .ZN(n6503) );
  OAI21_X1 U7441 ( .B1(n6505), .B2(n6504), .A(n6503), .ZN(U3461) );
  AOI21_X1 U7442 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6507) );
  AOI22_X1 U7443 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6507), .B2(n6506), .ZN(n6509) );
  AOI22_X1 U7444 ( .A1(n6510), .A2(n6509), .B1(n6508), .B2(n6513), .ZN(U3468)
         );
  NOR2_X1 U7445 ( .A1(n6513), .A2(REIP_REG_1__SCAN_IN), .ZN(n6511) );
  AOI22_X1 U7446 ( .A1(n6514), .A2(n6513), .B1(n6512), .B2(n6511), .ZN(U3469)
         );
  NAND2_X1 U7447 ( .A1(n6531), .A2(W_R_N_REG_SCAN_IN), .ZN(n6515) );
  OAI21_X1 U7448 ( .B1(n6531), .B2(READREQUEST_REG_SCAN_IN), .A(n6515), .ZN(
        U3470) );
  INV_X1 U7449 ( .A(MORE_REG_SCAN_IN), .ZN(n6517) );
  INV_X1 U7450 ( .A(n6519), .ZN(n6516) );
  AOI22_X1 U7451 ( .A1(n6519), .A2(n6518), .B1(n6517), .B2(n6516), .ZN(U3471)
         );
  AOI211_X1 U7452 ( .C1(n4378), .C2(n6572), .A(n6521), .B(n6520), .ZN(n6522)
         );
  AND2_X1 U7453 ( .A1(n6523), .A2(n6522), .ZN(n6530) );
  OAI211_X1 U7454 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6525), .A(n6524), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6527) );
  AOI21_X1 U7455 ( .B1(n6527), .B2(STATE2_REG_0__SCAN_IN), .A(n6526), .ZN(
        n6529) );
  NAND2_X1 U7456 ( .A1(n6530), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6528) );
  OAI21_X1 U7457 ( .B1(n6530), .B2(n6529), .A(n6528), .ZN(U3472) );
  MUX2_X1 U7458 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6531), .Z(U3473) );
  NAND3_X1 U7459 ( .A1(LWORD_REG_14__SCAN_IN), .A2(BE_N_REG_2__SCAN_IN), .A3(
        n6560), .ZN(n6553) );
  NOR4_X1 U7460 ( .A1(EBX_REG_22__SCAN_IN), .A2(EBX_REG_1__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A4(REIP_REG_11__SCAN_IN), .ZN(n6534) );
  NOR4_X1 U7461 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(
        INSTQUEUE_REG_1__6__SCAN_IN), .A3(INSTQUEUE_REG_15__3__SCAN_IN), .A4(
        REIP_REG_20__SCAN_IN), .ZN(n6533) );
  NOR4_X1 U7462 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(REIP_REG_23__SCAN_IN), 
        .A3(DATAI_12_), .A4(DATAI_23_), .ZN(n6532) );
  NAND3_X1 U7463 ( .A1(n6534), .A2(n6533), .A3(n6532), .ZN(n6552) );
  NOR4_X1 U7464 ( .A1(UWORD_REG_0__SCAN_IN), .A2(LWORD_REG_10__SCAN_IN), .A3(
        BE_N_REG_0__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6550) );
  NOR4_X1 U7465 ( .A1(LWORD_REG_3__SCAN_IN), .A2(DATAO_REG_10__SCAN_IN), .A3(
        DATAO_REG_5__SCAN_IN), .A4(DATAO_REG_1__SCAN_IN), .ZN(n6536) );
  NOR4_X1 U7466 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(UWORD_REG_14__SCAN_IN), .A3(DATAO_REG_18__SCAN_IN), .A4(DATAO_REG_17__SCAN_IN), .ZN(n6535) );
  AND4_X1 U7467 ( .A1(n6538), .A2(n6537), .A3(n6536), .A4(n6535), .ZN(n6549)
         );
  NAND4_X1 U7468 ( .A1(ADDRESS_REG_11__SCAN_IN), .A2(ADDRESS_REG_3__SCAN_IN), 
        .A3(ADDRESS_REG_7__SCAN_IN), .A4(ADDRESS_REG_23__SCAN_IN), .ZN(n6542)
         );
  NAND4_X1 U7469 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(D_C_N_REG_SCAN_IN), 
        .A3(BYTEENABLE_REG_3__SCAN_IN), .A4(ADDRESS_REG_1__SCAN_IN), .ZN(n6541) );
  NAND4_X1 U7470 ( .A1(STATE_REG_0__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .A3(EAX_REG_2__SCAN_IN), .A4(
        EAX_REG_5__SCAN_IN), .ZN(n6540) );
  NAND4_X1 U7471 ( .A1(UWORD_REG_3__SCAN_IN), .A2(DATAO_REG_30__SCAN_IN), .A3(
        DATAO_REG_3__SCAN_IN), .A4(DATAO_REG_2__SCAN_IN), .ZN(n6539) );
  NOR4_X1 U7472 ( .A1(n6542), .A2(n6541), .A3(n6540), .A4(n6539), .ZN(n6548)
         );
  NAND4_X1 U7473 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(
        INSTQUEUE_REG_14__2__SCAN_IN), .A3(PHYADDRPOINTER_REG_17__SCAN_IN), 
        .A4(EAX_REG_15__SCAN_IN), .ZN(n6546) );
  NAND4_X1 U7474 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(
        INSTQUEUE_REG_4__5__SCAN_IN), .A3(INSTQUEUE_REG_12__5__SCAN_IN), .A4(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6545) );
  NAND4_X1 U7475 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        INSTQUEUE_REG_3__5__SCAN_IN), .A3(INSTQUEUE_REG_8__6__SCAN_IN), .A4(
        INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6544) );
  NAND4_X1 U7476 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(
        INSTQUEUE_REG_0__7__SCAN_IN), .A3(REIP_REG_28__SCAN_IN), .A4(DATAI_31_), .ZN(n6543) );
  NOR4_X1 U7477 ( .A1(n6546), .A2(n6545), .A3(n6544), .A4(n6543), .ZN(n6547)
         );
  NAND4_X1 U7478 ( .A1(n6550), .A2(n6549), .A3(n6548), .A4(n6547), .ZN(n6551)
         );
  NOR4_X1 U7479 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n6553), .A3(n6552), 
        .A4(n6551), .ZN(n6687) );
  AOI22_X1 U7480 ( .A1(n3521), .A2(keyinput5), .B1(keyinput27), .B2(n6555), 
        .ZN(n6554) );
  OAI221_X1 U7481 ( .B1(n3521), .B2(keyinput5), .C1(n6555), .C2(keyinput27), 
        .A(n6554), .ZN(n6567) );
  INV_X1 U7482 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6557) );
  AOI22_X1 U7483 ( .A1(n3476), .A2(keyinput14), .B1(n6557), .B2(keyinput1), 
        .ZN(n6556) );
  OAI221_X1 U7484 ( .B1(n3476), .B2(keyinput14), .C1(n6557), .C2(keyinput1), 
        .A(n6556), .ZN(n6566) );
  INV_X1 U7485 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6559) );
  AOI22_X1 U7486 ( .A1(n6560), .A2(keyinput47), .B1(keyinput51), .B2(n6559), 
        .ZN(n6558) );
  OAI221_X1 U7487 ( .B1(n6560), .B2(keyinput47), .C1(n6559), .C2(keyinput51), 
        .A(n6558), .ZN(n6565) );
  INV_X1 U7488 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6562) );
  AOI22_X1 U7489 ( .A1(n6563), .A2(keyinput55), .B1(n6562), .B2(keyinput61), 
        .ZN(n6561) );
  OAI221_X1 U7490 ( .B1(n6563), .B2(keyinput55), .C1(n6562), .C2(keyinput61), 
        .A(n6561), .ZN(n6564) );
  NOR4_X1 U7491 ( .A1(n6567), .A2(n6566), .A3(n6565), .A4(n6564), .ZN(n6615)
         );
  AOI22_X1 U7492 ( .A1(n4998), .A2(keyinput39), .B1(n6569), .B2(keyinput33), 
        .ZN(n6568) );
  OAI221_X1 U7493 ( .B1(n4998), .B2(keyinput39), .C1(n6569), .C2(keyinput33), 
        .A(n6568), .ZN(n6581) );
  AOI22_X1 U7494 ( .A1(n6572), .A2(keyinput7), .B1(n6571), .B2(keyinput38), 
        .ZN(n6570) );
  OAI221_X1 U7495 ( .B1(n6572), .B2(keyinput7), .C1(n6571), .C2(keyinput38), 
        .A(n6570), .ZN(n6580) );
  INV_X1 U7496 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6575) );
  AOI22_X1 U7497 ( .A1(n6575), .A2(keyinput6), .B1(keyinput50), .B2(n6574), 
        .ZN(n6573) );
  OAI221_X1 U7498 ( .B1(n6575), .B2(keyinput6), .C1(n6574), .C2(keyinput50), 
        .A(n6573), .ZN(n6579) );
  AOI22_X1 U7499 ( .A1(n6577), .A2(keyinput56), .B1(n3554), .B2(keyinput36), 
        .ZN(n6576) );
  OAI221_X1 U7500 ( .B1(n6577), .B2(keyinput56), .C1(n3554), .C2(keyinput36), 
        .A(n6576), .ZN(n6578) );
  NOR4_X1 U7501 ( .A1(n6581), .A2(n6580), .A3(n6579), .A4(n6578), .ZN(n6614)
         );
  AOI22_X1 U7502 ( .A1(n6584), .A2(keyinput17), .B1(keyinput10), .B2(n6583), 
        .ZN(n6582) );
  OAI221_X1 U7503 ( .B1(n6584), .B2(keyinput17), .C1(n6583), .C2(keyinput10), 
        .A(n6582), .ZN(n6596) );
  INV_X1 U7504 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n6587) );
  AOI22_X1 U7505 ( .A1(n6587), .A2(keyinput21), .B1(n6586), .B2(keyinput42), 
        .ZN(n6585) );
  OAI221_X1 U7506 ( .B1(n6587), .B2(keyinput21), .C1(n6586), .C2(keyinput42), 
        .A(n6585), .ZN(n6595) );
  AOI22_X1 U7507 ( .A1(n6590), .A2(keyinput31), .B1(n6589), .B2(keyinput2), 
        .ZN(n6588) );
  OAI221_X1 U7508 ( .B1(n6590), .B2(keyinput31), .C1(n6589), .C2(keyinput2), 
        .A(n6588), .ZN(n6594) );
  INV_X1 U7509 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n6592) );
  AOI22_X1 U7510 ( .A1(n6592), .A2(keyinput46), .B1(keyinput28), .B2(n4988), 
        .ZN(n6591) );
  OAI221_X1 U7511 ( .B1(n6592), .B2(keyinput46), .C1(n4988), .C2(keyinput28), 
        .A(n6591), .ZN(n6593) );
  NOR4_X1 U7512 ( .A1(n6596), .A2(n6595), .A3(n6594), .A4(n6593), .ZN(n6613)
         );
  INV_X1 U7513 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n6598) );
  AOI22_X1 U7514 ( .A1(n4576), .A2(keyinput40), .B1(keyinput11), .B2(n6598), 
        .ZN(n6597) );
  OAI221_X1 U7515 ( .B1(n4576), .B2(keyinput40), .C1(n6598), .C2(keyinput11), 
        .A(n6597), .ZN(n6611) );
  INV_X1 U7516 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6601) );
  INV_X1 U7517 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n6600) );
  AOI22_X1 U7518 ( .A1(n6601), .A2(keyinput54), .B1(n6600), .B2(keyinput24), 
        .ZN(n6599) );
  OAI221_X1 U7519 ( .B1(n6601), .B2(keyinput54), .C1(n6600), .C2(keyinput24), 
        .A(n6599), .ZN(n6610) );
  INV_X1 U7520 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n6604) );
  INV_X1 U7521 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6603) );
  AOI22_X1 U7522 ( .A1(n6604), .A2(keyinput4), .B1(n6603), .B2(keyinput20), 
        .ZN(n6602) );
  OAI221_X1 U7523 ( .B1(n6604), .B2(keyinput4), .C1(n6603), .C2(keyinput20), 
        .A(n6602), .ZN(n6609) );
  INV_X1 U7524 ( .A(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n6607) );
  INV_X1 U7525 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n6606) );
  AOI22_X1 U7526 ( .A1(n6607), .A2(keyinput57), .B1(keyinput49), .B2(n6606), 
        .ZN(n6605) );
  OAI221_X1 U7527 ( .B1(n6607), .B2(keyinput57), .C1(n6606), .C2(keyinput49), 
        .A(n6605), .ZN(n6608) );
  NOR4_X1 U7528 ( .A1(n6611), .A2(n6610), .A3(n6609), .A4(n6608), .ZN(n6612)
         );
  NAND4_X1 U7529 ( .A1(n6615), .A2(n6614), .A3(n6613), .A4(n6612), .ZN(n6682)
         );
  INV_X1 U7530 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6617) );
  AOI22_X1 U7531 ( .A1(n6618), .A2(keyinput30), .B1(n6617), .B2(keyinput8), 
        .ZN(n6616) );
  OAI221_X1 U7532 ( .B1(n6618), .B2(keyinput30), .C1(n6617), .C2(keyinput8), 
        .A(n6616), .ZN(n6630) );
  AOI22_X1 U7533 ( .A1(n6621), .A2(keyinput25), .B1(n6620), .B2(keyinput62), 
        .ZN(n6619) );
  OAI221_X1 U7534 ( .B1(n6621), .B2(keyinput25), .C1(n6620), .C2(keyinput62), 
        .A(n6619), .ZN(n6629) );
  AOI22_X1 U7535 ( .A1(n6623), .A2(keyinput3), .B1(n4496), .B2(keyinput19), 
        .ZN(n6622) );
  OAI221_X1 U7536 ( .B1(n6623), .B2(keyinput3), .C1(n4496), .C2(keyinput19), 
        .A(n6622), .ZN(n6628) );
  NOR4_X1 U7537 ( .A1(n6630), .A2(n6629), .A3(n6628), .A4(n6627), .ZN(n6680)
         );
  INV_X1 U7538 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6633) );
  INV_X1 U7539 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n6632) );
  AOI22_X1 U7540 ( .A1(n6633), .A2(keyinput16), .B1(keyinput58), .B2(n6632), 
        .ZN(n6631) );
  OAI221_X1 U7541 ( .B1(n6633), .B2(keyinput16), .C1(n6632), .C2(keyinput58), 
        .A(n6631), .ZN(n6645) );
  INV_X1 U7542 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6636) );
  INV_X1 U7543 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6635) );
  AOI22_X1 U7544 ( .A1(n6636), .A2(keyinput13), .B1(n6635), .B2(keyinput60), 
        .ZN(n6634) );
  OAI221_X1 U7545 ( .B1(n6636), .B2(keyinput13), .C1(n6635), .C2(keyinput60), 
        .A(n6634), .ZN(n6644) );
  INV_X1 U7546 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n6638) );
  AOI22_X1 U7547 ( .A1(n3528), .A2(keyinput18), .B1(keyinput45), .B2(n6638), 
        .ZN(n6637) );
  OAI221_X1 U7548 ( .B1(n3528), .B2(keyinput18), .C1(n6638), .C2(keyinput45), 
        .A(n6637), .ZN(n6643) );
  INV_X1 U7549 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6641) );
  AOI22_X1 U7550 ( .A1(n6641), .A2(keyinput43), .B1(n6640), .B2(keyinput0), 
        .ZN(n6639) );
  OAI221_X1 U7551 ( .B1(n6641), .B2(keyinput43), .C1(n6640), .C2(keyinput0), 
        .A(n6639), .ZN(n6642) );
  NOR4_X1 U7552 ( .A1(n6645), .A2(n6644), .A3(n6643), .A4(n6642), .ZN(n6679)
         );
  INV_X1 U7553 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6648) );
  AOI22_X1 U7554 ( .A1(n6648), .A2(keyinput23), .B1(keyinput9), .B2(n6647), 
        .ZN(n6646) );
  OAI221_X1 U7555 ( .B1(n6648), .B2(keyinput23), .C1(n6647), .C2(keyinput9), 
        .A(n6646), .ZN(n6660) );
  AOI22_X1 U7556 ( .A1(n6651), .A2(keyinput59), .B1(n6650), .B2(keyinput48), 
        .ZN(n6649) );
  OAI221_X1 U7557 ( .B1(n6651), .B2(keyinput59), .C1(n6650), .C2(keyinput48), 
        .A(n6649), .ZN(n6659) );
  AOI22_X1 U7558 ( .A1(n3779), .A2(keyinput35), .B1(keyinput29), .B2(n6653), 
        .ZN(n6652) );
  OAI221_X1 U7559 ( .B1(n3779), .B2(keyinput35), .C1(n6653), .C2(keyinput29), 
        .A(n6652), .ZN(n6658) );
  INV_X1 U7560 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n6655) );
  AOI22_X1 U7561 ( .A1(n6656), .A2(keyinput37), .B1(n6655), .B2(keyinput26), 
        .ZN(n6654) );
  OAI221_X1 U7562 ( .B1(n6656), .B2(keyinput37), .C1(n6655), .C2(keyinput26), 
        .A(n6654), .ZN(n6657) );
  NOR4_X1 U7563 ( .A1(n6660), .A2(n6659), .A3(n6658), .A4(n6657), .ZN(n6678)
         );
  INV_X1 U7564 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6662) );
  AOI22_X1 U7565 ( .A1(n6663), .A2(keyinput15), .B1(n6662), .B2(keyinput53), 
        .ZN(n6661) );
  OAI221_X1 U7566 ( .B1(n6663), .B2(keyinput15), .C1(n6662), .C2(keyinput53), 
        .A(n6661), .ZN(n6676) );
  INV_X1 U7567 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6666) );
  INV_X1 U7568 ( .A(DATAI_23_), .ZN(n6665) );
  AOI22_X1 U7569 ( .A1(n6666), .A2(keyinput41), .B1(keyinput22), .B2(n6665), 
        .ZN(n6664) );
  OAI221_X1 U7570 ( .B1(n6666), .B2(keyinput41), .C1(n6665), .C2(keyinput22), 
        .A(n6664), .ZN(n6675) );
  INV_X1 U7571 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6669) );
  INV_X1 U7572 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6668) );
  AOI22_X1 U7573 ( .A1(n6669), .A2(keyinput44), .B1(keyinput32), .B2(n6668), 
        .ZN(n6667) );
  OAI221_X1 U7574 ( .B1(n6669), .B2(keyinput44), .C1(n6668), .C2(keyinput32), 
        .A(n6667), .ZN(n6674) );
  INV_X1 U7575 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n6672) );
  AOI22_X1 U7576 ( .A1(n6672), .A2(keyinput52), .B1(n6671), .B2(keyinput63), 
        .ZN(n6670) );
  OAI221_X1 U7577 ( .B1(n6672), .B2(keyinput52), .C1(n6671), .C2(keyinput63), 
        .A(n6670), .ZN(n6673) );
  NOR4_X1 U7578 ( .A1(n6676), .A2(n6675), .A3(n6674), .A4(n6673), .ZN(n6677)
         );
  NAND4_X1 U7579 ( .A1(n6680), .A2(n6679), .A3(n6678), .A4(n6677), .ZN(n6681)
         );
  NOR2_X1 U7580 ( .A1(n6682), .A2(n6681), .ZN(n6685) );
  NAND2_X1 U7581 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6683), .ZN(n6684) );
  XNOR2_X1 U7582 ( .A(n6685), .B(n6684), .ZN(n6686) );
  XOR2_X1 U7583 ( .A(n6687), .B(n6686), .Z(U3176) );
  AND2_X1 U3791 ( .A1(n4067), .A2(n2973), .ZN(n3316) );
  NAND4_X2 U3426 ( .A1(n3154), .A2(n3153), .A3(n3152), .A4(n3151), .ZN(n4497)
         );
  CLKBUF_X3 U3420 ( .A(n3323), .Z(n2955) );
  AND4_X1 U3434 ( .A1(n3150), .A2(n3149), .A3(n3148), .A4(n3147), .ZN(n3151)
         );
  CLKBUF_X1 U3439 ( .A(n3042), .Z(n3120) );
  CLKBUF_X1 U3440 ( .A(n5301), .Z(n5410) );
  CLKBUF_X1 U34600 ( .A(n3033), .Z(n5799) );
  CLKBUF_X1 U3564 ( .A(n5203), .Z(n5217) );
  CLKBUF_X1 U3624 ( .A(n5626), .Z(n6005) );
  CLKBUF_X1 U3640 ( .A(n3388), .Z(n5263) );
endmodule

