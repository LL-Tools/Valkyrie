

module b21_C_gen_AntiSAT_k_256_3 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67, 
        keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72, 
        keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77, 
        keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82, 
        keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87, 
        keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92, 
        keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97, 
        keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410;

  INV_X4 U4977 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NAND2_X1 U4978 ( .A1(n8432), .A2(n8435), .ZN(n8431) );
  INV_X1 U4979 ( .A(n5162), .ZN(n6491) );
  INV_X2 U4980 ( .A(n6309), .ZN(n6887) );
  CLKBUF_X2 U4981 ( .A(n5869), .Z(n8840) );
  CLKBUF_X1 U4982 ( .A(n8827), .Z(n4473) );
  NOR2_X1 U4983 ( .A1(n6386), .A2(n9632), .ZN(n8827) );
  NOR2_X1 U4984 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5032) );
  AND4_X1 U4985 ( .A1(n5030), .A2(n5029), .A3(n5028), .A4(n5027), .ZN(n5034)
         );
  INV_X1 U4986 ( .A(n9082), .ZN(n4673) );
  INV_X2 U4988 ( .A(n5167), .ZN(n6492) );
  AND2_X1 U4989 ( .A1(n4748), .A2(n4747), .ZN(n7301) );
  NAND2_X1 U4990 ( .A1(n4788), .A2(n5431), .ZN(n5676) );
  NAND2_X1 U4991 ( .A1(n4525), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5055) );
  INV_X1 U4992 ( .A(n5921), .ZN(n5866) );
  OAI21_X1 U4993 ( .B1(n8658), .B2(n8208), .A(n8431), .ZN(n8415) );
  NOR2_X1 U4994 ( .A1(n8710), .A2(n4500), .ZN(n8760) );
  XNOR2_X1 U4995 ( .A(n5777), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5784) );
  INV_X2 U4996 ( .A(n9751), .ZN(n9753) );
  OAI21_X2 U4997 ( .B1(n4993), .B2(n4996), .A(n4997), .ZN(n4992) );
  OAI22_X2 U4998 ( .A1(n7254), .A2(n6438), .B1(n7351), .B2(n6440), .ZN(n7364)
         );
  OAI222_X1 U4999 ( .A1(n8694), .A2(n6609), .B1(n8696), .B2(n6608), .C1(
        P2_U3152), .C2(n6797), .ZN(P2_U3350) );
  OAI222_X1 U5000 ( .A1(n9522), .A2(n6607), .B1(n9513), .B2(n6608), .C1(
        P1_U3084), .C2(n6606), .ZN(P1_U3345) );
  INV_X2 U5001 ( .A(n5665), .ZN(n5639) );
  NOR2_X2 U5002 ( .A1(n7518), .A2(n7523), .ZN(n7519) );
  OAI21_X2 U5003 ( .B1(n7630), .B2(n7629), .A(n8967), .ZN(n7646) );
  NAND2_X1 U5004 ( .A1(n9087), .A2(n8890), .ZN(n9052) );
  OAI21_X2 U5005 ( .B1(n5535), .B2(n4889), .A(n5539), .ZN(n5558) );
  NOR2_X2 U5006 ( .A1(n9230), .A2(n9233), .ZN(n9229) );
  AND2_X1 U5007 ( .A1(n5893), .A2(n6582), .ZN(n4474) );
  AND2_X1 U5008 ( .A1(n5893), .A2(n6582), .ZN(n5845) );
  OAI21_X2 U5009 ( .B1(n7643), .B2(n7627), .A(n7628), .ZN(n7780) );
  NAND2_X2 U5010 ( .A1(n7626), .A2(n7625), .ZN(n7643) );
  AND2_X4 U5011 ( .A1(n5792), .A2(n5776), .ZN(n5808) );
  INV_X4 U5012 ( .A(n5145), .ZN(n5161) );
  XNOR2_X2 U5013 ( .A(n5055), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8069) );
  AOI211_X2 U5014 ( .C1(n8016), .C2(n8015), .A(n8023), .B(n4722), .ZN(n8019)
         );
  AND2_X4 U5015 ( .A1(n4854), .A2(n4853), .ZN(n6582) );
  OAI21_X1 U5016 ( .B1(n8132), .B2(n4802), .A(n4800), .ZN(n8142) );
  NAND2_X1 U5017 ( .A1(n6298), .A2(n6297), .ZN(n9432) );
  AOI22_X1 U5018 ( .A1(n8485), .A2(n8480), .B1(n8256), .B2(n8487), .ZN(n8462)
         );
  OAI21_X1 U5019 ( .B1(n9390), .B2(n9176), .A(n9177), .ZN(n9386) );
  OAI21_X1 U5020 ( .B1(n9194), .B2(n4642), .A(n4640), .ZN(n9197) );
  NAND2_X1 U5021 ( .A1(n4837), .A2(n8989), .ZN(n9194) );
  NAND2_X1 U5022 ( .A1(n7645), .A2(n8973), .ZN(n7785) );
  NAND2_X1 U5023 ( .A1(n6974), .A2(n6976), .ZN(n6975) );
  NAND2_X1 U5024 ( .A1(n8788), .A2(n8790), .ZN(n8789) );
  INV_X1 U5025 ( .A(n7421), .ZN(n7500) );
  NAND2_X1 U5026 ( .A1(n7933), .A2(n7934), .ZN(n7040) );
  NAND2_X1 U5027 ( .A1(n9140), .A2(n6920), .ZN(n8890) );
  INV_X1 U5028 ( .A(n9141), .ZN(n6898) );
  INV_X1 U5029 ( .A(n8793), .ZN(n9766) );
  INV_X1 U5030 ( .A(n7054), .ZN(n6422) );
  BUF_X2 U5031 ( .A(n5854), .Z(n6405) );
  NAND2_X2 U5032 ( .A1(n6689), .A2(n6469), .ZN(n5199) );
  NOR2_X1 U5033 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5033) );
  OAI21_X1 U5034 ( .B1(n8073), .B2(n8066), .A(n8072), .ZN(n8067) );
  NAND2_X1 U5035 ( .A1(n6267), .A2(n6266), .ZN(n8778) );
  NAND2_X1 U5036 ( .A1(n8776), .A2(n8777), .ZN(n8775) );
  OAI211_X1 U5037 ( .C1(n8355), .C2(n4979), .A(n4976), .B(n4975), .ZN(n8093)
         );
  AOI21_X1 U5038 ( .B1(n4579), .B2(n9838), .A(n6501), .ZN(n8102) );
  NOR4_X1 U5039 ( .A1(n8058), .A2(n8057), .A3(n8356), .A4(n7921), .ZN(n7922)
         );
  AOI21_X1 U5040 ( .B1(n7879), .B2(n8051), .A(n7878), .ZN(n7896) );
  NAND2_X1 U5041 ( .A1(n8719), .A2(n6212), .ZN(n8769) );
  AOI21_X1 U5042 ( .B1(n8186), .B2(n5589), .A(n5026), .ZN(n5590) );
  NAND2_X1 U5043 ( .A1(n4680), .A2(n4678), .ZN(n8719) );
  AOI21_X1 U5044 ( .B1(n8415), .B2(n4991), .A(n4989), .ZN(n4988) );
  AND2_X1 U5045 ( .A1(n7881), .A2(n7880), .ZN(n8642) );
  XNOR2_X1 U5046 ( .A(n8569), .B(n8105), .ZN(n8356) );
  NAND2_X1 U5047 ( .A1(n6117), .A2(n6100), .ZN(n8699) );
  NAND2_X1 U5048 ( .A1(n4929), .A2(n4928), .ZN(n8700) );
  OR2_X1 U5049 ( .A1(n9437), .A2(n8911), .ZN(n9261) );
  OAI21_X1 U5050 ( .B1(n8255), .B2(n8604), .A(n6455), .ZN(n8448) );
  NAND2_X1 U5051 ( .A1(n5622), .A2(n5621), .ZN(n8577) );
  NAND2_X1 U5052 ( .A1(n6322), .A2(n6321), .ZN(n9426) );
  XNOR2_X1 U5053 ( .A(n6463), .B(n6462), .ZN(n9515) );
  NAND2_X1 U5054 ( .A1(n5601), .A2(n5600), .ZN(n8410) );
  NAND2_X1 U5055 ( .A1(n6272), .A2(n6271), .ZN(n9442) );
  NAND2_X1 U5056 ( .A1(n9175), .A2(n9174), .ZN(n9390) );
  AND2_X1 U5057 ( .A1(n4786), .A2(n8018), .ZN(n4782) );
  INV_X1 U5058 ( .A(n8468), .ZN(n8604) );
  AND2_X1 U5059 ( .A1(n5524), .A2(n5523), .ZN(n8468) );
  XNOR2_X1 U5060 ( .A(n5566), .B(n5565), .ZN(n7602) );
  OAI21_X1 U5061 ( .B1(n5558), .B2(n5557), .A(n5556), .ZN(n5566) );
  NAND2_X1 U5062 ( .A1(n5522), .A2(n5521), .ZN(n5535) );
  NAND2_X1 U5063 ( .A1(n4948), .A2(n4947), .ZN(n7624) );
  NAND2_X1 U5064 ( .A1(n6173), .A2(n6172), .ZN(n9475) );
  NAND2_X1 U5065 ( .A1(n5438), .A2(n5437), .ZN(n8535) );
  AND2_X1 U5066 ( .A1(n7999), .A2(n8000), .ZN(n8542) );
  AOI21_X1 U5067 ( .B1(n4954), .B2(n4952), .A(n4519), .ZN(n4951) );
  NAND2_X1 U5068 ( .A1(n5366), .A2(n5365), .ZN(n8120) );
  NAND2_X1 U5069 ( .A1(n5396), .A2(n5395), .ZN(n8550) );
  NOR2_X1 U5070 ( .A1(n5233), .A2(n4812), .ZN(n4811) );
  NAND2_X1 U5071 ( .A1(n6087), .A2(n6086), .ZN(n8875) );
  NAND2_X1 U5072 ( .A1(n6046), .A2(n6045), .ZN(n7745) );
  NAND2_X1 U5073 ( .A1(n6002), .A2(n6001), .ZN(n9587) );
  AND2_X1 U5074 ( .A1(n5273), .A2(n5272), .ZN(n7617) );
  OAI211_X1 U5075 ( .C1(n6689), .C2(n6797), .A(n5229), .B(n5228), .ZN(n7421)
         );
  INV_X1 U5076 ( .A(n6430), .ZN(n9929) );
  NAND4_X1 U5077 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n5146), .ZN(n8270)
         );
  AND4_X1 U5078 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n7046)
         );
  AND4_X1 U5079 ( .A1(n5108), .A2(n5107), .A3(n5106), .A4(n5105), .ZN(n9813)
         );
  NAND2_X1 U5080 ( .A1(n4750), .A2(n4498), .ZN(n7054) );
  OAI211_X1 U5081 ( .C1(n6689), .C2(n6721), .A(n5116), .B(n5115), .ZN(n9917)
         );
  NAND4_X1 U5082 ( .A1(n5829), .A2(n5828), .A3(n5827), .A4(n5826), .ZN(n9141)
         );
  NAND2_X1 U5083 ( .A1(n4712), .A2(n5132), .ZN(n5155) );
  NAND2_X1 U5084 ( .A1(n5049), .A2(n8689), .ZN(n5162) );
  OAI211_X1 U5085 ( .C1(n6689), .C2(n6593), .A(n5097), .B(n5096), .ZN(n7057)
         );
  NAND2_X1 U5086 ( .A1(n4673), .A2(n4672), .ZN(n6879) );
  INV_X2 U5087 ( .A(n5249), .ZN(n7890) );
  INV_X1 U5088 ( .A(n5852), .ZN(n6194) );
  AND2_X2 U5089 ( .A1(n5784), .A2(n8092), .ZN(n5921) );
  NAND2_X1 U5090 ( .A1(n6363), .A2(n9626), .ZN(n5893) );
  INV_X1 U5091 ( .A(n8530), .ZN(n7923) );
  XNOR2_X1 U5092 ( .A(n5042), .B(n5041), .ZN(n8689) );
  OR2_X1 U5093 ( .A1(n8679), .A2(n8680), .ZN(n5045) );
  MUX2_X1 U5094 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5779), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5780) );
  MUX2_X1 U5095 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5748), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5749) );
  OR2_X1 U5096 ( .A1(n4986), .A2(n8680), .ZN(n4749) );
  NAND2_X1 U5097 ( .A1(n4902), .A2(n5750), .ZN(n9626) );
  OR2_X1 U5098 ( .A1(n5061), .A2(n8680), .ZN(n5063) );
  NAND2_X1 U5099 ( .A1(n5778), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5777) );
  NOR2_X1 U5100 ( .A1(n5676), .A2(n4697), .ZN(n4986) );
  AND2_X1 U5101 ( .A1(n5017), .A2(n4789), .ZN(n4788) );
  INV_X2 U5102 ( .A(n6582), .ZN(n6469) );
  AND2_X1 U5103 ( .A1(n5018), .A2(n5038), .ZN(n5017) );
  NOR2_X1 U5104 ( .A1(n4790), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4789) );
  OAI21_X1 U5105 ( .B1(n4857), .B2(n4856), .A(n4855), .ZN(n5066) );
  AND3_X1 U5106 ( .A1(n5033), .A2(n5032), .A3(n5001), .ZN(n5000) );
  AND2_X1 U5107 ( .A1(n5037), .A2(n5036), .ZN(n5018) );
  INV_X1 U5108 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10072) );
  INV_X1 U5109 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4856) );
  NOR2_X1 U5110 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5830) );
  NOR2_X1 U5111 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P1_RD_REG_SCAN_IN), .ZN(
        n4710) );
  NOR2_X1 U5112 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5029) );
  NOR2_X1 U5113 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5028) );
  NOR2_X1 U5114 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5027) );
  NOR2_X1 U5115 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5088) );
  NOR3_X1 U5116 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5039) );
  NOR2_X1 U5117 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5031) );
  NOR2_X1 U5118 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5037) );
  NOR2_X1 U5119 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5737) );
  NOR2_X1 U5120 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5736) );
  NOR2_X1 U5121 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5738) );
  AND2_X1 U5122 ( .A1(n4854), .A2(n4853), .ZN(n4475) );
  NOR2_X2 U5123 ( .A1(n8523), .A2(n8514), .ZN(n4699) );
  NAND2_X1 U5124 ( .A1(n6689), .A2(n6469), .ZN(n4476) );
  INV_X1 U5125 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5244) );
  NAND2_X2 U5126 ( .A1(n6689), .A2(n6582), .ZN(n5249) );
  INV_X1 U5127 ( .A(n8001), .ZN(n4734) );
  OAI21_X1 U5128 ( .B1(n4731), .B2(n4478), .A(n4728), .ZN(n4727) );
  AND2_X1 U5129 ( .A1(n4735), .A2(n8059), .ZN(n4731) );
  NAND2_X1 U5130 ( .A1(n4600), .A2(n4597), .ZN(n9003) );
  NAND2_X1 U5131 ( .A1(n4601), .A2(n9032), .ZN(n4600) );
  NAND2_X1 U5132 ( .A1(n4598), .A2(n9030), .ZN(n4597) );
  NAND2_X1 U5133 ( .A1(n4604), .A2(n4602), .ZN(n4601) );
  INV_X1 U5134 ( .A(n7913), .ZN(n5011) );
  INV_X1 U5135 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5001) );
  AND2_X1 U5136 ( .A1(n6361), .A2(n6879), .ZN(n6309) );
  NAND2_X1 U5137 ( .A1(n9039), .A2(n8848), .ZN(n9081) );
  INV_X1 U5138 ( .A(n5536), .ZN(n4889) );
  NAND2_X1 U5139 ( .A1(n5356), .A2(n5355), .ZN(n5358) );
  BUF_X1 U5140 ( .A(n5162), .Z(n6663) );
  NAND2_X1 U5141 ( .A1(n4710), .A2(n4856), .ZN(n4854) );
  NAND2_X1 U5142 ( .A1(n5745), .A2(n4632), .ZN(n4631) );
  NAND2_X1 U5143 ( .A1(n7994), .A2(n7993), .ZN(n4736) );
  INV_X1 U5144 ( .A(n7995), .ZN(n4735) );
  NAND2_X1 U5145 ( .A1(n9003), .A2(n4596), .ZN(n8999) );
  AND2_X1 U5146 ( .A1(n9048), .A2(n8998), .ZN(n4596) );
  AND2_X1 U5147 ( .A1(n7274), .A2(n7951), .ZN(n7950) );
  NAND2_X1 U5148 ( .A1(n9127), .A2(n9745), .ZN(n6361) );
  INV_X1 U5149 ( .A(SI_9_), .ZN(n5245) );
  NAND2_X1 U5150 ( .A1(n4578), .A2(n4577), .ZN(n6489) );
  AND2_X1 U5151 ( .A1(n8388), .A2(n8040), .ZN(n4578) );
  NOR2_X1 U5152 ( .A1(n8496), .A2(n4785), .ZN(n4784) );
  INV_X1 U5153 ( .A(n7977), .ZN(n5012) );
  NAND2_X1 U5154 ( .A1(n7301), .A2(n8270), .ZN(n7951) );
  NAND2_X1 U5155 ( .A1(n7737), .A2(n4930), .ZN(n4929) );
  NOR2_X1 U5156 ( .A1(n7723), .A2(n4931), .ZN(n4930) );
  INV_X1 U5157 ( .A(n6064), .ZN(n4931) );
  AND2_X1 U5158 ( .A1(n7559), .A2(n4908), .ZN(n4907) );
  NAND2_X1 U5159 ( .A1(n4494), .A2(n6014), .ZN(n4908) );
  NAND2_X1 U5160 ( .A1(n9044), .A2(n9030), .ZN(n4615) );
  NAND2_X1 U5161 ( .A1(n4617), .A2(n9113), .ZN(n4616) );
  NOR2_X1 U5162 ( .A1(n9276), .A2(n4961), .ZN(n4960) );
  INV_X1 U5163 ( .A(n4963), .ZN(n4961) );
  NAND2_X1 U5164 ( .A1(n9186), .A2(n9187), .ZN(n4966) );
  OR2_X1 U5165 ( .A1(n7243), .A2(n7219), .ZN(n7187) );
  NAND2_X1 U5166 ( .A1(n4634), .A2(n9739), .ZN(n9089) );
  INV_X1 U5167 ( .A(n9138), .ZN(n4634) );
  AND2_X1 U5168 ( .A1(n5025), .A2(n5745), .ZN(n4845) );
  NAND2_X1 U5169 ( .A1(n5568), .A2(n5567), .ZN(n5596) );
  OAI21_X1 U5170 ( .B1(n5498), .B2(n5497), .A(n5499), .ZN(n5520) );
  OAI21_X1 U5171 ( .B1(n5457), .B2(n5456), .A(n5455), .ZN(n5476) );
  AND2_X1 U5172 ( .A1(n5428), .A2(n5392), .ZN(n5426) );
  OAI21_X1 U5173 ( .B1(n5286), .B2(n4885), .A(n4883), .ZN(n5356) );
  INV_X1 U5174 ( .A(n4884), .ZN(n4883) );
  OAI21_X1 U5175 ( .B1(n4887), .B2(n4885), .A(n5335), .ZN(n4884) );
  NAND2_X1 U5176 ( .A1(n4886), .A2(n5307), .ZN(n4885) );
  AND2_X1 U5177 ( .A1(n5357), .A2(n5338), .ZN(n5355) );
  NAND2_X1 U5178 ( .A1(n5265), .A2(n5264), .ZN(n5285) );
  INV_X1 U5179 ( .A(SI_10_), .ZN(n5264) );
  NAND2_X1 U5180 ( .A1(n5284), .A2(n5023), .ZN(n5286) );
  AOI21_X1 U5181 ( .B1(n4824), .B2(n7166), .A(n4823), .ZN(n4822) );
  INV_X1 U5182 ( .A(n5181), .ZN(n4823) );
  INV_X1 U5183 ( .A(n4811), .ZN(n4809) );
  AOI21_X1 U5184 ( .B1(n4811), .B2(n4808), .A(n4807), .ZN(n4806) );
  INV_X1 U5185 ( .A(n5259), .ZN(n4807) );
  INV_X1 U5186 ( .A(n7494), .ZN(n4808) );
  AND2_X1 U5187 ( .A1(n4825), .A2(n4826), .ZN(n4824) );
  INV_X1 U5188 ( .A(n7319), .ZN(n4825) );
  INV_X1 U5189 ( .A(n5161), .ZN(n6495) );
  AND4_X1 U5190 ( .A1(n5190), .A2(n5189), .A3(n5188), .A4(n5187), .ZN(n7345)
         );
  NAND2_X1 U5191 ( .A1(n5049), .A2(n5048), .ZN(n5163) );
  NOR2_X1 U5192 ( .A1(n8358), .A2(n4580), .ZN(n7879) );
  NOR2_X1 U5193 ( .A1(n8569), .A2(n8105), .ZN(n4580) );
  INV_X1 U5194 ( .A(n4992), .ZN(n4991) );
  OR2_X1 U5195 ( .A1(n8410), .A2(n8253), .ZN(n4997) );
  XNOR2_X1 U5196 ( .A(n8410), .B(n8253), .ZN(n8405) );
  OR2_X1 U5197 ( .A1(n8600), .A2(n8147), .ZN(n8434) );
  AOI22_X1 U5198 ( .A1(n8512), .A2(n6450), .B1(n8669), .B2(n6482), .ZN(n8493)
         );
  OR2_X1 U5199 ( .A1(n7771), .A2(n8263), .ZN(n5009) );
  INV_X1 U5200 ( .A(n7540), .ZN(n5004) );
  NAND2_X1 U5201 ( .A1(n5691), .A2(n9889), .ZN(n7008) );
  NAND2_X1 U5202 ( .A1(n7530), .A2(n7937), .ZN(n9897) );
  NAND2_X1 U5203 ( .A1(n5040), .A2(n4698), .ZN(n4697) );
  NAND2_X1 U5204 ( .A1(n6168), .A2(n4676), .ZN(n4680) );
  NOR2_X1 U5205 ( .A1(n4520), .A2(n4677), .ZN(n4676) );
  INV_X1 U5206 ( .A(n6167), .ZN(n4677) );
  AND2_X1 U5207 ( .A1(n4921), .A2(n4926), .ZN(n4920) );
  NAND2_X1 U5208 ( .A1(n4497), .A2(n4924), .ZN(n4921) );
  AND2_X1 U5209 ( .A1(n5843), .A2(n5844), .ZN(n8790) );
  INV_X1 U5210 ( .A(n5845), .ZN(n6190) );
  INV_X1 U5211 ( .A(n5846), .ZN(n6521) );
  OAI22_X1 U5212 ( .A1(n9241), .A2(n9248), .B1(n9265), .B2(n9426), .ZN(n9230)
         );
  INV_X1 U5213 ( .A(n4957), .ZN(n4952) );
  INV_X2 U5214 ( .A(n5834), .ZN(n8850) );
  NAND2_X1 U5215 ( .A1(n5019), .A2(n4509), .ZN(n7239) );
  INV_X1 U5216 ( .A(n6874), .ZN(n9054) );
  NAND2_X1 U5217 ( .A1(n6937), .A2(n6938), .ZN(n6936) );
  AND2_X1 U5218 ( .A1(n5025), .A2(n4974), .ZN(n4973) );
  NOR2_X1 U5219 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4974) );
  AND2_X1 U5220 ( .A1(n4935), .A2(n5753), .ZN(n4934) );
  AND2_X1 U5221 ( .A1(n10072), .A2(n5746), .ZN(n4935) );
  INV_X1 U5222 ( .A(n4751), .ZN(n4750) );
  NAND2_X1 U5223 ( .A1(n8811), .A2(n9140), .ZN(n4622) );
  INV_X1 U5224 ( .A(n4628), .ZN(n4627) );
  OAI21_X1 U5225 ( .B1(n9123), .B2(n9122), .A(n4629), .ZN(n4628) );
  INV_X1 U5226 ( .A(n9129), .ZN(n4629) );
  NAND2_X1 U5227 ( .A1(n9157), .A2(n9156), .ZN(n4567) );
  NAND2_X1 U5228 ( .A1(n4566), .A2(n4565), .ZN(n4564) );
  NAND2_X1 U5229 ( .A1(n9152), .A2(n9718), .ZN(n4566) );
  AOI21_X1 U5230 ( .B1(n9153), .B2(n9731), .A(n9156), .ZN(n4565) );
  XNOR2_X1 U5231 ( .A(n4588), .B(n8919), .ZN(n9409) );
  NAND2_X1 U5232 ( .A1(n4753), .A2(n4722), .ZN(n4721) );
  AOI21_X1 U5233 ( .B1(n7970), .B2(n7969), .A(n4765), .ZN(n4557) );
  OAI21_X1 U5234 ( .B1(n7986), .B2(n4478), .A(n4726), .ZN(n4730) );
  OAI21_X1 U5235 ( .B1(n7985), .B2(n7984), .A(n7983), .ZN(n7986) );
  INV_X1 U5236 ( .A(n4727), .ZN(n4726) );
  AND2_X1 U5237 ( .A1(n4735), .A2(n7987), .ZN(n4729) );
  NAND2_X1 U5238 ( .A1(n8996), .A2(n4605), .ZN(n4604) );
  AND2_X1 U5239 ( .A1(n9049), .A2(n9050), .ZN(n4605) );
  INV_X1 U5240 ( .A(n4611), .ZN(n4610) );
  AOI21_X1 U5241 ( .B1(n9000), .B2(n9047), .A(n4612), .ZN(n4611) );
  NAND2_X1 U5242 ( .A1(n9202), .A2(n9032), .ZN(n4612) );
  NAND2_X1 U5243 ( .A1(n8031), .A2(n8017), .ZN(n4718) );
  NAND2_X1 U5244 ( .A1(n8035), .A2(n8034), .ZN(n4716) );
  NAND2_X1 U5245 ( .A1(n8577), .A2(n8045), .ZN(n4746) );
  NAND2_X1 U5246 ( .A1(n7877), .A2(n7876), .ZN(n7883) );
  NAND2_X1 U5247 ( .A1(n7873), .A2(n7872), .ZN(n7877) );
  INV_X1 U5248 ( .A(n5426), .ZN(n4872) );
  NAND2_X1 U5249 ( .A1(n5390), .A2(n10323), .ZN(n5428) );
  NOR2_X1 U5250 ( .A1(n5403), .A2(n4878), .ZN(n4877) );
  INV_X1 U5251 ( .A(n5382), .ZN(n4878) );
  INV_X1 U5252 ( .A(SI_11_), .ZN(n10125) );
  INV_X1 U5253 ( .A(SI_14_), .ZN(n10113) );
  AND2_X1 U5254 ( .A1(n4819), .A2(n5419), .ZN(n4818) );
  NAND2_X1 U5255 ( .A1(n8114), .A2(n5379), .ZN(n4819) );
  NAND2_X1 U5256 ( .A1(n4818), .A2(n4816), .ZN(n4815) );
  INV_X1 U5257 ( .A(n5379), .ZN(n4816) );
  INV_X1 U5258 ( .A(n7614), .ZN(n4805) );
  NOR2_X1 U5259 ( .A1(n8439), .A2(n8442), .ZN(n8422) );
  OR2_X1 U5260 ( .A1(n8463), .A2(n8600), .ZN(n8439) );
  INV_X1 U5261 ( .A(n7991), .ZN(n4771) );
  INV_X1 U5262 ( .A(n6448), .ZN(n5006) );
  NOR2_X1 U5263 ( .A1(n8120), .A2(n7720), .ZN(n4704) );
  AND2_X1 U5264 ( .A1(n7976), .A2(n4764), .ZN(n4763) );
  NAND2_X1 U5265 ( .A1(n7967), .A2(n4765), .ZN(n4764) );
  NAND2_X1 U5266 ( .A1(n7923), .A2(n8079), .ZN(n8065) );
  OR2_X1 U5267 ( .A1(n7272), .A2(n7926), .ZN(n7225) );
  OR2_X1 U5268 ( .A1(n6477), .A2(n7950), .ZN(n7224) );
  NOR2_X1 U5269 ( .A1(n7088), .A2(n9917), .ZN(n9842) );
  INV_X1 U5270 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5062) );
  INV_X1 U5271 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U5272 ( .A1(n8775), .A2(n8778), .ZN(n6270) );
  NAND2_X1 U5273 ( .A1(n4684), .A2(n4480), .ZN(n7737) );
  INV_X1 U5274 ( .A(n7739), .ZN(n4683) );
  AOI21_X1 U5275 ( .B1(n4912), .B2(n4915), .A(n4518), .ZN(n4910) );
  INV_X1 U5276 ( .A(n8767), .ZN(n4915) );
  NAND2_X1 U5277 ( .A1(n8700), .A2(n8701), .ZN(n6123) );
  OR2_X1 U5278 ( .A1(n8919), .A2(n8916), .ZN(n9039) );
  OR2_X1 U5279 ( .A1(n9422), .A2(n8855), .ZN(n9209) );
  NOR2_X1 U5280 ( .A1(n9432), .A2(n9277), .ZN(n9189) );
  OR2_X1 U5281 ( .A1(n9458), .A2(n8861), .ZN(n9048) );
  INV_X1 U5282 ( .A(n9363), .ZN(n4641) );
  NOR2_X1 U5283 ( .A1(n4894), .A2(n9486), .ZN(n4591) );
  NAND2_X1 U5284 ( .A1(n4895), .A2(n9602), .ZN(n4894) );
  INV_X1 U5285 ( .A(n4896), .ZN(n4895) );
  OR2_X1 U5286 ( .A1(n9606), .A2(n8875), .ZN(n4896) );
  NOR2_X1 U5287 ( .A1(n9587), .A2(n7453), .ZN(n4590) );
  OR2_X1 U5288 ( .A1(n7436), .A2(n7217), .ZN(n8957) );
  INV_X1 U5289 ( .A(n8885), .ZN(n4606) );
  NAND2_X1 U5290 ( .A1(n8888), .A2(n9054), .ZN(n6904) );
  AND2_X1 U5291 ( .A1(n4845), .A2(n4844), .ZN(n4843) );
  INV_X1 U5292 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4844) );
  OR2_X1 U5293 ( .A1(n9346), .A2(n9199), .ZN(n9324) );
  XNOR2_X1 U5294 ( .A(n7883), .B(n7884), .ZN(n7882) );
  INV_X1 U5295 ( .A(n5615), .ZN(n4867) );
  INV_X1 U5296 ( .A(n5633), .ZN(n4866) );
  AND2_X1 U5297 ( .A1(n5631), .A2(n4863), .ZN(n4862) );
  NOR2_X1 U5298 ( .A1(n5616), .A2(n4864), .ZN(n4863) );
  INV_X1 U5299 ( .A(n5594), .ZN(n4864) );
  NOR2_X1 U5300 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5753) );
  AND2_X1 U5301 ( .A1(n5521), .A2(n5502), .ZN(n5519) );
  INV_X1 U5302 ( .A(n5474), .ZN(n5475) );
  AOI21_X1 U5303 ( .B1(n4875), .B2(n4877), .A(n4874), .ZN(n4873) );
  INV_X1 U5304 ( .A(n5389), .ZN(n4874) );
  INV_X1 U5305 ( .A(n4880), .ZN(n4875) );
  INV_X1 U5306 ( .A(n4877), .ZN(n4876) );
  NOR2_X1 U5307 ( .A1(n5308), .A2(n4888), .ZN(n4887) );
  INV_X1 U5308 ( .A(n5285), .ZN(n4888) );
  INV_X1 U5309 ( .A(n5305), .ZN(n5308) );
  XNOR2_X1 U5310 ( .A(n5306), .B(n10125), .ZN(n5305) );
  NAND2_X1 U5311 ( .A1(n5262), .A2(n5261), .ZN(n5284) );
  AND2_X1 U5312 ( .A1(n5285), .A2(n5267), .ZN(n5023) );
  NOR2_X1 U5313 ( .A1(n4851), .A2(n4848), .ZN(n4847) );
  INV_X1 U5314 ( .A(n5174), .ZN(n4848) );
  INV_X1 U5315 ( .A(n5196), .ZN(n4851) );
  INV_X1 U5316 ( .A(n5177), .ZN(n4850) );
  INV_X1 U5317 ( .A(SI_5_), .ZN(n10161) );
  OR2_X1 U5318 ( .A1(n5848), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U5319 ( .A1(n5081), .A2(n5795), .ZN(n5092) );
  INV_X1 U5320 ( .A(n8271), .ZN(n7168) );
  INV_X1 U5321 ( .A(n5233), .ZN(n4810) );
  INV_X1 U5322 ( .A(n7549), .ZN(n4812) );
  NAND2_X1 U5323 ( .A1(n5493), .A2(n5492), .ZN(n8132) );
  NAND2_X1 U5324 ( .A1(n5291), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5322) );
  OR2_X1 U5325 ( .A1(n5439), .A2(n8181), .ZN(n5462) );
  INV_X1 U5326 ( .A(n5369), .ZN(n5368) );
  AND2_X1 U5327 ( .A1(n5017), .A2(n5035), .ZN(n4787) );
  OR2_X1 U5328 ( .A1(n9942), .A2(n7923), .ZN(n7901) );
  AOI21_X1 U5329 ( .B1(n8378), .B2(n5718), .A(n5642), .ZN(n8227) );
  AND3_X1 U5330 ( .A1(n5584), .A2(n5583), .A3(n5582), .ZN(n8208) );
  AND4_X1 U5331 ( .A1(n5512), .A2(n5511), .A3(n5510), .A4(n5509), .ZN(n8146)
         );
  AND4_X1 U5332 ( .A1(n5215), .A2(n5214), .A3(n5213), .A4(n5212), .ZN(n7367)
         );
  AND4_X1 U5333 ( .A1(n5171), .A2(n5170), .A3(n5169), .A4(n5168), .ZN(n7261)
         );
  NAND2_X1 U5334 ( .A1(n8689), .A2(n5046), .ZN(n5145) );
  NOR2_X1 U5335 ( .A1(n9557), .A2(n9556), .ZN(n9555) );
  NOR2_X1 U5336 ( .A1(n6789), .A2(n4666), .ZN(n6792) );
  NOR2_X1 U5337 ( .A1(n6797), .A2(n4667), .ZN(n4666) );
  OR2_X1 U5338 ( .A1(n6792), .A2(n6791), .ZN(n4665) );
  NAND2_X1 U5339 ( .A1(n7202), .A2(n7203), .ZN(n7334) );
  INV_X1 U5340 ( .A(n4655), .ZN(n4653) );
  NOR2_X1 U5341 ( .A1(n4650), .A2(n8283), .ZN(n4654) );
  AND2_X1 U5342 ( .A1(n4657), .A2(n8283), .ZN(n4655) );
  NOR2_X1 U5343 ( .A1(n4657), .A2(n8283), .ZN(n4656) );
  NOR2_X1 U5344 ( .A1(n8320), .A2(n4671), .ZN(n8322) );
  AND2_X1 U5345 ( .A1(n8321), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U5346 ( .A1(n8322), .A2(n8323), .ZN(n8329) );
  NAND2_X1 U5347 ( .A1(n6490), .A2(n4982), .ZN(n4977) );
  NOR2_X1 U5348 ( .A1(n8356), .A2(n6461), .ZN(n4978) );
  NAND2_X1 U5349 ( .A1(n4773), .A2(n4496), .ZN(n8358) );
  NAND2_X1 U5350 ( .A1(n8401), .A2(n8405), .ZN(n4577) );
  NAND2_X1 U5351 ( .A1(n4995), .A2(n4994), .ZN(n4993) );
  NAND2_X1 U5352 ( .A1(n4996), .A2(n8417), .ZN(n4994) );
  INV_X1 U5353 ( .A(n8405), .ZN(n4995) );
  NAND2_X1 U5354 ( .A1(n8042), .A2(n6488), .ZN(n8393) );
  NOR2_X1 U5355 ( .A1(n8590), .A2(n4999), .ZN(n4998) );
  AND2_X1 U5356 ( .A1(n8036), .A2(n8035), .ZN(n8417) );
  NOR2_X1 U5357 ( .A1(n8415), .A2(n8417), .ZN(n8414) );
  AND2_X1 U5358 ( .A1(n6484), .A2(n4780), .ZN(n4779) );
  NAND2_X1 U5359 ( .A1(n4782), .A2(n4781), .ZN(n4780) );
  INV_X1 U5360 ( .A(n4784), .ZN(n4781) );
  NAND2_X1 U5361 ( .A1(n6483), .A2(n4784), .ZN(n4783) );
  NAND2_X1 U5362 ( .A1(n8507), .A2(n8012), .ZN(n6483) );
  OR2_X1 U5363 ( .A1(n5486), .A2(n10304), .ZN(n5507) );
  NAND2_X1 U5364 ( .A1(n4569), .A2(n8000), .ZN(n8525) );
  NAND2_X1 U5365 ( .A1(n8550), .A2(n8260), .ZN(n5015) );
  OR2_X1 U5366 ( .A1(n8539), .A2(n8542), .ZN(n5016) );
  OR2_X1 U5367 ( .A1(n5411), .A2(n5410), .ZN(n5413) );
  NAND2_X1 U5368 ( .A1(n7749), .A2(n7991), .ZN(n7821) );
  NAND2_X1 U5369 ( .A1(n5010), .A2(n5007), .ZN(n7713) );
  OR2_X1 U5370 ( .A1(n7366), .A2(n6478), .ZN(n7469) );
  OR2_X1 U5371 ( .A1(n7465), .A2(n7470), .ZN(n7467) );
  INV_X1 U5372 ( .A(n9838), .ZN(n8527) );
  AND2_X1 U5373 ( .A1(n7959), .A2(n7960), .ZN(n7957) );
  AOI21_X1 U5374 ( .B1(n7268), .B2(n6435), .A(n5021), .ZN(n7223) );
  NOR2_X1 U5375 ( .A1(n6434), .A2(n6433), .ZN(n5021) );
  NAND2_X1 U5376 ( .A1(n8065), .A2(n7900), .ZN(n9838) );
  NAND2_X1 U5377 ( .A1(n5460), .A2(n5459), .ZN(n8514) );
  NAND2_X1 U5378 ( .A1(n5320), .A2(n5319), .ZN(n7771) );
  NOR2_X1 U5379 ( .A1(n5688), .A2(n7864), .ZN(n9857) );
  AND2_X1 U5380 ( .A1(n7814), .A2(n5684), .ZN(n5688) );
  NAND2_X1 U5381 ( .A1(n5697), .A2(n5696), .ZN(n5699) );
  NAND2_X1 U5382 ( .A1(n6189), .A2(n8799), .ZN(n4679) );
  NAND2_X1 U5383 ( .A1(n5907), .A2(n5906), .ZN(n5908) );
  NAND2_X1 U5384 ( .A1(n5807), .A2(n5806), .ZN(n6808) );
  AND2_X1 U5385 ( .A1(n5812), .A2(n5811), .ZN(n6809) );
  AND2_X1 U5386 ( .A1(n4918), .A2(n8751), .ZN(n4917) );
  NAND2_X1 U5387 ( .A1(n8744), .A2(n6147), .ZN(n4918) );
  AOI21_X1 U5388 ( .B1(n4616), .B2(n9032), .A(n4614), .ZN(n4613) );
  NAND2_X1 U5389 ( .A1(n9116), .A2(n9118), .ZN(n9117) );
  INV_X1 U5390 ( .A(n8840), .ZN(n6323) );
  NAND4_X1 U5391 ( .A1(n5818), .A2(n5817), .A3(n5816), .A4(n5815), .ZN(n6872)
         );
  NAND2_X1 U5392 ( .A1(n5921), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5815) );
  OR2_X1 U5393 ( .A1(n9638), .A2(n4505), .ZN(n4563) );
  NAND2_X1 U5394 ( .A1(n9265), .A2(n9329), .ZN(n4840) );
  NAND2_X1 U5395 ( .A1(n9437), .A2(n8911), .ZN(n9205) );
  NAND2_X1 U5396 ( .A1(n4532), .A2(n4966), .ZN(n4963) );
  NAND2_X1 U5397 ( .A1(n9442), .A2(n9303), .ZN(n4967) );
  AND2_X1 U5398 ( .A1(n9261), .A2(n9205), .ZN(n9276) );
  NAND2_X1 U5399 ( .A1(n4966), .A2(n4965), .ZN(n4964) );
  INV_X1 U5400 ( .A(n9184), .ZN(n4965) );
  NAND2_X1 U5401 ( .A1(n9313), .A2(n4512), .ZN(n4646) );
  NAND2_X1 U5402 ( .A1(n4646), .A2(n4645), .ZN(n9283) );
  AND2_X1 U5403 ( .A1(n9285), .A2(n9203), .ZN(n4645) );
  AND2_X1 U5404 ( .A1(n9046), .A2(n9204), .ZN(n9285) );
  NAND2_X1 U5405 ( .A1(n4937), .A2(n4513), .ZN(n9294) );
  AND2_X1 U5406 ( .A1(n4940), .A2(n4533), .ZN(n4938) );
  NAND2_X1 U5407 ( .A1(n9314), .A2(n9315), .ZN(n9313) );
  NAND2_X1 U5408 ( .A1(n4531), .A2(n4941), .ZN(n4940) );
  INV_X1 U5409 ( .A(n4492), .ZN(n4941) );
  NAND2_X1 U5410 ( .A1(n9338), .A2(n4942), .ZN(n4939) );
  NOR2_X1 U5411 ( .A1(n4944), .A2(n4943), .ZN(n4942) );
  INV_X1 U5412 ( .A(n9181), .ZN(n4944) );
  INV_X1 U5413 ( .A(n4531), .ZN(n4943) );
  AND2_X1 U5414 ( .A1(n9047), .A2(n9202), .ZN(n9315) );
  OR2_X1 U5415 ( .A1(n9339), .A2(n9458), .ZN(n9321) );
  OR2_X1 U5416 ( .A1(n9391), .A2(n9475), .ZN(n9378) );
  AND2_X1 U5417 ( .A1(n8930), .A2(n9372), .ZN(n9398) );
  AOI21_X1 U5418 ( .B1(n4834), .B2(n7784), .A(n4833), .ZN(n4832) );
  AND2_X1 U5419 ( .A1(n7568), .A2(n7572), .ZN(n7653) );
  NAND2_X1 U5420 ( .A1(n7454), .A2(n4957), .ZN(n4956) );
  OR2_X1 U5421 ( .A1(n7453), .A2(n9577), .ZN(n4957) );
  NAND2_X1 U5422 ( .A1(n7395), .A2(n8957), .ZN(n9569) );
  NOR2_X1 U5423 ( .A1(n7187), .A2(n7436), .ZN(n7400) );
  NAND2_X1 U5424 ( .A1(n4648), .A2(n8954), .ZN(n7395) );
  INV_X1 U5425 ( .A(n7183), .ZN(n4648) );
  NAND2_X1 U5426 ( .A1(n7029), .A2(n9061), .ZN(n7178) );
  NAND2_X1 U5427 ( .A1(n4969), .A2(n7025), .ZN(n5019) );
  INV_X1 U5428 ( .A(n7024), .ZN(n4970) );
  CLKBUF_X1 U5429 ( .A(n6363), .Z(n9632) );
  NAND2_X1 U5430 ( .A1(n6940), .A2(n9053), .ZN(n6939) );
  CLKBUF_X1 U5431 ( .A(n9578), .Z(n9329) );
  NAND2_X1 U5432 ( .A1(n9040), .A2(n6892), .ZN(n9574) );
  CLKBUF_X1 U5433 ( .A(n9400), .Z(n9348) );
  INV_X1 U5434 ( .A(n9791), .ZN(n9487) );
  OR2_X1 U5435 ( .A1(n6882), .A2(n9122), .ZN(n9793) );
  NAND2_X1 U5436 ( .A1(n5650), .A2(n5649), .ZN(n6463) );
  NAND2_X1 U5437 ( .A1(n5648), .A2(n5647), .ZN(n5650) );
  AND2_X1 U5438 ( .A1(n5567), .A2(n5562), .ZN(n5565) );
  XNOR2_X1 U5439 ( .A(n5772), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9127) );
  NAND2_X1 U5440 ( .A1(n4879), .A2(n5382), .ZN(n5404) );
  NAND2_X1 U5441 ( .A1(n5358), .A2(n4880), .ZN(n4879) );
  OR2_X1 U5442 ( .A1(n5999), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6015) );
  OR2_X1 U5443 ( .A1(n6039), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U5444 ( .A1(n5222), .A2(n5221), .ZN(n5242) );
  NAND2_X1 U5445 ( .A1(n5915), .A2(n5914), .ZN(n6039) );
  INV_X1 U5446 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5914) );
  NOR2_X1 U5447 ( .A1(n5894), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U5448 ( .A1(n5695), .A2(n5694), .ZN(n6681) );
  NAND2_X1 U5449 ( .A1(n5207), .A2(n5206), .ZN(n7493) );
  NAND2_X1 U5450 ( .A1(n4821), .A2(n4508), .ZN(n5207) );
  XNOR2_X1 U5451 ( .A(n5553), .B(n5551), .ZN(n8205) );
  NAND2_X1 U5452 ( .A1(n4828), .A2(n4827), .ZN(n4826) );
  INV_X1 U5453 ( .A(n5159), .ZN(n4827) );
  INV_X1 U5454 ( .A(n5160), .ZN(n4828) );
  OR2_X1 U5455 ( .A1(n7167), .A2(n7166), .ZN(n4829) );
  NAND2_X1 U5456 ( .A1(n5722), .A2(n5709), .ZN(n8247) );
  AOI21_X1 U5457 ( .B1(n4759), .B2(n4756), .A(n7902), .ZN(n7899) );
  NAND2_X1 U5458 ( .A1(n7897), .A2(n8056), .ZN(n4759) );
  AOI21_X1 U5459 ( .B1(n4758), .B2(n4757), .A(n8058), .ZN(n4756) );
  NAND2_X1 U5460 ( .A1(n5610), .A2(n5609), .ZN(n8253) );
  AND2_X1 U5461 ( .A1(n5550), .A2(n5549), .ZN(n8147) );
  NAND2_X1 U5462 ( .A1(n7893), .A2(n7892), .ZN(n8560) );
  AOI21_X1 U5463 ( .B1(n8093), .B2(n9946), .A(n6502), .ZN(n6514) );
  OAI21_X1 U5464 ( .B1(n6601), .B2(n5249), .A(n4575), .ZN(n7312) );
  AND2_X1 U5465 ( .A1(n5178), .A2(n4501), .ZN(n4575) );
  NAND2_X1 U5466 ( .A1(n6514), .A2(n9949), .ZN(n4981) );
  INV_X1 U5467 ( .A(n6472), .ZN(n8072) );
  NAND2_X1 U5468 ( .A1(n5060), .A2(n5059), .ZN(n8530) );
  OR2_X1 U5469 ( .A1(n5058), .A2(n5057), .ZN(n5059) );
  NAND2_X1 U5470 ( .A1(n5944), .A2(n5943), .ZN(n7219) );
  INV_X1 U5471 ( .A(n4687), .ZN(n4693) );
  OAI21_X1 U5472 ( .B1(n8734), .B2(n4689), .A(n4688), .ZN(n4687) );
  NAND2_X1 U5473 ( .A1(n4695), .A2(n4692), .ZN(n4689) );
  AOI21_X1 U5474 ( .B1(n6316), .B2(n4695), .A(n4694), .ZN(n4688) );
  NAND2_X1 U5475 ( .A1(n6316), .A2(n4696), .ZN(n4690) );
  NAND2_X1 U5476 ( .A1(n4696), .A2(n4692), .ZN(n4691) );
  NOR2_X1 U5477 ( .A1(n6333), .A2(n6334), .ZN(n4696) );
  NAND2_X1 U5478 ( .A1(n6134), .A2(n6133), .ZN(n9173) );
  NAND2_X1 U5479 ( .A1(n6250), .A2(n6249), .ZN(n9451) );
  NAND2_X1 U5480 ( .A1(n4473), .A2(n4618), .ZN(n4623) );
  NAND3_X1 U5481 ( .A1(n5889), .A2(n4488), .A3(n5890), .ZN(n9138) );
  NAND4_X1 U5482 ( .A1(n5858), .A2(n5857), .A3(n5856), .A4(n5855), .ZN(n9140)
         );
  OR2_X1 U5483 ( .A1(n5866), .A2(n5853), .ZN(n5857) );
  NOR2_X1 U5484 ( .A1(n9664), .A2(n4568), .ZN(n9685) );
  AND2_X1 U5485 ( .A1(n9668), .A2(n7034), .ZN(n4568) );
  NOR2_X1 U5486 ( .A1(n9167), .A2(n9223), .ZN(n4585) );
  AND2_X1 U5487 ( .A1(n9422), .A2(n9250), .ZN(n9190) );
  NAND2_X1 U5488 ( .A1(n6936), .A2(n6873), .ZN(n6876) );
  OAI211_X1 U5489 ( .C1(n6594), .C2(n5834), .A(n5833), .B(n5832), .ZN(n8793)
         );
  AND2_X1 U5490 ( .A1(n5775), .A2(n4584), .ZN(n9156) );
  AOI21_X1 U5491 ( .B1(n9755), .B2(n6342), .A(n6341), .ZN(n6775) );
  AND2_X1 U5492 ( .A1(n4973), .A2(n4972), .ZN(n4971) );
  INV_X1 U5493 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4972) );
  NOR2_X1 U5494 ( .A1(n7954), .A2(n8059), .ZN(n4723) );
  INV_X1 U5495 ( .A(n8532), .ZN(n4733) );
  AOI21_X1 U5496 ( .B1(n7980), .B2(n7976), .A(n4762), .ZN(n7978) );
  NOR2_X1 U5497 ( .A1(n9199), .A2(n4603), .ZN(n4602) );
  INV_X1 U5498 ( .A(n9198), .ZN(n4603) );
  NAND2_X1 U5499 ( .A1(n4599), .A2(n8997), .ZN(n4598) );
  NAND2_X1 U5500 ( .A1(n8996), .A2(n8995), .ZN(n4599) );
  NAND2_X1 U5501 ( .A1(n9010), .A2(n9009), .ZN(n9019) );
  OAI211_X1 U5502 ( .C1(n9005), .C2(n9032), .A(n4610), .B(n9008), .ZN(n9009)
         );
  OAI21_X1 U5503 ( .B1(n8032), .B2(n8023), .A(n8031), .ZN(n8027) );
  AND2_X1 U5504 ( .A1(n8405), .A2(n8036), .ZN(n4713) );
  NAND2_X1 U5505 ( .A1(n6921), .A2(n8890), .ZN(n9086) );
  NAND2_X1 U5506 ( .A1(n4618), .A2(n4675), .ZN(n8882) );
  AND2_X1 U5507 ( .A1(n8726), .A2(n4913), .ZN(n4912) );
  NAND2_X1 U5508 ( .A1(n8767), .A2(n4914), .ZN(n4913) );
  INV_X1 U5509 ( .A(n8766), .ZN(n4914) );
  INV_X1 U5510 ( .A(n5333), .ZN(n4886) );
  INV_X1 U5511 ( .A(SI_12_), .ZN(n10159) );
  NAND2_X1 U5512 ( .A1(n7919), .A2(n4746), .ZN(n4745) );
  NOR2_X1 U5513 ( .A1(n8048), .A2(n8356), .ZN(n4744) );
  NAND2_X1 U5514 ( .A1(n8056), .A2(n4740), .ZN(n4739) );
  NOR2_X1 U5515 ( .A1(n4742), .A2(n4741), .ZN(n4740) );
  INV_X1 U5516 ( .A(n8054), .ZN(n4741) );
  INV_X1 U5517 ( .A(n8055), .ZN(n4742) );
  NAND2_X2 U5518 ( .A1(n8070), .A2(n7923), .ZN(n8059) );
  OR2_X1 U5519 ( .A1(n6495), .A2(n5211), .ZN(n5212) );
  NAND2_X1 U5520 ( .A1(n4990), .A2(n8393), .ZN(n4989) );
  NAND2_X1 U5521 ( .A1(n4991), .A2(n4993), .ZN(n4990) );
  NOR2_X1 U5522 ( .A1(n4776), .A2(n8368), .ZN(n4775) );
  INV_X1 U5523 ( .A(n6488), .ZN(n4776) );
  NOR2_X1 U5524 ( .A1(n8410), .A2(n8577), .ZN(n4708) );
  INV_X1 U5525 ( .A(n4998), .ZN(n4996) );
  OR2_X1 U5526 ( .A1(n8590), .A2(n8123), .ZN(n8036) );
  NAND2_X1 U5527 ( .A1(n7924), .A2(n7949), .ZN(n7944) );
  NAND2_X1 U5528 ( .A1(n8273), .A2(n9912), .ZN(n7940) );
  NAND2_X1 U5529 ( .A1(n8274), .A2(n6422), .ZN(n7933) );
  AND2_X1 U5530 ( .A1(n8423), .A2(n4706), .ZN(n8360) );
  AND2_X1 U5531 ( .A1(n4479), .A2(n8364), .ZN(n4706) );
  NAND2_X1 U5532 ( .A1(n5681), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5697) );
  OR2_X1 U5533 ( .A1(n5194), .A2(n5193), .ZN(n5216) );
  XNOR2_X1 U5534 ( .A(n4674), .B(n6309), .ZN(n5823) );
  NAND2_X1 U5535 ( .A1(n5820), .A2(n4559), .ZN(n4674) );
  NAND2_X1 U5536 ( .A1(n5792), .A2(n6948), .ZN(n4559) );
  NOR2_X1 U5537 ( .A1(n4925), .A2(n8712), .ZN(n4924) );
  NAND2_X1 U5538 ( .A1(n4925), .A2(n8712), .ZN(n4923) );
  NAND2_X1 U5539 ( .A1(n8759), .A2(n6285), .ZN(n4926) );
  NAND2_X1 U5540 ( .A1(n5958), .A2(n5957), .ZN(n5973) );
  NAND2_X1 U5541 ( .A1(n5797), .A2(n5770), .ZN(n5809) );
  NOR2_X1 U5542 ( .A1(n6089), .A2(n6088), .ZN(n6106) );
  NOR2_X1 U5543 ( .A1(n7071), .A2(n4561), .ZN(n6543) );
  AND2_X1 U5544 ( .A1(n6569), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4561) );
  NOR2_X1 U5545 ( .A1(n9442), .A2(n9447), .ZN(n4594) );
  AND2_X1 U5546 ( .A1(n6106), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6135) );
  NOR2_X1 U5547 ( .A1(n7848), .A2(n4835), .ZN(n4834) );
  INV_X1 U5548 ( .A(n8980), .ZN(n4835) );
  INV_X1 U5549 ( .A(n8986), .ZN(n4833) );
  OR2_X1 U5550 ( .A1(n7785), .A2(n7784), .ZN(n4836) );
  NAND2_X1 U5551 ( .A1(n4836), .A2(n4834), .ZN(n7845) );
  NAND2_X1 U5552 ( .A1(n7646), .A2(n9072), .ZN(n7645) );
  INV_X1 U5553 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6048) );
  OR2_X1 U5554 ( .A1(n7745), .A2(n7732), .ZN(n8968) );
  NAND2_X1 U5555 ( .A1(n6020), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6049) );
  INV_X1 U5556 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5962) );
  INV_X1 U5557 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U5558 ( .A1(n8885), .A2(n8886), .ZN(n6874) );
  NAND2_X1 U5559 ( .A1(n5749), .A2(n4633), .ZN(n6363) );
  NAND2_X1 U5560 ( .A1(n7400), .A2(n9792), .ZN(n9586) );
  NOR2_X1 U5561 ( .A1(n6919), .A2(n6968), .ZN(n7147) );
  NAND2_X1 U5562 ( .A1(n6468), .A2(n6467), .ZN(n7873) );
  INV_X1 U5563 ( .A(SI_17_), .ZN(n5430) );
  NAND2_X1 U5564 ( .A1(n5429), .A2(n5428), .ZN(n5457) );
  AOI21_X1 U5565 ( .B1(n4873), .B2(n4876), .A(n4872), .ZN(n4871) );
  NOR2_X1 U5566 ( .A1(n5383), .A2(n4881), .ZN(n4880) );
  INV_X1 U5567 ( .A(n5357), .ZN(n4881) );
  XNOR2_X1 U5568 ( .A(n5381), .B(n10113), .ZN(n5380) );
  NAND2_X1 U5569 ( .A1(n5336), .A2(n10303), .ZN(n5357) );
  OAI21_X1 U5570 ( .B1(n5242), .B2(n5241), .A(n5243), .ZN(n5260) );
  AND2_X1 U5571 ( .A1(n5261), .A2(n5248), .ZN(n5020) );
  NAND2_X1 U5572 ( .A1(n5830), .A2(n5742), .ZN(n5848) );
  OAI21_X1 U5573 ( .B1(n6582), .B2(n4738), .A(n4737), .ZN(n5112) );
  NAND2_X1 U5574 ( .A1(n4858), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4857) );
  OR2_X1 U5575 ( .A1(n8113), .A2(n8114), .ZN(n8111) );
  INV_X1 U5576 ( .A(n7407), .ZN(n4820) );
  NAND2_X1 U5577 ( .A1(n5073), .A2(n5072), .ZN(n4798) );
  INV_X1 U5578 ( .A(n4818), .ZN(n4817) );
  AND2_X1 U5579 ( .A1(n5425), .A2(n4815), .ZN(n4814) );
  NAND2_X1 U5580 ( .A1(n5572), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5604) );
  INV_X1 U5581 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U5582 ( .A1(n5505), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5525) );
  INV_X1 U5583 ( .A(n5507), .ZN(n5505) );
  NAND2_X1 U5584 ( .A1(n4804), .A2(n4803), .ZN(n6523) );
  AND2_X1 U5585 ( .A1(n5714), .A2(n6679), .ZN(n8228) );
  AND2_X1 U5586 ( .A1(n8560), .A2(n7898), .ZN(n7902) );
  NAND2_X1 U5587 ( .A1(n7896), .A2(n8642), .ZN(n4758) );
  NOR2_X1 U5588 ( .A1(n8347), .A2(n7937), .ZN(n4757) );
  AND2_X1 U5589 ( .A1(n9897), .A2(n8065), .ZN(n8070) );
  OR2_X1 U5590 ( .A1(n6503), .A2(P2_U3152), .ZN(n8078) );
  INV_X1 U5591 ( .A(n8228), .ZN(n9812) );
  AND4_X1 U5592 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n7824)
         );
  AND4_X1 U5593 ( .A1(n5374), .A2(n5373), .A3(n5372), .A4(n5371), .ZN(n7823)
         );
  AND4_X1 U5594 ( .A1(n5348), .A2(n5347), .A3(n5346), .A4(n5345), .ZN(n7753)
         );
  AND4_X1 U5595 ( .A1(n5327), .A2(n5326), .A3(n5325), .A4(n5324), .ZN(n7709)
         );
  AND4_X1 U5596 ( .A1(n5299), .A2(n5298), .A3(n5297), .A4(n5296), .ZN(n7535)
         );
  AND4_X1 U5597 ( .A1(n5240), .A2(n5239), .A3(n5238), .A4(n5237), .ZN(n7472)
         );
  OR2_X1 U5598 ( .A1(n5167), .A2(n5104), .ZN(n5105) );
  NOR2_X1 U5599 ( .A1(n9541), .A2(n4668), .ZN(n9539) );
  NAND2_X1 U5600 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n4668) );
  NOR2_X1 U5601 ( .A1(n9555), .A2(n4495), .ZN(n6713) );
  NOR2_X1 U5602 ( .A1(n6713), .A2(n6712), .ZN(n6711) );
  OR2_X1 U5603 ( .A1(n6752), .A2(n6751), .ZN(n4659) );
  NOR2_X1 U5604 ( .A1(n7106), .A2(n4662), .ZN(n7110) );
  AND2_X1 U5605 ( .A1(n7107), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4662) );
  NAND2_X1 U5606 ( .A1(n7110), .A2(n7109), .ZN(n7200) );
  NAND2_X1 U5607 ( .A1(n7200), .A2(n4661), .ZN(n7202) );
  OR2_X1 U5608 ( .A1(n7201), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4661) );
  NAND2_X1 U5609 ( .A1(n7336), .A2(n7337), .ZN(n7590) );
  NAND2_X1 U5610 ( .A1(n7339), .A2(n5367), .ZN(n4657) );
  OR2_X1 U5611 ( .A1(n5623), .A2(n10288), .ZN(n5656) );
  INV_X1 U5612 ( .A(n8047), .ZN(n4777) );
  NAND2_X1 U5613 ( .A1(n6489), .A2(n4775), .ZN(n4778) );
  NAND2_X1 U5614 ( .A1(n6489), .A2(n6488), .ZN(n8369) );
  NAND2_X1 U5615 ( .A1(n8423), .A2(n4708), .ZN(n8384) );
  NAND2_X1 U5616 ( .A1(n8423), .A2(n8653), .ZN(n8398) );
  NAND2_X1 U5617 ( .A1(n4573), .A2(n8024), .ZN(n4572) );
  INV_X1 U5618 ( .A(n6485), .ZN(n8450) );
  NAND2_X1 U5619 ( .A1(n8486), .A2(n8468), .ZN(n8463) );
  NAND2_X1 U5620 ( .A1(n4699), .A2(n6453), .ZN(n8500) );
  INV_X1 U5621 ( .A(n5462), .ZN(n5461) );
  AOI21_X1 U5622 ( .B1(n4477), .B2(n8542), .A(n4522), .ZN(n5014) );
  NAND2_X1 U5623 ( .A1(n5397), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U5624 ( .A1(n4570), .A2(n4767), .ZN(n8543) );
  INV_X1 U5625 ( .A(n4768), .ZN(n4767) );
  OAI21_X1 U5626 ( .B1(n7989), .B2(n4769), .A(n7996), .ZN(n4768) );
  AND2_X1 U5627 ( .A1(n7717), .A2(n4541), .ZN(n8549) );
  NAND2_X1 U5628 ( .A1(n5005), .A2(n5011), .ZN(n5003) );
  AOI21_X1 U5629 ( .B1(n5008), .B2(n5005), .A(n4483), .ZN(n5002) );
  NAND2_X1 U5630 ( .A1(n7717), .A2(n4704), .ZN(n7829) );
  NAND2_X1 U5631 ( .A1(n7717), .A2(n7979), .ZN(n7760) );
  INV_X1 U5632 ( .A(n7750), .ZN(n4772) );
  AOI21_X1 U5633 ( .B1(n4763), .B2(n4766), .A(n4762), .ZN(n4761) );
  INV_X1 U5634 ( .A(n7967), .ZN(n4766) );
  OR2_X1 U5635 ( .A1(n5343), .A2(n7205), .ZN(n5369) );
  NAND2_X1 U5636 ( .A1(n7513), .A2(n7967), .ZN(n7533) );
  NAND2_X1 U5637 ( .A1(n7469), .A2(n7966), .ZN(n7513) );
  OR2_X1 U5638 ( .A1(n5274), .A2(n10112), .ZN(n5293) );
  OR2_X1 U5639 ( .A1(n5235), .A2(n5234), .ZN(n5274) );
  NAND2_X1 U5640 ( .A1(n7364), .A2(n7910), .ZN(n7363) );
  AND2_X1 U5641 ( .A1(n6439), .A2(n7350), .ZN(n7351) );
  NAND2_X1 U5642 ( .A1(n4581), .A2(n7960), .ZN(n7344) );
  NAND2_X1 U5643 ( .A1(n4754), .A2(n4752), .ZN(n4581) );
  NOR2_X1 U5644 ( .A1(n4755), .A2(n4753), .ZN(n4752) );
  AND2_X1 U5645 ( .A1(n9842), .A2(n9929), .ZN(n9843) );
  OR2_X1 U5646 ( .A1(n9942), .A2(n8530), .ZN(n6505) );
  INV_X1 U5647 ( .A(n5199), .ZN(n5483) );
  INV_X1 U5648 ( .A(n6689), .ZN(n6666) );
  INV_X1 U5649 ( .A(n9940), .ZN(n9918) );
  OR2_X1 U5650 ( .A1(n9897), .A2(n5725), .ZN(n9940) );
  NAND2_X1 U5651 ( .A1(n5061), .A2(n5062), .ZN(n5043) );
  XNOR2_X1 U5652 ( .A(n4830), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6472) );
  NAND2_X1 U5653 ( .A1(n5060), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U5654 ( .A1(n5056), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5058) );
  INV_X1 U5655 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U5656 ( .A1(n5058), .A2(n5057), .ZN(n5060) );
  AND2_X1 U5657 ( .A1(n5287), .A2(n5271), .ZN(n6997) );
  NOR2_X1 U5658 ( .A1(n5216), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5251) );
  INV_X1 U5659 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5250) );
  INV_X1 U5660 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5191) );
  AND2_X1 U5661 ( .A1(n5172), .A2(n5153), .ZN(n6728) );
  INV_X1 U5662 ( .A(n6334), .ZN(n4694) );
  INV_X1 U5663 ( .A(n6333), .ZN(n4695) );
  AND2_X1 U5664 ( .A1(n6118), .A2(n7724), .ZN(n4928) );
  AOI21_X1 U5665 ( .B1(n4907), .B2(n4905), .A(n4510), .ZN(n4904) );
  INV_X1 U5666 ( .A(n6014), .ZN(n4905) );
  NAND2_X1 U5667 ( .A1(n7443), .A2(n4685), .ZN(n4684) );
  NOR2_X1 U5668 ( .A1(n4906), .A2(n4686), .ZN(n4685) );
  INV_X1 U5669 ( .A(n5996), .ZN(n4686) );
  INV_X1 U5670 ( .A(n4907), .ZN(n4906) );
  AND2_X1 U5671 ( .A1(n6135), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U5672 ( .A1(n6270), .A2(n6269), .ZN(n8711) );
  INV_X1 U5673 ( .A(n6270), .ZN(n4922) );
  AND2_X1 U5674 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5888) );
  OR2_X1 U5675 ( .A1(n5963), .A2(n5962), .ZN(n5982) );
  NOR2_X1 U5676 ( .A1(n5982), .A2(n7446), .ZN(n6003) );
  AND2_X1 U5677 ( .A1(n6196), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6236) );
  AND2_X1 U5678 ( .A1(n8720), .A2(n4679), .ZN(n4678) );
  NAND2_X1 U5679 ( .A1(n6236), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6254) );
  OR2_X1 U5680 ( .A1(n7485), .A2(n7484), .ZN(n6014) );
  OR2_X1 U5681 ( .A1(n8805), .A2(n8806), .ZN(n6316) );
  OR2_X1 U5682 ( .A1(n6803), .A2(n9754), .ZN(n6362) );
  OAI21_X1 U5683 ( .B1(n9081), .B2(n4890), .A(n9082), .ZN(n9118) );
  NAND2_X1 U5684 ( .A1(n9044), .A2(n4891), .ZN(n4890) );
  AND2_X1 U5685 ( .A1(n9045), .A2(n4504), .ZN(n4891) );
  NOR2_X1 U5686 ( .A1(n7073), .A2(n7072), .ZN(n7071) );
  OR2_X1 U5687 ( .A1(n7698), .A2(n7697), .ZN(n7695) );
  AND2_X1 U5688 ( .A1(n6548), .A2(n6520), .ZN(n6573) );
  NAND2_X1 U5689 ( .A1(n8843), .A2(n8842), .ZN(n9167) );
  NAND2_X1 U5690 ( .A1(n4636), .A2(n4635), .ZN(n9232) );
  AOI21_X1 U5691 ( .B1(n4482), .B2(n4637), .A(n9107), .ZN(n4635) );
  INV_X1 U5692 ( .A(n9233), .ZN(n4842) );
  AND2_X1 U5693 ( .A1(n9209), .A2(n9026), .ZN(n9233) );
  AOI21_X1 U5694 ( .B1(n9206), .B2(n4639), .A(n4638), .ZN(n4637) );
  INV_X1 U5695 ( .A(n9205), .ZN(n4639) );
  NOR2_X1 U5696 ( .A1(n9271), .A2(n9432), .ZN(n9256) );
  OR2_X1 U5697 ( .A1(n9189), .A2(n9078), .ZN(n9264) );
  AOI21_X1 U5698 ( .B1(n4960), .B2(n4964), .A(n4521), .ZN(n4959) );
  NAND2_X1 U5699 ( .A1(n9309), .A2(n4592), .ZN(n9271) );
  NOR2_X1 U5700 ( .A1(n9437), .A2(n4593), .ZN(n4592) );
  INV_X1 U5701 ( .A(n4594), .ZN(n4593) );
  NOR2_X1 U5702 ( .A1(n6274), .A2(n8761), .ZN(n6289) );
  NAND2_X1 U5703 ( .A1(n9309), .A2(n9301), .ZN(n9295) );
  NOR2_X1 U5704 ( .A1(n9321), .A2(n9451), .ZN(n9309) );
  NAND2_X1 U5705 ( .A1(n9338), .A2(n9181), .ZN(n4946) );
  OR2_X1 U5706 ( .A1(n9325), .A2(n9199), .ZN(n9347) );
  AOI21_X1 U5707 ( .B1(n9196), .B2(n4643), .A(n4641), .ZN(n4640) );
  INV_X1 U5708 ( .A(n9196), .ZN(n4642) );
  NAND2_X1 U5709 ( .A1(n9373), .A2(n9196), .ZN(n9364) );
  AND2_X1 U5710 ( .A1(n9049), .A2(n9198), .ZN(n9361) );
  NAND2_X1 U5711 ( .A1(n9194), .A2(n8873), .ZN(n9373) );
  NAND2_X1 U5712 ( .A1(n7653), .A2(n4481), .ZN(n9391) );
  NOR2_X1 U5713 ( .A1(n7655), .A2(n4896), .ZN(n7854) );
  NAND2_X1 U5714 ( .A1(n4836), .A2(n8980), .ZN(n7847) );
  OR2_X1 U5715 ( .A1(n6070), .A2(n6069), .ZN(n6089) );
  NAND2_X1 U5716 ( .A1(n7653), .A2(n7656), .ZN(n7655) );
  AOI21_X1 U5717 ( .B1(n4949), .B2(n4955), .A(n4507), .ZN(n4947) );
  AND2_X1 U5718 ( .A1(n7400), .A2(n4486), .ZN(n7568) );
  NAND2_X1 U5719 ( .A1(n7400), .A2(n4590), .ZN(n9588) );
  NOR2_X1 U5720 ( .A1(n5925), .A2(n5924), .ZN(n5945) );
  NAND2_X1 U5721 ( .A1(n7148), .A2(n7147), .ZN(n7241) );
  NAND2_X1 U5722 ( .A1(n4582), .A2(n9779), .ZN(n7243) );
  INV_X1 U5723 ( .A(n7241), .ZN(n4582) );
  INV_X1 U5724 ( .A(n8890), .ZN(n4609) );
  AND2_X1 U5725 ( .A1(n4608), .A2(n9087), .ZN(n4607) );
  NAND2_X1 U5726 ( .A1(n9767), .A2(n6920), .ZN(n6919) );
  NAND2_X1 U5727 ( .A1(n6904), .A2(n8885), .ZN(n6921) );
  NAND2_X1 U5728 ( .A1(n4618), .A2(n6948), .ZN(n6873) );
  INV_X1 U5729 ( .A(n9053), .ZN(n6938) );
  OAI21_X1 U5730 ( .B1(n4584), .B2(n4583), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4903) );
  OR2_X1 U5731 ( .A1(n9490), .A2(n4673), .ZN(n6770) );
  NAND2_X1 U5732 ( .A1(n6193), .A2(n6192), .ZN(n9468) );
  INV_X1 U5733 ( .A(n9788), .ZN(n9484) );
  NAND2_X1 U5734 ( .A1(n7025), .A2(n7024), .ZN(n7145) );
  INV_X1 U5735 ( .A(n9793), .ZN(n9764) );
  INV_X1 U5736 ( .A(n6933), .ZN(n6945) );
  XNOR2_X1 U5737 ( .A(n7873), .B(n7872), .ZN(n8851) );
  NAND2_X1 U5738 ( .A1(n4861), .A2(n4859), .ZN(n5648) );
  AND2_X1 U5739 ( .A1(n4860), .A2(n4865), .ZN(n4859) );
  AOI21_X1 U5740 ( .B1(n5631), .B2(n4867), .A(n4866), .ZN(n4865) );
  AND2_X1 U5741 ( .A1(n5649), .A2(n5636), .ZN(n5647) );
  NAND2_X1 U5742 ( .A1(n4868), .A2(n5615), .ZN(n5632) );
  NAND2_X1 U5743 ( .A1(n4869), .A2(n4863), .ZN(n4868) );
  NAND2_X1 U5744 ( .A1(n4936), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5756) );
  INV_X1 U5745 ( .A(n5763), .ZN(n5764) );
  AND2_X1 U5746 ( .A1(n6169), .A2(n6153), .ZN(n9145) );
  OAI21_X1 U5747 ( .B1(n5358), .B2(n4876), .A(n4873), .ZN(n5427) );
  OR2_X1 U5748 ( .A1(n6039), .A2(n6038), .ZN(n6042) );
  OR2_X1 U5749 ( .A1(n6042), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U5750 ( .A1(n4882), .A2(n5307), .ZN(n5334) );
  NAND2_X1 U5751 ( .A1(n5286), .A2(n4887), .ZN(n4882) );
  NAND2_X1 U5752 ( .A1(n5286), .A2(n5285), .ZN(n5309) );
  AOI21_X1 U5753 ( .B1(n4850), .B2(n5196), .A(n4527), .ZN(n4849) );
  AND2_X1 U5754 ( .A1(n5897), .A2(n5896), .ZN(n5915) );
  XNOR2_X1 U5755 ( .A(n5819), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U5756 ( .A1(n4821), .A2(n4822), .ZN(n7408) );
  NAND2_X1 U5757 ( .A1(n5564), .A2(n5563), .ZN(n8442) );
  OAI21_X1 U5758 ( .B1(n7493), .B2(n4809), .A(n4806), .ZN(n7613) );
  NAND2_X1 U5759 ( .A1(n6854), .A2(n5103), .ZN(n6868) );
  NAND2_X1 U5760 ( .A1(n5710), .A2(n8247), .ZN(n4792) );
  INV_X1 U5761 ( .A(n4801), .ZN(n4800) );
  OAI21_X1 U5762 ( .B1(n4493), .B2(n4802), .A(n8143), .ZN(n4801) );
  INV_X1 U5763 ( .A(n5518), .ZN(n4802) );
  NAND2_X1 U5764 ( .A1(n8198), .A2(n5518), .ZN(n8144) );
  NOR2_X1 U5765 ( .A1(n5022), .A2(n4795), .ZN(n4794) );
  INV_X1 U5766 ( .A(n9811), .ZN(n4795) );
  INV_X1 U5767 ( .A(n7377), .ZN(n9933) );
  NAND2_X1 U5768 ( .A1(n4813), .A2(n4811), .ZN(n7548) );
  AND2_X1 U5769 ( .A1(n4813), .A2(n4810), .ZN(n7550) );
  NAND2_X1 U5770 ( .A1(n7493), .A2(n7494), .ZN(n4813) );
  NAND2_X1 U5771 ( .A1(n8132), .A2(n4493), .ZN(n8198) );
  NAND2_X1 U5772 ( .A1(n5544), .A2(n5543), .ZN(n8600) );
  AND2_X1 U5773 ( .A1(n5704), .A2(n9845), .ZN(n9819) );
  INV_X1 U5774 ( .A(n8247), .ZN(n9821) );
  INV_X1 U5775 ( .A(n9819), .ZN(n8244) );
  NAND2_X1 U5776 ( .A1(n5127), .A2(n5126), .ZN(n8271) );
  NAND2_X1 U5777 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  NOR2_X1 U5778 ( .A1(n6711), .A2(n4663), .ZN(n6762) );
  AND2_X1 U5779 ( .A1(n6697), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4663) );
  NOR2_X1 U5780 ( .A1(n6726), .A2(n6725), .ZN(n6735) );
  NOR2_X1 U5781 ( .A1(n6735), .A2(n4660), .ZN(n6752) );
  NOR2_X1 U5782 ( .A1(n6743), .A2(n6724), .ZN(n4660) );
  INV_X1 U5783 ( .A(n4659), .ZN(n6750) );
  AND2_X1 U5784 ( .A1(n4659), .A2(n4658), .ZN(n6738) );
  NAND2_X1 U5785 ( .A1(n6740), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4658) );
  INV_X1 U5786 ( .A(n4665), .ZN(n6840) );
  NOR2_X1 U5787 ( .A1(n6843), .A2(n6842), .ZN(n6996) );
  AND2_X1 U5788 ( .A1(n4665), .A2(n4664), .ZN(n6843) );
  NAND2_X1 U5789 ( .A1(n6845), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4664) );
  AOI21_X1 U5790 ( .B1(n4655), .B2(n4650), .A(n4656), .ZN(n4649) );
  OR2_X1 U5791 ( .A1(n7336), .A2(n4653), .ZN(n4652) );
  XNOR2_X1 U5792 ( .A(n4670), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U5793 ( .A1(n8329), .A2(n4555), .ZN(n4670) );
  INV_X1 U5794 ( .A(n9830), .ZN(n9825) );
  NAND2_X1 U5795 ( .A1(n4514), .A2(n9841), .ZN(n8561) );
  NAND2_X1 U5796 ( .A1(n6500), .A2(n6499), .ZN(n6501) );
  XNOR2_X1 U5797 ( .A(n7879), .B(n8051), .ZN(n4579) );
  NAND2_X1 U5798 ( .A1(n8051), .A2(n4982), .ZN(n4979) );
  OAI21_X1 U5799 ( .B1(n6490), .B2(n4978), .A(n4977), .ZN(n4976) );
  NAND2_X1 U5800 ( .A1(n8355), .A2(n4499), .ZN(n4975) );
  NAND2_X1 U5801 ( .A1(n4577), .A2(n8040), .ZN(n8389) );
  OAI21_X1 U5802 ( .B1(n8415), .B2(n4993), .A(n4991), .ZN(n8394) );
  NOR2_X1 U5803 ( .A1(n8414), .A2(n4998), .ZN(n8406) );
  NAND2_X1 U5804 ( .A1(n4779), .A2(n4574), .ZN(n8471) );
  NAND2_X1 U5805 ( .A1(n4783), .A2(n8018), .ZN(n8479) );
  NAND2_X1 U5806 ( .A1(n6483), .A2(n8007), .ZN(n8497) );
  NAND2_X1 U5807 ( .A1(n5016), .A2(n4477), .ZN(n8531) );
  AND2_X1 U5808 ( .A1(n5016), .A2(n5015), .ZN(n8533) );
  NAND2_X1 U5809 ( .A1(n7713), .A2(n6448), .ZN(n7758) );
  NAND2_X1 U5810 ( .A1(n5010), .A2(n5009), .ZN(n7715) );
  NAND2_X1 U5811 ( .A1(n7467), .A2(n6444), .ZN(n7512) );
  INV_X1 U5812 ( .A(n7617), .ZN(n7481) );
  NAND2_X1 U5813 ( .A1(n4754), .A2(n7958), .ZN(n7260) );
  OR2_X1 U5814 ( .A1(n9855), .A2(n7017), .ZN(n9851) );
  INV_X1 U5815 ( .A(n8506), .ZN(n9853) );
  OR2_X1 U5816 ( .A1(n5249), .A2(n6583), .ZN(n5115) );
  OR2_X1 U5817 ( .A1(n5249), .A2(n6594), .ZN(n5096) );
  OR2_X1 U5818 ( .A1(n4476), .A2(n6595), .ZN(n5097) );
  OR2_X1 U5819 ( .A1(n7042), .A2(n7923), .ZN(n9847) );
  INV_X1 U5820 ( .A(n9851), .ZN(n8534) );
  AND2_X1 U5821 ( .A1(n8561), .A2(n8563), .ZN(n8635) );
  INV_X1 U5822 ( .A(n8442), .ZN(n8658) );
  INV_X1 U5823 ( .A(n8514), .ZN(n8669) );
  INV_X1 U5824 ( .A(n7771), .ZN(n7669) );
  AND2_X2 U5825 ( .A1(n7011), .A2(n6513), .ZN(n9949) );
  NOR2_X1 U5826 ( .A1(n6582), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8683) );
  INV_X1 U5827 ( .A(n4986), .ZN(n5686) );
  XNOR2_X1 U5828 ( .A(n5683), .B(n5682), .ZN(n7694) );
  NAND2_X1 U5829 ( .A1(n5699), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5683) );
  INV_X1 U5830 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7531) );
  INV_X1 U5831 ( .A(n8079), .ZN(n7530) );
  INV_X1 U5832 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7464) );
  INV_X1 U5833 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7441) );
  INV_X1 U5834 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7306) );
  INV_X1 U5835 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6986) );
  INV_X1 U5836 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6833) );
  INV_X1 U5837 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6786) );
  INV_X1 U5838 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6671) );
  INV_X1 U5839 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6646) );
  INV_X1 U5840 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6602) );
  XNOR2_X1 U5841 ( .A(n4669), .B(n5065), .ZN(n9546) );
  NAND2_X1 U5842 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4669) );
  NAND2_X1 U5843 ( .A1(n7443), .A2(n5996), .ZN(n7487) );
  NAND2_X1 U5844 ( .A1(n5961), .A2(n5960), .ZN(n7436) );
  AOI22_X1 U5845 ( .A1(n6397), .A2(n6948), .B1(n6872), .B2(n5808), .ZN(n6862)
         );
  NAND2_X1 U5846 ( .A1(n4911), .A2(n8767), .ZN(n8725) );
  NAND2_X1 U5847 ( .A1(n8769), .A2(n8766), .ZN(n4911) );
  INV_X1 U5848 ( .A(n4933), .ZN(n4932) );
  NAND2_X1 U5849 ( .A1(n5912), .A2(n5908), .ZN(n7080) );
  NAND2_X1 U5850 ( .A1(n8741), .A2(n6147), .ZN(n8752) );
  NAND2_X1 U5851 ( .A1(n6975), .A2(n5865), .ZN(n6965) );
  INV_X1 U5852 ( .A(n8811), .ZN(n8824) );
  AND2_X1 U5853 ( .A1(n5977), .A2(n7429), .ZN(n7442) );
  NAND2_X1 U5854 ( .A1(n6214), .A2(n6213), .ZN(n9464) );
  NAND2_X1 U5855 ( .A1(n7737), .A2(n6064), .ZN(n7727) );
  OAI21_X1 U5856 ( .B1(n7487), .B2(n4494), .A(n6014), .ZN(n7560) );
  NAND2_X1 U5857 ( .A1(n4682), .A2(n6188), .ZN(n8797) );
  NAND2_X1 U5858 ( .A1(n6105), .A2(n6104), .ZN(n9606) );
  NAND4_X1 U5859 ( .A1(n6329), .A2(n6328), .A3(n6327), .A4(n6326), .ZN(n9265)
         );
  NAND4_X1 U5860 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5871), .ZN(n9139)
         );
  OR2_X1 U5861 ( .A1(n5854), .A2(n6931), .ZN(n5802) );
  NAND2_X1 U5862 ( .A1(n4563), .A2(n4562), .ZN(n9530) );
  INV_X1 U5863 ( .A(n9527), .ZN(n4562) );
  INV_X1 U5864 ( .A(n4563), .ZN(n9528) );
  OAI21_X1 U5865 ( .B1(n9685), .B2(n6540), .A(n9684), .ZN(n9693) );
  AOI21_X1 U5866 ( .B1(n4841), .B2(n9574), .A(n4838), .ZN(n9424) );
  NAND2_X1 U5867 ( .A1(n4840), .A2(n4839), .ZN(n4838) );
  XNOR2_X1 U5868 ( .A(n9232), .B(n4842), .ZN(n4841) );
  NAND2_X1 U5869 ( .A1(n9234), .A2(n9400), .ZN(n4839) );
  NAND2_X1 U5870 ( .A1(n6393), .A2(n6392), .ZN(n9422) );
  NAND2_X1 U5871 ( .A1(n4962), .A2(n4963), .ZN(n9270) );
  OR2_X1 U5872 ( .A1(n9185), .A2(n4964), .ZN(n4962) );
  AND2_X1 U5873 ( .A1(n4646), .A2(n9203), .ZN(n9284) );
  NAND2_X1 U5874 ( .A1(n4968), .A2(n4491), .ZN(n9282) );
  OR2_X1 U5875 ( .A1(n9185), .A2(n9184), .ZN(n4968) );
  NAND2_X1 U5876 ( .A1(n9313), .A2(n9202), .ZN(n9302) );
  NAND2_X1 U5877 ( .A1(n4939), .A2(n4940), .ZN(n9308) );
  NAND2_X1 U5878 ( .A1(n6234), .A2(n6233), .ZN(n9458) );
  NAND2_X1 U5879 ( .A1(n9194), .A2(n9193), .ZN(n9399) );
  NAND2_X1 U5880 ( .A1(n4950), .A2(n4951), .ZN(n7567) );
  OR2_X1 U5881 ( .A1(n7455), .A2(n4955), .ZN(n4950) );
  NAND2_X1 U5882 ( .A1(n4953), .A2(n4957), .ZN(n9567) );
  OR2_X1 U5883 ( .A1(n7455), .A2(n7454), .ZN(n4953) );
  NAND2_X1 U5884 ( .A1(n7178), .A2(n7177), .ZN(n7180) );
  INV_X1 U5885 ( .A(n9585), .ZN(n9396) );
  AND2_X1 U5886 ( .A1(n5019), .A2(n7026), .ZN(n7240) );
  OR2_X1 U5887 ( .A1(n9257), .A2(n9793), .ZN(n9225) );
  AOI21_X1 U5888 ( .B1(n9329), .B2(n4618), .A(n4551), .ZN(n6895) );
  OR2_X1 U5889 ( .A1(n9754), .A2(n6770), .ZN(n9743) );
  AND2_X1 U5890 ( .A1(n4621), .A2(n4552), .ZN(n6930) );
  NAND2_X1 U5891 ( .A1(n9348), .A2(n4618), .ZN(n4621) );
  AND2_X1 U5892 ( .A1(n9751), .A2(n9738), .ZN(n9585) );
  INV_X1 U5893 ( .A(n9225), .ZN(n9406) );
  AND3_X2 U5894 ( .A1(n6782), .A2(n6781), .A3(n6805), .ZN(n9809) );
  OAI21_X1 U5895 ( .B1(n9409), .B2(n9793), .A(n4586), .ZN(n9494) );
  NOR2_X1 U5896 ( .A1(n4503), .A2(n4587), .ZN(n4586) );
  INV_X1 U5897 ( .A(n9411), .ZN(n4587) );
  NOR2_X1 U5898 ( .A1(n9418), .A2(n9417), .ZN(n9419) );
  AND2_X2 U5899 ( .A1(n6782), .A2(n6878), .ZN(n9800) );
  AOI21_X1 U5900 ( .B1(n9755), .B2(n6354), .A(n6353), .ZN(n6877) );
  NAND2_X1 U5901 ( .A1(n4633), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5779) );
  XNOR2_X1 U5902 ( .A(n5648), .B(n5647), .ZN(n9519) );
  INV_X1 U5903 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U5904 ( .A1(n6355), .A2(n10072), .ZN(n5759) );
  INV_X1 U5905 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10122) );
  INV_X1 U5906 ( .A(n9127), .ZN(n9042) );
  INV_X1 U5907 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7452) );
  INV_X1 U5908 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7427) );
  INV_X1 U5909 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7308) );
  INV_X1 U5910 ( .A(n9156), .ZN(n9745) );
  INV_X1 U5911 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10097) );
  INV_X1 U5912 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10321) );
  AND2_X1 U5913 ( .A1(n6015), .A2(n6000), .ZN(n6816) );
  INV_X1 U5914 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6607) );
  INV_X1 U5915 ( .A(n9681), .ZN(n6606) );
  INV_X1 U5916 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6600) );
  XNOR2_X1 U5917 ( .A(n4576), .B(n5196), .ZN(n6601) );
  NAND2_X1 U5918 ( .A1(n4852), .A2(n5177), .ZN(n4576) );
  XNOR2_X1 U5919 ( .A(n5175), .B(n5174), .ZN(n6589) );
  NAND2_X1 U5920 ( .A1(n4829), .A2(n4826), .ZN(n7318) );
  OR2_X1 U5921 ( .A1(n8081), .A2(n8080), .ZN(n4556) );
  OAI21_X1 U5922 ( .B1(n8635), .B2(n9958), .A(n4700), .ZN(P2_U3551) );
  INV_X1 U5923 ( .A(n4701), .ZN(n4700) );
  OAI21_X1 U5924 ( .B1(n8638), .B2(n8634), .A(n4702), .ZN(n4701) );
  OR2_X1 U5925 ( .A1(n9960), .A2(n8562), .ZN(n4702) );
  NAND2_X1 U5926 ( .A1(n4981), .A2(n4980), .ZN(n6518) );
  OAI21_X1 U5927 ( .B1(n6403), .B2(n4693), .A(n8808), .ZN(n6391) );
  AOI22_X1 U5928 ( .A1(n8811), .A2(n4618), .B1(n8828), .B2(n6933), .ZN(n6811)
         );
  AND2_X1 U5929 ( .A1(n4623), .A2(n4622), .ZN(n8794) );
  NAND2_X1 U5930 ( .A1(n4553), .A2(n4625), .ZN(n4624) );
  NAND2_X1 U5931 ( .A1(n4630), .A2(n4627), .ZN(n4626) );
  INV_X1 U5932 ( .A(n9128), .ZN(n4625) );
  NAND2_X1 U5933 ( .A1(n4620), .A2(n4619), .ZN(P1_U3556) );
  NAND2_X1 U5934 ( .A1(P1_U4006), .A2(n4618), .ZN(n4619) );
  OR2_X1 U5935 ( .A1(P1_U4006), .A2(n6597), .ZN(n4620) );
  INV_X1 U5936 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U5937 ( .A1(n4567), .A2(n4564), .ZN(n9160) );
  INV_X1 U5938 ( .A(n5893), .ZN(n5846) );
  INV_X1 U5939 ( .A(n7470), .ZN(n6443) );
  AND2_X1 U5940 ( .A1(n6479), .A2(n7971), .ZN(n7470) );
  INV_X1 U5941 ( .A(n8733), .ZN(n4692) );
  AND2_X1 U5942 ( .A1(n8532), .A2(n5015), .ZN(n4477) );
  NAND2_X1 U5943 ( .A1(n5785), .A2(n5782), .ZN(n5869) );
  INV_X1 U5944 ( .A(n8356), .ZN(n4774) );
  XNOR2_X1 U5945 ( .A(n5769), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9122) );
  INV_X1 U5946 ( .A(n9122), .ZN(n4672) );
  NAND2_X1 U5947 ( .A1(n5570), .A2(n5569), .ZN(n8590) );
  OR2_X1 U5948 ( .A1(n4736), .A2(n4734), .ZN(n4478) );
  INV_X1 U5949 ( .A(n4955), .ZN(n4954) );
  NAND2_X1 U5950 ( .A1(n9572), .A2(n4956), .ZN(n4955) );
  AND2_X1 U5951 ( .A1(n4708), .A2(n4707), .ZN(n4479) );
  AND2_X1 U5952 ( .A1(n4904), .A2(n4683), .ZN(n4480) );
  AND2_X1 U5953 ( .A1(n4591), .A2(n9397), .ZN(n4481) );
  NAND2_X1 U5954 ( .A1(n9309), .A2(n4594), .ZN(n4595) );
  OR2_X1 U5955 ( .A1(n8487), .A2(n8146), .ZN(n8017) );
  INV_X1 U5956 ( .A(n8105), .ZN(n8250) );
  AND2_X1 U5957 ( .A1(n5664), .A2(n5663), .ZN(n8105) );
  AND2_X1 U5958 ( .A1(n9106), .A2(n9248), .ZN(n4482) );
  NOR2_X1 U5959 ( .A1(n8120), .A2(n8261), .ZN(n4483) );
  AND2_X1 U5960 ( .A1(n4704), .A2(n4703), .ZN(n4484) );
  AND2_X1 U5961 ( .A1(n5283), .A2(n5282), .ZN(n4485) );
  AND2_X1 U5962 ( .A1(n4590), .A2(n4589), .ZN(n4486) );
  NAND2_X1 U5963 ( .A1(n4684), .A2(n4904), .ZN(n7736) );
  NAND2_X1 U5964 ( .A1(n4772), .A2(n7989), .ZN(n7749) );
  AND2_X1 U5965 ( .A1(n4796), .A2(n4797), .ZN(n4487) );
  NAND2_X1 U5966 ( .A1(n6168), .A2(n6167), .ZN(n4682) );
  AND2_X1 U5967 ( .A1(n8053), .A2(n8052), .ZN(n8051) );
  AND2_X1 U5968 ( .A1(n5891), .A2(n5892), .ZN(n4488) );
  NAND4_X1 U5969 ( .A1(n5805), .A2(n5804), .A3(n5803), .A4(n5802), .ZN(n6776)
         );
  NAND2_X1 U5970 ( .A1(n6335), .A2(n5762), .ZN(n5797) );
  INV_X1 U5971 ( .A(n6269), .ZN(n4925) );
  AND2_X1 U5972 ( .A1(n4783), .A2(n4782), .ZN(n4489) );
  INV_X1 U5973 ( .A(n4584), .ZN(n5768) );
  OR2_X1 U5974 ( .A1(n9464), .A2(n9367), .ZN(n4490) );
  INV_X1 U5975 ( .A(n9293), .ZN(n4647) );
  OR2_X1 U5976 ( .A1(n9301), .A2(n9183), .ZN(n4491) );
  XNOR2_X1 U5977 ( .A(n8377), .B(n8227), .ZN(n8368) );
  AND2_X1 U5978 ( .A1(n9334), .A2(n4490), .ZN(n4492) );
  NAND2_X1 U5979 ( .A1(n4973), .A2(n5763), .ZN(n4633) );
  AND2_X1 U5980 ( .A1(n8199), .A2(n5496), .ZN(n4493) );
  AND2_X1 U5981 ( .A1(n6320), .A2(n6319), .ZN(n6333) );
  AND2_X1 U5982 ( .A1(n7485), .A2(n7484), .ZN(n4494) );
  AND2_X1 U5983 ( .A1(n9559), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4495) );
  INV_X1 U5984 ( .A(n7958), .ZN(n4753) );
  NAND2_X1 U5985 ( .A1(n5752), .A2(n5751), .ZN(n9447) );
  OR2_X1 U5986 ( .A1(n8356), .A2(n4777), .ZN(n4496) );
  AND2_X1 U5987 ( .A1(n6285), .A2(n4923), .ZN(n4497) );
  OR2_X1 U5988 ( .A1(n5249), .A2(n6596), .ZN(n4498) );
  NAND2_X1 U5989 ( .A1(n5485), .A2(n5484), .ZN(n8614) );
  NAND2_X1 U5990 ( .A1(n8835), .A2(n8834), .ZN(n8919) );
  AND2_X1 U5991 ( .A1(n6490), .A2(n8356), .ZN(n4499) );
  INV_X1 U5992 ( .A(n8007), .ZN(n4785) );
  NAND2_X1 U5993 ( .A1(n5408), .A2(n5407), .ZN(n8245) );
  INV_X1 U5994 ( .A(n8245), .ZN(n4703) );
  AND2_X1 U5995 ( .A1(n8711), .A2(n8712), .ZN(n4500) );
  NAND2_X1 U5996 ( .A1(n5638), .A2(n5637), .ZN(n8377) );
  INV_X1 U5997 ( .A(n8377), .ZN(n4707) );
  INV_X1 U5998 ( .A(n8480), .ZN(n4786) );
  INV_X1 U5999 ( .A(n7982), .ZN(n4762) );
  OR2_X1 U6000 ( .A1(n6689), .A2(n6743), .ZN(n4501) );
  OR3_X1 U6001 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4502) );
  AND2_X1 U6002 ( .A1(n8919), .A2(n9487), .ZN(n4503) );
  INV_X1 U6003 ( .A(n7514), .ZN(n4985) );
  INV_X1 U6004 ( .A(n9207), .ZN(n4638) );
  AND3_X1 U6005 ( .A1(n9211), .A2(n9233), .A3(n9080), .ZN(n4504) );
  AND2_X1 U6006 ( .A1(n6557), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4505) );
  AND2_X1 U6007 ( .A1(n4806), .A2(n4805), .ZN(n4506) );
  AND2_X1 U6008 ( .A1(n7574), .A2(n9576), .ZN(n4507) );
  AND2_X1 U6009 ( .A1(n4822), .A2(n4820), .ZN(n4508) );
  AND2_X1 U6010 ( .A1(n7964), .A2(n7963), .ZN(n7962) );
  AND2_X1 U6011 ( .A1(n8932), .A2(n7026), .ZN(n4509) );
  NAND2_X1 U6012 ( .A1(n5431), .A2(n4787), .ZN(n5054) );
  INV_X1 U6013 ( .A(n7966), .ZN(n4765) );
  AND2_X1 U6014 ( .A1(n6033), .A2(n6032), .ZN(n4510) );
  AND3_X1 U6015 ( .A1(n8165), .A2(n5422), .A3(n8166), .ZN(n4511) );
  AND2_X1 U6016 ( .A1(n4647), .A2(n9202), .ZN(n4512) );
  OR2_X1 U6017 ( .A1(n9312), .A2(n9182), .ZN(n4513) );
  NAND2_X1 U6018 ( .A1(n6068), .A2(n6067), .ZN(n9486) );
  INV_X1 U6019 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8680) );
  INV_X1 U6020 ( .A(n4897), .ZN(n9235) );
  NOR2_X1 U6021 ( .A1(n9242), .A2(n9422), .ZN(n4897) );
  NAND2_X1 U6022 ( .A1(n5778), .A2(n5780), .ZN(n8092) );
  NAND2_X1 U6023 ( .A1(n8423), .A2(n4479), .ZN(n4709) );
  XOR2_X1 U6024 ( .A(n8350), .B(n8560), .Z(n4514) );
  NOR2_X1 U6025 ( .A1(n8760), .A2(n8759), .ZN(n4515) );
  AND2_X1 U6026 ( .A1(n5121), .A2(n5103), .ZN(n4516) );
  INV_X1 U6027 ( .A(n7720), .ZN(n7979) );
  NAND2_X1 U6028 ( .A1(n5341), .A2(n5340), .ZN(n7720) );
  NAND2_X1 U6029 ( .A1(n4778), .A2(n4777), .ZN(n4517) );
  AND4_X1 U6030 ( .A1(n5053), .A2(n5052), .A3(n5051), .A4(n5050), .ZN(n6420)
         );
  OR2_X1 U6031 ( .A1(n9195), .A2(n4644), .ZN(n4643) );
  NAND2_X1 U6032 ( .A1(n8853), .A2(n8852), .ZN(n9223) );
  NAND2_X1 U6033 ( .A1(n6155), .A2(n6154), .ZN(n9480) );
  AND2_X1 U6034 ( .A1(n6248), .A2(n6247), .ZN(n4518) );
  INV_X1 U6035 ( .A(n8550), .ZN(n8678) );
  NOR2_X1 U6036 ( .A1(n9587), .A2(n9134), .ZN(n4519) );
  AND2_X1 U6037 ( .A1(n6188), .A2(n4681), .ZN(n4520) );
  NOR2_X1 U6038 ( .A1(n9437), .A2(n9286), .ZN(n4521) );
  NOR2_X1 U6039 ( .A1(n8535), .A2(n8259), .ZN(n4522) );
  OR2_X1 U6040 ( .A1(n4682), .A2(n6188), .ZN(n4523) );
  AND2_X1 U6041 ( .A1(n7998), .A2(n8542), .ZN(n4524) );
  NAND2_X1 U6042 ( .A1(n5435), .A2(n5018), .ZN(n4525) );
  AND2_X1 U6043 ( .A1(n7149), .A2(n9089), .ZN(n4526) );
  INV_X1 U6044 ( .A(n4927), .ZN(n8710) );
  NAND2_X1 U6045 ( .A1(n4922), .A2(n4925), .ZN(n4927) );
  INV_X1 U6046 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5035) );
  AND2_X1 U6047 ( .A1(n5198), .A2(SI_6_), .ZN(n4527) );
  AND2_X1 U6048 ( .A1(n4809), .A2(n4805), .ZN(n4528) );
  OR2_X1 U6049 ( .A1(n8732), .A2(n6316), .ZN(n4529) );
  NOR2_X1 U6050 ( .A1(n7989), .A2(n5006), .ZN(n5005) );
  INV_X1 U6051 ( .A(n5008), .ZN(n5007) );
  NAND2_X1 U6052 ( .A1(n5012), .A2(n5009), .ZN(n5008) );
  OR2_X1 U6053 ( .A1(n7574), .A2(n9576), .ZN(n4530) );
  INV_X1 U6054 ( .A(n5792), .ZN(n5835) );
  OAI21_X1 U6055 ( .B1(n4524), .B2(n4734), .A(n4733), .ZN(n4732) );
  INV_X1 U6056 ( .A(n4732), .ZN(n4728) );
  OR2_X1 U6057 ( .A1(n7895), .A2(n7894), .ZN(n8056) );
  AND2_X1 U6058 ( .A1(n8957), .A2(n8954), .ZN(n9063) );
  NAND2_X1 U6059 ( .A1(n9458), .A2(n9349), .ZN(n4531) );
  INV_X1 U6060 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5745) );
  INV_X1 U6061 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U6062 ( .A1(n4967), .A2(n4491), .ZN(n4532) );
  OR2_X1 U6063 ( .A1(n9426), .A2(n8856), .ZN(n9208) );
  OR2_X1 U6064 ( .A1(n9451), .A2(n9330), .ZN(n4533) );
  AND3_X1 U6065 ( .A1(n8051), .A2(n8050), .A3(n8049), .ZN(n4534) );
  AND2_X1 U6066 ( .A1(n4637), .A2(n9248), .ZN(n4535) );
  AND2_X1 U6067 ( .A1(n8025), .A2(n8024), .ZN(n4536) );
  AND2_X1 U6068 ( .A1(n8024), .A2(n8012), .ZN(n4537) );
  AND2_X1 U6069 ( .A1(n4775), .A2(n4774), .ZN(n4538) );
  OR2_X1 U6070 ( .A1(n6689), .A2(n6710), .ZN(n4539) );
  AND2_X1 U6071 ( .A1(n9208), .A2(n9023), .ZN(n9248) );
  INV_X1 U6072 ( .A(n9248), .ZN(n4560) );
  AND2_X1 U6073 ( .A1(n7957), .A2(n4721), .ZN(n4540) );
  INV_X1 U6074 ( .A(n8569), .ZN(n8364) );
  NAND2_X1 U6075 ( .A1(n5652), .A2(n5651), .ZN(n8569) );
  AND2_X1 U6076 ( .A1(n4484), .A2(n8678), .ZN(n4541) );
  AND2_X1 U6077 ( .A1(n7182), .A2(n7177), .ZN(n4542) );
  INV_X1 U6078 ( .A(n4770), .ZN(n4769) );
  NOR2_X1 U6079 ( .A1(n6481), .A2(n4771), .ZN(n4770) );
  AND2_X1 U6080 ( .A1(n4680), .A2(n4679), .ZN(n4543) );
  INV_X1 U6081 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5064) );
  INV_X1 U6082 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4632) );
  INV_X1 U6083 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4698) );
  AND2_X1 U6084 ( .A1(n4946), .A2(n4490), .ZN(n4544) );
  INV_X1 U6085 ( .A(n8059), .ZN(n4722) );
  NAND2_X1 U6086 ( .A1(n5004), .A2(n5011), .ZN(n5010) );
  AND3_X1 U6087 ( .A1(n5576), .A2(n5575), .A3(n5574), .ZN(n8123) );
  INV_X1 U6088 ( .A(n8123), .ZN(n4999) );
  NAND2_X1 U6089 ( .A1(n8111), .A2(n5379), .ZN(n8164) );
  INV_X1 U6090 ( .A(n8069), .ZN(n7937) );
  NAND2_X1 U6091 ( .A1(n7653), .A2(n4591), .ZN(n4545) );
  INV_X1 U6092 ( .A(n8099), .ZN(n6515) );
  NAND2_X1 U6093 ( .A1(n6471), .A2(n6470), .ZN(n8099) );
  AND2_X1 U6094 ( .A1(n5431), .A2(n5035), .ZN(n5435) );
  INV_X1 U6095 ( .A(n9193), .ZN(n4644) );
  INV_X1 U6096 ( .A(n9437), .ZN(n4898) );
  OR2_X1 U6097 ( .A1(n8743), .A2(n8744), .ZN(n8741) );
  AOI21_X1 U6098 ( .B1(n8386), .B2(n5718), .A(n5627), .ZN(n8157) );
  INV_X1 U6099 ( .A(n4699), .ZN(n8513) );
  NAND2_X1 U6100 ( .A1(n7717), .A2(n4484), .ZN(n4705) );
  INV_X1 U6101 ( .A(n8799), .ZN(n4681) );
  OR2_X1 U6102 ( .A1(n7655), .A2(n8875), .ZN(n4546) );
  INV_X1 U6103 ( .A(n4945), .ZN(n9461) );
  NAND2_X1 U6104 ( .A1(n4946), .A2(n4492), .ZN(n4945) );
  AND2_X1 U6105 ( .A1(n8132), .A2(n5496), .ZN(n4547) );
  INV_X1 U6106 ( .A(n7337), .ZN(n4650) );
  OAI211_X2 U6107 ( .C1(n5834), .C2(n6596), .A(n4901), .B(n4900), .ZN(n6948)
         );
  INV_X1 U6108 ( .A(n6948), .ZN(n4675) );
  NAND2_X1 U6109 ( .A1(n5767), .A2(n5771), .ZN(n9082) );
  NAND2_X1 U6110 ( .A1(n6437), .A2(n6436), .ZN(n7254) );
  INV_X1 U6111 ( .A(n9587), .ZN(n4893) );
  NAND2_X1 U6112 ( .A1(n4933), .A2(n5912), .ZN(n7134) );
  NAND2_X1 U6113 ( .A1(n4558), .A2(n5881), .ZN(n6963) );
  AND2_X1 U6114 ( .A1(n4932), .A2(n5912), .ZN(n4548) );
  OR2_X1 U6115 ( .A1(n5676), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4549) );
  AND2_X1 U6116 ( .A1(n5633), .A2(n5620), .ZN(n5631) );
  AND2_X1 U6117 ( .A1(n4829), .A2(n4824), .ZN(n4550) );
  AND2_X1 U6118 ( .A1(n5405), .A2(n5364), .ZN(n7592) );
  INV_X1 U6119 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n4667) );
  AND2_X1 U6120 ( .A1(n9140), .A2(n9400), .ZN(n4551) );
  NAND2_X1 U6121 ( .A1(n6018), .A2(n6017), .ZN(n7574) );
  INV_X1 U6122 ( .A(n7574), .ZN(n4589) );
  OR3_X1 U6123 ( .A1(n9056), .A2(n9125), .A3(n6777), .ZN(n4552) );
  OR2_X1 U6124 ( .A1(n9754), .A2(n9126), .ZN(n4553) );
  AND2_X1 U6125 ( .A1(n4798), .A2(n4799), .ZN(n4554) );
  INV_X1 U6126 ( .A(n5022), .ZN(n4797) );
  OR2_X1 U6127 ( .A1(n8332), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4555) );
  NOR2_X1 U6128 ( .A1(n5043), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8679) );
  INV_X1 U6129 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4738) );
  OAI21_X1 U6130 ( .B1(n8083), .B2(n8082), .A(n4556), .ZN(P2_U3244) );
  OAI21_X1 U6131 ( .B1(n4557), .B2(n7973), .A(n7972), .ZN(n7974) );
  OR2_X1 U6132 ( .A1(n8006), .A2(n8005), .ZN(n8013) );
  MUX2_X1 U6133 ( .A(n7926), .B(n7925), .S(n8059), .Z(n7952) );
  NAND2_X1 U6134 ( .A1(n5435), .A2(n5036), .ZN(n5056) );
  OAI21_X1 U6135 ( .B1(n4724), .B2(n4723), .A(n4540), .ZN(n4720) );
  AOI21_X1 U6136 ( .B1(n4743), .B2(n4534), .A(n4739), .ZN(n8064) );
  NOR2_X2 U6137 ( .A1(n5741), .A2(n5740), .ZN(n5744) );
  INV_X1 U6138 ( .A(n6965), .ZN(n4558) );
  NAND2_X1 U6139 ( .A1(n8816), .A2(n8819), .ZN(n6126) );
  NOR2_X2 U6140 ( .A1(n8734), .A2(n8733), .ZN(n8732) );
  OAI21_X1 U6141 ( .B1(n8113), .B2(n4817), .A(n4814), .ZN(n8178) );
  NAND2_X1 U6142 ( .A1(n4711), .A2(n5157), .ZN(n5175) );
  NAND2_X1 U6143 ( .A1(n4846), .A2(n4849), .ZN(n5219) );
  NAND2_X1 U6144 ( .A1(n5479), .A2(n5478), .ZN(n5498) );
  OR2_X1 U6145 ( .A1(n9019), .A2(n4560), .ZN(n9011) );
  NAND2_X1 U6146 ( .A1(n5114), .A2(n5113), .ZN(n5130) );
  NAND2_X1 U6147 ( .A1(n4626), .A2(n4624), .ZN(P1_U3240) );
  NAND2_X1 U6148 ( .A1(n5520), .A2(n5519), .ZN(n5522) );
  NAND2_X1 U6149 ( .A1(n5260), .A2(n5020), .ZN(n5262) );
  AOI21_X1 U6150 ( .B1(n9029), .B2(n9111), .A(n4615), .ZN(n4614) );
  NAND2_X1 U6151 ( .A1(n4869), .A2(n5594), .ZN(n5617) );
  NAND2_X1 U6152 ( .A1(n9038), .A2(n4613), .ZN(n9043) );
  XNOR2_X1 U6153 ( .A(n5092), .B(n5069), .ZN(n5091) );
  INV_X1 U6154 ( .A(n4715), .ZN(n4714) );
  NAND2_X1 U6155 ( .A1(n4714), .A2(n4713), .ZN(n8037) );
  OAI21_X1 U6156 ( .B1(n8032), .B2(n4718), .A(n4536), .ZN(n4717) );
  NOR2_X1 U6157 ( .A1(n7956), .A2(n7955), .ZN(n4724) );
  OAI21_X1 U6158 ( .B1(n8044), .B2(n4745), .A(n4744), .ZN(n4743) );
  NOR2_X1 U6159 ( .A1(n7386), .A2(n6544), .ZN(n7683) );
  NAND2_X1 U6160 ( .A1(n4796), .A2(n4794), .ZN(n9810) );
  INV_X1 U6161 ( .A(n6867), .ZN(n5121) );
  AND2_X4 U6162 ( .A1(n8070), .A2(n7900), .ZN(n5665) );
  NAND2_X1 U6163 ( .A1(n8543), .A2(n7999), .ZN(n4569) );
  NAND2_X1 U6164 ( .A1(n7750), .A2(n4770), .ZN(n4570) );
  NAND2_X1 U6165 ( .A1(n8449), .A2(n8450), .ZN(n8433) );
  NAND2_X1 U6166 ( .A1(n4572), .A2(n4571), .ZN(n8449) );
  NAND3_X1 U6167 ( .A1(n4782), .A2(n8507), .A3(n4537), .ZN(n4571) );
  INV_X1 U6168 ( .A(n4779), .ZN(n4573) );
  NAND3_X1 U6169 ( .A1(n8507), .A2(n4782), .A3(n8012), .ZN(n4574) );
  NAND3_X1 U6170 ( .A1(n4858), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4853) );
  INV_X2 U6171 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4858) );
  NAND3_X1 U6172 ( .A1(n7908), .A2(n7225), .A3(n7224), .ZN(n4754) );
  NAND3_X1 U6173 ( .A1(n9632), .A2(n9626), .A3(n6578), .ZN(n4900) );
  INV_X1 U6174 ( .A(n4845), .ZN(n4583) );
  NAND2_X1 U6175 ( .A1(n5744), .A2(n5743), .ZN(n5773) );
  NAND3_X1 U6176 ( .A1(n5744), .A2(n4632), .A3(n5743), .ZN(n4584) );
  NAND2_X1 U6177 ( .A1(n4897), .A2(n4585), .ZN(n4588) );
  NAND2_X1 U6178 ( .A1(n4897), .A2(n9415), .ZN(n9219) );
  INV_X1 U6179 ( .A(n4595), .ZN(n4899) );
  NAND2_X1 U6180 ( .A1(n8890), .A2(n4606), .ZN(n4608) );
  OAI21_X2 U6181 ( .B1(n6904), .B2(n4609), .A(n4607), .ZN(n7151) );
  NAND3_X1 U6182 ( .A1(n9033), .A2(n9111), .A3(n9234), .ZN(n4617) );
  INV_X1 U6183 ( .A(n6872), .ZN(n6890) );
  CLKBUF_X1 U6184 ( .A(n6872), .Z(n4618) );
  NAND4_X1 U6185 ( .A1(n9121), .A2(n9120), .A3(n9122), .A4(n9119), .ZN(n4630)
         );
  NOR2_X4 U6186 ( .A1(n5773), .A2(n4631), .ZN(n5763) );
  OAI21_X1 U6187 ( .B1(n9275), .B2(n9106), .A(n4637), .ZN(n9249) );
  NAND2_X1 U6188 ( .A1(n9275), .A2(n4535), .ZN(n4636) );
  NAND2_X1 U6189 ( .A1(n9275), .A2(n9205), .ZN(n9262) );
  OAI21_X1 U6190 ( .B1(n7181), .B2(n9061), .A(n8940), .ZN(n7183) );
  NAND2_X1 U6191 ( .A1(n7336), .A2(n4654), .ZN(n4651) );
  NAND3_X1 U6192 ( .A1(n4652), .A2(n4651), .A3(n4649), .ZN(n7591) );
  NAND2_X1 U6193 ( .A1(n7590), .A2(n4657), .ZN(n8276) );
  NOR2_X1 U6194 ( .A1(n7591), .A2(n7870), .ZN(n8278) );
  MUX2_X1 U6195 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6683), .S(n9546), .Z(n9541)
         );
  OAI21_X1 U6196 ( .B1(n8734), .B2(n4691), .A(n4690), .ZN(n6403) );
  NAND3_X1 U6197 ( .A1(n8699), .A2(n6123), .A3(n6116), .ZN(n8816) );
  NOR2_X2 U6198 ( .A1(n5676), .A2(n4987), .ZN(n5061) );
  NOR2_X2 U6199 ( .A1(n8500), .A2(n8487), .ZN(n8486) );
  INV_X1 U6200 ( .A(n4705), .ZN(n8548) );
  INV_X1 U6201 ( .A(n4709), .ZN(n8376) );
  NAND2_X1 U6202 ( .A1(n4710), .A2(n4856), .ZN(n4855) );
  NAND2_X1 U6203 ( .A1(n5155), .A2(n5154), .ZN(n4711) );
  NAND2_X1 U6204 ( .A1(n5130), .A2(n5129), .ZN(n4712) );
  AOI21_X1 U6205 ( .B1(n4717), .B2(n8033), .A(n4716), .ZN(n4715) );
  NAND3_X1 U6206 ( .A1(n4719), .A2(n7965), .A3(n7969), .ZN(n7970) );
  NAND3_X1 U6207 ( .A1(n4720), .A2(n7961), .A3(n7962), .ZN(n4719) );
  NAND2_X1 U6208 ( .A1(n4725), .A2(n4730), .ZN(n8006) );
  NAND3_X1 U6209 ( .A1(n7988), .A2(n4728), .A3(n4729), .ZN(n4725) );
  NAND2_X1 U6210 ( .A1(n6582), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4737) );
  MUX2_X1 U6211 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6582), .Z(n5131) );
  MUX2_X1 U6212 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n6582), .Z(n5156) );
  MUX2_X1 U6213 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6582), .Z(n5176) );
  MUX2_X1 U6214 ( .A(n6600), .B(n6602), .S(n6582), .Z(n5197) );
  MUX2_X1 U6215 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6582), .Z(n5220) );
  MUX2_X1 U6216 ( .A(n6607), .B(n6609), .S(n6582), .Z(n5224) );
  MUX2_X1 U6217 ( .A(n5244), .B(n6646), .S(n6582), .Z(n5246) );
  MUX2_X1 U6218 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n6582), .Z(n5306) );
  MUX2_X1 U6219 ( .A(n6788), .B(n6786), .S(n6582), .Z(n5310) );
  MUX2_X1 U6220 ( .A(n5263), .B(n6671), .S(n6582), .Z(n5265) );
  MUX2_X1 U6221 ( .A(n10321), .B(n6833), .S(n6582), .Z(n5336) );
  INV_X1 U6222 ( .A(n7301), .ZN(n7283) );
  AND2_X1 U6223 ( .A1(n5158), .A2(n4539), .ZN(n4747) );
  OR2_X1 U6224 ( .A1(n6589), .A2(n5249), .ZN(n4748) );
  XNOR2_X2 U6225 ( .A(n4749), .B(n5064), .ZN(n6496) );
  OAI22_X1 U6226 ( .A1(n5199), .A2(n6597), .B1(n6689), .B2(n9546), .ZN(n4751)
         );
  INV_X1 U6227 ( .A(n7959), .ZN(n4755) );
  NAND2_X1 U6228 ( .A1(n7469), .A2(n4763), .ZN(n4760) );
  NAND2_X1 U6229 ( .A1(n4760), .A2(n4761), .ZN(n7708) );
  NAND2_X1 U6230 ( .A1(n6489), .A2(n4538), .ZN(n4773) );
  INV_X1 U6231 ( .A(n4778), .ZN(n8372) );
  INV_X1 U6232 ( .A(n5039), .ZN(n4790) );
  NAND2_X1 U6233 ( .A1(n4791), .A2(n5732), .ZN(P2_U3222) );
  OAI211_X1 U6234 ( .C1(n5712), .C2(n5706), .A(n4793), .B(n4792), .ZN(n4791)
         );
  NAND2_X1 U6235 ( .A1(n5712), .A2(n5711), .ZN(n4793) );
  NAND2_X1 U6236 ( .A1(n6854), .A2(n4516), .ZN(n4796) );
  NAND2_X1 U6237 ( .A1(n5071), .A2(n5070), .ZN(n4799) );
  NAND3_X1 U6238 ( .A1(n4798), .A2(n8085), .A3(n4799), .ZN(n8084) );
  NAND2_X1 U6239 ( .A1(n8084), .A2(n4799), .ZN(n6855) );
  NAND2_X1 U6240 ( .A1(n7493), .A2(n4506), .ZN(n4804) );
  AOI21_X1 U6241 ( .B1(n4528), .B2(n4806), .A(n4485), .ZN(n4803) );
  NAND2_X1 U6242 ( .A1(n7167), .A2(n4824), .ZN(n4821) );
  NAND2_X1 U6243 ( .A1(n7785), .A2(n4834), .ZN(n4831) );
  NAND2_X1 U6244 ( .A1(n4831), .A2(n4832), .ZN(n4837) );
  OAI21_X2 U6245 ( .B1(n9569), .B2(n8963), .A(n8877), .ZN(n7575) );
  XNOR2_X2 U6246 ( .A(n6948), .B(n6872), .ZN(n9053) );
  NAND2_X1 U6247 ( .A1(n4843), .A2(n5768), .ZN(n5750) );
  NAND2_X1 U6248 ( .A1(n5175), .A2(n5174), .ZN(n4852) );
  NAND2_X1 U6249 ( .A1(n5175), .A2(n4847), .ZN(n4846) );
  NAND2_X1 U6250 ( .A1(n5596), .A2(n4862), .ZN(n4861) );
  NAND3_X1 U6251 ( .A1(n5631), .A2(n4863), .A3(n5595), .ZN(n4860) );
  OR2_X1 U6252 ( .A1(n5596), .A2(n5595), .ZN(n4869) );
  NAND2_X1 U6253 ( .A1(n5358), .A2(n4873), .ZN(n4870) );
  NAND2_X1 U6254 ( .A1(n4870), .A2(n4871), .ZN(n5429) );
  NAND2_X1 U6255 ( .A1(n5358), .A2(n5357), .ZN(n5384) );
  XNOR2_X1 U6256 ( .A(n4892), .B(n7889), .ZN(n8833) );
  OAI21_X1 U6257 ( .B1(n7882), .B2(n10098), .A(n7887), .ZN(n4892) );
  NAND2_X1 U6258 ( .A1(n4474), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4901) );
  MUX2_X1 U6259 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4903), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n4902) );
  NAND2_X1 U6260 ( .A1(n8769), .A2(n4912), .ZN(n4909) );
  NAND2_X1 U6261 ( .A1(n4909), .A2(n4910), .ZN(n6264) );
  NAND2_X1 U6262 ( .A1(n4916), .A2(n4917), .ZN(n6168) );
  NAND2_X1 U6263 ( .A1(n8743), .A2(n6147), .ZN(n4916) );
  NAND2_X1 U6264 ( .A1(n6270), .A2(n4497), .ZN(n4919) );
  NAND2_X1 U6265 ( .A1(n4919), .A2(n4920), .ZN(n8734) );
  NAND2_X1 U6266 ( .A1(n4929), .A2(n7724), .ZN(n6117) );
  NAND2_X1 U6267 ( .A1(n5908), .A2(n5911), .ZN(n4933) );
  NAND2_X1 U6268 ( .A1(n5763), .A2(n4934), .ZN(n4936) );
  AND2_X1 U6269 ( .A1(n5763), .A2(n5753), .ZN(n6355) );
  NAND3_X1 U6270 ( .A1(n5977), .A2(n7429), .A3(n7444), .ZN(n7443) );
  NAND2_X1 U6271 ( .A1(n4938), .A2(n4939), .ZN(n4937) );
  NAND2_X1 U6272 ( .A1(n7455), .A2(n4949), .ZN(n4948) );
  AND2_X1 U6273 ( .A1(n4951), .A2(n4530), .ZN(n4949) );
  NAND2_X1 U6274 ( .A1(n7178), .A2(n4542), .ZN(n7394) );
  NAND2_X1 U6275 ( .A1(n9185), .A2(n4960), .ZN(n4958) );
  NAND2_X1 U6276 ( .A1(n4958), .A2(n4959), .ZN(n9255) );
  NOR2_X1 U6277 ( .A1(n7144), .A2(n4970), .ZN(n4969) );
  NAND3_X1 U6278 ( .A1(n6874), .A2(n6936), .A3(n6873), .ZN(n6900) );
  OR2_X2 U6279 ( .A1(n9386), .A2(n9385), .ZN(n9474) );
  OAI22_X2 U6280 ( .A1(n7780), .A2(n7779), .B1(n8874), .B2(n9614), .ZN(n7849)
         );
  NAND2_X1 U6281 ( .A1(n5763), .A2(n4971), .ZN(n5778) );
  OR2_X1 U6282 ( .A1(n9949), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4980) );
  INV_X1 U6283 ( .A(n6461), .ZN(n4982) );
  NAND2_X1 U6284 ( .A1(n4983), .A2(n4984), .ZN(n6446) );
  NAND2_X1 U6285 ( .A1(n7465), .A2(n6444), .ZN(n4983) );
  AOI21_X1 U6286 ( .B1(n7470), .B2(n6444), .A(n4985), .ZN(n4984) );
  NAND3_X1 U6287 ( .A1(n5040), .A2(n4698), .A3(n5064), .ZN(n4987) );
  INV_X1 U6288 ( .A(n4988), .ZN(n6458) );
  AND3_X2 U6289 ( .A1(n5034), .A2(n5151), .A3(n5000), .ZN(n5431) );
  NAND4_X1 U6290 ( .A1(n5034), .A2(n5151), .A3(n5033), .A4(n5032), .ZN(n5393)
         );
  OAI21_X1 U6291 ( .B1(n5003), .B2(n7540), .A(n5002), .ZN(n7820) );
  NAND2_X1 U6292 ( .A1(n8539), .A2(n4477), .ZN(n5013) );
  NAND2_X1 U6293 ( .A1(n5013), .A2(n5014), .ZN(n8512) );
  INV_X1 U6294 ( .A(n5016), .ZN(n8541) );
  OAI21_X1 U6295 ( .B1(n7905), .B2(n7058), .A(n7938), .ZN(n7094) );
  NAND2_X1 U6296 ( .A1(n6463), .A2(n6462), .ZN(n6468) );
  AOI22_X1 U6297 ( .A1(n5808), .A2(n9141), .B1(n6397), .B2(n8793), .ZN(n5841)
         );
  NOR2_X2 U6298 ( .A1(n7355), .A2(n7421), .ZN(n7374) );
  NAND4_X1 U6299 ( .A1(n5078), .A2(n5077), .A3(n5076), .A4(n5075), .ZN(n6475)
         );
  NAND2_X1 U6300 ( .A1(n8274), .A2(n7901), .ZN(n5071) );
  NAND2_X2 U6301 ( .A1(n6460), .A2(n6459), .ZN(n8355) );
  NAND2_X1 U6302 ( .A1(n5976), .A2(n5975), .ZN(n7429) );
  INV_X1 U6303 ( .A(n6264), .ZN(n6267) );
  XNOR2_X1 U6304 ( .A(n5632), .B(n5631), .ZN(n7817) );
  INV_X1 U6305 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10234) );
  INV_X1 U6306 ( .A(n5973), .ZN(n5976) );
  OR2_X1 U6307 ( .A1(n5797), .A2(n6519), .ZN(n6548) );
  NAND2_X1 U6308 ( .A1(n5797), .A2(n6358), .ZN(n9754) );
  INV_X1 U6309 ( .A(n5797), .ZN(n5798) );
  NAND2_X1 U6310 ( .A1(n5893), .A2(n6469), .ZN(n5834) );
  XNOR2_X1 U6311 ( .A(n7882), .B(SI_30_), .ZN(n8841) );
  OAI21_X1 U6312 ( .B1(n7344), .B2(n6439), .A(n7964), .ZN(n7366) );
  NAND2_X1 U6313 ( .A1(n5566), .A2(n5565), .ZN(n5568) );
  XNOR2_X1 U6314 ( .A(n5617), .B(n5616), .ZN(n7813) );
  NAND2_X1 U6315 ( .A1(n8126), .A2(n5585), .ZN(n5591) );
  NAND2_X1 U6316 ( .A1(n5782), .A2(n5784), .ZN(n5854) );
  OAI21_X1 U6317 ( .B1(n9255), .B2(n9189), .A(n9188), .ZN(n9241) );
  NAND2_X1 U6318 ( .A1(n5047), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5085) );
  INV_X1 U6319 ( .A(n8689), .ZN(n5048) );
  NAND2_X1 U6320 ( .A1(n6420), .A2(n7054), .ZN(n7934) );
  AOI22_X1 U6321 ( .A1(n8448), .A2(n6485), .B1(n8147), .B2(n8458), .ZN(n8432)
         );
  NAND2_X2 U6322 ( .A1(n7035), .A2(n9743), .ZN(n9751) );
  AND2_X1 U6323 ( .A1(n5120), .A2(n5119), .ZN(n5022) );
  INV_X1 U6324 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10293) );
  NAND2_X2 U6325 ( .A1(n7042), .A2(n9845), .ZN(n8553) );
  INV_X1 U6326 ( .A(n8634), .ZN(n6508) );
  AND2_X1 U6327 ( .A1(n6492), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5024) );
  AND4_X1 U6328 ( .A1(n5530), .A2(n5529), .A3(n5528), .A4(n5527), .ZN(n8207)
         );
  AND4_X1 U6329 ( .A1(n5753), .A2(n5747), .A3(n5746), .A4(n10072), .ZN(n5025)
         );
  NOR2_X1 U6330 ( .A1(n8189), .A2(n8188), .ZN(n5026) );
  INV_X1 U6331 ( .A(n8577), .ZN(n6456) );
  INV_X1 U6332 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5746) );
  INV_X1 U6333 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5036) );
  NOR2_X1 U6334 ( .A1(n5848), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5743) );
  INV_X1 U6335 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5038) );
  INV_X1 U6336 ( .A(n6188), .ZN(n6189) );
  INV_X1 U6337 ( .A(n7081), .ZN(n5911) );
  INV_X1 U6338 ( .A(n6175), .ZN(n5783) );
  INV_X1 U6339 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5263) );
  INV_X1 U6340 ( .A(n5071), .ZN(n5073) );
  INV_X1 U6341 ( .A(n5581), .ZN(n5572) );
  OR2_X1 U6342 ( .A1(n5579), .A2(n5571), .ZN(n5581) );
  INV_X1 U6343 ( .A(n5413), .ZN(n5397) );
  OAI22_X1 U6344 ( .A1(n5809), .A2(n6945), .B1(n5797), .B2(n10275), .ZN(n5810)
         );
  AND2_X1 U6345 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(n5783), .ZN(n6174) );
  AND2_X1 U6346 ( .A1(n6174), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6196) );
  INV_X1 U6347 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6069) );
  INV_X1 U6348 ( .A(SI_20_), .ZN(n10306) );
  INV_X1 U6349 ( .A(SI_16_), .ZN(n10323) );
  INV_X1 U6350 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6036) );
  INV_X1 U6351 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5742) );
  INV_X1 U6352 ( .A(n5293), .ZN(n5291) );
  OR2_X1 U6353 ( .A1(n5525), .A2(n10176), .ZN(n5579) );
  NAND2_X1 U6354 ( .A1(n6456), .A2(n8157), .ZN(n6457) );
  NAND2_X1 U6355 ( .A1(n8604), .A2(n8255), .ZN(n6454) );
  NAND2_X1 U6356 ( .A1(n5461), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6357 ( .A1(n5368), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5411) );
  INV_X1 U6358 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U6359 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n6301), .ZN(n6368) );
  INV_X1 U6360 ( .A(n6300), .ZN(n6301) );
  OR2_X1 U6361 ( .A1(n6049), .A2(n6048), .ZN(n6070) );
  AND2_X1 U6362 ( .A1(n6003), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U6363 ( .A1(n9042), .A2(n9156), .ZN(n9030) );
  OR2_X1 U6364 ( .A1(n6889), .A2(n6378), .ZN(n6779) );
  NAND2_X1 U6365 ( .A1(n5476), .A2(n5475), .ZN(n5479) );
  INV_X1 U6366 ( .A(n5380), .ZN(n5383) );
  NAND2_X1 U6367 ( .A1(n5310), .A2(n10159), .ZN(n5335) );
  INV_X1 U6368 ( .A(n6475), .ZN(n7047) );
  AND2_X1 U6369 ( .A1(n8072), .A2(n8530), .ZN(n5725) );
  AND2_X1 U6370 ( .A1(n5656), .A2(n5624), .ZN(n8386) );
  NAND2_X1 U6371 ( .A1(n5047), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5051) );
  INV_X1 U6372 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10112) );
  INV_X1 U6373 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7205) );
  INV_X1 U6374 ( .A(n8590), .ZN(n8428) );
  AND2_X1 U6375 ( .A1(n7990), .A2(n6447), .ZN(n7977) );
  AND2_X1 U6376 ( .A1(n7983), .A2(n7982), .ZN(n7913) );
  INV_X1 U6377 ( .A(n8218), .ZN(n9814) );
  AND2_X1 U6378 ( .A1(n5689), .A2(n9857), .ZN(n6504) );
  NOR2_X1 U6379 ( .A1(n6254), .A2(n8782), .ZN(n6253) );
  NAND2_X1 U6380 ( .A1(n6156), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6175) );
  INV_X1 U6381 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7446) );
  NOR2_X1 U6382 ( .A1(n9447), .A2(n9316), .ZN(n9184) );
  AND2_X1 U6383 ( .A1(n9464), .A2(n8865), .ZN(n9199) );
  AND2_X1 U6384 ( .A1(n9050), .A2(n9363), .ZN(n9385) );
  AND2_X1 U6385 ( .A1(n8948), .A2(n8973), .ZN(n9072) );
  AND2_X1 U6386 ( .A1(n4672), .A2(n9745), .ZN(n6378) );
  INV_X1 U6387 ( .A(n9171), .ZN(n8989) );
  INV_X1 U6388 ( .A(n9065), .ZN(n9568) );
  INV_X1 U6389 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5765) );
  INV_X1 U6390 ( .A(SI_7_), .ZN(n10175) );
  OAI21_X1 U6391 ( .B1(n8357), .B2(n8233), .A(n5730), .ZN(n5731) );
  INV_X1 U6392 ( .A(n8233), .ZN(n9817) );
  NOR2_X1 U6393 ( .A1(n6504), .A2(n5703), .ZN(n5722) );
  INV_X1 U6394 ( .A(n5658), .ZN(n5718) );
  AND4_X1 U6395 ( .A1(n5444), .A2(n5443), .A3(n5442), .A4(n5441), .ZN(n8217)
         );
  INV_X1 U6396 ( .A(n9827), .ZN(n9554) );
  AND2_X1 U6397 ( .A1(n6691), .A2(n6690), .ZN(n9827) );
  INV_X1 U6398 ( .A(n9847), .ZN(n8556) );
  INV_X1 U6399 ( .A(n9946), .ZN(n9898) );
  NAND2_X1 U6400 ( .A1(n8547), .A2(n9921), .ZN(n9946) );
  NOR2_X1 U6401 ( .A1(n6504), .A2(n8078), .ZN(n7011) );
  NAND2_X1 U6402 ( .A1(n6681), .A2(n5700), .ZN(n9856) );
  INV_X1 U6403 ( .A(n8810), .ZN(n8822) );
  INV_X1 U6404 ( .A(n8831), .ZN(n8808) );
  OR2_X1 U6405 ( .A1(n8840), .A2(n6302), .ZN(n6303) );
  INV_X1 U6406 ( .A(n9724), .ZN(n9705) );
  INV_X1 U6407 ( .A(n9718), .ZN(n9690) );
  AND2_X1 U6408 ( .A1(n6570), .A2(n9162), .ZN(n9718) );
  AND2_X1 U6409 ( .A1(n6888), .A2(n6887), .ZN(n9735) );
  AND2_X1 U6410 ( .A1(n6775), .A2(n6772), .ZN(n6781) );
  OR2_X1 U6411 ( .A1(n6882), .A2(n6378), .ZN(n9791) );
  NOR2_X1 U6412 ( .A1(n6775), .A2(n6774), .ZN(n6878) );
  AND3_X1 U6413 ( .A1(n6335), .A2(n6340), .A3(n6339), .ZN(n9755) );
  AND2_X1 U6414 ( .A1(n6085), .A2(n6101), .ZN(n7389) );
  NAND2_X1 U6415 ( .A1(n6665), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9892) );
  INV_X1 U6416 ( .A(n5731), .ZN(n5732) );
  NAND2_X1 U6417 ( .A1(n5729), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9824) );
  AND4_X1 U6418 ( .A1(n5418), .A2(n5417), .A3(n5416), .A4(n5415), .ZN(n8170)
         );
  INV_X2 U6419 ( .A(P2_U3966), .ZN(n8275) );
  OR2_X1 U6420 ( .A1(n8541), .A2(n8540), .ZN(n8628) );
  INV_X1 U6421 ( .A(n8553), .ZN(n9849) );
  INV_X1 U6422 ( .A(n8553), .ZN(n9855) );
  OR2_X1 U6423 ( .A1(n9855), .A2(n7012), .ZN(n8506) );
  NAND2_X1 U6424 ( .A1(n9960), .A2(n9918), .ZN(n8634) );
  AND2_X2 U6425 ( .A1(n7011), .A2(n6506), .ZN(n9960) );
  INV_X1 U6426 ( .A(n8410), .ZN(n8653) );
  INV_X1 U6427 ( .A(n8535), .ZN(n8673) );
  NAND2_X1 U6428 ( .A1(n9949), .A2(n9918), .ZN(n8677) );
  INV_X1 U6429 ( .A(n9949), .ZN(n9948) );
  NOR2_X1 U6430 ( .A1(n9857), .A2(n9856), .ZN(n9872) );
  CLKBUF_X1 U6431 ( .A(n9872), .Z(n9893) );
  INV_X1 U6432 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7604) );
  INV_X1 U6433 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6984) );
  INV_X1 U6434 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6609) );
  INV_X1 U6435 ( .A(n8875), .ZN(n9614) );
  OR2_X1 U6436 ( .A1(n6403), .A2(n6401), .ZN(n6419) );
  OR2_X1 U6437 ( .A1(n6362), .A2(n6377), .ZN(n8831) );
  NAND4_X1 U6438 ( .A1(n6306), .A2(n6305), .A3(n6304), .A4(n6303), .ZN(n9277)
         );
  INV_X1 U6439 ( .A(n9730), .ZN(n9717) );
  NAND2_X1 U6440 ( .A1(n9751), .A2(n9735), .ZN(n9408) );
  INV_X1 U6441 ( .A(n9592), .ZN(n7661) );
  INV_X1 U6442 ( .A(n9809), .ZN(n9806) );
  OR2_X1 U6443 ( .A1(n9493), .A2(n9492), .ZN(n9509) );
  INV_X1 U6444 ( .A(n9800), .ZN(n9799) );
  OR2_X1 U6445 ( .A1(n9755), .A2(n9754), .ZN(n9757) );
  INV_X1 U6446 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10244) );
  INV_X1 U6447 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10107) );
  INV_X1 U6448 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6788) );
  OR2_X1 U6449 ( .A1(n5917), .A2(n5916), .ZN(n6623) );
  NOR2_X2 U6450 ( .A1(n6681), .A2(n9892), .ZN(P2_U3966) );
  NOR2_X2 U6451 ( .A1(n6548), .A2(P1_U3084), .ZN(P1_U4006) );
  NOR2_X1 U6452 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5030) );
  AND2_X2 U6453 ( .A1(n5088), .A2(n5031), .ZN(n5151) );
  NAND2_X1 U6454 ( .A1(n5043), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5042) );
  INV_X1 U6455 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5041) );
  INV_X1 U6456 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5044) );
  XNOR2_X2 U6457 ( .A(n5045), .B(n5044), .ZN(n5046) );
  NAND2_X1 U6458 ( .A1(n5161), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5053) );
  INV_X1 U6459 ( .A(n5046), .ZN(n5049) );
  INV_X1 U6460 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7049) );
  OR2_X1 U6461 ( .A1(n5162), .A2(n7049), .ZN(n5052) );
  NAND2_X2 U6462 ( .A1(n5046), .A2(n5048), .ZN(n5167) );
  INV_X1 U6463 ( .A(n5167), .ZN(n5047) );
  INV_X1 U6464 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10120) );
  OR2_X1 U6465 ( .A1(n5163), .A2(n10120), .ZN(n5050) );
  NAND2_X1 U6466 ( .A1(n5054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5680) );
  XNOR2_X1 U6467 ( .A(n5680), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8079) );
  OR2_X4 U6468 ( .A1(n9897), .A2(n6472), .ZN(n9942) );
  INV_X2 U6469 ( .A(n7901), .ZN(n7018) );
  XNOR2_X2 U6470 ( .A(n5063), .B(n5062), .ZN(n5713) );
  NAND2_X4 U6471 ( .A1(n5713), .A2(n6496), .ZN(n6689) );
  INV_X1 U6472 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5065) );
  INV_X1 U6473 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6597) );
  AND2_X1 U6474 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U6475 ( .A1(n5066), .A2(n5067), .ZN(n5795) );
  AND2_X1 U6476 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U6477 ( .A1(n4475), .A2(n5068), .ZN(n5081) );
  INV_X1 U6478 ( .A(SI_1_), .ZN(n5069) );
  MUX2_X1 U6479 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5066), .Z(n5090) );
  XNOR2_X1 U6480 ( .A(n5091), .B(n5090), .ZN(n6596) );
  NAND2_X1 U6481 ( .A1(n6472), .A2(n8069), .ZN(n7900) );
  XNOR2_X1 U6482 ( .A(n7054), .B(n5665), .ZN(n5072) );
  INV_X1 U6483 ( .A(n5072), .ZN(n5070) );
  NAND2_X1 U6484 ( .A1(n6491), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5078) );
  INV_X1 U6485 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9826) );
  OR2_X1 U6486 ( .A1(n5167), .A2(n9826), .ZN(n5077) );
  INV_X1 U6487 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5074) );
  OR2_X1 U6488 ( .A1(n5145), .A2(n5074), .ZN(n5076) );
  INV_X1 U6489 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10273) );
  OR2_X1 U6490 ( .A1(n5163), .A2(n10273), .ZN(n5075) );
  NAND2_X1 U6491 ( .A1(n6582), .A2(SI_0_), .ZN(n5080) );
  INV_X1 U6492 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6493 ( .A1(n5080), .A2(n5079), .ZN(n5082) );
  AND2_X1 U6494 ( .A1(n5082), .A2(n5081), .ZN(n8698) );
  MUX2_X1 U6495 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8698), .S(n6689), .Z(n7053) );
  NAND2_X1 U6496 ( .A1(n6475), .A2(n7053), .ZN(n6421) );
  INV_X1 U6497 ( .A(n6421), .ZN(n7041) );
  NOR2_X1 U6498 ( .A1(n7053), .A2(n5665), .ZN(n5083) );
  AOI21_X1 U6499 ( .B1(n7041), .B2(n7901), .A(n5083), .ZN(n8085) );
  NAND2_X1 U6500 ( .A1(n5161), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5087) );
  INV_X1 U6501 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7061) );
  OR2_X1 U6502 ( .A1(n5162), .A2(n7061), .ZN(n5086) );
  INV_X1 U6503 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10319) );
  OR2_X1 U6504 ( .A1(n5163), .A2(n10319), .ZN(n5084) );
  NOR2_X1 U6505 ( .A1(n7046), .A2(n7018), .ZN(n5098) );
  OR2_X1 U6506 ( .A1(n5088), .A2(n8680), .ZN(n5089) );
  XNOR2_X1 U6507 ( .A(n5089), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9559) );
  INV_X1 U6508 ( .A(n9559), .ZN(n6593) );
  INV_X1 U6509 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U6510 ( .A1(n5091), .A2(n5090), .ZN(n5094) );
  NAND2_X1 U6511 ( .A1(n5092), .A2(SI_1_), .ZN(n5093) );
  NAND2_X1 U6512 ( .A1(n5094), .A2(n5093), .ZN(n5111) );
  INV_X1 U6513 ( .A(SI_2_), .ZN(n5095) );
  XNOR2_X1 U6514 ( .A(n5112), .B(n5095), .ZN(n5110) );
  XNOR2_X1 U6515 ( .A(n5111), .B(n5110), .ZN(n6594) );
  XNOR2_X1 U6516 ( .A(n7057), .B(n5665), .ZN(n5099) );
  NAND2_X1 U6517 ( .A1(n5098), .A2(n5099), .ZN(n5102) );
  INV_X1 U6518 ( .A(n5098), .ZN(n5101) );
  INV_X1 U6519 ( .A(n5099), .ZN(n5100) );
  NAND2_X1 U6520 ( .A1(n5101), .A2(n5100), .ZN(n5103) );
  AND2_X1 U6521 ( .A1(n5102), .A2(n5103), .ZN(n6856) );
  NAND2_X1 U6522 ( .A1(n6855), .A2(n6856), .ZN(n6854) );
  NAND2_X1 U6523 ( .A1(n5161), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5108) );
  OR2_X1 U6524 ( .A1(n5163), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5107) );
  INV_X1 U6525 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6698) );
  OR2_X1 U6526 ( .A1(n5162), .A2(n6698), .ZN(n5106) );
  INV_X1 U6527 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5104) );
  OR2_X1 U6528 ( .A1(n9813), .A2(n7018), .ZN(n5117) );
  NAND2_X1 U6529 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4502), .ZN(n5109) );
  XNOR2_X1 U6530 ( .A(n5109), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6697) );
  INV_X1 U6531 ( .A(n6697), .ZN(n6721) );
  INV_X1 U6532 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6584) );
  OR2_X1 U6533 ( .A1(n5199), .A2(n6584), .ZN(n5116) );
  NAND2_X1 U6534 ( .A1(n5111), .A2(n5110), .ZN(n5114) );
  NAND2_X1 U6535 ( .A1(n5112), .A2(SI_2_), .ZN(n5113) );
  INV_X1 U6536 ( .A(SI_3_), .ZN(n10324) );
  XNOR2_X1 U6537 ( .A(n5131), .B(n10324), .ZN(n5129) );
  XNOR2_X1 U6538 ( .A(n5130), .B(n5129), .ZN(n6583) );
  XNOR2_X1 U6539 ( .A(n9917), .B(n5639), .ZN(n5118) );
  XNOR2_X1 U6540 ( .A(n5117), .B(n5118), .ZN(n6867) );
  INV_X1 U6541 ( .A(n5117), .ZN(n5120) );
  INV_X1 U6542 ( .A(n5118), .ZN(n5119) );
  INV_X1 U6543 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5122) );
  OR2_X1 U6544 ( .A1(n5145), .A2(n5122), .ZN(n5127) );
  XNOR2_X1 U6545 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9846) );
  OR2_X1 U6546 ( .A1(n5163), .A2(n9846), .ZN(n5124) );
  INV_X1 U6547 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6696) );
  OR2_X1 U6548 ( .A1(n5162), .A2(n6696), .ZN(n5123) );
  NOR2_X1 U6549 ( .A1(n5024), .A2(n5125), .ZN(n5126) );
  NOR2_X1 U6550 ( .A1(n7168), .A2(n7018), .ZN(n5135) );
  OR2_X1 U6551 ( .A1(n5151), .A2(n8680), .ZN(n5128) );
  XNOR2_X1 U6552 ( .A(n5128), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6695) );
  INV_X1 U6553 ( .A(n6695), .ZN(n6769) );
  NAND2_X1 U6554 ( .A1(n5131), .A2(SI_3_), .ZN(n5132) );
  INV_X1 U6555 ( .A(SI_4_), .ZN(n10307) );
  XNOR2_X1 U6556 ( .A(n5156), .B(n10307), .ZN(n5154) );
  XNOR2_X1 U6557 ( .A(n5155), .B(n5154), .ZN(n6591) );
  OR2_X1 U6558 ( .A1(n5249), .A2(n6591), .ZN(n5134) );
  INV_X1 U6559 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6592) );
  OR2_X1 U6560 ( .A1(n4476), .A2(n6592), .ZN(n5133) );
  OAI211_X1 U6561 ( .C1(n6689), .C2(n6769), .A(n5134), .B(n5133), .ZN(n6430)
         );
  XNOR2_X1 U6562 ( .A(n6430), .B(n5665), .ZN(n5136) );
  NAND2_X1 U6563 ( .A1(n5135), .A2(n5136), .ZN(n5139) );
  INV_X1 U6564 ( .A(n5135), .ZN(n5138) );
  INV_X1 U6565 ( .A(n5136), .ZN(n5137) );
  NAND2_X1 U6566 ( .A1(n5138), .A2(n5137), .ZN(n5140) );
  AND2_X1 U6567 ( .A1(n5139), .A2(n5140), .ZN(n9811) );
  NAND2_X1 U6568 ( .A1(n9810), .A2(n5140), .ZN(n7167) );
  NAND2_X1 U6569 ( .A1(n6492), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5149) );
  INV_X1 U6570 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6703) );
  OR2_X1 U6571 ( .A1(n5162), .A2(n6703), .ZN(n5148) );
  NAND3_X1 U6572 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5165) );
  INV_X1 U6573 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U6574 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5141) );
  NAND2_X1 U6575 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  NAND2_X1 U6576 ( .A1(n5165), .A2(n5143), .ZN(n7280) );
  OR2_X1 U6577 ( .A1(n5163), .A2(n7280), .ZN(n5147) );
  INV_X1 U6578 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5144) );
  OR2_X1 U6579 ( .A1(n5145), .A2(n5144), .ZN(n5146) );
  NAND2_X1 U6580 ( .A1(n8270), .A2(n7901), .ZN(n5159) );
  INV_X1 U6581 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6582 ( .A1(n5151), .A2(n5150), .ZN(n5194) );
  NAND2_X1 U6583 ( .A1(n5194), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6584 ( .A1(n5152), .A2(n5192), .ZN(n5172) );
  OR2_X1 U6585 ( .A1(n5152), .A2(n5192), .ZN(n5153) );
  INV_X1 U6586 ( .A(n6728), .ZN(n6710) );
  NAND2_X1 U6587 ( .A1(n5156), .A2(SI_4_), .ZN(n5157) );
  XNOR2_X1 U6588 ( .A(n5176), .B(n10161), .ZN(n5174) );
  INV_X1 U6589 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6590) );
  OR2_X1 U6590 ( .A1(n5199), .A2(n6590), .ZN(n5158) );
  XNOR2_X1 U6591 ( .A(n7283), .B(n5639), .ZN(n5160) );
  XNOR2_X1 U6592 ( .A(n5159), .B(n5160), .ZN(n7166) );
  NAND2_X1 U6593 ( .A1(n5161), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5171) );
  INV_X1 U6594 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7233) );
  OR2_X1 U6595 ( .A1(n6663), .A2(n7233), .ZN(n5170) );
  INV_X1 U6596 ( .A(n5165), .ZN(n5164) );
  NAND2_X1 U6597 ( .A1(n5164), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5184) );
  INV_X1 U6598 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6722) );
  NAND2_X1 U6599 ( .A1(n5165), .A2(n6722), .ZN(n5166) );
  NAND2_X1 U6600 ( .A1(n5184), .A2(n5166), .ZN(n7320) );
  OR2_X1 U6601 ( .A1(n5658), .A2(n7320), .ZN(n5169) );
  INV_X1 U6602 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6724) );
  OR2_X1 U6603 ( .A1(n5167), .A2(n6724), .ZN(n5168) );
  OR2_X1 U6604 ( .A1(n7261), .A2(n7018), .ZN(n5180) );
  NAND2_X1 U6605 ( .A1(n5172), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5173) );
  XNOR2_X1 U6606 ( .A(n5173), .B(n5191), .ZN(n6743) );
  NAND2_X1 U6607 ( .A1(n5176), .A2(SI_5_), .ZN(n5177) );
  XNOR2_X1 U6608 ( .A(n5197), .B(SI_6_), .ZN(n5196) );
  OR2_X1 U6609 ( .A1(n4476), .A2(n6602), .ZN(n5178) );
  XNOR2_X1 U6610 ( .A(n7312), .B(n5639), .ZN(n5179) );
  NAND2_X1 U6611 ( .A1(n5180), .A2(n5179), .ZN(n5181) );
  OAI21_X1 U6612 ( .B1(n5180), .B2(n5179), .A(n5181), .ZN(n7319) );
  NAND2_X1 U6613 ( .A1(n5161), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5190) );
  INV_X1 U6614 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7265) );
  OR2_X1 U6615 ( .A1(n6663), .A2(n7265), .ZN(n5189) );
  INV_X1 U6616 ( .A(n5184), .ZN(n5182) );
  NAND2_X1 U6617 ( .A1(n5182), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5209) );
  INV_X1 U6618 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6619 ( .A1(n5184), .A2(n5183), .ZN(n5185) );
  NAND2_X1 U6620 ( .A1(n5209), .A2(n5185), .ZN(n7414) );
  OR2_X1 U6621 ( .A1(n5658), .A2(n7414), .ZN(n5188) );
  INV_X1 U6622 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5186) );
  OR2_X1 U6623 ( .A1(n5167), .A2(n5186), .ZN(n5187) );
  OR2_X1 U6624 ( .A1(n7345), .A2(n7018), .ZN(n5202) );
  NAND2_X1 U6625 ( .A1(n5192), .A2(n5191), .ZN(n5193) );
  NAND2_X1 U6626 ( .A1(n5216), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5195) );
  XNOR2_X1 U6627 ( .A(n5195), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6740) );
  INV_X1 U6628 ( .A(n6740), .ZN(n6759) );
  INV_X1 U6629 ( .A(n5197), .ZN(n5198) );
  XNOR2_X1 U6630 ( .A(n5220), .B(n10175), .ZN(n5218) );
  XNOR2_X1 U6631 ( .A(n5219), .B(n5218), .ZN(n6604) );
  OR2_X1 U6632 ( .A1(n5249), .A2(n6604), .ZN(n5201) );
  INV_X1 U6633 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6603) );
  OR2_X1 U6634 ( .A1(n4476), .A2(n6603), .ZN(n5200) );
  OAI211_X1 U6635 ( .C1(n6689), .C2(n6759), .A(n5201), .B(n5200), .ZN(n7255)
         );
  XNOR2_X1 U6636 ( .A(n7255), .B(n5639), .ZN(n5203) );
  XNOR2_X1 U6637 ( .A(n5202), .B(n5203), .ZN(n7407) );
  INV_X1 U6638 ( .A(n5202), .ZN(n5205) );
  INV_X1 U6639 ( .A(n5203), .ZN(n5204) );
  NAND2_X1 U6640 ( .A1(n5205), .A2(n5204), .ZN(n5206) );
  NAND2_X1 U6641 ( .A1(n6492), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5215) );
  INV_X1 U6642 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6745) );
  OR2_X1 U6643 ( .A1(n6663), .A2(n6745), .ZN(n5214) );
  INV_X1 U6644 ( .A(n5209), .ZN(n5208) );
  NAND2_X1 U6645 ( .A1(n5208), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5235) );
  INV_X1 U6646 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10318) );
  NAND2_X1 U6647 ( .A1(n5209), .A2(n10318), .ZN(n5210) );
  NAND2_X1 U6648 ( .A1(n5235), .A2(n5210), .ZN(n7497) );
  OR2_X1 U6649 ( .A1(n5658), .A2(n7497), .ZN(n5213) );
  INV_X1 U6650 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5211) );
  OR2_X1 U6651 ( .A1(n7367), .A2(n7018), .ZN(n5232) );
  OR2_X1 U6652 ( .A1(n5251), .A2(n8680), .ZN(n5217) );
  XNOR2_X1 U6653 ( .A(n5217), .B(n5250), .ZN(n6797) );
  NAND2_X1 U6654 ( .A1(n5219), .A2(n5218), .ZN(n5222) );
  NAND2_X1 U6655 ( .A1(n5220), .A2(SI_7_), .ZN(n5221) );
  INV_X1 U6656 ( .A(SI_8_), .ZN(n5223) );
  NAND2_X1 U6657 ( .A1(n5224), .A2(n5223), .ZN(n5243) );
  INV_X1 U6658 ( .A(n5224), .ZN(n5225) );
  NAND2_X1 U6659 ( .A1(n5225), .A2(SI_8_), .ZN(n5226) );
  NAND2_X1 U6660 ( .A1(n5243), .A2(n5226), .ZN(n5241) );
  INV_X1 U6661 ( .A(n5241), .ZN(n5227) );
  XNOR2_X1 U6662 ( .A(n5242), .B(n5227), .ZN(n6608) );
  OR2_X1 U6663 ( .A1(n6608), .A2(n5249), .ZN(n5229) );
  OR2_X1 U6664 ( .A1(n5199), .A2(n6609), .ZN(n5228) );
  XNOR2_X1 U6665 ( .A(n7421), .B(n5665), .ZN(n5230) );
  XNOR2_X1 U6666 ( .A(n5232), .B(n5230), .ZN(n7494) );
  INV_X1 U6667 ( .A(n5230), .ZN(n5231) );
  NOR2_X1 U6668 ( .A1(n5232), .A2(n5231), .ZN(n5233) );
  NAND2_X1 U6669 ( .A1(n5161), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5240) );
  INV_X1 U6670 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7375) );
  OR2_X1 U6671 ( .A1(n6663), .A2(n7375), .ZN(n5239) );
  NAND2_X1 U6672 ( .A1(n5235), .A2(n5234), .ZN(n5236) );
  NAND2_X1 U6673 ( .A1(n5274), .A2(n5236), .ZN(n7554) );
  OR2_X1 U6674 ( .A1(n5658), .A2(n7554), .ZN(n5238) );
  INV_X1 U6675 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6790) );
  OR2_X1 U6676 ( .A1(n5167), .A2(n6790), .ZN(n5237) );
  NOR2_X1 U6677 ( .A1(n7472), .A2(n7018), .ZN(n5254) );
  NAND2_X1 U6678 ( .A1(n5246), .A2(n5245), .ZN(n5261) );
  INV_X1 U6679 ( .A(n5246), .ZN(n5247) );
  NAND2_X1 U6680 ( .A1(n5247), .A2(SI_9_), .ZN(n5248) );
  XNOR2_X1 U6681 ( .A(n5260), .B(n5020), .ZN(n6632) );
  NAND2_X1 U6682 ( .A1(n6632), .A2(n7890), .ZN(n5253) );
  NAND2_X1 U6683 ( .A1(n5251), .A2(n5250), .ZN(n5317) );
  NAND2_X1 U6684 ( .A1(n5317), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5268) );
  XNOR2_X1 U6685 ( .A(n5268), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6845) );
  AOI22_X1 U6686 ( .A1(n5483), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6666), .B2(
        n6845), .ZN(n5252) );
  NAND2_X1 U6687 ( .A1(n5253), .A2(n5252), .ZN(n7377) );
  XNOR2_X1 U6688 ( .A(n7377), .B(n5665), .ZN(n5255) );
  NAND2_X1 U6689 ( .A1(n5254), .A2(n5255), .ZN(n5258) );
  INV_X1 U6690 ( .A(n5254), .ZN(n5257) );
  INV_X1 U6691 ( .A(n5255), .ZN(n5256) );
  NAND2_X1 U6692 ( .A1(n5257), .A2(n5256), .ZN(n5259) );
  AND2_X1 U6693 ( .A1(n5258), .A2(n5259), .ZN(n7549) );
  INV_X1 U6694 ( .A(n5265), .ZN(n5266) );
  NAND2_X1 U6695 ( .A1(n5266), .A2(SI_10_), .ZN(n5267) );
  XNOR2_X1 U6696 ( .A(n5284), .B(n5023), .ZN(n6659) );
  NAND2_X1 U6697 ( .A1(n6659), .A2(n7890), .ZN(n5273) );
  INV_X1 U6698 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6699 ( .A1(n5268), .A2(n5314), .ZN(n5269) );
  NAND2_X1 U6700 ( .A1(n5269), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5270) );
  INV_X1 U6701 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6702 ( .A1(n5270), .A2(n5315), .ZN(n5287) );
  OR2_X1 U6703 ( .A1(n5270), .A2(n5315), .ZN(n5271) );
  AOI22_X1 U6704 ( .A1(n5483), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6666), .B2(
        n6997), .ZN(n5272) );
  XNOR2_X1 U6705 ( .A(n7617), .B(n5665), .ZN(n5280) );
  NAND2_X1 U6706 ( .A1(n6492), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U6707 ( .A1(n5161), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5278) );
  INV_X1 U6708 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7476) );
  OR2_X1 U6709 ( .A1(n6663), .A2(n7476), .ZN(n5277) );
  NAND2_X1 U6710 ( .A1(n5274), .A2(n10112), .ZN(n5275) );
  NAND2_X1 U6711 ( .A1(n5293), .A2(n5275), .ZN(n7620) );
  OR2_X1 U6712 ( .A1(n5658), .A2(n7620), .ZN(n5276) );
  NAND4_X1 U6713 ( .A1(n5279), .A2(n5278), .A3(n5277), .A4(n5276), .ZN(n8265)
         );
  NAND2_X1 U6714 ( .A1(n8265), .A2(n7901), .ZN(n5281) );
  XNOR2_X1 U6715 ( .A(n5280), .B(n5281), .ZN(n7614) );
  INV_X1 U6716 ( .A(n5280), .ZN(n5283) );
  INV_X1 U6717 ( .A(n5281), .ZN(n5282) );
  XNOR2_X1 U6718 ( .A(n5309), .B(n5305), .ZN(n6673) );
  NAND2_X1 U6719 ( .A1(n6673), .A2(n7890), .ZN(n5290) );
  NAND2_X1 U6720 ( .A1(n5287), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5288) );
  XNOR2_X1 U6721 ( .A(n5288), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7107) );
  AOI22_X1 U6722 ( .A1(n5483), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6666), .B2(
        n7107), .ZN(n5289) );
  NAND2_X1 U6723 ( .A1(n5290), .A2(n5289), .ZN(n7523) );
  XNOR2_X1 U6724 ( .A(n7523), .B(n5639), .ZN(n5300) );
  NAND2_X1 U6725 ( .A1(n6492), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5299) );
  INV_X1 U6726 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6991) );
  OR2_X1 U6727 ( .A1(n6663), .A2(n6991), .ZN(n5298) );
  INV_X1 U6728 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6729 ( .A1(n5293), .A2(n5292), .ZN(n5294) );
  NAND2_X1 U6730 ( .A1(n5322), .A2(n5294), .ZN(n7521) );
  OR2_X1 U6731 ( .A1(n5658), .A2(n7521), .ZN(n5297) );
  INV_X1 U6732 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5295) );
  OR2_X1 U6733 ( .A1(n6495), .A2(n5295), .ZN(n5296) );
  NOR2_X1 U6734 ( .A1(n7535), .A2(n7018), .ZN(n5301) );
  XNOR2_X1 U6735 ( .A(n5300), .B(n5301), .ZN(n6522) );
  NAND2_X1 U6736 ( .A1(n6523), .A2(n6522), .ZN(n5304) );
  INV_X1 U6737 ( .A(n5300), .ZN(n5302) );
  NAND2_X1 U6738 ( .A1(n5302), .A2(n5301), .ZN(n5303) );
  NAND2_X1 U6739 ( .A1(n5304), .A2(n5303), .ZN(n7770) );
  NAND2_X1 U6740 ( .A1(n5306), .A2(SI_11_), .ZN(n5307) );
  INV_X1 U6741 ( .A(n5310), .ZN(n5311) );
  NAND2_X1 U6742 ( .A1(n5311), .A2(SI_12_), .ZN(n5312) );
  NAND2_X1 U6743 ( .A1(n5335), .A2(n5312), .ZN(n5333) );
  XNOR2_X1 U6744 ( .A(n5334), .B(n5333), .ZN(n6785) );
  NAND2_X1 U6745 ( .A1(n6785), .A2(n7890), .ZN(n5320) );
  INV_X1 U6746 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5313) );
  NAND3_X1 U6747 ( .A1(n5315), .A2(n5314), .A3(n5313), .ZN(n5316) );
  OR2_X1 U6748 ( .A1(n5317), .A2(n5316), .ZN(n5339) );
  NAND2_X1 U6749 ( .A1(n5339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5318) );
  XNOR2_X1 U6750 ( .A(n5318), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7201) );
  AOI22_X1 U6751 ( .A1(n5483), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6666), .B2(
        n7201), .ZN(n5319) );
  XNOR2_X1 U6752 ( .A(n7771), .B(n5639), .ZN(n5328) );
  NAND2_X1 U6753 ( .A1(n5161), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5327) );
  INV_X1 U6754 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7108) );
  OR2_X1 U6755 ( .A1(n5167), .A2(n7108), .ZN(n5326) );
  INV_X1 U6756 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7542) );
  OR2_X1 U6757 ( .A1(n6663), .A2(n7542), .ZN(n5325) );
  INV_X1 U6758 ( .A(n5322), .ZN(n5321) );
  NAND2_X1 U6759 ( .A1(n5321), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5343) );
  INV_X1 U6760 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10257) );
  NAND2_X1 U6761 ( .A1(n5322), .A2(n10257), .ZN(n5323) );
  NAND2_X1 U6762 ( .A1(n5343), .A2(n5323), .ZN(n7775) );
  OR2_X1 U6763 ( .A1(n5658), .A2(n7775), .ZN(n5324) );
  OR2_X1 U6764 ( .A1(n7709), .A2(n7018), .ZN(n5329) );
  NAND2_X1 U6765 ( .A1(n5328), .A2(n5329), .ZN(n7767) );
  NAND2_X1 U6766 ( .A1(n7770), .A2(n7767), .ZN(n5332) );
  INV_X1 U6767 ( .A(n5328), .ZN(n5331) );
  INV_X1 U6768 ( .A(n5329), .ZN(n5330) );
  NAND2_X1 U6769 ( .A1(n5331), .A2(n5330), .ZN(n7768) );
  NAND2_X1 U6770 ( .A1(n5332), .A2(n7768), .ZN(n7838) );
  INV_X1 U6771 ( .A(n5336), .ZN(n5337) );
  NAND2_X1 U6772 ( .A1(n5337), .A2(SI_13_), .ZN(n5338) );
  XNOR2_X1 U6773 ( .A(n5356), .B(n5355), .ZN(n6824) );
  NAND2_X1 U6774 ( .A1(n6824), .A2(n7890), .ZN(n5341) );
  OAI21_X1 U6775 ( .B1(n5339), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5360) );
  XNOR2_X1 U6776 ( .A(n5360), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7335) );
  AOI22_X1 U6777 ( .A1(n5483), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6666), .B2(
        n7335), .ZN(n5340) );
  XNOR2_X1 U6778 ( .A(n7720), .B(n5665), .ZN(n5349) );
  NAND2_X1 U6779 ( .A1(n5161), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5348) );
  INV_X1 U6780 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5342) );
  OR2_X1 U6781 ( .A1(n5167), .A2(n5342), .ZN(n5347) );
  INV_X1 U6782 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7716) );
  OR2_X1 U6783 ( .A1(n6663), .A2(n7716), .ZN(n5346) );
  NAND2_X1 U6784 ( .A1(n5343), .A2(n7205), .ZN(n5344) );
  NAND2_X1 U6785 ( .A1(n5369), .A2(n5344), .ZN(n7839) );
  OR2_X1 U6786 ( .A1(n5658), .A2(n7839), .ZN(n5345) );
  NOR2_X1 U6787 ( .A1(n7753), .A2(n7018), .ZN(n5350) );
  NAND2_X1 U6788 ( .A1(n5349), .A2(n5350), .ZN(n5354) );
  INV_X1 U6789 ( .A(n5349), .ZN(n5352) );
  INV_X1 U6790 ( .A(n5350), .ZN(n5351) );
  NAND2_X1 U6791 ( .A1(n5352), .A2(n5351), .ZN(n5353) );
  AND2_X1 U6792 ( .A1(n5354), .A2(n5353), .ZN(n7837) );
  NAND2_X1 U6793 ( .A1(n7838), .A2(n7837), .ZN(n7836) );
  NAND2_X1 U6794 ( .A1(n7836), .A2(n5354), .ZN(n8113) );
  MUX2_X1 U6795 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6469), .Z(n5381) );
  XNOR2_X1 U6796 ( .A(n5384), .B(n5380), .ZN(n6834) );
  NAND2_X1 U6797 ( .A1(n6834), .A2(n7890), .ZN(n5366) );
  INV_X1 U6798 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6799 ( .A1(n5360), .A2(n5359), .ZN(n5361) );
  NAND2_X1 U6800 ( .A1(n5361), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5363) );
  INV_X1 U6801 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6802 ( .A1(n5363), .A2(n5362), .ZN(n5405) );
  OR2_X1 U6803 ( .A1(n5363), .A2(n5362), .ZN(n5364) );
  AOI22_X1 U6804 ( .A1(n5483), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6666), .B2(
        n7592), .ZN(n5365) );
  XNOR2_X1 U6805 ( .A(n8120), .B(n5665), .ZN(n5375) );
  NAND2_X1 U6806 ( .A1(n5161), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5374) );
  INV_X1 U6807 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5367) );
  OR2_X1 U6808 ( .A1(n5167), .A2(n5367), .ZN(n5373) );
  INV_X1 U6809 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7761) );
  OR2_X1 U6810 ( .A1(n6663), .A2(n7761), .ZN(n5372) );
  INV_X1 U6811 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10260) );
  NAND2_X1 U6812 ( .A1(n5369), .A2(n10260), .ZN(n5370) );
  NAND2_X1 U6813 ( .A1(n5411), .A2(n5370), .ZN(n8118) );
  OR2_X1 U6814 ( .A1(n5658), .A2(n8118), .ZN(n5371) );
  NOR2_X1 U6815 ( .A1(n7823), .A2(n7018), .ZN(n5376) );
  XNOR2_X1 U6816 ( .A(n5375), .B(n5376), .ZN(n8114) );
  INV_X1 U6817 ( .A(n5375), .ZN(n5378) );
  INV_X1 U6818 ( .A(n5376), .ZN(n5377) );
  NAND2_X1 U6819 ( .A1(n5378), .A2(n5377), .ZN(n5379) );
  NAND2_X1 U6820 ( .A1(n5381), .A2(SI_14_), .ZN(n5382) );
  MUX2_X1 U6821 ( .A(n6984), .B(n10097), .S(n6469), .Z(n5386) );
  INV_X1 U6822 ( .A(SI_15_), .ZN(n5385) );
  NAND2_X1 U6823 ( .A1(n5386), .A2(n5385), .ZN(n5389) );
  INV_X1 U6824 ( .A(n5386), .ZN(n5387) );
  NAND2_X1 U6825 ( .A1(n5387), .A2(SI_15_), .ZN(n5388) );
  NAND2_X1 U6826 ( .A1(n5389), .A2(n5388), .ZN(n5403) );
  MUX2_X1 U6827 ( .A(n6986), .B(n10107), .S(n6469), .Z(n5390) );
  INV_X1 U6828 ( .A(n5390), .ZN(n5391) );
  NAND2_X1 U6829 ( .A1(n5391), .A2(SI_16_), .ZN(n5392) );
  XNOR2_X1 U6830 ( .A(n5427), .B(n5426), .ZN(n6985) );
  NAND2_X1 U6831 ( .A1(n6985), .A2(n7890), .ZN(n5396) );
  NAND2_X1 U6832 ( .A1(n5393), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5394) );
  XNOR2_X1 U6833 ( .A(n5394), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8304) );
  AOI22_X1 U6834 ( .A1(n5483), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6666), .B2(
        n8304), .ZN(n5395) );
  XNOR2_X1 U6835 ( .A(n8550), .B(n5665), .ZN(n8167) );
  NAND2_X1 U6836 ( .A1(n5161), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5402) );
  INV_X1 U6837 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8632) );
  OR2_X1 U6838 ( .A1(n5167), .A2(n8632), .ZN(n5401) );
  INV_X1 U6839 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8552) );
  OR2_X1 U6840 ( .A1(n6663), .A2(n8552), .ZN(n5400) );
  INV_X1 U6841 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5410) );
  INV_X1 U6842 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8171) );
  NAND2_X1 U6843 ( .A1(n5413), .A2(n8171), .ZN(n5398) );
  NAND2_X1 U6844 ( .A1(n5439), .A2(n5398), .ZN(n8551) );
  OR2_X1 U6845 ( .A1(n5658), .A2(n8551), .ZN(n5399) );
  NOR2_X1 U6846 ( .A1(n7824), .A2(n7018), .ZN(n5421) );
  XNOR2_X1 U6847 ( .A(n5404), .B(n5403), .ZN(n6982) );
  NAND2_X1 U6848 ( .A1(n6982), .A2(n7890), .ZN(n5408) );
  NAND2_X1 U6849 ( .A1(n5405), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5406) );
  XNOR2_X1 U6850 ( .A(n5406), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8283) );
  AOI22_X1 U6851 ( .A1(n5483), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6666), .B2(
        n8283), .ZN(n5407) );
  XNOR2_X1 U6852 ( .A(n8245), .B(n5665), .ZN(n5420) );
  NAND2_X1 U6853 ( .A1(n6492), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5418) );
  INV_X1 U6854 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5409) );
  OR2_X1 U6855 ( .A1(n6663), .A2(n5409), .ZN(n5417) );
  NAND2_X1 U6856 ( .A1(n5411), .A2(n5410), .ZN(n5412) );
  NAND2_X1 U6857 ( .A1(n5413), .A2(n5412), .ZN(n8242) );
  OR2_X1 U6858 ( .A1(n5658), .A2(n8242), .ZN(n5416) );
  INV_X1 U6859 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5414) );
  OR2_X1 U6860 ( .A1(n6495), .A2(n5414), .ZN(n5415) );
  NOR2_X1 U6861 ( .A1(n8170), .A2(n7018), .ZN(n8239) );
  AOI22_X1 U6862 ( .A1(n8167), .A2(n5421), .B1(n5420), .B2(n8239), .ZN(n5419)
         );
  INV_X1 U6863 ( .A(n8167), .ZN(n5424) );
  OAI21_X1 U6864 ( .B1(n5420), .B2(n8239), .A(n5421), .ZN(n5423) );
  INV_X1 U6865 ( .A(n5420), .ZN(n8165) );
  INV_X1 U6866 ( .A(n8239), .ZN(n5422) );
  INV_X1 U6867 ( .A(n5421), .ZN(n8166) );
  AOI21_X1 U6868 ( .B1(n5424), .B2(n5423), .A(n4511), .ZN(n5425) );
  INV_X1 U6869 ( .A(n8178), .ZN(n5451) );
  MUX2_X1 U6870 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n6469), .Z(n5454) );
  XNOR2_X1 U6871 ( .A(n5454), .B(n5430), .ZN(n5453) );
  XNOR2_X1 U6872 ( .A(n5457), .B(n5453), .ZN(n7064) );
  NAND2_X1 U6873 ( .A1(n7064), .A2(n7890), .ZN(n5438) );
  INV_X1 U6874 ( .A(n5431), .ZN(n5432) );
  NAND2_X1 U6875 ( .A1(n5432), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5433) );
  MUX2_X1 U6876 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5433), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5434) );
  INV_X1 U6877 ( .A(n5434), .ZN(n5436) );
  NOR2_X1 U6878 ( .A1(n5436), .A2(n5435), .ZN(n8321) );
  AOI22_X1 U6879 ( .A1(n5483), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6666), .B2(
        n8321), .ZN(n5437) );
  XNOR2_X1 U6880 ( .A(n8535), .B(n5665), .ZN(n5445) );
  NAND2_X1 U6881 ( .A1(n6492), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5444) );
  OR2_X1 U6882 ( .A1(n6663), .A2(n8299), .ZN(n5443) );
  INV_X1 U6883 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U6884 ( .A1(n5439), .A2(n8181), .ZN(n5440) );
  NAND2_X1 U6885 ( .A1(n5462), .A2(n5440), .ZN(n8524) );
  OR2_X1 U6886 ( .A1(n5658), .A2(n8524), .ZN(n5442) );
  INV_X1 U6887 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8671) );
  OR2_X1 U6888 ( .A1(n6495), .A2(n8671), .ZN(n5441) );
  NOR2_X1 U6889 ( .A1(n8217), .A2(n7018), .ZN(n5446) );
  NAND2_X1 U6890 ( .A1(n5445), .A2(n5446), .ZN(n5452) );
  INV_X1 U6891 ( .A(n5445), .ZN(n5448) );
  INV_X1 U6892 ( .A(n5446), .ZN(n5447) );
  NAND2_X1 U6893 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  NAND2_X1 U6894 ( .A1(n5452), .A2(n5449), .ZN(n8177) );
  INV_X1 U6895 ( .A(n8177), .ZN(n5450) );
  NAND2_X1 U6896 ( .A1(n5451), .A2(n5450), .ZN(n8179) );
  NAND2_X1 U6897 ( .A1(n8179), .A2(n5452), .ZN(n8216) );
  INV_X1 U6898 ( .A(n5453), .ZN(n5456) );
  NAND2_X1 U6899 ( .A1(n5454), .A2(SI_17_), .ZN(n5455) );
  MUX2_X1 U6900 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6469), .Z(n5477) );
  XNOR2_X1 U6901 ( .A(n5477), .B(SI_18_), .ZN(n5474) );
  XNOR2_X1 U6902 ( .A(n5476), .B(n5474), .ZN(n7210) );
  NAND2_X1 U6903 ( .A1(n7210), .A2(n7890), .ZN(n5460) );
  OR2_X1 U6904 ( .A1(n5435), .A2(n8680), .ZN(n5458) );
  XNOR2_X1 U6905 ( .A(n5458), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8332) );
  AOI22_X1 U6906 ( .A1(n5483), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6666), .B2(
        n8332), .ZN(n5459) );
  XNOR2_X1 U6907 ( .A(n8514), .B(n5665), .ZN(n5468) );
  NAND2_X1 U6908 ( .A1(n5161), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5467) );
  INV_X1 U6909 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8621) );
  OR2_X1 U6910 ( .A1(n5167), .A2(n8621), .ZN(n5466) );
  INV_X1 U6911 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8516) );
  OR2_X1 U6912 ( .A1(n6663), .A2(n8516), .ZN(n5465) );
  INV_X1 U6913 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U6914 ( .A1(n5462), .A2(n8317), .ZN(n5463) );
  NAND2_X1 U6915 ( .A1(n5486), .A2(n5463), .ZN(n8515) );
  OR2_X1 U6916 ( .A1(n5658), .A2(n8515), .ZN(n5464) );
  NAND4_X1 U6917 ( .A1(n5467), .A2(n5466), .A3(n5465), .A4(n5464), .ZN(n8258)
         );
  AND2_X1 U6918 ( .A1(n8258), .A2(n7901), .ZN(n5469) );
  NAND2_X1 U6919 ( .A1(n5468), .A2(n5469), .ZN(n5473) );
  INV_X1 U6920 ( .A(n5468), .ZN(n5471) );
  INV_X1 U6921 ( .A(n5469), .ZN(n5470) );
  NAND2_X1 U6922 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  AND2_X1 U6923 ( .A1(n5473), .A2(n5472), .ZN(n8215) );
  NAND2_X1 U6924 ( .A1(n8216), .A2(n8215), .ZN(n8214) );
  NAND2_X1 U6925 ( .A1(n8214), .A2(n5473), .ZN(n8134) );
  INV_X1 U6926 ( .A(n8134), .ZN(n5493) );
  NAND2_X1 U6927 ( .A1(n5477), .A2(SI_18_), .ZN(n5478) );
  MUX2_X1 U6928 ( .A(n7306), .B(n7308), .S(n6469), .Z(n5480) );
  INV_X1 U6929 ( .A(SI_19_), .ZN(n10071) );
  NAND2_X1 U6930 ( .A1(n5480), .A2(n10071), .ZN(n5499) );
  INV_X1 U6931 ( .A(n5480), .ZN(n5481) );
  NAND2_X1 U6932 ( .A1(n5481), .A2(SI_19_), .ZN(n5482) );
  NAND2_X1 U6933 ( .A1(n5499), .A2(n5482), .ZN(n5497) );
  XNOR2_X1 U6934 ( .A(n5498), .B(n5497), .ZN(n7305) );
  NAND2_X1 U6935 ( .A1(n7305), .A2(n7890), .ZN(n5485) );
  AOI22_X1 U6936 ( .A1(n5483), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7923), .B2(
        n6666), .ZN(n5484) );
  XNOR2_X1 U6937 ( .A(n8614), .B(n5639), .ZN(n5495) );
  NAND2_X1 U6938 ( .A1(n5161), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5491) );
  INV_X1 U6939 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8330) );
  OR2_X1 U6940 ( .A1(n5167), .A2(n8330), .ZN(n5490) );
  INV_X1 U6941 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8495) );
  OR2_X1 U6942 ( .A1(n6663), .A2(n8495), .ZN(n5489) );
  INV_X1 U6943 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U6944 ( .A1(n5486), .A2(n10304), .ZN(n5487) );
  NAND2_X1 U6945 ( .A1(n5507), .A2(n5487), .ZN(n8494) );
  OR2_X1 U6946 ( .A1(n5658), .A2(n8494), .ZN(n5488) );
  NAND4_X1 U6947 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5488), .ZN(n8257)
         );
  NAND2_X1 U6948 ( .A1(n8257), .A2(n7901), .ZN(n5494) );
  XNOR2_X1 U6949 ( .A(n5495), .B(n5494), .ZN(n8135) );
  INV_X1 U6950 ( .A(n8135), .ZN(n5492) );
  NAND2_X1 U6951 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  MUX2_X1 U6952 ( .A(n7441), .B(n7427), .S(n6469), .Z(n5500) );
  NAND2_X1 U6953 ( .A1(n5500), .A2(n10306), .ZN(n5521) );
  INV_X1 U6954 ( .A(n5500), .ZN(n5501) );
  NAND2_X1 U6955 ( .A1(n5501), .A2(SI_20_), .ZN(n5502) );
  XNOR2_X1 U6956 ( .A(n5520), .B(n5519), .ZN(n7426) );
  NAND2_X1 U6957 ( .A1(n7426), .A2(n7890), .ZN(n5504) );
  OR2_X1 U6958 ( .A1(n5199), .A2(n7441), .ZN(n5503) );
  NAND2_X2 U6959 ( .A1(n5504), .A2(n5503), .ZN(n8487) );
  XNOR2_X1 U6960 ( .A(n8487), .B(n5665), .ZN(n5513) );
  NAND2_X1 U6961 ( .A1(n6492), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5512) );
  INV_X1 U6962 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8488) );
  OR2_X1 U6963 ( .A1(n6663), .A2(n8488), .ZN(n5511) );
  INV_X1 U6964 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U6965 ( .A1(n5507), .A2(n5506), .ZN(n5508) );
  NAND2_X1 U6966 ( .A1(n5525), .A2(n5508), .ZN(n8478) );
  OR2_X1 U6967 ( .A1(n5658), .A2(n8478), .ZN(n5510) );
  INV_X1 U6968 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8662) );
  OR2_X1 U6969 ( .A1(n6495), .A2(n8662), .ZN(n5509) );
  NOR2_X1 U6970 ( .A1(n8146), .A2(n7018), .ZN(n5514) );
  NAND2_X1 U6971 ( .A1(n5513), .A2(n5514), .ZN(n5518) );
  INV_X1 U6972 ( .A(n5513), .ZN(n5516) );
  INV_X1 U6973 ( .A(n5514), .ZN(n5515) );
  NAND2_X1 U6974 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  AND2_X1 U6975 ( .A1(n5518), .A2(n5517), .ZN(n8199) );
  MUX2_X1 U6976 ( .A(n7464), .B(n7452), .S(n6469), .Z(n5537) );
  XNOR2_X1 U6977 ( .A(n5537), .B(SI_21_), .ZN(n5536) );
  XNOR2_X1 U6978 ( .A(n5535), .B(n5536), .ZN(n7451) );
  NAND2_X1 U6979 ( .A1(n7451), .A2(n7890), .ZN(n5524) );
  OR2_X1 U6980 ( .A1(n4476), .A2(n7464), .ZN(n5523) );
  XNOR2_X1 U6981 ( .A(n8468), .B(n5639), .ZN(n5533) );
  INV_X1 U6982 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10176) );
  NAND2_X1 U6983 ( .A1(n5525), .A2(n10176), .ZN(n5526) );
  NAND2_X1 U6984 ( .A1(n5579), .A2(n5526), .ZN(n8145) );
  OR2_X1 U6985 ( .A1(n8145), .A2(n5658), .ZN(n5530) );
  NAND2_X1 U6986 ( .A1(n6492), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U6987 ( .A1(n6491), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U6988 ( .A1(n5161), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5527) );
  INV_X1 U6989 ( .A(n8207), .ZN(n8255) );
  NAND2_X1 U6990 ( .A1(n8255), .A2(n7901), .ZN(n5531) );
  XNOR2_X1 U6991 ( .A(n5533), .B(n5531), .ZN(n8143) );
  INV_X1 U6992 ( .A(n5531), .ZN(n5532) );
  NAND2_X1 U6993 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  NAND2_X1 U6994 ( .A1(n8142), .A2(n5534), .ZN(n5553) );
  INV_X1 U6995 ( .A(n5537), .ZN(n5538) );
  NAND2_X1 U6996 ( .A1(n5538), .A2(SI_21_), .ZN(n5539) );
  MUX2_X1 U6997 ( .A(n7531), .B(n10122), .S(n6469), .Z(n5540) );
  INV_X1 U6998 ( .A(SI_22_), .ZN(n10261) );
  NAND2_X1 U6999 ( .A1(n5540), .A2(n10261), .ZN(n5556) );
  INV_X1 U7000 ( .A(n5540), .ZN(n5541) );
  NAND2_X1 U7001 ( .A1(n5541), .A2(SI_22_), .ZN(n5542) );
  NAND2_X1 U7002 ( .A1(n5556), .A2(n5542), .ZN(n5557) );
  XNOR2_X1 U7003 ( .A(n5558), .B(n5557), .ZN(n7529) );
  NAND2_X1 U7004 ( .A1(n7529), .A2(n7890), .ZN(n5544) );
  OR2_X1 U7005 ( .A1(n5199), .A2(n7531), .ZN(n5543) );
  XNOR2_X1 U7006 ( .A(n8600), .B(n5639), .ZN(n5551) );
  XNOR2_X1 U7007 ( .A(n5579), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U7008 ( .A1(n8455), .A2(n5718), .ZN(n5550) );
  INV_X1 U7009 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U7010 ( .A1(n6492), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7011 ( .A1(n6491), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5545) );
  OAI211_X1 U7012 ( .C1(n5547), .C2(n6495), .A(n5546), .B(n5545), .ZN(n5548)
         );
  INV_X1 U7013 ( .A(n5548), .ZN(n5549) );
  OR2_X1 U7014 ( .A1(n8147), .A2(n7018), .ZN(n8206) );
  NAND2_X1 U7015 ( .A1(n8205), .A2(n8206), .ZN(n5555) );
  INV_X1 U7016 ( .A(n5551), .ZN(n5552) );
  OR2_X1 U7017 ( .A1(n5553), .A2(n5552), .ZN(n5554) );
  NAND2_X1 U7018 ( .A1(n5555), .A2(n5554), .ZN(n5588) );
  INV_X1 U7019 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5559) );
  MUX2_X1 U7020 ( .A(n7604), .B(n5559), .S(n6469), .Z(n5560) );
  INV_X1 U7021 ( .A(SI_23_), .ZN(n10287) );
  NAND2_X1 U7022 ( .A1(n5560), .A2(n10287), .ZN(n5567) );
  INV_X1 U7023 ( .A(n5560), .ZN(n5561) );
  NAND2_X1 U7024 ( .A1(n5561), .A2(SI_23_), .ZN(n5562) );
  NAND2_X1 U7025 ( .A1(n7602), .A2(n7890), .ZN(n5564) );
  OR2_X1 U7026 ( .A1(n4476), .A2(n7604), .ZN(n5563) );
  XNOR2_X1 U7027 ( .A(n8442), .B(n5665), .ZN(n5586) );
  XNOR2_X1 U7028 ( .A(n5588), .B(n5586), .ZN(n8126) );
  MUX2_X1 U7029 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n6469), .Z(n5593) );
  INV_X1 U7030 ( .A(SI_24_), .ZN(n10274) );
  XNOR2_X1 U7031 ( .A(n5593), .B(n10274), .ZN(n5592) );
  XNOR2_X1 U7032 ( .A(n5596), .B(n5592), .ZN(n7641) );
  NAND2_X1 U7033 ( .A1(n7641), .A2(n7890), .ZN(n5570) );
  INV_X1 U7034 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7692) );
  OR2_X1 U7035 ( .A1(n5199), .A2(n7692), .ZN(n5569) );
  XNOR2_X1 U7036 ( .A(n8590), .B(n5639), .ZN(n8189) );
  NAND2_X1 U7037 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5571) );
  INV_X1 U7038 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U7039 ( .A1(n5581), .A2(n10315), .ZN(n5573) );
  NAND2_X1 U7040 ( .A1(n5604), .A2(n5573), .ZN(n8424) );
  OR2_X1 U7041 ( .A1(n8424), .A2(n5658), .ZN(n5576) );
  AOI22_X1 U7042 ( .A1(n6491), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n6492), .B2(
        P2_REG1_REG_24__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7043 ( .A1(n5161), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5574) );
  INV_X1 U7044 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5578) );
  INV_X1 U7045 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5577) );
  OAI21_X1 U7046 ( .B1(n5579), .B2(n5578), .A(n5577), .ZN(n5580) );
  AND2_X1 U7047 ( .A1(n5581), .A2(n5580), .ZN(n8441) );
  NAND2_X1 U7048 ( .A1(n8441), .A2(n5718), .ZN(n5584) );
  AOI22_X1 U7049 ( .A1(n6491), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n6492), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7050 ( .A1(n5161), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5582) );
  INV_X1 U7051 ( .A(n8208), .ZN(n8254) );
  NAND2_X1 U7052 ( .A1(n8254), .A2(n7901), .ZN(n8127) );
  AOI21_X1 U7053 ( .B1(n8189), .B2(n8123), .A(n8127), .ZN(n5585) );
  INV_X1 U7054 ( .A(n5586), .ZN(n5587) );
  NOR2_X1 U7055 ( .A1(n5588), .A2(n5587), .ZN(n8186) );
  NAND2_X1 U7056 ( .A1(n4999), .A2(n7901), .ZN(n8188) );
  NAND2_X1 U7057 ( .A1(n8189), .A2(n8188), .ZN(n5589) );
  NAND2_X1 U7058 ( .A1(n5591), .A2(n5590), .ZN(n8156) );
  INV_X1 U7059 ( .A(n5592), .ZN(n5595) );
  NAND2_X1 U7060 ( .A1(n5593), .A2(SI_24_), .ZN(n5594) );
  INV_X1 U7061 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7816) );
  MUX2_X1 U7062 ( .A(n7816), .B(n10301), .S(n6469), .Z(n5597) );
  INV_X1 U7063 ( .A(SI_25_), .ZN(n10110) );
  NAND2_X1 U7064 ( .A1(n5597), .A2(n10110), .ZN(n5615) );
  INV_X1 U7065 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7066 ( .A1(n5598), .A2(SI_25_), .ZN(n5599) );
  NAND2_X1 U7067 ( .A1(n5615), .A2(n5599), .ZN(n5616) );
  NAND2_X1 U7068 ( .A1(n7813), .A2(n7890), .ZN(n5601) );
  OR2_X1 U7069 ( .A1(n4476), .A2(n7816), .ZN(n5600) );
  XNOR2_X1 U7070 ( .A(n8410), .B(n5665), .ZN(n5611) );
  INV_X1 U7071 ( .A(n5604), .ZN(n5602) );
  NAND2_X1 U7072 ( .A1(n5602), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5623) );
  INV_X1 U7073 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U7074 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  NAND2_X1 U7075 ( .A1(n5623), .A2(n5605), .ZN(n8407) );
  OR2_X1 U7076 ( .A1(n8407), .A2(n5658), .ZN(n5610) );
  INV_X1 U7077 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U7078 ( .A1(n6491), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U7079 ( .A1(n6492), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5606) );
  OAI211_X1 U7080 ( .C1(n6495), .C2(n8651), .A(n5607), .B(n5606), .ZN(n5608)
         );
  INV_X1 U7081 ( .A(n5608), .ZN(n5609) );
  AND2_X1 U7082 ( .A1(n8253), .A2(n7901), .ZN(n5612) );
  AND2_X1 U7083 ( .A1(n5611), .A2(n5612), .ZN(n8153) );
  INV_X1 U7084 ( .A(n5611), .ZN(n5614) );
  INV_X1 U7085 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U7086 ( .A1(n5614), .A2(n5613), .ZN(n8152) );
  OAI21_X2 U7087 ( .B1(n8156), .B2(n8153), .A(n8152), .ZN(n8226) );
  INV_X1 U7088 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7862) );
  INV_X1 U7089 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10124) );
  MUX2_X1 U7090 ( .A(n7862), .B(n10124), .S(n6469), .Z(n5618) );
  INV_X1 U7091 ( .A(SI_26_), .ZN(n10095) );
  NAND2_X1 U7092 ( .A1(n5618), .A2(n10095), .ZN(n5633) );
  INV_X1 U7093 ( .A(n5618), .ZN(n5619) );
  NAND2_X1 U7094 ( .A1(n5619), .A2(SI_26_), .ZN(n5620) );
  NAND2_X1 U7095 ( .A1(n7817), .A2(n7890), .ZN(n5622) );
  OR2_X1 U7096 ( .A1(n5199), .A2(n7862), .ZN(n5621) );
  XNOR2_X1 U7097 ( .A(n8577), .B(n5665), .ZN(n5629) );
  INV_X1 U7098 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10288) );
  NAND2_X1 U7099 ( .A1(n5623), .A2(n10288), .ZN(n5624) );
  INV_X1 U7100 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U7101 ( .A1(n6492), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7102 ( .A1(n6491), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5625) );
  OAI211_X1 U7103 ( .C1(n8648), .C2(n6495), .A(n5626), .B(n5625), .ZN(n5627)
         );
  NOR2_X1 U7104 ( .A1(n8157), .A2(n7018), .ZN(n5628) );
  XNOR2_X1 U7105 ( .A(n5629), .B(n5628), .ZN(n8225) );
  NAND2_X1 U7106 ( .A1(n5629), .A2(n5628), .ZN(n5630) );
  OAI21_X2 U7107 ( .B1(n8226), .B2(n8225), .A(n5630), .ZN(n8104) );
  INV_X1 U7108 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8697) );
  MUX2_X1 U7109 ( .A(n8697), .B(n10244), .S(n6469), .Z(n5634) );
  INV_X1 U7110 ( .A(SI_27_), .ZN(n10106) );
  NAND2_X1 U7111 ( .A1(n5634), .A2(n10106), .ZN(n5649) );
  INV_X1 U7112 ( .A(n5634), .ZN(n5635) );
  NAND2_X1 U7113 ( .A1(n5635), .A2(SI_27_), .ZN(n5636) );
  NAND2_X1 U7114 ( .A1(n9519), .A2(n7890), .ZN(n5638) );
  OR2_X1 U7115 ( .A1(n5199), .A2(n8697), .ZN(n5637) );
  XNOR2_X1 U7116 ( .A(n8377), .B(n5639), .ZN(n5643) );
  XNOR2_X1 U7117 ( .A(n5656), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8378) );
  INV_X1 U7118 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U7119 ( .A1(n6491), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7120 ( .A1(n6492), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5640) );
  OAI211_X1 U7121 ( .C1(n8645), .C2(n6495), .A(n5641), .B(n5640), .ZN(n5642)
         );
  NOR2_X1 U7122 ( .A1(n8227), .A2(n7018), .ZN(n5644) );
  XNOR2_X1 U7123 ( .A(n5643), .B(n5644), .ZN(n8103) );
  INV_X1 U7124 ( .A(n5643), .ZN(n5645) );
  AND2_X1 U7125 ( .A1(n5645), .A2(n5644), .ZN(n5646) );
  AOI21_X1 U7126 ( .B1(n8104), .B2(n8103), .A(n5646), .ZN(n5712) );
  MUX2_X1 U7127 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6469), .Z(n6464) );
  INV_X1 U7128 ( .A(SI_28_), .ZN(n6465) );
  XNOR2_X1 U7129 ( .A(n6464), .B(n6465), .ZN(n6462) );
  NAND2_X1 U7130 ( .A1(n9515), .A2(n7890), .ZN(n5652) );
  INV_X1 U7131 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8693) );
  OR2_X1 U7132 ( .A1(n5199), .A2(n8693), .ZN(n5651) );
  INV_X1 U7133 ( .A(n5656), .ZN(n5654) );
  AND2_X1 U7134 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5653) );
  NAND2_X1 U7135 ( .A1(n5654), .A2(n5653), .ZN(n8094) );
  INV_X1 U7136 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10255) );
  INV_X1 U7137 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5655) );
  OAI21_X1 U7138 ( .B1(n5656), .B2(n10255), .A(n5655), .ZN(n5657) );
  NAND2_X1 U7139 ( .A1(n8094), .A2(n5657), .ZN(n5723) );
  OR2_X1 U7140 ( .A1(n5723), .A2(n5658), .ZN(n5664) );
  INV_X1 U7141 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7142 ( .A1(n6492), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U7143 ( .A1(n6491), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5659) );
  OAI211_X1 U7144 ( .C1(n5661), .C2(n6495), .A(n5660), .B(n5659), .ZN(n5662)
         );
  INV_X1 U7145 ( .A(n5662), .ZN(n5663) );
  NOR2_X1 U7146 ( .A1(n8105), .A2(n7018), .ZN(n5666) );
  XNOR2_X1 U7147 ( .A(n5666), .B(n5665), .ZN(n5708) );
  NOR4_X1 U7148 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5675) );
  INV_X1 U7149 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9888) );
  INV_X1 U7150 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9887) );
  INV_X1 U7151 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9886) );
  INV_X1 U7152 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9885) );
  NAND4_X1 U7153 ( .A1(n9888), .A2(n9887), .A3(n9886), .A4(n9885), .ZN(n5672)
         );
  NOR4_X1 U7154 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5670) );
  NOR4_X1 U7155 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5669) );
  NOR4_X1 U7156 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5668) );
  NOR4_X1 U7157 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5667) );
  NAND4_X1 U7158 ( .A1(n5670), .A2(n5669), .A3(n5668), .A4(n5667), .ZN(n5671)
         );
  NOR4_X1 U7159 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n5672), .A4(n5671), .ZN(n5674) );
  NOR4_X1 U7160 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5673) );
  NAND3_X1 U7161 ( .A1(n5675), .A2(n5674), .A3(n5673), .ZN(n5689) );
  NAND2_X1 U7162 ( .A1(n5676), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5677) );
  MUX2_X1 U7163 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5677), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5678) );
  NAND2_X1 U7164 ( .A1(n5678), .A2(n4549), .ZN(n7814) );
  INV_X1 U7165 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7166 ( .A1(n5680), .A2(n5679), .ZN(n5681) );
  INV_X1 U7167 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5682) );
  INV_X1 U7168 ( .A(P2_B_REG_SCAN_IN), .ZN(n10148) );
  XOR2_X1 U7169 ( .A(n7694), .B(n10148), .Z(n5684) );
  NAND2_X1 U7170 ( .A1(n4549), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5685) );
  MUX2_X1 U7171 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5685), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5687) );
  NAND2_X1 U7172 ( .A1(n5687), .A2(n5686), .ZN(n7864) );
  INV_X1 U7173 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U7174 ( .A1(n9857), .A2(n5690), .ZN(n5691) );
  NAND2_X1 U7175 ( .A1(n7694), .A2(n7864), .ZN(n9889) );
  INV_X1 U7176 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U7177 ( .A1(n9857), .A2(n5692), .ZN(n5693) );
  NAND2_X1 U7178 ( .A1(n7864), .A2(n7814), .ZN(n9891) );
  NAND2_X1 U7179 ( .A1(n5693), .A2(n9891), .ZN(n7007) );
  OR2_X1 U7180 ( .A1(n7008), .A2(n7007), .ZN(n5724) );
  INV_X1 U7181 ( .A(n5724), .ZN(n5702) );
  INV_X1 U7182 ( .A(n7694), .ZN(n5695) );
  NOR2_X1 U7183 ( .A1(n7864), .A2(n7814), .ZN(n5694) );
  OR2_X1 U7184 ( .A1(n5697), .A2(n5696), .ZN(n5698) );
  NAND2_X1 U7185 ( .A1(n5699), .A2(n5698), .ZN(n6665) );
  INV_X1 U7186 ( .A(n9892), .ZN(n5700) );
  INV_X1 U7187 ( .A(n9856), .ZN(n5701) );
  NAND2_X1 U7188 ( .A1(n5702), .A2(n5701), .ZN(n5703) );
  NOR2_X1 U7189 ( .A1(n9897), .A2(n8072), .ZN(n7016) );
  NAND2_X1 U7190 ( .A1(n5722), .A2(n7016), .ZN(n5704) );
  OR2_X2 U7191 ( .A1(n9856), .A2(n6505), .ZN(n9845) );
  NOR3_X1 U7192 ( .A1(n8364), .A2(n5708), .A3(n8244), .ZN(n5705) );
  AOI21_X1 U7193 ( .B1(n8364), .B2(n5708), .A(n5705), .ZN(n5706) );
  NAND3_X1 U7194 ( .A1(n8569), .A2(n9819), .A3(n5708), .ZN(n5707) );
  OAI21_X1 U7195 ( .B1(n8569), .B2(n5708), .A(n5707), .ZN(n5711) );
  NAND2_X1 U7196 ( .A1(n8079), .A2(n8069), .ZN(n6668) );
  AND2_X1 U7197 ( .A1(n9940), .A2(n6668), .ZN(n5709) );
  NAND2_X1 U7198 ( .A1(n8569), .A2(n8244), .ZN(n5710) );
  INV_X1 U7199 ( .A(n5713), .ZN(n5714) );
  INV_X1 U7200 ( .A(n6668), .ZN(n6679) );
  OR2_X1 U7201 ( .A1(n8227), .A2(n9812), .ZN(n5721) );
  INV_X1 U7202 ( .A(n8094), .ZN(n5719) );
  INV_X1 U7203 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U7204 ( .A1(n6491), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U7205 ( .A1(n5161), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5715) );
  OAI211_X1 U7206 ( .C1(n6507), .C2(n5167), .A(n5716), .B(n5715), .ZN(n5717)
         );
  AOI21_X1 U7207 ( .B1(n5719), .B2(n5718), .A(n5717), .ZN(n6839) );
  AND2_X1 U7208 ( .A1(n5713), .A2(n6679), .ZN(n8218) );
  OR2_X1 U7209 ( .A1(n6839), .A2(n9814), .ZN(n5720) );
  AND2_X1 U7210 ( .A1(n5721), .A2(n5720), .ZN(n8357) );
  NAND2_X1 U7211 ( .A1(n5722), .A2(n5725), .ZN(n8233) );
  INV_X1 U7212 ( .A(n5723), .ZN(n8361) );
  OAI21_X1 U7213 ( .B1(n6504), .B2(n5724), .A(n6505), .ZN(n6826) );
  OAI21_X1 U7214 ( .B1(n6668), .B2(n5725), .A(n6665), .ZN(n5726) );
  INV_X1 U7215 ( .A(n5726), .ZN(n5727) );
  NAND2_X1 U7216 ( .A1(n6681), .A2(n5727), .ZN(n6503) );
  INV_X1 U7217 ( .A(n6503), .ZN(n5728) );
  NAND2_X1 U7218 ( .A1(n6826), .A2(n5728), .ZN(n5729) );
  INV_X1 U7219 ( .A(n9824), .ZN(n8231) );
  AOI22_X1 U7220 ( .A1(n8361), .A2(n8231), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5730) );
  INV_X2 U7221 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U7222 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5735) );
  NOR2_X1 U7223 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5734) );
  NOR2_X1 U7224 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5733) );
  NAND4_X1 U7225 ( .A1(n5735), .A2(n5734), .A3(n5733), .A4(n6036), .ZN(n5741)
         );
  NOR2_X1 U7226 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5739) );
  NAND4_X1 U7227 ( .A1(n5739), .A2(n5738), .A3(n5737), .A4(n5736), .ZN(n5740)
         );
  NOR2_X1 U7228 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5747) );
  NAND2_X1 U7229 ( .A1(n5750), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U7230 ( .A1(n7602), .A2(n8850), .ZN(n5752) );
  NAND2_X1 U7231 ( .A1(n4474), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5751) );
  INV_X1 U7232 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7233 ( .A1(n5756), .A2(n10293), .ZN(n5757) );
  NAND2_X1 U7234 ( .A1(n5757), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5755) );
  XNOR2_X1 U7235 ( .A(n5755), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6335) );
  OR2_X1 U7236 ( .A1(n5756), .A2(n10293), .ZN(n5758) );
  NAND2_X1 U7237 ( .A1(n5758), .A2(n5757), .ZN(n6336) );
  NAND2_X1 U7238 ( .A1(n5759), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5760) );
  MUX2_X1 U7239 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5760), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5761) );
  NAND2_X1 U7240 ( .A1(n5761), .A2(n4936), .ZN(n7642) );
  NOR2_X1 U7241 ( .A1(n6336), .A2(n7642), .ZN(n5762) );
  NAND2_X1 U7242 ( .A1(n5764), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5766) );
  OR2_X1 U7243 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  NAND2_X1 U7244 ( .A1(n5766), .A2(n5765), .ZN(n5771) );
  NAND2_X1 U7245 ( .A1(n4584), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5769) );
  INV_X1 U7246 ( .A(n6879), .ZN(n5770) );
  INV_X4 U7247 ( .A(n5809), .ZN(n6397) );
  AND2_X2 U7248 ( .A1(n5797), .A2(n6879), .ZN(n5792) );
  NAND2_X1 U7249 ( .A1(n5771), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U7250 ( .A1(n5773), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5774) );
  MUX2_X1 U7251 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5774), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5775) );
  NAND2_X1 U7252 ( .A1(n9042), .A2(n6378), .ZN(n5776) );
  NAND2_X1 U7253 ( .A1(n6323), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5790) );
  INV_X1 U7254 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5781) );
  OR2_X1 U7255 ( .A1(n5866), .A2(n5781), .ZN(n5789) );
  INV_X1 U7256 ( .A(n8092), .ZN(n5782) );
  NAND2_X1 U7257 ( .A1(n5888), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7258 ( .A1(n5945), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5963) );
  INV_X1 U7259 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6088) );
  INV_X1 U7260 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8782) );
  NAND2_X1 U7261 ( .A1(n6253), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6274) );
  OAI21_X1 U7262 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n6253), .A(n6274), .ZN(
        n9298) );
  OR2_X1 U7263 ( .A1(n6405), .A2(n9298), .ZN(n5788) );
  INV_X1 U7264 ( .A(n5784), .ZN(n5785) );
  NAND2_X2 U7265 ( .A1(n5785), .A2(n8092), .ZN(n5852) );
  INV_X1 U7266 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n5786) );
  OR2_X1 U7267 ( .A1(n5852), .A2(n5786), .ZN(n5787) );
  NAND4_X1 U7268 ( .A1(n5790), .A2(n5789), .A3(n5788), .A4(n5787), .ZN(n9316)
         );
  AND2_X1 U7269 ( .A1(n5808), .A2(n9316), .ZN(n5791) );
  AOI21_X1 U7270 ( .B1(n9447), .B2(n6397), .A(n5791), .ZN(n8712) );
  NAND2_X1 U7271 ( .A1(n6469), .A2(SI_0_), .ZN(n5794) );
  INV_X1 U7272 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7273 ( .A1(n5794), .A2(n5793), .ZN(n5796) );
  AND2_X1 U7274 ( .A1(n5796), .A2(n5795), .ZN(n9523) );
  MUX2_X1 U7275 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9523), .S(n5893), .Z(n6933) );
  NAND2_X1 U7276 ( .A1(n5798), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5799) );
  OAI21_X1 U7277 ( .B1(n5835), .B2(n6945), .A(n5799), .ZN(n5800) );
  INV_X1 U7278 ( .A(n5800), .ZN(n5807) );
  NAND2_X1 U7279 ( .A1(n5921), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5805) );
  INV_X1 U7280 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6556) );
  OR2_X1 U7281 ( .A1(n5869), .A2(n6556), .ZN(n5804) );
  INV_X1 U7282 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5801) );
  OR2_X1 U7283 ( .A1(n5852), .A2(n5801), .ZN(n5803) );
  INV_X1 U7284 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U7285 ( .A1(n6776), .A2(n6397), .ZN(n5806) );
  NAND2_X1 U7286 ( .A1(n6776), .A2(n5808), .ZN(n5812) );
  INV_X1 U7287 ( .A(n5810), .ZN(n5811) );
  NAND2_X1 U7288 ( .A1(n6809), .A2(n6808), .ZN(n6807) );
  OAI21_X1 U7289 ( .B1(n6808), .B2(n6309), .A(n6807), .ZN(n5824) );
  INV_X1 U7290 ( .A(n5824), .ZN(n5822) );
  INV_X1 U7291 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5813) );
  OR2_X1 U7292 ( .A1(n5869), .A2(n5813), .ZN(n5818) );
  INV_X1 U7293 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6946) );
  OR2_X1 U7294 ( .A1(n5854), .A2(n6946), .ZN(n5817) );
  INV_X1 U7295 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5814) );
  OR2_X1 U7296 ( .A1(n5852), .A2(n5814), .ZN(n5816) );
  NAND2_X1 U7297 ( .A1(n6872), .A2(n6397), .ZN(n5820) );
  NAND2_X1 U7298 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5819) );
  INV_X1 U7299 ( .A(n5823), .ZN(n5821) );
  NAND2_X1 U7300 ( .A1(n5822), .A2(n5821), .ZN(n6860) );
  NAND2_X1 U7301 ( .A1(n6860), .A2(n6862), .ZN(n5825) );
  NAND2_X1 U7302 ( .A1(n5824), .A2(n5823), .ZN(n6861) );
  NAND2_X1 U7303 ( .A1(n5825), .A2(n6861), .ZN(n8788) );
  NAND2_X1 U7304 ( .A1(n5921), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5829) );
  INV_X1 U7305 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6558) );
  OR2_X1 U7306 ( .A1(n5869), .A2(n6558), .ZN(n5828) );
  INV_X1 U7307 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9623) );
  OR2_X1 U7308 ( .A1(n5854), .A2(n9623), .ZN(n5827) );
  OR2_X1 U7309 ( .A1(n5852), .A2(n9772), .ZN(n5826) );
  NAND2_X1 U7310 ( .A1(n5845), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5833) );
  OR2_X1 U7311 ( .A1(n5830), .A2(n5754), .ZN(n5831) );
  XNOR2_X1 U7312 ( .A(n5831), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U7313 ( .A1(n5846), .A2(n6557), .ZN(n5832) );
  INV_X1 U7314 ( .A(n5841), .ZN(n5839) );
  NAND2_X1 U7315 ( .A1(n9141), .A2(n6397), .ZN(n5837) );
  INV_X2 U7316 ( .A(n5835), .ZN(n6398) );
  NAND2_X1 U7317 ( .A1(n8793), .A2(n6398), .ZN(n5836) );
  NAND2_X1 U7318 ( .A1(n5837), .A2(n5836), .ZN(n5840) );
  XNOR2_X1 U7319 ( .A(n5840), .B(n6887), .ZN(n5838) );
  NAND2_X1 U7320 ( .A1(n5839), .A2(n5838), .ZN(n5843) );
  XNOR2_X1 U7321 ( .A(n5840), .B(n6309), .ZN(n5842) );
  NAND2_X1 U7322 ( .A1(n5842), .A2(n5841), .ZN(n5844) );
  NAND2_X1 U7323 ( .A1(n8789), .A2(n5844), .ZN(n6974) );
  NAND2_X1 U7324 ( .A1(n5845), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U7325 ( .A1(n5848), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5847) );
  MUX2_X1 U7326 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5847), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n5849) );
  AND2_X1 U7327 ( .A1(n5849), .A2(n5894), .ZN(n6580) );
  NAND2_X1 U7328 ( .A1(n5846), .A2(n6580), .ZN(n5850) );
  OAI211_X1 U7329 ( .C1(n6583), .C2(n5834), .A(n5851), .B(n5850), .ZN(n7119)
         );
  NAND2_X1 U7330 ( .A1(n6398), .A2(n7119), .ZN(n5860) );
  NAND2_X1 U7331 ( .A1(n6194), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5858) );
  INV_X1 U7332 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5853) );
  INV_X1 U7333 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6559) );
  OR2_X1 U7334 ( .A1(n8840), .A2(n6559), .ZN(n5856) );
  OR2_X1 U7335 ( .A1(n5854), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U7336 ( .A1(n9140), .A2(n6397), .ZN(n5859) );
  NAND2_X1 U7337 ( .A1(n5860), .A2(n5859), .ZN(n5861) );
  XNOR2_X1 U7338 ( .A(n5861), .B(n6887), .ZN(n5862) );
  AOI22_X1 U7339 ( .A1(n5808), .A2(n9140), .B1(n6397), .B2(n7119), .ZN(n5863)
         );
  XNOR2_X1 U7340 ( .A(n5862), .B(n5863), .ZN(n6976) );
  INV_X1 U7341 ( .A(n5862), .ZN(n5864) );
  NAND2_X1 U7342 ( .A1(n5864), .A2(n5863), .ZN(n5865) );
  NAND2_X1 U7343 ( .A1(n6194), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5874) );
  INV_X1 U7344 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6909) );
  OR2_X1 U7345 ( .A1(n5866), .A2(n6909), .ZN(n5873) );
  INV_X1 U7346 ( .A(n5888), .ZN(n5868) );
  INV_X1 U7347 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7118) );
  INV_X1 U7348 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6967) );
  NAND2_X1 U7349 ( .A1(n7118), .A2(n6967), .ZN(n5867) );
  NAND2_X1 U7350 ( .A1(n5868), .A2(n5867), .ZN(n6971) );
  OR2_X1 U7351 ( .A1(n6405), .A2(n6971), .ZN(n5872) );
  INV_X1 U7352 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5870) );
  OR2_X1 U7353 ( .A1(n8840), .A2(n5870), .ZN(n5871) );
  NAND2_X1 U7354 ( .A1(n9139), .A2(n6397), .ZN(n5879) );
  NAND2_X1 U7355 ( .A1(n4474), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7356 ( .A1(n5894), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5875) );
  XNOR2_X1 U7357 ( .A(n5875), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9654) );
  NAND2_X1 U7358 ( .A1(n5846), .A2(n9654), .ZN(n5876) );
  OAI211_X1 U7359 ( .C1(n6591), .C2(n5834), .A(n5877), .B(n5876), .ZN(n6968)
         );
  NAND2_X1 U7360 ( .A1(n6398), .A2(n6968), .ZN(n5878) );
  NAND2_X1 U7361 ( .A1(n5879), .A2(n5878), .ZN(n5880) );
  XNOR2_X1 U7362 ( .A(n5880), .B(n6309), .ZN(n5882) );
  AOI22_X1 U7363 ( .A1(n5808), .A2(n9139), .B1(n6397), .B2(n6968), .ZN(n5883)
         );
  XNOR2_X1 U7364 ( .A(n5882), .B(n5883), .ZN(n6966) );
  INV_X1 U7365 ( .A(n6966), .ZN(n5881) );
  INV_X1 U7366 ( .A(n5882), .ZN(n5885) );
  INV_X1 U7367 ( .A(n5883), .ZN(n5884) );
  NAND2_X1 U7368 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  NAND2_X1 U7369 ( .A1(n6963), .A2(n5886), .ZN(n5907) );
  INV_X1 U7370 ( .A(n5907), .ZN(n5904) );
  NAND2_X1 U7371 ( .A1(n6194), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5892) );
  INV_X1 U7372 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5887) );
  OR2_X1 U7373 ( .A1(n5866), .A2(n5887), .ZN(n5891) );
  INV_X1 U7374 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6555) );
  OR2_X1 U7375 ( .A1(n8840), .A2(n6555), .ZN(n5890) );
  OAI21_X1 U7376 ( .B1(n5888), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5925), .ZN(
        n9742) );
  OR2_X1 U7377 ( .A1(n6405), .A2(n9742), .ZN(n5889) );
  NAND2_X1 U7378 ( .A1(n9138), .A2(n6397), .ZN(n5902) );
  INV_X1 U7379 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6588) );
  NOR2_X1 U7380 ( .A1(n5897), .A2(n5754), .ZN(n5895) );
  MUX2_X1 U7381 ( .A(n5754), .B(n5895), .S(P1_IR_REG_5__SCAN_IN), .Z(n5898) );
  INV_X1 U7382 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5896) );
  OR2_X1 U7383 ( .A1(n5898), .A2(n5915), .ZN(n6587) );
  OAI22_X1 U7384 ( .A1(n6190), .A2(n6588), .B1(n6521), .B2(n6587), .ZN(n5899)
         );
  INV_X1 U7385 ( .A(n5899), .ZN(n5900) );
  OAI21_X1 U7386 ( .B1(n6589), .B2(n5834), .A(n5900), .ZN(n9739) );
  NAND2_X1 U7387 ( .A1(n6398), .A2(n9739), .ZN(n5901) );
  NAND2_X1 U7388 ( .A1(n5902), .A2(n5901), .ZN(n5903) );
  XNOR2_X1 U7389 ( .A(n5903), .B(n6309), .ZN(n5905) );
  NAND2_X1 U7390 ( .A1(n5904), .A2(n5905), .ZN(n5912) );
  INV_X1 U7391 ( .A(n5905), .ZN(n5906) );
  NAND2_X1 U7392 ( .A1(n5808), .A2(n9138), .ZN(n5910) );
  NAND2_X1 U7393 ( .A1(n6397), .A2(n9739), .ZN(n5909) );
  NAND2_X1 U7394 ( .A1(n5910), .A2(n5909), .ZN(n7081) );
  OR2_X1 U7395 ( .A1(n5834), .A2(n6601), .ZN(n5920) );
  NOR2_X1 U7396 ( .A1(n5915), .A2(n5754), .ZN(n5913) );
  MUX2_X1 U7397 ( .A(n5754), .B(n5913), .S(P1_IR_REG_6__SCAN_IN), .Z(n5917) );
  INV_X1 U7398 ( .A(n6039), .ZN(n5916) );
  OAI22_X1 U7399 ( .A1(n6190), .A2(n6600), .B1(n6521), .B2(n6623), .ZN(n5918)
         );
  INV_X1 U7400 ( .A(n5918), .ZN(n5919) );
  NAND2_X1 U7401 ( .A1(n5920), .A2(n5919), .ZN(n7246) );
  NAND2_X1 U7402 ( .A1(n7246), .A2(n6398), .ZN(n5932) );
  NAND2_X1 U7403 ( .A1(n5921), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5930) );
  INV_X1 U7404 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5922) );
  OR2_X1 U7405 ( .A1(n8840), .A2(n5922), .ZN(n5929) );
  INV_X1 U7406 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5923) );
  OR2_X1 U7407 ( .A1(n5852), .A2(n5923), .ZN(n5928) );
  AND2_X1 U7408 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  OR2_X1 U7409 ( .A1(n5926), .A2(n5945), .ZN(n7244) );
  OR2_X1 U7410 ( .A1(n6405), .A2(n7244), .ZN(n5927) );
  NAND4_X1 U7411 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(n9137)
         );
  NAND2_X1 U7412 ( .A1(n9137), .A2(n6397), .ZN(n5931) );
  NAND2_X1 U7413 ( .A1(n5932), .A2(n5931), .ZN(n5933) );
  XNOR2_X1 U7414 ( .A(n5933), .B(n6887), .ZN(n5936) );
  NAND2_X1 U7415 ( .A1(n5808), .A2(n9137), .ZN(n5935) );
  NAND2_X1 U7416 ( .A1(n7246), .A2(n6397), .ZN(n5934) );
  NAND2_X1 U7417 ( .A1(n5935), .A2(n5934), .ZN(n5937) );
  NAND2_X1 U7418 ( .A1(n5936), .A2(n5937), .ZN(n7136) );
  NAND2_X1 U7419 ( .A1(n7134), .A2(n7136), .ZN(n5940) );
  INV_X1 U7420 ( .A(n5936), .ZN(n5939) );
  INV_X1 U7421 ( .A(n5937), .ZN(n5938) );
  NAND2_X1 U7422 ( .A1(n5939), .A2(n5938), .ZN(n7135) );
  NAND2_X1 U7423 ( .A1(n5940), .A2(n7135), .ZN(n7213) );
  OR2_X1 U7424 ( .A1(n6604), .A2(n5834), .ZN(n5944) );
  INV_X1 U7425 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U7426 ( .A1(n6039), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5941) );
  INV_X1 U7427 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6035) );
  XNOR2_X1 U7428 ( .A(n5941), .B(n6035), .ZN(n9668) );
  OAI22_X1 U7429 ( .A1(n6190), .A2(n6605), .B1(n6521), .B2(n9668), .ZN(n5942)
         );
  INV_X1 U7430 ( .A(n5942), .ZN(n5943) );
  NAND2_X1 U7431 ( .A1(n7219), .A2(n6398), .ZN(n5952) );
  NAND2_X1 U7432 ( .A1(n6194), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5950) );
  INV_X1 U7433 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7034) );
  OR2_X1 U7434 ( .A1(n5866), .A2(n7034), .ZN(n5949) );
  OR2_X1 U7435 ( .A1(n5945), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7436 ( .A1(n5963), .A2(n5946), .ZN(n7216) );
  OR2_X1 U7437 ( .A1(n6405), .A2(n7216), .ZN(n5948) );
  INV_X1 U7438 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6564) );
  OR2_X1 U7439 ( .A1(n8840), .A2(n6564), .ZN(n5947) );
  NAND4_X1 U7440 ( .A1(n5950), .A2(n5949), .A3(n5948), .A4(n5947), .ZN(n9136)
         );
  NAND2_X1 U7441 ( .A1(n9136), .A2(n6397), .ZN(n5951) );
  NAND2_X1 U7442 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  XNOR2_X1 U7443 ( .A(n5953), .B(n6887), .ZN(n5954) );
  AOI22_X1 U7444 ( .A1(n7219), .A2(n6397), .B1(n5808), .B2(n9136), .ZN(n5955)
         );
  XNOR2_X1 U7445 ( .A(n5954), .B(n5955), .ZN(n7214) );
  NAND2_X1 U7446 ( .A1(n7213), .A2(n7214), .ZN(n5958) );
  INV_X1 U7447 ( .A(n5954), .ZN(n5956) );
  NAND2_X1 U7448 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  OR2_X1 U7449 ( .A1(n6608), .A2(n5834), .ZN(n5961) );
  NAND2_X1 U7450 ( .A1(n5959), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5998) );
  XNOR2_X1 U7451 ( .A(n5998), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9681) );
  AOI22_X1 U7452 ( .A1(n4474), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5846), .B2(
        n9681), .ZN(n5960) );
  NAND2_X1 U7453 ( .A1(n6194), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5968) );
  INV_X1 U7454 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6554) );
  OR2_X1 U7455 ( .A1(n8840), .A2(n6554), .ZN(n5967) );
  INV_X1 U7456 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7190) );
  OR2_X1 U7457 ( .A1(n5866), .A2(n7190), .ZN(n5966) );
  NAND2_X1 U7458 ( .A1(n5963), .A2(n5962), .ZN(n5964) );
  NAND2_X1 U7459 ( .A1(n5982), .A2(n5964), .ZN(n7432) );
  OR2_X1 U7460 ( .A1(n6405), .A2(n7432), .ZN(n5965) );
  NAND4_X1 U7461 ( .A1(n5968), .A2(n5967), .A3(n5966), .A4(n5965), .ZN(n9135)
         );
  AND2_X1 U7462 ( .A1(n5808), .A2(n9135), .ZN(n5969) );
  AOI21_X1 U7463 ( .B1(n7436), .B2(n6397), .A(n5969), .ZN(n5974) );
  NAND2_X1 U7464 ( .A1(n5973), .A2(n5974), .ZN(n7428) );
  NAND2_X1 U7465 ( .A1(n7436), .A2(n5792), .ZN(n5971) );
  NAND2_X1 U7466 ( .A1(n9135), .A2(n6397), .ZN(n5970) );
  NAND2_X1 U7467 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  XNOR2_X1 U7468 ( .A(n5972), .B(n6887), .ZN(n7431) );
  NAND2_X1 U7469 ( .A1(n7428), .A2(n7431), .ZN(n5977) );
  INV_X1 U7470 ( .A(n5974), .ZN(n5975) );
  NAND2_X1 U7471 ( .A1(n6632), .A2(n8850), .ZN(n5981) );
  INV_X1 U7472 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7473 ( .A1(n5998), .A2(n6034), .ZN(n5978) );
  NAND2_X1 U7474 ( .A1(n5978), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5979) );
  XNOR2_X1 U7475 ( .A(n5979), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9696) );
  AOI22_X1 U7476 ( .A1(n5845), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5846), .B2(
        n9696), .ZN(n5980) );
  NAND2_X1 U7477 ( .A1(n5981), .A2(n5980), .ZN(n7453) );
  NAND2_X1 U7478 ( .A1(n7453), .A2(n6398), .ZN(n5990) );
  NAND2_X1 U7479 ( .A1(n5921), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5988) );
  AND2_X1 U7480 ( .A1(n5982), .A2(n7446), .ZN(n5983) );
  OR2_X1 U7481 ( .A1(n5983), .A2(n6003), .ZN(n7447) );
  OR2_X1 U7482 ( .A1(n6405), .A2(n7447), .ZN(n5987) );
  INV_X1 U7483 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5984) );
  OR2_X1 U7484 ( .A1(n5852), .A2(n5984), .ZN(n5986) );
  OR2_X1 U7485 ( .A1(n8840), .A2(n9807), .ZN(n5985) );
  NAND4_X1 U7486 ( .A1(n5988), .A2(n5987), .A3(n5986), .A4(n5985), .ZN(n9577)
         );
  NAND2_X1 U7487 ( .A1(n9577), .A2(n6397), .ZN(n5989) );
  NAND2_X1 U7488 ( .A1(n5990), .A2(n5989), .ZN(n5991) );
  XNOR2_X1 U7489 ( .A(n5991), .B(n6887), .ZN(n5993) );
  AND2_X1 U7490 ( .A1(n5808), .A2(n9577), .ZN(n5992) );
  AOI21_X1 U7491 ( .B1(n7453), .B2(n6397), .A(n5992), .ZN(n5994) );
  XNOR2_X1 U7492 ( .A(n5993), .B(n5994), .ZN(n7444) );
  INV_X1 U7493 ( .A(n5993), .ZN(n5995) );
  NAND2_X1 U7494 ( .A1(n5995), .A2(n5994), .ZN(n5996) );
  NAND2_X1 U7495 ( .A1(n6659), .A2(n8850), .ZN(n6002) );
  OAI21_X1 U7496 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7497 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  NAND2_X1 U7498 ( .A1(n5999), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6000) );
  AOI22_X1 U7499 ( .A1(n5845), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5846), .B2(
        n6816), .ZN(n6001) );
  NAND2_X1 U7500 ( .A1(n9587), .A2(n5792), .ZN(n6011) );
  NAND2_X1 U7501 ( .A1(n5921), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6009) );
  INV_X1 U7502 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6552) );
  OR2_X1 U7503 ( .A1(n8840), .A2(n6552), .ZN(n6008) );
  NOR2_X1 U7504 ( .A1(n6003), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6004) );
  OR2_X1 U7505 ( .A1(n6020), .A2(n6004), .ZN(n9582) );
  OR2_X1 U7506 ( .A1(n6405), .A2(n9582), .ZN(n6007) );
  INV_X1 U7507 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6005) );
  OR2_X1 U7508 ( .A1(n5852), .A2(n6005), .ZN(n6006) );
  NAND4_X1 U7509 ( .A1(n6009), .A2(n6008), .A3(n6007), .A4(n6006), .ZN(n9134)
         );
  NAND2_X1 U7510 ( .A1(n9134), .A2(n6397), .ZN(n6010) );
  NAND2_X1 U7511 ( .A1(n6011), .A2(n6010), .ZN(n6012) );
  XNOR2_X1 U7512 ( .A(n6012), .B(n6309), .ZN(n7485) );
  AND2_X1 U7513 ( .A1(n5808), .A2(n9134), .ZN(n6013) );
  AOI21_X1 U7514 ( .B1(n9587), .B2(n6397), .A(n6013), .ZN(n7484) );
  NAND2_X1 U7515 ( .A1(n6673), .A2(n8850), .ZN(n6018) );
  NAND2_X1 U7516 ( .A1(n6015), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6016) );
  XNOR2_X1 U7517 ( .A(n6016), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9704) );
  AOI22_X1 U7518 ( .A1(n4474), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5846), .B2(
        n9704), .ZN(n6017) );
  NAND2_X1 U7519 ( .A1(n7574), .A2(n6398), .ZN(n6028) );
  NAND2_X1 U7520 ( .A1(n6194), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6026) );
  INV_X1 U7521 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6019) );
  OR2_X1 U7522 ( .A1(n5866), .A2(n6019), .ZN(n6025) );
  OR2_X1 U7523 ( .A1(n6020), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7524 ( .A1(n6049), .A2(n6021), .ZN(n7562) );
  OR2_X1 U7525 ( .A1(n6405), .A2(n7562), .ZN(n6024) );
  INV_X1 U7526 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6022) );
  OR2_X1 U7527 ( .A1(n8840), .A2(n6022), .ZN(n6023) );
  NAND4_X1 U7528 ( .A1(n6026), .A2(n6025), .A3(n6024), .A4(n6023), .ZN(n9576)
         );
  NAND2_X1 U7529 ( .A1(n9576), .A2(n6397), .ZN(n6027) );
  NAND2_X1 U7530 ( .A1(n6028), .A2(n6027), .ZN(n6029) );
  XNOR2_X1 U7531 ( .A(n6029), .B(n6887), .ZN(n6033) );
  AND2_X1 U7532 ( .A1(n5808), .A2(n9576), .ZN(n6030) );
  AOI21_X1 U7533 ( .B1(n7574), .B2(n6397), .A(n6030), .ZN(n6031) );
  XNOR2_X1 U7534 ( .A(n6033), .B(n6031), .ZN(n7559) );
  INV_X1 U7535 ( .A(n6031), .ZN(n6032) );
  NAND2_X1 U7536 ( .A1(n6785), .A2(n8850), .ZN(n6046) );
  NOR2_X1 U7537 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6037) );
  NAND4_X1 U7538 ( .A1(n6037), .A2(n6036), .A3(n6035), .A4(n6034), .ZN(n6038)
         );
  NAND2_X1 U7539 ( .A1(n6042), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6041) );
  INV_X1 U7540 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6040) );
  MUX2_X1 U7541 ( .A(n6041), .B(P1_IR_REG_31__SCAN_IN), .S(n6040), .Z(n6043)
         );
  NAND2_X1 U7542 ( .A1(n6043), .A2(n6127), .ZN(n6955) );
  OAI22_X1 U7543 ( .A1(n6190), .A2(n6788), .B1(n6521), .B2(n6955), .ZN(n6044)
         );
  INV_X1 U7544 ( .A(n6044), .ZN(n6045) );
  NAND2_X1 U7545 ( .A1(n7745), .A2(n5792), .ZN(n6056) );
  NAND2_X1 U7546 ( .A1(n5921), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6054) );
  INV_X1 U7547 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6047) );
  OR2_X1 U7548 ( .A1(n5852), .A2(n6047), .ZN(n6053) );
  NAND2_X1 U7549 ( .A1(n6049), .A2(n6048), .ZN(n6050) );
  NAND2_X1 U7550 ( .A1(n6070), .A2(n6050), .ZN(n7741) );
  OR2_X1 U7551 ( .A1(n6405), .A2(n7741), .ZN(n6052) );
  INV_X1 U7552 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6566) );
  OR2_X1 U7553 ( .A1(n8840), .A2(n6566), .ZN(n6051) );
  NAND4_X1 U7554 ( .A1(n6054), .A2(n6053), .A3(n6052), .A4(n6051), .ZN(n9133)
         );
  NAND2_X1 U7555 ( .A1(n9133), .A2(n6397), .ZN(n6055) );
  NAND2_X1 U7556 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  XNOR2_X1 U7557 ( .A(n6057), .B(n6309), .ZN(n6059) );
  AND2_X1 U7558 ( .A1(n5808), .A2(n9133), .ZN(n6058) );
  AOI21_X1 U7559 ( .B1(n7745), .B2(n6397), .A(n6058), .ZN(n6060) );
  NAND2_X1 U7560 ( .A1(n6059), .A2(n6060), .ZN(n6064) );
  INV_X1 U7561 ( .A(n6059), .ZN(n6062) );
  INV_X1 U7562 ( .A(n6060), .ZN(n6061) );
  NAND2_X1 U7563 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  NAND2_X1 U7564 ( .A1(n6064), .A2(n6063), .ZN(n7739) );
  NAND2_X1 U7565 ( .A1(n6824), .A2(n8850), .ZN(n6068) );
  NAND2_X1 U7566 ( .A1(n6127), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6065) );
  XNOR2_X1 U7567 ( .A(n6065), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6569) );
  INV_X1 U7568 ( .A(n6569), .ZN(n7070) );
  OAI22_X1 U7569 ( .A1(n6190), .A2(n10321), .B1(n6521), .B2(n7070), .ZN(n6066)
         );
  INV_X1 U7570 ( .A(n6066), .ZN(n6067) );
  NAND2_X1 U7571 ( .A1(n9486), .A2(n6398), .ZN(n6077) );
  NAND2_X1 U7572 ( .A1(n6194), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6075) );
  INV_X1 U7573 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6568) );
  OR2_X1 U7574 ( .A1(n8840), .A2(n6568), .ZN(n6074) );
  INV_X1 U7575 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6542) );
  OR2_X1 U7576 ( .A1(n5866), .A2(n6542), .ZN(n6073) );
  NAND2_X1 U7577 ( .A1(n6070), .A2(n6069), .ZN(n6071) );
  NAND2_X1 U7578 ( .A1(n6089), .A2(n6071), .ZN(n7728) );
  OR2_X1 U7579 ( .A1(n6405), .A2(n7728), .ZN(n6072) );
  NAND4_X1 U7580 ( .A1(n6075), .A2(n6074), .A3(n6073), .A4(n6072), .ZN(n9132)
         );
  NAND2_X1 U7581 ( .A1(n9132), .A2(n6397), .ZN(n6076) );
  NAND2_X1 U7582 ( .A1(n6077), .A2(n6076), .ZN(n6078) );
  XNOR2_X1 U7583 ( .A(n6078), .B(n6309), .ZN(n6080) );
  AND2_X1 U7584 ( .A1(n5808), .A2(n9132), .ZN(n6079) );
  AOI21_X1 U7585 ( .B1(n9486), .B2(n6397), .A(n6079), .ZN(n6081) );
  AND2_X1 U7586 ( .A1(n6080), .A2(n6081), .ZN(n7723) );
  INV_X1 U7587 ( .A(n6080), .ZN(n6083) );
  INV_X1 U7588 ( .A(n6081), .ZN(n6082) );
  NAND2_X1 U7589 ( .A1(n6083), .A2(n6082), .ZN(n7724) );
  NAND2_X1 U7590 ( .A1(n6834), .A2(n8850), .ZN(n6087) );
  OAI21_X1 U7591 ( .B1(n6127), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6084) );
  INV_X1 U7592 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10379) );
  OR2_X1 U7593 ( .A1(n6084), .A2(n10379), .ZN(n6085) );
  NAND2_X1 U7594 ( .A1(n6084), .A2(n10379), .ZN(n6101) );
  AOI22_X1 U7595 ( .A1(n5845), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5846), .B2(
        n7389), .ZN(n6086) );
  NAND2_X1 U7596 ( .A1(n8875), .A2(n6398), .ZN(n6098) );
  INV_X1 U7597 ( .A(n6405), .ZN(n6108) );
  AND2_X1 U7598 ( .A1(n6089), .A2(n6088), .ZN(n6090) );
  NOR2_X1 U7599 ( .A1(n6106), .A2(n6090), .ZN(n7635) );
  NAND2_X1 U7600 ( .A1(n6108), .A2(n7635), .ZN(n6096) );
  INV_X1 U7601 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6091) );
  OR2_X1 U7602 ( .A1(n5866), .A2(n6091), .ZN(n6095) );
  INV_X1 U7603 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6092) );
  OR2_X1 U7604 ( .A1(n5852), .A2(n6092), .ZN(n6094) );
  INV_X1 U7605 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6551) );
  OR2_X1 U7606 ( .A1(n8840), .A2(n6551), .ZN(n6093) );
  NAND4_X1 U7607 ( .A1(n6096), .A2(n6095), .A3(n6094), .A4(n6093), .ZN(n9131)
         );
  NAND2_X1 U7608 ( .A1(n9131), .A2(n6397), .ZN(n6097) );
  NAND2_X1 U7609 ( .A1(n6098), .A2(n6097), .ZN(n6099) );
  XNOR2_X1 U7610 ( .A(n6099), .B(n6309), .ZN(n6118) );
  INV_X1 U7611 ( .A(n6118), .ZN(n6100) );
  NAND2_X1 U7612 ( .A1(n6982), .A2(n8850), .ZN(n6105) );
  NAND2_X1 U7613 ( .A1(n6101), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6102) );
  INV_X1 U7614 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6128) );
  XNOR2_X1 U7615 ( .A(n6102), .B(n6128), .ZN(n7682) );
  OAI22_X1 U7616 ( .A1(n7682), .A2(n6521), .B1(n6190), .B2(n10097), .ZN(n6103)
         );
  INV_X1 U7617 ( .A(n6103), .ZN(n6104) );
  NAND2_X1 U7618 ( .A1(n9606), .A2(n6398), .ZN(n6114) );
  NOR2_X1 U7619 ( .A1(n6106), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6107) );
  OR2_X1 U7620 ( .A1(n6135), .A2(n6107), .ZN(n8821) );
  INV_X1 U7621 ( .A(n8821), .ZN(n7856) );
  NAND2_X1 U7622 ( .A1(n7856), .A2(n6108), .ZN(n6112) );
  NAND2_X1 U7623 ( .A1(n5921), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7624 ( .A1(n6194), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7625 ( .A1(n6323), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6109) );
  NAND4_X1 U7626 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n9130)
         );
  NAND2_X1 U7627 ( .A1(n9130), .A2(n6397), .ZN(n6113) );
  NAND2_X1 U7628 ( .A1(n6114), .A2(n6113), .ZN(n6115) );
  XNOR2_X1 U7629 ( .A(n6115), .B(n6887), .ZN(n6124) );
  INV_X1 U7630 ( .A(n6124), .ZN(n6116) );
  NAND2_X1 U7631 ( .A1(n8875), .A2(n6397), .ZN(n6120) );
  NAND2_X1 U7632 ( .A1(n5808), .A2(n9131), .ZN(n6119) );
  NAND2_X1 U7633 ( .A1(n6120), .A2(n6119), .ZN(n8701) );
  NAND2_X1 U7634 ( .A1(n9606), .A2(n6397), .ZN(n6122) );
  NAND2_X1 U7635 ( .A1(n5808), .A2(n9130), .ZN(n6121) );
  NAND2_X1 U7636 ( .A1(n6122), .A2(n6121), .ZN(n8819) );
  NAND2_X1 U7637 ( .A1(n6123), .A2(n8699), .ZN(n6125) );
  NAND2_X1 U7638 ( .A1(n6125), .A2(n6124), .ZN(n8817) );
  NAND2_X1 U7639 ( .A1(n6126), .A2(n8817), .ZN(n8743) );
  NAND2_X1 U7640 ( .A1(n6985), .A2(n8850), .ZN(n6134) );
  INV_X1 U7641 ( .A(n6127), .ZN(n6131) );
  INV_X1 U7642 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6129) );
  AND3_X1 U7643 ( .A1(n6129), .A2(n6128), .A3(n10379), .ZN(n6130) );
  NAND2_X1 U7644 ( .A1(n6131), .A2(n6130), .ZN(n6148) );
  NAND2_X1 U7645 ( .A1(n6148), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6132) );
  XNOR2_X1 U7646 ( .A(n6132), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7702) );
  AOI22_X1 U7647 ( .A1(n4474), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5846), .B2(
        n7702), .ZN(n6133) );
  NAND2_X1 U7648 ( .A1(n9173), .A2(n6398), .ZN(n6142) );
  NOR2_X1 U7649 ( .A1(n6135), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6136) );
  OR2_X1 U7650 ( .A1(n6156), .A2(n6136), .ZN(n8745) );
  NAND2_X1 U7651 ( .A1(n5921), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7652 ( .A1(n6194), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6137) );
  AND2_X1 U7653 ( .A1(n6138), .A2(n6137), .ZN(n6140) );
  NAND2_X1 U7654 ( .A1(n6323), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6139) );
  OAI211_X1 U7655 ( .C1(n8745), .C2(n6405), .A(n6140), .B(n6139), .ZN(n9402)
         );
  NAND2_X1 U7656 ( .A1(n9402), .A2(n6397), .ZN(n6141) );
  NAND2_X1 U7657 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  XNOR2_X1 U7658 ( .A(n6143), .B(n6309), .ZN(n6146) );
  AND2_X1 U7659 ( .A1(n9402), .A2(n5808), .ZN(n6144) );
  AOI21_X1 U7660 ( .B1(n9173), .B2(n6397), .A(n6144), .ZN(n6145) );
  XNOR2_X1 U7661 ( .A(n6146), .B(n6145), .ZN(n8744) );
  NAND2_X1 U7662 ( .A1(n6146), .A2(n6145), .ZN(n6147) );
  NAND2_X1 U7663 ( .A1(n7064), .A2(n8850), .ZN(n6155) );
  INV_X1 U7664 ( .A(n6148), .ZN(n6150) );
  INV_X1 U7665 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7666 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  NAND2_X1 U7667 ( .A1(n6151), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6152) );
  INV_X1 U7668 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10294) );
  NAND2_X1 U7669 ( .A1(n6152), .A2(n10294), .ZN(n6169) );
  OR2_X1 U7670 ( .A1(n6152), .A2(n10294), .ZN(n6153) );
  AOI22_X1 U7671 ( .A1(n5845), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9145), .B2(
        n5846), .ZN(n6154) );
  NAND2_X1 U7672 ( .A1(n9480), .A2(n5792), .ZN(n6161) );
  OR2_X1 U7673 ( .A1(n6156), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7674 ( .A1(n6157), .A2(n6175), .ZN(n9393) );
  AOI22_X1 U7675 ( .A1(n6323), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n5921), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7676 ( .A1(n6194), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6158) );
  OAI211_X1 U7677 ( .C1(n9393), .C2(n6405), .A(n6159), .B(n6158), .ZN(n9376)
         );
  NAND2_X1 U7678 ( .A1(n9376), .A2(n6397), .ZN(n6160) );
  NAND2_X1 U7679 ( .A1(n6161), .A2(n6160), .ZN(n6162) );
  XNOR2_X1 U7680 ( .A(n6162), .B(n6887), .ZN(n6164) );
  AND2_X1 U7681 ( .A1(n9376), .A2(n5808), .ZN(n6163) );
  AOI21_X1 U7682 ( .B1(n9480), .B2(n6397), .A(n6163), .ZN(n6165) );
  XNOR2_X1 U7683 ( .A(n6164), .B(n6165), .ZN(n8751) );
  INV_X1 U7684 ( .A(n6164), .ZN(n6166) );
  NAND2_X1 U7685 ( .A1(n6166), .A2(n6165), .ZN(n6167) );
  NAND2_X1 U7686 ( .A1(n7210), .A2(n8850), .ZN(n6173) );
  NAND2_X1 U7687 ( .A1(n6169), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6170) );
  XNOR2_X1 U7688 ( .A(n6170), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9148) );
  INV_X1 U7689 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10149) );
  NOR2_X1 U7690 ( .A1(n6190), .A2(n10149), .ZN(n6171) );
  AOI21_X1 U7691 ( .B1(n9148), .B2(n5846), .A(n6171), .ZN(n6172) );
  NAND2_X1 U7692 ( .A1(n9475), .A2(n6398), .ZN(n6184) );
  NAND2_X1 U7693 ( .A1(n5921), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6182) );
  INV_X1 U7694 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9143) );
  OR2_X1 U7695 ( .A1(n8840), .A2(n9143), .ZN(n6181) );
  INV_X1 U7696 ( .A(n6174), .ZN(n6198) );
  INV_X1 U7697 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7698 ( .A1(n6176), .A2(n6175), .ZN(n6177) );
  NAND2_X1 U7699 ( .A1(n6198), .A2(n6177), .ZN(n9380) );
  OR2_X1 U7700 ( .A1(n6405), .A2(n9380), .ZN(n6180) );
  INV_X1 U7701 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n6178) );
  OR2_X1 U7702 ( .A1(n5852), .A2(n6178), .ZN(n6179) );
  NAND4_X1 U7703 ( .A1(n6182), .A2(n6181), .A3(n6180), .A4(n6179), .ZN(n9401)
         );
  NAND2_X1 U7704 ( .A1(n9401), .A2(n6397), .ZN(n6183) );
  NAND2_X1 U7705 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  XNOR2_X1 U7706 ( .A(n6185), .B(n6309), .ZN(n6188) );
  NAND2_X1 U7707 ( .A1(n9475), .A2(n6397), .ZN(n6187) );
  NAND2_X1 U7708 ( .A1(n5808), .A2(n9401), .ZN(n6186) );
  NAND2_X1 U7709 ( .A1(n6187), .A2(n6186), .ZN(n8799) );
  NAND2_X1 U7710 ( .A1(n7305), .A2(n8850), .ZN(n6193) );
  OAI22_X1 U7711 ( .A1(n6190), .A2(n7308), .B1(n9745), .B2(n6521), .ZN(n6191)
         );
  INV_X1 U7712 ( .A(n6191), .ZN(n6192) );
  NAND2_X1 U7713 ( .A1(n9468), .A2(n6398), .ZN(n6206) );
  NAND2_X1 U7714 ( .A1(n6194), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6204) );
  INV_X1 U7715 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6195) );
  OR2_X1 U7716 ( .A1(n5866), .A2(n6195), .ZN(n6203) );
  INV_X1 U7717 ( .A(n6196), .ZN(n6217) );
  INV_X1 U7718 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7719 ( .A1(n6198), .A2(n6197), .ZN(n6199) );
  NAND2_X1 U7720 ( .A1(n6217), .A2(n6199), .ZN(n9357) );
  OR2_X1 U7721 ( .A1(n6405), .A2(n9357), .ZN(n6202) );
  INV_X1 U7722 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6200) );
  OR2_X1 U7723 ( .A1(n8840), .A2(n6200), .ZN(n6201) );
  NAND4_X1 U7724 ( .A1(n6204), .A2(n6203), .A3(n6202), .A4(n6201), .ZN(n9375)
         );
  NAND2_X1 U7725 ( .A1(n9375), .A2(n6397), .ZN(n6205) );
  NAND2_X1 U7726 ( .A1(n6206), .A2(n6205), .ZN(n6207) );
  XNOR2_X1 U7727 ( .A(n6207), .B(n6887), .ZN(n6209) );
  AND2_X1 U7728 ( .A1(n5808), .A2(n9375), .ZN(n6208) );
  AOI21_X1 U7729 ( .B1(n9468), .B2(n6397), .A(n6208), .ZN(n6210) );
  XNOR2_X1 U7730 ( .A(n6209), .B(n6210), .ZN(n8720) );
  INV_X1 U7731 ( .A(n6209), .ZN(n6211) );
  NAND2_X1 U7732 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  NAND2_X1 U7733 ( .A1(n7426), .A2(n8850), .ZN(n6214) );
  NAND2_X1 U7734 ( .A1(n4474), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7735 ( .A1(n9464), .A2(n6398), .ZN(n6225) );
  NAND2_X1 U7736 ( .A1(n6323), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6223) );
  INV_X1 U7737 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6215) );
  OR2_X1 U7738 ( .A1(n5866), .A2(n6215), .ZN(n6222) );
  INV_X1 U7739 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n6216) );
  OR2_X1 U7740 ( .A1(n5852), .A2(n6216), .ZN(n6221) );
  INV_X1 U7741 ( .A(n6236), .ZN(n6219) );
  INV_X1 U7742 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U7743 ( .A1(n6217), .A2(n8770), .ZN(n6218) );
  NAND2_X1 U7744 ( .A1(n6219), .A2(n6218), .ZN(n9342) );
  OR2_X1 U7745 ( .A1(n6405), .A2(n9342), .ZN(n6220) );
  NAND4_X1 U7746 ( .A1(n6223), .A2(n6222), .A3(n6221), .A4(n6220), .ZN(n9367)
         );
  NAND2_X1 U7747 ( .A1(n9367), .A2(n6397), .ZN(n6224) );
  NAND2_X1 U7748 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  XNOR2_X1 U7749 ( .A(n6226), .B(n6887), .ZN(n6229) );
  NAND2_X1 U7750 ( .A1(n9464), .A2(n6397), .ZN(n6228) );
  NAND2_X1 U7751 ( .A1(n5808), .A2(n9367), .ZN(n6227) );
  NAND2_X1 U7752 ( .A1(n6228), .A2(n6227), .ZN(n6230) );
  NAND2_X1 U7753 ( .A1(n6229), .A2(n6230), .ZN(n8766) );
  INV_X1 U7754 ( .A(n6229), .ZN(n6232) );
  INV_X1 U7755 ( .A(n6230), .ZN(n6231) );
  NAND2_X1 U7756 ( .A1(n6232), .A2(n6231), .ZN(n8767) );
  NAND2_X1 U7757 ( .A1(n7451), .A2(n8850), .ZN(n6234) );
  NAND2_X1 U7758 ( .A1(n5845), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U7759 ( .A1(n9458), .A2(n6398), .ZN(n6243) );
  NAND2_X1 U7760 ( .A1(n5921), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6241) );
  INV_X1 U7761 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n6235) );
  OR2_X1 U7762 ( .A1(n5852), .A2(n6235), .ZN(n6240) );
  OAI21_X1 U7763 ( .B1(n6236), .B2(P1_REG3_REG_21__SCAN_IN), .A(n6254), .ZN(
        n9323) );
  OR2_X1 U7764 ( .A1(n6405), .A2(n9323), .ZN(n6239) );
  INV_X1 U7765 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6237) );
  OR2_X1 U7766 ( .A1(n8840), .A2(n6237), .ZN(n6238) );
  NAND4_X1 U7767 ( .A1(n6241), .A2(n6240), .A3(n6239), .A4(n6238), .ZN(n9349)
         );
  NAND2_X1 U7768 ( .A1(n9349), .A2(n6397), .ZN(n6242) );
  NAND2_X1 U7769 ( .A1(n6243), .A2(n6242), .ZN(n6244) );
  XNOR2_X1 U7770 ( .A(n6244), .B(n6887), .ZN(n6246) );
  AND2_X1 U7771 ( .A1(n5808), .A2(n9349), .ZN(n6245) );
  AOI21_X1 U7772 ( .B1(n9458), .B2(n6397), .A(n6245), .ZN(n6247) );
  XNOR2_X1 U7773 ( .A(n6246), .B(n6247), .ZN(n8726) );
  INV_X1 U7774 ( .A(n6246), .ZN(n6248) );
  NAND2_X1 U7775 ( .A1(n7529), .A2(n8850), .ZN(n6250) );
  NAND2_X1 U7776 ( .A1(n5845), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7777 ( .A1(n5921), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6259) );
  INV_X1 U7778 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6251) );
  OR2_X1 U7779 ( .A1(n8840), .A2(n6251), .ZN(n6258) );
  INV_X1 U7780 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n6252) );
  OR2_X1 U7781 ( .A1(n5852), .A2(n6252), .ZN(n6257) );
  AOI21_X1 U7782 ( .B1(n6254), .B2(n8782), .A(n6253), .ZN(n9310) );
  INV_X1 U7783 ( .A(n9310), .ZN(n6255) );
  OR2_X1 U7784 ( .A1(n6405), .A2(n6255), .ZN(n6256) );
  NAND4_X1 U7785 ( .A1(n6259), .A2(n6258), .A3(n6257), .A4(n6256), .ZN(n9330)
         );
  AND2_X1 U7786 ( .A1(n5808), .A2(n9330), .ZN(n6260) );
  AOI21_X1 U7787 ( .B1(n9451), .B2(n6397), .A(n6260), .ZN(n6265) );
  NAND2_X1 U7788 ( .A1(n6264), .A2(n6265), .ZN(n8776) );
  NAND2_X1 U7789 ( .A1(n9451), .A2(n5792), .ZN(n6262) );
  NAND2_X1 U7790 ( .A1(n9330), .A2(n6397), .ZN(n6261) );
  NAND2_X1 U7791 ( .A1(n6262), .A2(n6261), .ZN(n6263) );
  XNOR2_X1 U7792 ( .A(n6263), .B(n6887), .ZN(n8777) );
  INV_X1 U7793 ( .A(n6265), .ZN(n6266) );
  AOI22_X1 U7794 ( .A1(n9447), .A2(n6398), .B1(n6397), .B2(n9316), .ZN(n6268)
         );
  XOR2_X1 U7795 ( .A(n6887), .B(n6268), .Z(n6269) );
  NAND2_X1 U7796 ( .A1(n7641), .A2(n8850), .ZN(n6272) );
  NAND2_X1 U7797 ( .A1(n5845), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7798 ( .A1(n5921), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6281) );
  INV_X1 U7799 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6273) );
  OR2_X1 U7800 ( .A1(n5852), .A2(n6273), .ZN(n6280) );
  INV_X1 U7801 ( .A(n6274), .ZN(n6276) );
  INV_X1 U7802 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8761) );
  INV_X1 U7803 ( .A(n6289), .ZN(n6275) );
  OAI21_X1 U7804 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n6276), .A(n6275), .ZN(
        n9289) );
  OR2_X1 U7805 ( .A1(n6405), .A2(n9289), .ZN(n6279) );
  INV_X1 U7806 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6277) );
  OR2_X1 U7807 ( .A1(n8840), .A2(n6277), .ZN(n6278) );
  NAND4_X1 U7808 ( .A1(n6281), .A2(n6280), .A3(n6279), .A4(n6278), .ZN(n9303)
         );
  AOI22_X1 U7809 ( .A1(n9442), .A2(n6398), .B1(n6397), .B2(n9303), .ZN(n6282)
         );
  XNOR2_X1 U7810 ( .A(n6282), .B(n6887), .ZN(n6284) );
  AOI22_X1 U7811 ( .A1(n9442), .A2(n6397), .B1(n5808), .B2(n9303), .ZN(n6283)
         );
  NAND2_X1 U7812 ( .A1(n6284), .A2(n6283), .ZN(n6285) );
  OAI21_X1 U7813 ( .B1(n6284), .B2(n6283), .A(n6285), .ZN(n8759) );
  NAND2_X1 U7814 ( .A1(n7813), .A2(n8850), .ZN(n6287) );
  NAND2_X1 U7815 ( .A1(n4474), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6286) );
  NAND2_X2 U7816 ( .A1(n6287), .A2(n6286), .ZN(n9437) );
  NAND2_X1 U7817 ( .A1(n6323), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6294) );
  INV_X1 U7818 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6288) );
  OR2_X1 U7819 ( .A1(n5866), .A2(n6288), .ZN(n6293) );
  NAND2_X1 U7820 ( .A1(n6289), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6300) );
  OAI21_X1 U7821 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n6289), .A(n6300), .ZN(
        n8736) );
  OR2_X1 U7822 ( .A1(n6405), .A2(n8736), .ZN(n6292) );
  INV_X1 U7823 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n6290) );
  OR2_X1 U7824 ( .A1(n5852), .A2(n6290), .ZN(n6291) );
  NAND4_X1 U7825 ( .A1(n6294), .A2(n6293), .A3(n6292), .A4(n6291), .ZN(n9286)
         );
  AOI22_X1 U7826 ( .A1(n9437), .A2(n6398), .B1(n6397), .B2(n9286), .ZN(n6295)
         );
  XNOR2_X1 U7827 ( .A(n6295), .B(n6887), .ZN(n6312) );
  AND2_X1 U7828 ( .A1(n5808), .A2(n9286), .ZN(n6296) );
  AOI21_X1 U7829 ( .B1(n9437), .B2(n6397), .A(n6296), .ZN(n6313) );
  XNOR2_X1 U7830 ( .A(n6312), .B(n6313), .ZN(n8733) );
  NAND2_X1 U7831 ( .A1(n7817), .A2(n8850), .ZN(n6298) );
  NAND2_X1 U7832 ( .A1(n4474), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U7833 ( .A1(n9432), .A2(n5792), .ZN(n6308) );
  NAND2_X1 U7834 ( .A1(n5921), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6306) );
  INV_X1 U7835 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6299) );
  OR2_X1 U7836 ( .A1(n5852), .A2(n6299), .ZN(n6305) );
  OAI21_X1 U7837 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n6301), .A(n6368), .ZN(
        n8809) );
  OR2_X1 U7838 ( .A1(n6405), .A2(n8809), .ZN(n6304) );
  INV_X1 U7839 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7840 ( .A1(n9277), .A2(n6397), .ZN(n6307) );
  NAND2_X1 U7841 ( .A1(n6308), .A2(n6307), .ZN(n6310) );
  XNOR2_X1 U7842 ( .A(n6310), .B(n6309), .ZN(n6317) );
  AND2_X1 U7843 ( .A1(n5808), .A2(n9277), .ZN(n6311) );
  AOI21_X1 U7844 ( .B1(n9432), .B2(n6397), .A(n6311), .ZN(n6318) );
  XNOR2_X1 U7845 ( .A(n6317), .B(n6318), .ZN(n8805) );
  INV_X1 U7846 ( .A(n6312), .ZN(n6315) );
  INV_X1 U7847 ( .A(n6313), .ZN(n6314) );
  NOR2_X1 U7848 ( .A1(n6315), .A2(n6314), .ZN(n8806) );
  INV_X1 U7849 ( .A(n6317), .ZN(n6320) );
  INV_X1 U7850 ( .A(n6318), .ZN(n6319) );
  NAND2_X1 U7851 ( .A1(n9519), .A2(n8850), .ZN(n6322) );
  NAND2_X1 U7852 ( .A1(n5845), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U7853 ( .A1(n6323), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6329) );
  INV_X1 U7854 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6324) );
  OR2_X1 U7855 ( .A1(n5866), .A2(n6324), .ZN(n6328) );
  INV_X1 U7856 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6367) );
  XNOR2_X1 U7857 ( .A(n6368), .B(n6367), .ZN(n6376) );
  OR2_X1 U7858 ( .A1(n6405), .A2(n6376), .ZN(n6327) );
  INV_X1 U7859 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6325) );
  OR2_X1 U7860 ( .A1(n5852), .A2(n6325), .ZN(n6326) );
  AOI22_X1 U7861 ( .A1(n9426), .A2(n6398), .B1(n6397), .B2(n9265), .ZN(n6330)
         );
  XNOR2_X1 U7862 ( .A(n6330), .B(n6887), .ZN(n6332) );
  AOI22_X1 U7863 ( .A1(n9426), .A2(n6397), .B1(n5808), .B2(n9265), .ZN(n6331)
         );
  NAND2_X1 U7864 ( .A1(n6332), .A2(n6331), .ZN(n6413) );
  OAI21_X1 U7865 ( .B1(n6332), .B2(n6331), .A(n6413), .ZN(n6334) );
  NAND3_X1 U7866 ( .A1(n7642), .A2(P1_B_REG_SCAN_IN), .A3(n6336), .ZN(n6340)
         );
  INV_X1 U7867 ( .A(n7642), .ZN(n6338) );
  INV_X1 U7868 ( .A(P1_B_REG_SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7869 ( .A1(n6338), .A2(n6337), .ZN(n6339) );
  INV_X1 U7870 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6342) );
  INV_X1 U7871 ( .A(n6335), .ZN(n7818) );
  AND2_X1 U7872 ( .A1(n7818), .A2(n7642), .ZN(n6341) );
  NOR4_X1 U7873 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6351) );
  NOR4_X1 U7874 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6350) );
  OR4_X1 U7875 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6348) );
  NOR4_X1 U7876 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6346) );
  NOR4_X1 U7877 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6345) );
  NOR4_X1 U7878 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6344) );
  NOR4_X1 U7879 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6343) );
  NAND4_X1 U7880 ( .A1(n6346), .A2(n6345), .A3(n6344), .A4(n6343), .ZN(n6347)
         );
  NOR4_X1 U7881 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6348), .A4(n6347), .ZN(n6349) );
  NAND3_X1 U7882 ( .A1(n6351), .A2(n6350), .A3(n6349), .ZN(n6352) );
  NAND2_X1 U7883 ( .A1(n9755), .A2(n6352), .ZN(n6772) );
  INV_X1 U7884 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6354) );
  AND2_X1 U7885 ( .A1(n7818), .A2(n6336), .ZN(n6353) );
  NAND2_X1 U7886 ( .A1(n6781), .A2(n6877), .ZN(n6803) );
  INV_X1 U7887 ( .A(n6355), .ZN(n6356) );
  NAND2_X1 U7888 ( .A1(n6356), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6357) );
  XNOR2_X1 U7889 ( .A(n6357), .B(n10072), .ZN(n7587) );
  AND2_X1 U7890 ( .A1(n7587), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6358) );
  NAND2_X1 U7891 ( .A1(n9042), .A2(n9082), .ZN(n6882) );
  NAND2_X1 U7892 ( .A1(n9127), .A2(n4673), .ZN(n6889) );
  NAND2_X1 U7893 ( .A1(n9791), .A2(n6889), .ZN(n6377) );
  INV_X1 U7894 ( .A(n6362), .ZN(n6359) );
  INV_X1 U7895 ( .A(n6882), .ZN(n6777) );
  AND2_X1 U7896 ( .A1(n6777), .A2(n9122), .ZN(n9738) );
  NAND2_X1 U7897 ( .A1(n6359), .A2(n9738), .ZN(n6360) );
  OR2_X1 U7898 ( .A1(n9030), .A2(n9122), .ZN(n9490) );
  NAND2_X2 U7899 ( .A1(n6360), .A2(n9743), .ZN(n8828) );
  NAND2_X1 U7900 ( .A1(n9426), .A2(n8828), .ZN(n6390) );
  OR2_X1 U7901 ( .A1(n6361), .A2(n6879), .ZN(n6888) );
  OR2_X1 U7902 ( .A1(n6362), .A2(n6888), .ZN(n6386) );
  INV_X1 U7903 ( .A(n9632), .ZN(n9124) );
  NOR2_X2 U7904 ( .A1(n6386), .A2(n9124), .ZN(n8811) );
  NAND2_X1 U7905 ( .A1(n5921), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6375) );
  INV_X1 U7906 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6364) );
  OR2_X1 U7907 ( .A1(n8840), .A2(n6364), .ZN(n6374) );
  INV_X1 U7908 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6365) );
  OR2_X1 U7909 ( .A1(n5852), .A2(n6365), .ZN(n6373) );
  INV_X1 U7910 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6366) );
  OAI21_X1 U7911 ( .B1(n6368), .B2(n6367), .A(n6366), .ZN(n6371) );
  INV_X1 U7912 ( .A(n6368), .ZN(n6370) );
  AND2_X1 U7913 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6369) );
  NAND2_X1 U7914 ( .A1(n6370), .A2(n6369), .ZN(n9220) );
  NAND2_X1 U7915 ( .A1(n6371), .A2(n9220), .ZN(n9237) );
  OR2_X1 U7916 ( .A1(n6405), .A2(n9237), .ZN(n6372) );
  NAND4_X1 U7917 ( .A1(n6375), .A2(n6374), .A3(n6373), .A4(n6372), .ZN(n9250)
         );
  INV_X1 U7918 ( .A(n6376), .ZN(n9245) );
  INV_X1 U7919 ( .A(n6377), .ZN(n6380) );
  NAND3_X1 U7920 ( .A1(n5797), .A2(n7587), .A3(n6779), .ZN(n6379) );
  AOI21_X1 U7921 ( .B1(n6803), .B2(n6380), .A(n6379), .ZN(n6381) );
  OR2_X1 U7922 ( .A1(n6381), .A2(P1_U3084), .ZN(n6385) );
  INV_X1 U7923 ( .A(n9738), .ZN(n6382) );
  AND2_X1 U7924 ( .A1(n6382), .A2(n6888), .ZN(n6383) );
  NOR2_X1 U7925 ( .A1(n9754), .A2(n6383), .ZN(n6384) );
  NAND2_X1 U7926 ( .A1(n6803), .A2(n6384), .ZN(n6804) );
  NAND2_X1 U7927 ( .A1(n6385), .A2(n6804), .ZN(n8810) );
  AOI22_X1 U7928 ( .A1(n8811), .A2(n9250), .B1(n9245), .B2(n8810), .ZN(n6388)
         );
  AOI22_X1 U7929 ( .A1(n4473), .A2(n9277), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n6387) );
  AND2_X1 U7930 ( .A1(n6388), .A2(n6387), .ZN(n6389) );
  NAND3_X1 U7931 ( .A1(n6391), .A2(n6390), .A3(n6389), .ZN(P1_U3212) );
  NAND2_X1 U7932 ( .A1(n9515), .A2(n8850), .ZN(n6393) );
  NAND2_X1 U7933 ( .A1(n4474), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U7934 ( .A1(n9422), .A2(n6397), .ZN(n6395) );
  NAND2_X1 U7935 ( .A1(n5808), .A2(n9250), .ZN(n6394) );
  NAND2_X1 U7936 ( .A1(n6395), .A2(n6394), .ZN(n6396) );
  XNOR2_X1 U7937 ( .A(n6396), .B(n6887), .ZN(n6400) );
  AOI22_X1 U7938 ( .A1(n9422), .A2(n6398), .B1(n6397), .B2(n9250), .ZN(n6399)
         );
  XNOR2_X1 U7939 ( .A(n6400), .B(n6399), .ZN(n6402) );
  INV_X1 U7940 ( .A(n6402), .ZN(n6414) );
  NAND3_X1 U7941 ( .A1(n6414), .A2(n8808), .A3(n6413), .ZN(n6401) );
  NAND3_X1 U7942 ( .A1(n6403), .A2(n6402), .A3(n8808), .ZN(n6418) );
  NAND2_X1 U7943 ( .A1(n5921), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6410) );
  INV_X1 U7944 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6404) );
  OR2_X1 U7945 ( .A1(n8840), .A2(n6404), .ZN(n6409) );
  OR2_X1 U7946 ( .A1(n6405), .A2(n9220), .ZN(n6408) );
  INV_X1 U7947 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6406) );
  OR2_X1 U7948 ( .A1(n5852), .A2(n6406), .ZN(n6407) );
  NAND4_X1 U7949 ( .A1(n6410), .A2(n6409), .A3(n6408), .A4(n6407), .ZN(n9234)
         );
  AOI22_X1 U7950 ( .A1(n8811), .A2(n9234), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6412) );
  NAND2_X1 U7951 ( .A1(n4473), .A2(n9265), .ZN(n6411) );
  OAI211_X1 U7952 ( .C1(n8822), .C2(n9237), .A(n6412), .B(n6411), .ZN(n6416)
         );
  NOR3_X1 U7953 ( .A1(n6414), .A2(n8831), .A3(n6413), .ZN(n6415) );
  AOI211_X1 U7954 ( .C1(n9422), .C2(n8828), .A(n6416), .B(n6415), .ZN(n6417)
         );
  NAND3_X1 U7955 ( .A1(n6419), .A2(n6418), .A3(n6417), .ZN(P1_U3218) );
  INV_X1 U7956 ( .A(n8614), .ZN(n6453) );
  INV_X1 U7957 ( .A(n8257), .ZN(n8200) );
  INV_X1 U7958 ( .A(n7824), .ZN(n8260) );
  INV_X1 U7959 ( .A(n6420), .ZN(n8274) );
  NAND2_X1 U7960 ( .A1(n7040), .A2(n6421), .ZN(n6424) );
  NAND2_X1 U7961 ( .A1(n6420), .A2(n6422), .ZN(n6423) );
  NAND2_X1 U7962 ( .A1(n6424), .A2(n6423), .ZN(n7052) );
  INV_X1 U7963 ( .A(n7046), .ZN(n8273) );
  INV_X1 U7964 ( .A(n7057), .ZN(n9912) );
  NAND2_X1 U7965 ( .A1(n7046), .A2(n7057), .ZN(n7938) );
  NAND2_X1 U7966 ( .A1(n7940), .A2(n7938), .ZN(n7905) );
  NAND2_X1 U7967 ( .A1(n7052), .A2(n7905), .ZN(n6426) );
  NAND2_X1 U7968 ( .A1(n7046), .A2(n9912), .ZN(n6425) );
  NAND2_X1 U7969 ( .A1(n6426), .A2(n6425), .ZN(n7087) );
  NAND2_X1 U7970 ( .A1(n9813), .A2(n9917), .ZN(n7924) );
  INV_X1 U7971 ( .A(n9813), .ZN(n8272) );
  INV_X1 U7972 ( .A(n9917), .ZN(n6427) );
  NAND2_X1 U7973 ( .A1(n8272), .A2(n6427), .ZN(n7949) );
  NAND2_X1 U7974 ( .A1(n7087), .A2(n7944), .ZN(n6429) );
  NAND2_X1 U7975 ( .A1(n9813), .A2(n6427), .ZN(n6428) );
  NAND2_X1 U7976 ( .A1(n6429), .A2(n6428), .ZN(n7268) );
  NAND2_X1 U7977 ( .A1(n7168), .A2(n6430), .ZN(n7273) );
  NAND2_X1 U7978 ( .A1(n8271), .A2(n9929), .ZN(n7274) );
  NAND2_X1 U7979 ( .A1(n7273), .A2(n7274), .ZN(n9840) );
  NAND2_X1 U7980 ( .A1(n8270), .A2(n7283), .ZN(n6431) );
  AND2_X1 U7981 ( .A1(n9840), .A2(n6431), .ZN(n6435) );
  INV_X1 U7982 ( .A(n6431), .ZN(n6434) );
  NAND2_X1 U7983 ( .A1(n7168), .A2(n9929), .ZN(n7269) );
  OR2_X1 U7984 ( .A1(n8270), .A2(n7283), .ZN(n6432) );
  AND2_X1 U7985 ( .A1(n7269), .A2(n6432), .ZN(n6433) );
  NAND2_X1 U7986 ( .A1(n7261), .A2(n7312), .ZN(n7958) );
  INV_X1 U7987 ( .A(n7261), .ZN(n8269) );
  INV_X1 U7988 ( .A(n7312), .ZN(n7325) );
  NAND2_X1 U7989 ( .A1(n8269), .A2(n7325), .ZN(n7948) );
  NAND2_X1 U7990 ( .A1(n7958), .A2(n7948), .ZN(n7226) );
  NAND2_X1 U7991 ( .A1(n7223), .A2(n7226), .ZN(n6437) );
  NAND2_X1 U7992 ( .A1(n8269), .A2(n7312), .ZN(n6436) );
  NAND2_X1 U7993 ( .A1(n7345), .A2(n7255), .ZN(n7959) );
  INV_X1 U7994 ( .A(n7345), .ZN(n8268) );
  INV_X1 U7995 ( .A(n7255), .ZN(n7411) );
  NAND2_X1 U7996 ( .A1(n8268), .A2(n7411), .ZN(n7960) );
  INV_X1 U7997 ( .A(n7367), .ZN(n8267) );
  AND2_X1 U7998 ( .A1(n8267), .A2(n7421), .ZN(n6440) );
  OR2_X1 U7999 ( .A1(n7957), .A2(n6440), .ZN(n6438) );
  NAND2_X1 U8000 ( .A1(n7345), .A2(n7411), .ZN(n7350) );
  NAND2_X1 U8001 ( .A1(n7367), .A2(n7421), .ZN(n7964) );
  NAND2_X1 U8002 ( .A1(n8267), .A2(n7500), .ZN(n7963) );
  INV_X1 U8003 ( .A(n7962), .ZN(n6439) );
  NAND2_X1 U8004 ( .A1(n7472), .A2(n7377), .ZN(n7969) );
  INV_X1 U8005 ( .A(n7472), .ZN(n8266) );
  NAND2_X1 U8006 ( .A1(n8266), .A2(n9933), .ZN(n7468) );
  NAND2_X1 U8007 ( .A1(n7969), .A2(n7468), .ZN(n7910) );
  NAND2_X1 U8008 ( .A1(n7472), .A2(n9933), .ZN(n6441) );
  NAND2_X1 U8009 ( .A1(n7363), .A2(n6441), .ZN(n7465) );
  NAND2_X1 U8010 ( .A1(n7617), .A2(n8265), .ZN(n6479) );
  INV_X1 U8011 ( .A(n8265), .ZN(n6442) );
  NAND2_X1 U8012 ( .A1(n6442), .A2(n7481), .ZN(n7971) );
  NAND2_X1 U8013 ( .A1(n7481), .A2(n8265), .ZN(n6444) );
  OR2_X1 U8014 ( .A1(n7523), .A2(n7535), .ZN(n7972) );
  NAND2_X1 U8015 ( .A1(n7523), .A2(n7535), .ZN(n7981) );
  NAND2_X1 U8016 ( .A1(n7972), .A2(n7981), .ZN(n7514) );
  INV_X1 U8017 ( .A(n7535), .ZN(n8264) );
  NAND2_X1 U8018 ( .A1(n7523), .A2(n8264), .ZN(n6445) );
  NAND2_X1 U8019 ( .A1(n6446), .A2(n6445), .ZN(n7540) );
  OR2_X1 U8020 ( .A1(n7771), .A2(n7709), .ZN(n7983) );
  NAND2_X1 U8021 ( .A1(n7771), .A2(n7709), .ZN(n7982) );
  INV_X1 U8022 ( .A(n7709), .ZN(n8263) );
  NAND2_X1 U8023 ( .A1(n7720), .A2(n7753), .ZN(n7990) );
  OR2_X1 U8024 ( .A1(n7720), .A2(n7753), .ZN(n6447) );
  INV_X1 U8025 ( .A(n7753), .ZN(n8262) );
  NAND2_X1 U8026 ( .A1(n7720), .A2(n8262), .ZN(n6448) );
  OR2_X1 U8027 ( .A1(n8120), .A2(n7823), .ZN(n7991) );
  NAND2_X1 U8028 ( .A1(n8120), .A2(n7823), .ZN(n7992) );
  INV_X1 U8030 ( .A(n7823), .ZN(n8261) );
  OR2_X1 U8031 ( .A1(n8245), .A2(n8170), .ZN(n7997) );
  NAND2_X1 U8032 ( .A1(n8245), .A2(n8170), .ZN(n7996) );
  NAND2_X1 U8033 ( .A1(n7997), .A2(n7996), .ZN(n7903) );
  NAND2_X1 U8034 ( .A1(n7820), .A2(n7903), .ZN(n7819) );
  NAND2_X1 U8035 ( .A1(n4703), .A2(n8170), .ZN(n6449) );
  NAND2_X1 U8036 ( .A1(n7819), .A2(n6449), .ZN(n8539) );
  OR2_X1 U8037 ( .A1(n8550), .A2(n7824), .ZN(n7999) );
  NAND2_X1 U8038 ( .A1(n8550), .A2(n7824), .ZN(n8000) );
  XNOR2_X1 U8039 ( .A(n8535), .B(n8217), .ZN(n8532) );
  INV_X1 U8040 ( .A(n8217), .ZN(n8259) );
  NAND2_X1 U8041 ( .A1(n8514), .A2(n8258), .ZN(n6450) );
  INV_X1 U8042 ( .A(n8258), .ZN(n6482) );
  OR2_X1 U8043 ( .A1(n8614), .A2(n8257), .ZN(n6451) );
  NAND2_X1 U8044 ( .A1(n8493), .A2(n6451), .ZN(n6452) );
  OAI21_X1 U8045 ( .B1(n6453), .B2(n8200), .A(n6452), .ZN(n8485) );
  NAND2_X1 U8046 ( .A1(n8487), .A2(n8146), .ZN(n8014) );
  NAND2_X1 U8047 ( .A1(n8017), .A2(n8014), .ZN(n8480) );
  INV_X1 U8048 ( .A(n8146), .ZN(n8256) );
  NAND2_X1 U8049 ( .A1(n8462), .A2(n6454), .ZN(n6455) );
  NAND2_X1 U8050 ( .A1(n8600), .A2(n8147), .ZN(n8025) );
  NAND2_X1 U8051 ( .A1(n8434), .A2(n8025), .ZN(n6485) );
  INV_X1 U8052 ( .A(n8600), .ZN(n8458) );
  OR2_X1 U8053 ( .A1(n8442), .A2(n8208), .ZN(n8028) );
  NAND2_X1 U8054 ( .A1(n8442), .A2(n8208), .ZN(n8034) );
  NAND2_X1 U8055 ( .A1(n8028), .A2(n8034), .ZN(n8435) );
  NAND2_X1 U8056 ( .A1(n8590), .A2(n8123), .ZN(n8035) );
  OR2_X1 U8057 ( .A1(n8577), .A2(n8157), .ZN(n8042) );
  NAND2_X1 U8058 ( .A1(n8577), .A2(n8157), .ZN(n6488) );
  INV_X1 U8059 ( .A(n8157), .ZN(n8252) );
  NAND2_X1 U8060 ( .A1(n6458), .A2(n6457), .ZN(n8367) );
  NAND2_X1 U8061 ( .A1(n8367), .A2(n8368), .ZN(n6460) );
  NAND2_X1 U8062 ( .A1(n4707), .A2(n8227), .ZN(n6459) );
  NOR2_X1 U8063 ( .A1(n8569), .A2(n8250), .ZN(n6461) );
  INV_X1 U8064 ( .A(n6464), .ZN(n6466) );
  NAND2_X1 U8065 ( .A1(n6466), .A2(n6465), .ZN(n6467) );
  MUX2_X1 U8066 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6469), .Z(n7874) );
  INV_X1 U8067 ( .A(SI_29_), .ZN(n10172) );
  XNOR2_X1 U8068 ( .A(n7874), .B(n10172), .ZN(n7872) );
  NAND2_X1 U8069 ( .A1(n8851), .A2(n7890), .ZN(n6471) );
  INV_X1 U8070 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8687) );
  OR2_X1 U8071 ( .A1(n4476), .A2(n8687), .ZN(n6470) );
  OR2_X1 U8072 ( .A1(n8099), .A2(n6839), .ZN(n8053) );
  NAND2_X1 U8073 ( .A1(n8099), .A2(n6839), .ZN(n8052) );
  NAND2_X1 U8074 ( .A1(n7530), .A2(n6472), .ZN(n6473) );
  NAND4_X1 U8075 ( .A1(n6668), .A2(n9897), .A3(n8530), .A4(n6473), .ZN(n8547)
         );
  AND2_X1 U8076 ( .A1(n8072), .A2(n7923), .ZN(n6474) );
  NAND2_X1 U8077 ( .A1(n7530), .A2(n6474), .ZN(n9921) );
  NAND2_X1 U8078 ( .A1(n7047), .A2(n7053), .ZN(n7045) );
  NAND2_X1 U8079 ( .A1(n7045), .A2(n7934), .ZN(n6476) );
  NAND2_X1 U8080 ( .A1(n6476), .A2(n7933), .ZN(n7058) );
  INV_X1 U8081 ( .A(n7944), .ZN(n7095) );
  NAND2_X1 U8082 ( .A1(n7094), .A2(n7095), .ZN(n7093) );
  NAND2_X1 U8083 ( .A1(n7093), .A2(n7924), .ZN(n7272) );
  INV_X1 U8084 ( .A(n8270), .ZN(n9815) );
  NAND2_X1 U8085 ( .A1(n9815), .A2(n7283), .ZN(n7930) );
  NAND2_X1 U8086 ( .A1(n7273), .A2(n7930), .ZN(n7926) );
  INV_X1 U8087 ( .A(n7930), .ZN(n6477) );
  INV_X1 U8088 ( .A(n7226), .ZN(n7908) );
  INV_X1 U8089 ( .A(n7969), .ZN(n6478) );
  AND2_X1 U8090 ( .A1(n6479), .A2(n7468), .ZN(n7966) );
  AND2_X1 U8091 ( .A1(n7981), .A2(n7971), .ZN(n7967) );
  AND2_X1 U8092 ( .A1(n7983), .A2(n7972), .ZN(n7976) );
  NAND2_X1 U8093 ( .A1(n7708), .A2(n7977), .ZN(n6480) );
  NAND2_X1 U8094 ( .A1(n6480), .A2(n7990), .ZN(n7750) );
  INV_X1 U8095 ( .A(n7989), .ZN(n7751) );
  INV_X1 U8096 ( .A(n7997), .ZN(n6481) );
  OR2_X1 U8097 ( .A1(n8535), .A2(n8217), .ZN(n8002) );
  OAI21_X1 U8098 ( .B1(n8525), .B2(n8532), .A(n8002), .ZN(n8507) );
  NAND2_X1 U8099 ( .A1(n8514), .A2(n6482), .ZN(n8012) );
  OR2_X1 U8100 ( .A1(n8514), .A2(n6482), .ZN(n8007) );
  OR2_X1 U8101 ( .A1(n8614), .A2(n8200), .ZN(n8015) );
  NAND2_X1 U8102 ( .A1(n8614), .A2(n8200), .ZN(n8018) );
  NAND2_X1 U8103 ( .A1(n8015), .A2(n8018), .ZN(n8496) );
  OR2_X1 U8104 ( .A1(n8604), .A2(n8207), .ZN(n8031) );
  NAND2_X1 U8105 ( .A1(n8604), .A2(n8207), .ZN(n8024) );
  NAND2_X1 U8106 ( .A1(n8031), .A2(n8024), .ZN(n8469) );
  INV_X1 U8107 ( .A(n8017), .ZN(n8470) );
  NOR2_X1 U8108 ( .A1(n8469), .A2(n8470), .ZN(n6484) );
  INV_X1 U8109 ( .A(n8434), .ZN(n8026) );
  NOR2_X1 U8110 ( .A1(n8435), .A2(n8026), .ZN(n8033) );
  INV_X1 U8111 ( .A(n8034), .ZN(n6486) );
  AOI21_X1 U8112 ( .B1(n8433), .B2(n8033), .A(n6486), .ZN(n8418) );
  NAND2_X1 U8113 ( .A1(n8418), .A2(n8417), .ZN(n8416) );
  NAND2_X1 U8114 ( .A1(n8416), .A2(n8036), .ZN(n8401) );
  INV_X1 U8115 ( .A(n8253), .ZN(n6487) );
  OR2_X1 U8116 ( .A1(n8410), .A2(n6487), .ZN(n8040) );
  NOR2_X1 U8117 ( .A1(n8377), .A2(n8227), .ZN(n8047) );
  INV_X1 U8118 ( .A(n8051), .ZN(n6490) );
  NAND2_X1 U8119 ( .A1(n8250), .A2(n8228), .ZN(n6500) );
  INV_X1 U8120 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U8121 ( .A1(n6491), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U8122 ( .A1(n6492), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6493) );
  OAI211_X1 U8123 ( .C1(n6495), .C2(n8640), .A(n6494), .B(n6493), .ZN(n8249)
         );
  INV_X1 U8124 ( .A(n6496), .ZN(n6497) );
  NAND2_X1 U8125 ( .A1(n6497), .A2(P2_B_REG_SCAN_IN), .ZN(n6498) );
  AND2_X1 U8126 ( .A1(n8218), .A2(n6498), .ZN(n8346) );
  NAND2_X1 U8127 ( .A1(n8249), .A2(n8346), .ZN(n6499) );
  INV_X1 U8128 ( .A(n7053), .ZN(n9896) );
  NAND3_X1 U8129 ( .A1(n6422), .A2(n9912), .A3(n9896), .ZN(n7088) );
  NAND2_X1 U8130 ( .A1(n9843), .A2(n7301), .ZN(n7279) );
  OR2_X1 U8131 ( .A1(n7279), .A2(n7312), .ZN(n7256) );
  OR2_X2 U8132 ( .A1(n7256), .A2(n7255), .ZN(n7355) );
  NAND2_X1 U8133 ( .A1(n7374), .A2(n9933), .ZN(n7477) );
  OR2_X2 U8134 ( .A1(n7477), .A2(n7481), .ZN(n7518) );
  AND2_X2 U8135 ( .A1(n7519), .A2(n7669), .ZN(n7717) );
  NAND2_X1 U8136 ( .A1(n8549), .A2(n8673), .ZN(n8523) );
  AND2_X2 U8137 ( .A1(n8422), .A2(n8428), .ZN(n8423) );
  INV_X1 U8138 ( .A(n9942), .ZN(n9841) );
  NAND2_X1 U8139 ( .A1(n8360), .A2(n6515), .ZN(n8344) );
  OAI211_X1 U8140 ( .C1(n8360), .C2(n6515), .A(n9841), .B(n8344), .ZN(n8096)
         );
  NAND2_X1 U8141 ( .A1(n8102), .A2(n8096), .ZN(n6502) );
  NAND2_X1 U8142 ( .A1(n7007), .A2(n6505), .ZN(n6511) );
  NOR2_X1 U8143 ( .A1(n6511), .A2(n7008), .ZN(n6506) );
  MUX2_X1 U8144 ( .A(n6507), .B(n6514), .S(n9960), .Z(n6510) );
  NAND2_X1 U8145 ( .A1(n8099), .A2(n6508), .ZN(n6509) );
  NAND2_X1 U8146 ( .A1(n6510), .A2(n6509), .ZN(P2_U3549) );
  INV_X1 U8147 ( .A(n7008), .ZN(n6512) );
  NOR2_X1 U8148 ( .A1(n6512), .A2(n6511), .ZN(n6513) );
  INV_X1 U8149 ( .A(n8677), .ZN(n6516) );
  NAND2_X1 U8150 ( .A1(n8099), .A2(n6516), .ZN(n6517) );
  NAND2_X1 U8151 ( .A1(n6518), .A2(n6517), .ZN(P2_U3517) );
  INV_X1 U8152 ( .A(n7587), .ZN(n6519) );
  OR2_X1 U8153 ( .A1(n6889), .A2(n6519), .ZN(n6520) );
  NAND2_X1 U8154 ( .A1(n6573), .A2(n6521), .ZN(n6615) );
  NAND2_X1 U8155 ( .A1(n6615), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  XNOR2_X1 U8156 ( .A(n6523), .B(n6522), .ZN(n6524) );
  NOR2_X1 U8157 ( .A1(n6524), .A2(n8247), .ZN(n6530) );
  INV_X1 U8158 ( .A(n7523), .ZN(n9941) );
  NOR2_X1 U8159 ( .A1(n9819), .A2(n9941), .ZN(n6529) );
  NOR2_X1 U8160 ( .A1(n9824), .A2(n7521), .ZN(n6528) );
  OR2_X1 U8161 ( .A1(n7709), .A2(n9814), .ZN(n6526) );
  NAND2_X1 U8162 ( .A1(n8265), .A2(n8228), .ZN(n6525) );
  AND2_X1 U8163 ( .A1(n6526), .A2(n6525), .ZN(n7516) );
  OAI22_X1 U8164 ( .A1(n7516), .A2(n8233), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5292), .ZN(n6527) );
  OR4_X1 U8165 ( .A1(n6530), .A2(n6529), .A3(n6528), .A4(n6527), .ZN(P2_U3238)
         );
  INV_X1 U8166 ( .A(n6955), .ZN(n6567) );
  NOR2_X1 U8167 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n9704), .ZN(n6531) );
  AOI21_X1 U8168 ( .B1(n9704), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6531), .ZN(
        n9708) );
  NAND2_X1 U8169 ( .A1(n9696), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6532) );
  OAI21_X1 U8170 ( .B1(n9696), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6532), .ZN(
        n9692) );
  NOR2_X1 U8171 ( .A1(n6606), .A2(n7190), .ZN(n6540) );
  MUX2_X1 U8172 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7034), .S(n9668), .Z(n9665)
         );
  INV_X1 U8173 ( .A(n6587), .ZN(n6653) );
  NOR2_X1 U8174 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6653), .ZN(n6536) );
  NOR2_X1 U8175 ( .A1(n9654), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U8176 ( .A1(n6580), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6534) );
  INV_X1 U8177 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6533) );
  MUX2_X1 U8178 ( .A(n6533), .B(P1_REG2_REG_1__SCAN_IN), .S(n6578), .Z(n6635)
         );
  INV_X1 U8179 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6610) );
  INV_X1 U8180 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10275) );
  NOR3_X1 U8181 ( .A1(n6635), .A2(n6610), .A3(n10275), .ZN(n6634) );
  AOI21_X1 U8182 ( .B1(n6578), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6634), .ZN(
        n9640) );
  INV_X1 U8183 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6881) );
  MUX2_X1 U8184 ( .A(n6881), .B(P1_REG2_REG_2__SCAN_IN), .S(n6557), .Z(n9639)
         );
  NOR2_X1 U8185 ( .A1(n9640), .A2(n9639), .ZN(n9638) );
  MUX2_X1 U8186 ( .A(n5853), .B(P1_REG2_REG_3__SCAN_IN), .S(n6580), .Z(n9527)
         );
  NAND2_X1 U8187 ( .A1(n6534), .A2(n9530), .ZN(n9650) );
  INV_X1 U8188 ( .A(n9654), .ZN(n6585) );
  AOI22_X1 U8189 ( .A1(n9654), .A2(n6909), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n6585), .ZN(n9649) );
  NOR2_X1 U8190 ( .A1(n9650), .A2(n9649), .ZN(n9648) );
  NOR2_X1 U8191 ( .A1(n6535), .A2(n9648), .ZN(n6649) );
  AOI22_X1 U8192 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6587), .B1(n6653), .B2(
        n5887), .ZN(n6648) );
  NOR2_X1 U8193 ( .A1(n6649), .A2(n6648), .ZN(n6647) );
  NOR2_X1 U8194 ( .A1(n6536), .A2(n6647), .ZN(n6628) );
  INV_X1 U8195 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6537) );
  MUX2_X1 U8196 ( .A(n6537), .B(P1_REG2_REG_6__SCAN_IN), .S(n6623), .Z(n6627)
         );
  NAND2_X1 U8197 ( .A1(n6628), .A2(n6627), .ZN(n6626) );
  INV_X1 U8198 ( .A(n6623), .ZN(n6538) );
  NAND2_X1 U8199 ( .A1(n6538), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U8200 ( .A1(n6626), .A2(n6539), .ZN(n9666) );
  NOR2_X1 U8201 ( .A1(n9665), .A2(n9666), .ZN(n9664) );
  NAND2_X1 U8202 ( .A1(n6606), .A2(n7190), .ZN(n9684) );
  NOR2_X1 U8203 ( .A1(n9692), .A2(n9693), .ZN(n9691) );
  AOI21_X1 U8204 ( .B1(n9696), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9691), .ZN(
        n6814) );
  NAND2_X1 U8205 ( .A1(n6816), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6541) );
  OAI21_X1 U8206 ( .B1(n6816), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6541), .ZN(
        n6813) );
  NOR2_X1 U8207 ( .A1(n6814), .A2(n6813), .ZN(n6812) );
  AOI21_X1 U8208 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6816), .A(n6812), .ZN(
        n9707) );
  NAND2_X1 U8209 ( .A1(n9708), .A2(n9707), .ZN(n9706) );
  OAI21_X1 U8210 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9704), .A(n9706), .ZN(
        n6957) );
  XOR2_X1 U8211 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n6955), .Z(n6958) );
  NOR2_X1 U8212 ( .A1(n6957), .A2(n6958), .ZN(n6956) );
  AOI21_X1 U8213 ( .B1(n6567), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6956), .ZN(
        n7073) );
  MUX2_X1 U8214 ( .A(n6542), .B(P1_REG2_REG_13__SCAN_IN), .S(n6569), .Z(n7072)
         );
  INV_X1 U8215 ( .A(n7389), .ZN(n6835) );
  NOR2_X1 U8216 ( .A1(n6543), .A2(n6835), .ZN(n6544) );
  XNOR2_X1 U8217 ( .A(n6835), .B(n6543), .ZN(n7387) );
  NOR2_X1 U8218 ( .A1(n6091), .A2(n7387), .ZN(n7386) );
  XNOR2_X1 U8219 ( .A(n7683), .B(n7682), .ZN(n6547) );
  INV_X1 U8220 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6546) );
  NOR2_X1 U8221 ( .A1(n6546), .A2(n6547), .ZN(n7684) );
  INV_X1 U8222 ( .A(n6573), .ZN(n6545) );
  NAND2_X1 U8223 ( .A1(n9124), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9516) );
  NOR2_X1 U8224 ( .A1(n6545), .A2(n9516), .ZN(n6570) );
  INV_X1 U8225 ( .A(n9626), .ZN(n9162) );
  AOI211_X1 U8226 ( .C1(n6547), .C2(n6546), .A(n7684), .B(n9690), .ZN(n6577)
         );
  INV_X1 U8227 ( .A(n6548), .ZN(n6549) );
  NOR2_X1 U8228 ( .A1(P1_U3083), .A2(n6549), .ZN(n9730) );
  INV_X1 U8229 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n6550) );
  NOR2_X1 U8230 ( .A1(n9717), .A2(n6550), .ZN(n6576) );
  MUX2_X1 U8231 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n6551), .S(n7389), .Z(n7383)
         );
  INV_X1 U8232 ( .A(n9704), .ZN(n6674) );
  AOI22_X1 U8233 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n9704), .B1(n6674), .B2(
        n6022), .ZN(n9711) );
  MUX2_X1 U8234 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6552), .S(n6816), .Z(n6818)
         );
  NOR2_X1 U8235 ( .A1(n9696), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6553) );
  AOI21_X1 U8236 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9696), .A(n6553), .ZN(
        n9699) );
  NOR2_X1 U8237 ( .A1(n6606), .A2(n6554), .ZN(n6565) );
  NAND2_X1 U8238 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6653), .ZN(n6562) );
  MUX2_X1 U8239 ( .A(n6555), .B(P1_REG1_REG_5__SCAN_IN), .S(n6587), .Z(n6651)
         );
  NOR2_X1 U8240 ( .A1(n9654), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6561) );
  AOI22_X1 U8241 ( .A1(n9654), .A2(n5870), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n6585), .ZN(n9647) );
  NAND2_X1 U8242 ( .A1(n6580), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6560) );
  INV_X1 U8243 ( .A(n6557), .ZN(n9624) );
  MUX2_X1 U8244 ( .A(n5813), .B(P1_REG1_REG_1__SCAN_IN), .S(n6578), .Z(n6638)
         );
  NOR3_X1 U8245 ( .A1(n6638), .A2(n6556), .A3(n10275), .ZN(n6636) );
  AOI21_X1 U8246 ( .B1(n6578), .B2(P1_REG1_REG_1__SCAN_IN), .A(n6636), .ZN(
        n9635) );
  MUX2_X1 U8247 ( .A(n6558), .B(P1_REG1_REG_2__SCAN_IN), .S(n6557), .Z(n9634)
         );
  OR2_X1 U8248 ( .A1(n9635), .A2(n9634), .ZN(n9637) );
  OAI21_X1 U8249 ( .B1(n9624), .B2(n6558), .A(n9637), .ZN(n9533) );
  MUX2_X1 U8250 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6559), .S(n6580), .Z(n9532)
         );
  NAND2_X1 U8251 ( .A1(n9533), .A2(n9532), .ZN(n9531) );
  NAND2_X1 U8252 ( .A1(n6560), .A2(n9531), .ZN(n9646) );
  NOR2_X1 U8253 ( .A1(n9647), .A2(n9646), .ZN(n9645) );
  NOR2_X1 U8254 ( .A1(n6561), .A2(n9645), .ZN(n6652) );
  NAND2_X1 U8255 ( .A1(n6651), .A2(n6652), .ZN(n6650) );
  AND2_X1 U8256 ( .A1(n6562), .A2(n6650), .ZN(n6621) );
  MUX2_X1 U8257 ( .A(n5922), .B(P1_REG1_REG_6__SCAN_IN), .S(n6623), .Z(n6622)
         );
  NAND2_X1 U8258 ( .A1(n6621), .A2(n6622), .ZN(n6620) );
  NAND2_X1 U8259 ( .A1(n6623), .A2(n5922), .ZN(n6563) );
  AND2_X1 U8260 ( .A1(n6620), .A2(n6563), .ZN(n9663) );
  MUX2_X1 U8261 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6564), .S(n9668), .Z(n9662)
         );
  NOR2_X1 U8262 ( .A1(n9663), .A2(n9662), .ZN(n9661) );
  AOI21_X1 U8263 ( .B1(n9668), .B2(n6564), .A(n9661), .ZN(n9683) );
  NAND2_X1 U8264 ( .A1(n6606), .A2(n6554), .ZN(n9682) );
  OAI21_X1 U8265 ( .B1(n6565), .B2(n9683), .A(n9682), .ZN(n9698) );
  NAND2_X1 U8266 ( .A1(n9699), .A2(n9698), .ZN(n9697) );
  OAI21_X1 U8267 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9696), .A(n9697), .ZN(
        n6819) );
  NAND2_X1 U8268 ( .A1(n6818), .A2(n6819), .ZN(n6817) );
  OAI21_X1 U8269 ( .B1(n6816), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6817), .ZN(
        n9710) );
  NAND2_X1 U8270 ( .A1(n9711), .A2(n9710), .ZN(n9709) );
  OAI21_X1 U8271 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9704), .A(n9709), .ZN(
        n6952) );
  MUX2_X1 U8272 ( .A(n6566), .B(P1_REG1_REG_12__SCAN_IN), .S(n6955), .Z(n6953)
         );
  NAND2_X1 U8273 ( .A1(n6952), .A2(n6953), .ZN(n6951) );
  OAI21_X1 U8274 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n6567), .A(n6951), .ZN(
        n7067) );
  MUX2_X1 U8275 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6568), .S(n6569), .Z(n7068)
         );
  NAND2_X1 U8276 ( .A1(n7067), .A2(n7068), .ZN(n7066) );
  OAI21_X1 U8277 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n6569), .A(n7066), .ZN(
        n7384) );
  NAND2_X1 U8278 ( .A1(n7383), .A2(n7384), .ZN(n7382) );
  OAI21_X1 U8279 ( .B1(n7389), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7382), .ZN(
        n7672) );
  XNOR2_X1 U8280 ( .A(n7682), .B(n7672), .ZN(n6571) );
  INV_X1 U8281 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9612) );
  NOR2_X1 U8282 ( .A1(n9612), .A2(n6571), .ZN(n7673) );
  NAND2_X1 U8283 ( .A1(n6570), .A2(n9626), .ZN(n9673) );
  AOI211_X1 U8284 ( .C1(n6571), .C2(n9612), .A(n7673), .B(n9673), .ZN(n6575)
         );
  NAND2_X1 U8285 ( .A1(n9162), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9520) );
  NOR2_X1 U8286 ( .A1(n9124), .A2(n9520), .ZN(n6572) );
  NAND2_X1 U8287 ( .A1(n6573), .A2(n6572), .ZN(n9724) );
  NAND2_X1 U8288 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8820) );
  OAI21_X1 U8289 ( .B1(n9724), .B2(n7682), .A(n8820), .ZN(n6574) );
  OR4_X1 U8290 ( .A1(n6577), .A2(n6576), .A3(n6575), .A4(n6574), .ZN(P1_U3256)
         );
  NOR2_X1 U8291 ( .A1(n6469), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9511) );
  INV_X2 U8292 ( .A(n9511), .ZN(n9522) );
  INV_X1 U8293 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6579) );
  AND2_X1 U8294 ( .A1(n6469), .A2(P1_U3084), .ZN(n9518) );
  INV_X2 U8295 ( .A(n9518), .ZN(n9513) );
  INV_X1 U8296 ( .A(n6578), .ZN(n6639) );
  OAI222_X1 U8297 ( .A1(n9522), .A2(n6579), .B1(n9513), .B2(n6596), .C1(
        P1_U3084), .C2(n6639), .ZN(P1_U3352) );
  OAI222_X1 U8298 ( .A1(n9522), .A2(n4738), .B1(n9513), .B2(n6594), .C1(
        P1_U3084), .C2(n9624), .ZN(P1_U3351) );
  INV_X1 U8299 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6581) );
  INV_X1 U8300 ( .A(n6580), .ZN(n9524) );
  OAI222_X1 U8301 ( .A1(n9522), .A2(n6581), .B1(n9513), .B2(n6583), .C1(
        P1_U3084), .C2(n9524), .ZN(P1_U3350) );
  INV_X2 U8302 ( .A(n8683), .ZN(n8694) );
  AND2_X1 U8303 ( .A1(n6582), .A2(P2_U3152), .ZN(n8690) );
  INV_X2 U8304 ( .A(n8690), .ZN(n8696) );
  OAI222_X1 U8305 ( .A1(n8694), .A2(n6584), .B1(n8696), .B2(n6583), .C1(
        P2_U3152), .C2(n6721), .ZN(P2_U3355) );
  INV_X1 U8306 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6586) );
  OAI222_X1 U8307 ( .A1(n9522), .A2(n6586), .B1(n9513), .B2(n6591), .C1(
        P1_U3084), .C2(n6585), .ZN(P1_U3349) );
  OAI222_X1 U8308 ( .A1(n9522), .A2(n6588), .B1(n9513), .B2(n6589), .C1(
        P1_U3084), .C2(n6587), .ZN(P1_U3348) );
  OAI222_X1 U8309 ( .A1(n8694), .A2(n6590), .B1(n8696), .B2(n6589), .C1(
        P2_U3152), .C2(n6710), .ZN(P2_U3353) );
  OAI222_X1 U8310 ( .A1(n8694), .A2(n6592), .B1(n8696), .B2(n6591), .C1(
        P2_U3152), .C2(n6769), .ZN(P2_U3354) );
  OAI222_X1 U8311 ( .A1(n8694), .A2(n6595), .B1(n8696), .B2(n6594), .C1(
        P2_U3152), .C2(n6593), .ZN(P2_U3356) );
  OAI222_X1 U8312 ( .A1(n8694), .A2(n6597), .B1(n8696), .B2(n6596), .C1(
        P2_U3152), .C2(n9546), .ZN(P2_U3357) );
  INV_X1 U8313 ( .A(n9754), .ZN(n6773) );
  NAND2_X1 U8314 ( .A1(n6775), .A2(n6773), .ZN(n6598) );
  OAI21_X1 U8315 ( .B1(n6773), .B2(n6342), .A(n6598), .ZN(P1_U3440) );
  NAND2_X1 U8316 ( .A1(n6877), .A2(n6773), .ZN(n6599) );
  OAI21_X1 U8317 ( .B1(n6773), .B2(n6354), .A(n6599), .ZN(P1_U3441) );
  OAI222_X1 U8318 ( .A1(n9522), .A2(n6600), .B1(n9513), .B2(n6601), .C1(
        P1_U3084), .C2(n6623), .ZN(P1_U3347) );
  OAI222_X1 U8319 ( .A1(n8694), .A2(n6602), .B1(n8696), .B2(n6601), .C1(
        P2_U3152), .C2(n6743), .ZN(P2_U3352) );
  OAI222_X1 U8320 ( .A1(n8694), .A2(n6603), .B1(n8696), .B2(n6604), .C1(
        P2_U3152), .C2(n6759), .ZN(P2_U3351) );
  OAI222_X1 U8321 ( .A1(n9522), .A2(n6605), .B1(n9513), .B2(n6604), .C1(
        P1_U3084), .C2(n9668), .ZN(P1_U3346) );
  INV_X1 U8322 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U8323 ( .A1(n9162), .A2(n6610), .ZN(n6611) );
  NAND2_X1 U8324 ( .A1(n9124), .A2(n6611), .ZN(n9629) );
  INV_X1 U8325 ( .A(n9629), .ZN(n6613) );
  OAI21_X1 U8326 ( .B1(n9162), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6613), .ZN(
        n6612) );
  MUX2_X1 U8327 ( .A(n6613), .B(n6612), .S(n10275), .Z(n6614) );
  NOR3_X1 U8328 ( .A1(n6615), .A2(n6614), .A3(P1_U3084), .ZN(n6616) );
  AOI21_X1 U8329 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .A(n6616), .ZN(
        n6618) );
  INV_X1 U8330 ( .A(n9673), .ZN(n9731) );
  NAND3_X1 U8331 ( .A1(n9731), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6556), .ZN(
        n6617) );
  OAI211_X1 U8332 ( .C1(n9717), .C2(n6619), .A(n6618), .B(n6617), .ZN(P1_U3241) );
  INV_X1 U8333 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6631) );
  OAI21_X1 U8334 ( .B1(n6622), .B2(n6621), .A(n6620), .ZN(n6625) );
  AND2_X1 U8335 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7140) );
  NOR2_X1 U8336 ( .A1(n9724), .A2(n6623), .ZN(n6624) );
  AOI211_X1 U8337 ( .C1(n9731), .C2(n6625), .A(n7140), .B(n6624), .ZN(n6630)
         );
  OAI211_X1 U8338 ( .C1(n6628), .C2(n6627), .A(n9718), .B(n6626), .ZN(n6629)
         );
  OAI211_X1 U8339 ( .C1(n6631), .C2(n9717), .A(n6630), .B(n6629), .ZN(P1_U3247) );
  INV_X1 U8340 ( .A(n6632), .ZN(n6645) );
  AOI22_X1 U8341 ( .A1(n9696), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9511), .ZN(n6633) );
  OAI21_X1 U8342 ( .B1(n6645), .B2(n9513), .A(n6633), .ZN(P1_U3344) );
  INV_X1 U8343 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U8344 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9628) );
  AOI211_X1 U8345 ( .C1(n9628), .C2(n6635), .A(n6634), .B(n9690), .ZN(n6642)
         );
  NAND2_X1 U8346 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6637) );
  AOI211_X1 U8347 ( .C1(n6638), .C2(n6637), .A(n6636), .B(n9673), .ZN(n6641)
         );
  OAI22_X1 U8348 ( .A1(n9724), .A2(n6639), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6946), .ZN(n6640) );
  NOR3_X1 U8349 ( .A1(n6642), .A2(n6641), .A3(n6640), .ZN(n6643) );
  OAI21_X1 U8350 ( .B1(n9717), .B2(n6644), .A(n6643), .ZN(P1_U3242) );
  INV_X1 U8351 ( .A(n6845), .ZN(n6802) );
  OAI222_X1 U8352 ( .A1(n8694), .A2(n6646), .B1(n8696), .B2(n6645), .C1(n6802), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  AOI21_X1 U8353 ( .B1(n6649), .B2(n6648), .A(n6647), .ZN(n6656) );
  OAI211_X1 U8354 ( .C1(n6652), .C2(n6651), .A(n9731), .B(n6650), .ZN(n6655)
         );
  AND2_X1 U8355 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7083) );
  AOI21_X1 U8356 ( .B1(n9705), .B2(n6653), .A(n7083), .ZN(n6654) );
  OAI211_X1 U8357 ( .C1(n9690), .C2(n6656), .A(n6655), .B(n6654), .ZN(n6657)
         );
  AOI21_X1 U8358 ( .B1(n9730), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6657), .ZN(
        n6658) );
  INV_X1 U8359 ( .A(n6658), .ZN(P1_U3246) );
  INV_X1 U8360 ( .A(n6659), .ZN(n6672) );
  AOI22_X1 U8361 ( .A1(n6816), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9511), .ZN(n6660) );
  OAI21_X1 U8362 ( .B1(n6672), .B2(n9513), .A(n6660), .ZN(P1_U3343) );
  INV_X1 U8363 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10083) );
  INV_X1 U8364 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8345) );
  INV_X1 U8365 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8562) );
  OR2_X1 U8366 ( .A1(n5167), .A2(n8562), .ZN(n6662) );
  NAND2_X1 U8367 ( .A1(n5161), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6661) );
  OAI211_X1 U8368 ( .C1(n6663), .C2(n8345), .A(n6662), .B(n6661), .ZN(n8347)
         );
  NAND2_X1 U8369 ( .A1(n8347), .A2(P2_U3966), .ZN(n6664) );
  OAI21_X1 U8370 ( .B1(P2_U3966), .B2(n10083), .A(n6664), .ZN(P2_U3583) );
  OR2_X1 U8371 ( .A1(n6665), .A2(P2_U3152), .ZN(n8082) );
  NAND2_X1 U8372 ( .A1(n9856), .A2(n8082), .ZN(n6667) );
  NAND2_X1 U8373 ( .A1(n6667), .A2(n6666), .ZN(n6670) );
  OR2_X1 U8374 ( .A1(n9856), .A2(n6668), .ZN(n6669) );
  AND2_X1 U8375 ( .A1(n6670), .A2(n6669), .ZN(n9537) );
  INV_X1 U8376 ( .A(n9537), .ZN(n9832) );
  NOR2_X1 U8377 ( .A1(n9832), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8378 ( .A(n6997), .ZN(n6853) );
  OAI222_X1 U8379 ( .A1(P2_U3152), .A2(n6853), .B1(n8696), .B2(n6672), .C1(
        n6671), .C2(n8694), .ZN(P2_U3348) );
  INV_X1 U8380 ( .A(n6673), .ZN(n6677) );
  INV_X1 U8381 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10158) );
  OAI222_X1 U8382 ( .A1(n9513), .A2(n6677), .B1(n6674), .B2(P1_U3084), .C1(
        n10158), .C2(n9522), .ZN(P1_U3342) );
  NAND2_X1 U8383 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n8275), .ZN(n6675) );
  OAI21_X1 U8384 ( .B1(n8170), .B2(n8275), .A(n6675), .ZN(P2_U3567) );
  INV_X1 U8385 ( .A(n7107), .ZN(n7003) );
  INV_X1 U8386 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6676) );
  OAI222_X1 U8387 ( .A1(P2_U3152), .A2(n7003), .B1(n8696), .B2(n6677), .C1(
        n6676), .C2(n8694), .ZN(P2_U3347) );
  NAND2_X1 U8388 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n8275), .ZN(n6678) );
  OAI21_X1 U8389 ( .B1(n8147), .B2(n8275), .A(n6678), .ZN(P2_U3574) );
  OR2_X1 U8390 ( .A1(n5713), .A2(P2_U3152), .ZN(n8691) );
  OR2_X1 U8391 ( .A1(n9856), .A2(n6679), .ZN(n6680) );
  OAI211_X1 U8392 ( .C1(n6681), .C2(n8691), .A(n6680), .B(n8082), .ZN(n6691)
         );
  NAND2_X1 U8393 ( .A1(n6691), .A2(n6689), .ZN(n6682) );
  NAND2_X1 U8394 ( .A1(n6682), .A2(n8275), .ZN(n6705) );
  NAND2_X1 U8395 ( .A1(n6705), .A2(n5713), .ZN(n9828) );
  NOR2_X1 U8396 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5142), .ZN(n7171) );
  INV_X1 U8397 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9835) );
  INV_X1 U8398 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6683) );
  NOR2_X1 U8399 ( .A1(n9546), .A2(n6683), .ZN(n6684) );
  NOR2_X1 U8400 ( .A1(n9539), .A2(n6684), .ZN(n9557) );
  NAND2_X1 U8401 ( .A1(P2_REG1_REG_2__SCAN_IN), .A2(n9559), .ZN(n6685) );
  OAI21_X1 U8402 ( .B1(n9559), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6685), .ZN(
        n9556) );
  NAND2_X1 U8403 ( .A1(n6697), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6686) );
  OAI21_X1 U8404 ( .B1(n6697), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6686), .ZN(
        n6712) );
  NAND2_X1 U8405 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n6695), .ZN(n6687) );
  OAI21_X1 U8406 ( .B1(n6695), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6687), .ZN(
        n6761) );
  NOR2_X1 U8407 ( .A1(n6762), .A2(n6761), .ZN(n6760) );
  AOI21_X1 U8408 ( .B1(n6695), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6760), .ZN(
        n6693) );
  NAND2_X1 U8409 ( .A1(n6728), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6688) );
  OAI21_X1 U8410 ( .B1(n6728), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6688), .ZN(
        n6692) );
  NOR2_X1 U8411 ( .A1(n6693), .A2(n6692), .ZN(n6723) );
  AND2_X1 U8412 ( .A1(n6689), .A2(n6496), .ZN(n6690) );
  AOI211_X1 U8413 ( .C1(n6693), .C2(n6692), .A(n6723), .B(n9554), .ZN(n6694)
         );
  AOI211_X1 U8414 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9832), .A(n7171), .B(
        n6694), .ZN(n6709) );
  NAND2_X1 U8415 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n6695), .ZN(n6702) );
  MUX2_X1 U8416 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6696), .S(n6695), .Z(n6765)
         );
  NAND2_X1 U8417 ( .A1(n6697), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6701) );
  MUX2_X1 U8418 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6698), .S(n6697), .Z(n6717)
         );
  NAND2_X1 U8419 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(n9559), .ZN(n6700) );
  MUX2_X1 U8420 ( .A(n7061), .B(P2_REG2_REG_2__SCAN_IN), .S(n9559), .Z(n6699)
         );
  INV_X1 U8421 ( .A(n6699), .ZN(n9562) );
  MUX2_X1 U8422 ( .A(n7049), .B(P2_REG2_REG_1__SCAN_IN), .S(n9546), .Z(n9550)
         );
  NAND3_X1 U8423 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9550), .ZN(n9549) );
  OAI21_X1 U8424 ( .B1(n9546), .B2(n7049), .A(n9549), .ZN(n9563) );
  NAND2_X1 U8425 ( .A1(n9562), .A2(n9563), .ZN(n9561) );
  NAND2_X1 U8426 ( .A1(n6700), .A2(n9561), .ZN(n6718) );
  NAND2_X1 U8427 ( .A1(n6717), .A2(n6718), .ZN(n6716) );
  NAND2_X1 U8428 ( .A1(n6701), .A2(n6716), .ZN(n6766) );
  NAND2_X1 U8429 ( .A1(n6765), .A2(n6766), .ZN(n6764) );
  NAND2_X1 U8430 ( .A1(n6702), .A2(n6764), .ZN(n6707) );
  MUX2_X1 U8431 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6703), .S(n6728), .Z(n6706)
         );
  NOR2_X1 U8432 ( .A1(n5713), .A2(n6496), .ZN(n6704) );
  NAND2_X1 U8433 ( .A1(n6705), .A2(n6704), .ZN(n9830) );
  NAND2_X1 U8434 ( .A1(n6706), .A2(n6707), .ZN(n6729) );
  OAI211_X1 U8435 ( .C1(n6707), .C2(n6706), .A(n9825), .B(n6729), .ZN(n6708)
         );
  OAI211_X1 U8436 ( .C1(n9828), .C2(n6710), .A(n6709), .B(n6708), .ZN(P2_U3250) );
  INV_X1 U8437 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10300) );
  NOR2_X1 U8438 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10300), .ZN(n6715) );
  AOI211_X1 U8439 ( .C1(n6713), .C2(n6712), .A(n6711), .B(n9554), .ZN(n6714)
         );
  AOI211_X1 U8440 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9832), .A(n6715), .B(
        n6714), .ZN(n6720) );
  OAI211_X1 U8441 ( .C1(n6718), .C2(n6717), .A(n9825), .B(n6716), .ZN(n6719)
         );
  OAI211_X1 U8442 ( .C1(n9828), .C2(n6721), .A(n6720), .B(n6719), .ZN(P2_U3248) );
  NOR2_X1 U8443 ( .A1(n6722), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7321) );
  AOI21_X1 U8444 ( .B1(n6728), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6723), .ZN(
        n6726) );
  MUX2_X1 U8445 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6724), .S(n6743), .Z(n6725)
         );
  AOI211_X1 U8446 ( .C1(n6726), .C2(n6725), .A(n6735), .B(n9554), .ZN(n6727)
         );
  AOI211_X1 U8447 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9832), .A(n7321), .B(
        n6727), .ZN(n6734) );
  NAND2_X1 U8448 ( .A1(n6728), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6730) );
  NAND2_X1 U8449 ( .A1(n6730), .A2(n6729), .ZN(n6732) );
  MUX2_X1 U8450 ( .A(n7233), .B(P2_REG2_REG_6__SCAN_IN), .S(n6743), .Z(n6731)
         );
  NAND2_X1 U8451 ( .A1(n6731), .A2(n6732), .ZN(n6742) );
  OAI211_X1 U8452 ( .C1(n6732), .C2(n6731), .A(n9825), .B(n6742), .ZN(n6733)
         );
  OAI211_X1 U8453 ( .C1(n9828), .C2(n6743), .A(n6734), .B(n6733), .ZN(P2_U3251) );
  NOR2_X1 U8454 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10318), .ZN(n7495) );
  NAND2_X1 U8455 ( .A1(n6740), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6736) );
  OAI21_X1 U8456 ( .B1(n6740), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6736), .ZN(
        n6751) );
  MUX2_X1 U8457 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n4667), .S(n6797), .Z(n6737)
         );
  NOR2_X1 U8458 ( .A1(n6738), .A2(n6737), .ZN(n6789) );
  AOI211_X1 U8459 ( .C1(n6738), .C2(n6737), .A(n6789), .B(n9554), .ZN(n6739)
         );
  AOI211_X1 U8460 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9832), .A(n7495), .B(
        n6739), .ZN(n6749) );
  NAND2_X1 U8461 ( .A1(n6740), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6744) );
  MUX2_X1 U8462 ( .A(n7265), .B(P2_REG2_REG_7__SCAN_IN), .S(n6740), .Z(n6741)
         );
  INV_X1 U8463 ( .A(n6741), .ZN(n6756) );
  OAI21_X1 U8464 ( .B1(n6743), .B2(n7233), .A(n6742), .ZN(n6755) );
  NAND2_X1 U8465 ( .A1(n6756), .A2(n6755), .ZN(n6754) );
  NAND2_X1 U8466 ( .A1(n6744), .A2(n6754), .ZN(n6747) );
  MUX2_X1 U8467 ( .A(n6745), .B(P2_REG2_REG_8__SCAN_IN), .S(n6797), .Z(n6746)
         );
  NAND2_X1 U8468 ( .A1(n6746), .A2(n6747), .ZN(n6796) );
  OAI211_X1 U8469 ( .C1(n6747), .C2(n6746), .A(n9825), .B(n6796), .ZN(n6748)
         );
  OAI211_X1 U8470 ( .C1(n9828), .C2(n6797), .A(n6749), .B(n6748), .ZN(P2_U3253) );
  NOR2_X1 U8471 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5183), .ZN(n7409) );
  AOI211_X1 U8472 ( .C1(n6752), .C2(n6751), .A(n6750), .B(n9554), .ZN(n6753)
         );
  AOI211_X1 U8473 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9832), .A(n7409), .B(
        n6753), .ZN(n6758) );
  OAI211_X1 U8474 ( .C1(n6756), .C2(n6755), .A(n9825), .B(n6754), .ZN(n6757)
         );
  OAI211_X1 U8475 ( .C1(n9828), .C2(n6759), .A(n6758), .B(n6757), .ZN(P2_U3252) );
  INV_X1 U8476 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10170) );
  NOR2_X1 U8477 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10170), .ZN(n9816) );
  AOI211_X1 U8478 ( .C1(n6762), .C2(n6761), .A(n6760), .B(n9554), .ZN(n6763)
         );
  AOI211_X1 U8479 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9832), .A(n9816), .B(
        n6763), .ZN(n6768) );
  OAI211_X1 U8480 ( .C1(n6766), .C2(n6765), .A(n9825), .B(n6764), .ZN(n6767)
         );
  OAI211_X1 U8481 ( .C1(n9828), .C2(n6769), .A(n6768), .B(n6767), .ZN(P2_U3249) );
  INV_X1 U8482 ( .A(n6770), .ZN(n6771) );
  NOR2_X1 U8483 ( .A1(n6877), .A2(n6771), .ZN(n6782) );
  NAND3_X1 U8484 ( .A1(n6773), .A2(n6772), .A3(n6779), .ZN(n6774) );
  NOR2_X2 U8485 ( .A1(n9124), .A2(n6889), .ZN(n9400) );
  NOR2_X1 U8486 ( .A1(n6776), .A2(n6945), .ZN(n6940) );
  AND2_X1 U8487 ( .A1(n6945), .A2(n6776), .ZN(n8881) );
  NOR2_X1 U8488 ( .A1(n6940), .A2(n8881), .ZN(n9056) );
  INV_X1 U8489 ( .A(n6888), .ZN(n9125) );
  OAI21_X1 U8490 ( .B1(n6945), .B2(n6882), .A(n6930), .ZN(n6783) );
  NAND2_X1 U8491 ( .A1(n6783), .A2(n9800), .ZN(n6778) );
  OAI21_X1 U8492 ( .B1(n9800), .B2(n5801), .A(n6778), .ZN(P1_U3454) );
  INV_X1 U8493 ( .A(n6779), .ZN(n6780) );
  NOR2_X1 U8494 ( .A1(n9754), .A2(n6780), .ZN(n6805) );
  NAND2_X1 U8495 ( .A1(n6783), .A2(n9809), .ZN(n6784) );
  OAI21_X1 U8496 ( .B1(n9809), .B2(n6556), .A(n6784), .ZN(P1_U3523) );
  INV_X1 U8497 ( .A(n6785), .ZN(n6787) );
  INV_X1 U8498 ( .A(n7201), .ZN(n7117) );
  OAI222_X1 U8499 ( .A1(n8694), .A2(n6786), .B1(n8696), .B2(n6787), .C1(
        P2_U3152), .C2(n7117), .ZN(P2_U3346) );
  OAI222_X1 U8500 ( .A1(n9522), .A2(n6788), .B1(n9513), .B2(n6787), .C1(
        P1_U3084), .C2(n6955), .ZN(P1_U3341) );
  NAND2_X1 U8501 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7552) );
  INV_X1 U8502 ( .A(n7552), .ZN(n6794) );
  MUX2_X1 U8503 ( .A(n6790), .B(P2_REG1_REG_9__SCAN_IN), .S(n6845), .Z(n6791)
         );
  AOI211_X1 U8504 ( .C1(n6792), .C2(n6791), .A(n6840), .B(n9554), .ZN(n6793)
         );
  AOI211_X1 U8505 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9832), .A(n6794), .B(
        n6793), .ZN(n6801) );
  MUX2_X1 U8506 ( .A(n7375), .B(P2_REG2_REG_9__SCAN_IN), .S(n6845), .Z(n6795)
         );
  INV_X1 U8507 ( .A(n6795), .ZN(n6799) );
  OAI21_X1 U8508 ( .B1(n6797), .B2(n6745), .A(n6796), .ZN(n6798) );
  NAND2_X1 U8509 ( .A1(n6799), .A2(n6798), .ZN(n6846) );
  OAI211_X1 U8510 ( .C1(n6799), .C2(n6798), .A(n9825), .B(n6846), .ZN(n6800)
         );
  OAI211_X1 U8511 ( .C1(n9828), .C2(n6802), .A(n6801), .B(n6800), .ZN(P2_U3254) );
  INV_X1 U8512 ( .A(n6803), .ZN(n6806) );
  OAI211_X1 U8513 ( .C1(n6806), .C2(n9487), .A(n6805), .B(n6804), .ZN(n8792)
         );
  OAI21_X1 U8514 ( .B1(n6809), .B2(n6808), .A(n6807), .ZN(n9627) );
  AOI22_X1 U8515 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n8792), .B1(n8808), .B2(
        n9627), .ZN(n6810) );
  NAND2_X1 U8516 ( .A1(n6811), .A2(n6810), .ZN(P1_U3230) );
  INV_X1 U8517 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6823) );
  AND2_X1 U8518 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7489) );
  AOI211_X1 U8519 ( .C1(n6814), .C2(n6813), .A(n6812), .B(n9690), .ZN(n6815)
         );
  AOI211_X1 U8520 ( .C1(n9705), .C2(n6816), .A(n7489), .B(n6815), .ZN(n6822)
         );
  OAI21_X1 U8521 ( .B1(n6819), .B2(n6818), .A(n6817), .ZN(n6820) );
  NAND2_X1 U8522 ( .A1(n6820), .A2(n9731), .ZN(n6821) );
  OAI211_X1 U8523 ( .C1(n9717), .C2(n6823), .A(n6822), .B(n6821), .ZN(P1_U3251) );
  INV_X1 U8524 ( .A(n6824), .ZN(n6832) );
  OAI222_X1 U8525 ( .A1(n9513), .A2(n6832), .B1(n7070), .B2(P1_U3084), .C1(
        n10321), .C2(n9522), .ZN(P1_U3340) );
  NOR2_X1 U8526 ( .A1(n6420), .A2(n9814), .ZN(n7013) );
  INV_X1 U8527 ( .A(n8078), .ZN(n6825) );
  NAND2_X1 U8528 ( .A1(n6826), .A2(n6825), .ZN(n8087) );
  AOI22_X1 U8529 ( .A1(n9817), .A2(n7013), .B1(n8087), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n6831) );
  NAND2_X1 U8530 ( .A1(n6475), .A2(n9896), .ZN(n7932) );
  INV_X1 U8531 ( .A(n7932), .ZN(n6827) );
  MUX2_X1 U8532 ( .A(n6827), .B(n7053), .S(n7018), .Z(n6829) );
  INV_X1 U8533 ( .A(n7045), .ZN(n6828) );
  OAI21_X1 U8534 ( .B1(n6829), .B2(n6828), .A(n9821), .ZN(n6830) );
  OAI211_X1 U8535 ( .C1(n9819), .C2(n9896), .A(n6831), .B(n6830), .ZN(P2_U3234) );
  INV_X1 U8536 ( .A(n7335), .ZN(n7331) );
  OAI222_X1 U8537 ( .A1(n8694), .A2(n6833), .B1(n8696), .B2(n6832), .C1(n7331), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8538 ( .A(n6834), .ZN(n6836) );
  INV_X1 U8539 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10316) );
  OAI222_X1 U8540 ( .A1(n9513), .A2(n6836), .B1(n6835), .B2(P1_U3084), .C1(
        n10316), .C2(n9522), .ZN(P1_U3339) );
  INV_X1 U8541 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6837) );
  INV_X1 U8542 ( .A(n7592), .ZN(n7339) );
  OAI222_X1 U8543 ( .A1(n8694), .A2(n6837), .B1(n8696), .B2(n6836), .C1(n7339), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NAND2_X1 U8544 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8275), .ZN(n6838) );
  OAI21_X1 U8545 ( .B1(n6839), .B2(n8275), .A(n6838), .ZN(P2_U3581) );
  NOR2_X1 U8546 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10112), .ZN(n7615) );
  INV_X1 U8547 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6841) );
  MUX2_X1 U8548 ( .A(n6841), .B(P2_REG1_REG_10__SCAN_IN), .S(n6997), .Z(n6842)
         );
  AOI211_X1 U8549 ( .C1(n6843), .C2(n6842), .A(n6996), .B(n9554), .ZN(n6844)
         );
  AOI211_X1 U8550 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9832), .A(n7615), .B(
        n6844), .ZN(n6852) );
  NAND2_X1 U8551 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n6845), .ZN(n6847) );
  NAND2_X1 U8552 ( .A1(n6847), .A2(n6846), .ZN(n6850) );
  MUX2_X1 U8553 ( .A(n7476), .B(P2_REG2_REG_10__SCAN_IN), .S(n6997), .Z(n6848)
         );
  INV_X1 U8554 ( .A(n6848), .ZN(n6849) );
  NAND2_X1 U8555 ( .A1(n6849), .A2(n6850), .ZN(n6989) );
  OAI211_X1 U8556 ( .C1(n6850), .C2(n6849), .A(n9825), .B(n6989), .ZN(n6851)
         );
  OAI211_X1 U8557 ( .C1(n9828), .C2(n6853), .A(n6852), .B(n6851), .ZN(P2_U3255) );
  OAI21_X1 U8558 ( .B1(n6856), .B2(n6855), .A(n6854), .ZN(n6857) );
  NAND2_X1 U8559 ( .A1(n6857), .A2(n9821), .ZN(n6859) );
  OAI22_X1 U8560 ( .A1(n6420), .A2(n9812), .B1(n9813), .B2(n9814), .ZN(n7059)
         );
  AOI22_X1 U8561 ( .A1(n9817), .A2(n7059), .B1(n8087), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6858) );
  OAI211_X1 U8562 ( .C1(n9912), .C2(n9819), .A(n6859), .B(n6858), .ZN(P2_U3239) );
  NAND2_X1 U8563 ( .A1(n6860), .A2(n6861), .ZN(n6863) );
  XNOR2_X1 U8564 ( .A(n6863), .B(n6862), .ZN(n6866) );
  AOI22_X1 U8565 ( .A1(n4473), .A2(n6776), .B1(n8811), .B2(n9141), .ZN(n6865)
         );
  AOI22_X1 U8566 ( .A1(n6948), .A2(n8828), .B1(n8792), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6864) );
  OAI211_X1 U8567 ( .C1(n6866), .C2(n8831), .A(n6865), .B(n6864), .ZN(P1_U3220) );
  XNOR2_X1 U8568 ( .A(n6868), .B(n6867), .ZN(n6871) );
  OAI22_X1 U8569 ( .A1(n7046), .A2(n9812), .B1(n7168), .B2(n9814), .ZN(n7096)
         );
  AOI22_X1 U8570 ( .A1(n8244), .A2(n9917), .B1(n9817), .B2(n7096), .ZN(n6870)
         );
  MUX2_X1 U8571 ( .A(n9824), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6869) );
  OAI211_X1 U8572 ( .C1(n6871), .C2(n8247), .A(n6870), .B(n6869), .ZN(P2_U3220) );
  NAND2_X1 U8573 ( .A1(n6898), .A2(n8793), .ZN(n8885) );
  NAND2_X1 U8574 ( .A1(n9141), .A2(n9766), .ZN(n8886) );
  AND2_X1 U8575 ( .A1(n6776), .A2(n6933), .ZN(n6937) );
  INV_X1 U8576 ( .A(n6900), .ZN(n6875) );
  AOI21_X1 U8577 ( .B1(n9054), .B2(n6876), .A(n6875), .ZN(n9763) );
  NAND2_X1 U8578 ( .A1(n6878), .A2(n6877), .ZN(n7035) );
  NOR2_X1 U8579 ( .A1(n6879), .A2(n9745), .ZN(n6880) );
  AND2_X1 U8580 ( .A1(n9751), .A2(n6880), .ZN(n9592) );
  OAI22_X1 U8581 ( .A1(n9743), .A2(n9623), .B1(n6881), .B2(n9751), .ZN(n6886)
         );
  NAND2_X1 U8582 ( .A1(n9751), .A2(n9745), .ZN(n9257) );
  NOR2_X1 U8583 ( .A1(n6948), .A2(n6933), .ZN(n6883) );
  AND2_X1 U8584 ( .A1(n6883), .A2(n9766), .ZN(n9767) );
  INV_X1 U8585 ( .A(n6883), .ZN(n6944) );
  NAND2_X1 U8586 ( .A1(n6944), .A2(n8793), .ZN(n9765) );
  INV_X1 U8587 ( .A(n9765), .ZN(n6884) );
  NOR3_X1 U8588 ( .A1(n9225), .A2(n9767), .A3(n6884), .ZN(n6885) );
  AOI211_X1 U8589 ( .C1(n9585), .C2(n8793), .A(n6886), .B(n6885), .ZN(n6897)
         );
  NAND2_X1 U8590 ( .A1(n9735), .A2(n9745), .ZN(n7127) );
  NOR2_X1 U8591 ( .A1(n6889), .A2(n9632), .ZN(n9578) );
  NAND2_X1 U8592 ( .A1(n6890), .A2(n6948), .ZN(n6891) );
  NAND2_X1 U8593 ( .A1(n6939), .A2(n6891), .ZN(n8888) );
  OAI21_X1 U8594 ( .B1(n9054), .B2(n8888), .A(n6904), .ZN(n6893) );
  OR2_X1 U8595 ( .A1(n9042), .A2(n9745), .ZN(n9040) );
  NAND2_X1 U8596 ( .A1(n4673), .A2(n9122), .ZN(n6892) );
  NAND2_X1 U8597 ( .A1(n6893), .A2(n9574), .ZN(n6894) );
  OAI211_X1 U8598 ( .C1(n9763), .C2(n7127), .A(n6895), .B(n6894), .ZN(n9769)
         );
  NAND2_X1 U8599 ( .A1(n9769), .A2(n9751), .ZN(n6896) );
  OAI211_X1 U8600 ( .C1(n9763), .C2(n7661), .A(n6897), .B(n6896), .ZN(P1_U3289) );
  NAND2_X1 U8601 ( .A1(n6898), .A2(n9766), .ZN(n6899) );
  NAND2_X1 U8602 ( .A1(n6900), .A2(n6899), .ZN(n6918) );
  INV_X1 U8603 ( .A(n9140), .ZN(n6901) );
  NAND2_X1 U8604 ( .A1(n6901), .A2(n7119), .ZN(n9087) );
  INV_X1 U8605 ( .A(n7119), .ZN(n6920) );
  NAND2_X1 U8606 ( .A1(n6918), .A2(n9052), .ZN(n6917) );
  NAND2_X1 U8607 ( .A1(n6901), .A2(n6920), .ZN(n6902) );
  NAND2_X1 U8608 ( .A1(n6917), .A2(n6902), .ZN(n6903) );
  INV_X1 U8609 ( .A(n9139), .ZN(n7023) );
  NAND2_X1 U8610 ( .A1(n7023), .A2(n6968), .ZN(n7149) );
  INV_X1 U8611 ( .A(n6968), .ZN(n9773) );
  NAND2_X1 U8612 ( .A1(n9139), .A2(n9773), .ZN(n9083) );
  NAND2_X1 U8613 ( .A1(n7149), .A2(n9083), .ZN(n6905) );
  NAND2_X1 U8614 ( .A1(n6903), .A2(n6905), .ZN(n7025) );
  OAI21_X1 U8615 ( .B1(n6903), .B2(n6905), .A(n7025), .ZN(n9777) );
  INV_X1 U8616 ( .A(n9777), .ZN(n6916) );
  XNOR2_X1 U8617 ( .A(n7151), .B(n6905), .ZN(n6908) );
  INV_X1 U8618 ( .A(n9574), .ZN(n7853) );
  INV_X1 U8619 ( .A(n7127), .ZN(n9581) );
  NAND2_X1 U8620 ( .A1(n9777), .A2(n9581), .ZN(n6907) );
  AOI22_X1 U8621 ( .A1(n9329), .A2(n9140), .B1(n9138), .B2(n9400), .ZN(n6906)
         );
  OAI211_X1 U8622 ( .C1(n6908), .C2(n7853), .A(n6907), .B(n6906), .ZN(n9775)
         );
  NAND2_X1 U8623 ( .A1(n9775), .A2(n9751), .ZN(n6915) );
  OAI22_X1 U8624 ( .A1(n9751), .A2(n6909), .B1(n6971), .B2(n9743), .ZN(n6913)
         );
  INV_X1 U8625 ( .A(n6919), .ZN(n6911) );
  INV_X1 U8626 ( .A(n7147), .ZN(n6910) );
  OAI21_X1 U8627 ( .B1(n9773), .B2(n6911), .A(n6910), .ZN(n9774) );
  NOR2_X1 U8628 ( .A1(n9225), .A2(n9774), .ZN(n6912) );
  AOI211_X1 U8629 ( .C1(n9585), .C2(n6968), .A(n6913), .B(n6912), .ZN(n6914)
         );
  OAI211_X1 U8630 ( .C1(n6916), .C2(n7661), .A(n6915), .B(n6914), .ZN(P1_U3287) );
  INV_X1 U8631 ( .A(n9490), .ZN(n9798) );
  OAI21_X1 U8632 ( .B1(n6918), .B2(n9052), .A(n6917), .ZN(n7125) );
  OAI21_X1 U8633 ( .B1(n9767), .B2(n6920), .A(n6919), .ZN(n7121) );
  OAI22_X1 U8634 ( .A1(n7121), .A2(n9793), .B1(n6920), .B2(n9791), .ZN(n6925)
         );
  XNOR2_X1 U8635 ( .A(n6921), .B(n9052), .ZN(n6924) );
  NAND2_X1 U8636 ( .A1(n7125), .A2(n9581), .ZN(n6923) );
  AOI22_X1 U8637 ( .A1(n9329), .A2(n9141), .B1(n9139), .B2(n9348), .ZN(n6922)
         );
  OAI211_X1 U8638 ( .C1(n7853), .C2(n6924), .A(n6923), .B(n6922), .ZN(n7122)
         );
  AOI211_X1 U8639 ( .C1(n9798), .C2(n7125), .A(n6925), .B(n7122), .ZN(n6927)
         );
  OR2_X1 U8640 ( .A1(n6927), .A2(n9806), .ZN(n6926) );
  OAI21_X1 U8641 ( .B1(n9809), .B2(n6559), .A(n6926), .ZN(P1_U3526) );
  INV_X1 U8642 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6929) );
  OR2_X1 U8643 ( .A1(n6927), .A2(n9799), .ZN(n6928) );
  OAI21_X1 U8644 ( .B1(n9800), .B2(n6929), .A(n6928), .ZN(P1_U3463) );
  OAI21_X1 U8645 ( .B1(n6931), .B2(n9743), .A(n6930), .ZN(n6932) );
  NAND2_X1 U8646 ( .A1(n6932), .A2(n9751), .ZN(n6935) );
  OAI21_X1 U8647 ( .B1(n9406), .B2(n9585), .A(n6933), .ZN(n6934) );
  OAI211_X1 U8648 ( .C1(n6610), .C2(n9751), .A(n6935), .B(n6934), .ZN(P1_U3291) );
  OAI21_X1 U8649 ( .B1(n6938), .B2(n6937), .A(n6936), .ZN(n9758) );
  AOI22_X1 U8650 ( .A1(n9329), .A2(n6776), .B1(n9141), .B2(n9400), .ZN(n6943)
         );
  OAI21_X1 U8651 ( .B1(n9053), .B2(n6940), .A(n6939), .ZN(n6941) );
  NAND2_X1 U8652 ( .A1(n6941), .A2(n9574), .ZN(n6942) );
  OAI211_X1 U8653 ( .C1(n9758), .C2(n7127), .A(n6943), .B(n6942), .ZN(n9760)
         );
  OAI211_X1 U8654 ( .C1(n4675), .C2(n6945), .A(n6944), .B(n9764), .ZN(n9759)
         );
  OAI22_X1 U8655 ( .A1(n9759), .A2(n9156), .B1(n9743), .B2(n6946), .ZN(n6947)
         );
  OAI21_X1 U8656 ( .B1(n9760), .B2(n6947), .A(n9751), .ZN(n6950) );
  AOI22_X1 U8657 ( .A1(n9585), .A2(n6948), .B1(n9753), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6949) );
  OAI211_X1 U8658 ( .C1(n9758), .C2(n7661), .A(n6950), .B(n6949), .ZN(P1_U3290) );
  OAI21_X1 U8659 ( .B1(n6953), .B2(n6952), .A(n6951), .ZN(n6961) );
  NAND2_X1 U8660 ( .A1(n9730), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U8661 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7740) );
  OAI211_X1 U8662 ( .C1(n9724), .C2(n6955), .A(n6954), .B(n7740), .ZN(n6960)
         );
  AOI211_X1 U8663 ( .C1(n6958), .C2(n6957), .A(n9690), .B(n6956), .ZN(n6959)
         );
  AOI211_X1 U8664 ( .C1(n9731), .C2(n6961), .A(n6960), .B(n6959), .ZN(n6962)
         );
  INV_X1 U8665 ( .A(n6962), .ZN(P1_U3253) );
  INV_X1 U8666 ( .A(n6963), .ZN(n6964) );
  AOI211_X1 U8667 ( .C1(n6966), .C2(n6965), .A(n8831), .B(n6964), .ZN(n6973)
         );
  AOI22_X1 U8668 ( .A1(n4473), .A2(n9140), .B1(n8811), .B2(n9138), .ZN(n6970)
         );
  NOR2_X1 U8669 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6967), .ZN(n9653) );
  AOI21_X1 U8670 ( .B1(n8828), .B2(n6968), .A(n9653), .ZN(n6969) );
  OAI211_X1 U8671 ( .C1(n8822), .C2(n6971), .A(n6970), .B(n6969), .ZN(n6972)
         );
  OR2_X1 U8672 ( .A1(n6973), .A2(n6972), .ZN(P1_U3228) );
  OAI21_X1 U8673 ( .B1(n6976), .B2(n6974), .A(n6975), .ZN(n6980) );
  AOI22_X1 U8674 ( .A1(n4473), .A2(n9141), .B1(n8811), .B2(n9139), .ZN(n6978)
         );
  NOR2_X1 U8675 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7118), .ZN(n9526) );
  AOI21_X1 U8676 ( .B1(n8828), .B2(n7119), .A(n9526), .ZN(n6977) );
  OAI211_X1 U8677 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8822), .A(n6978), .B(
        n6977), .ZN(n6979) );
  AOI21_X1 U8678 ( .B1(n8808), .B2(n6980), .A(n6979), .ZN(n6981) );
  INV_X1 U8679 ( .A(n6981), .ZN(P1_U3216) );
  INV_X1 U8680 ( .A(n6982), .ZN(n6983) );
  OAI222_X1 U8681 ( .A1(n9522), .A2(n10097), .B1(n9513), .B2(n6983), .C1(
        P1_U3084), .C2(n7682), .ZN(P1_U3338) );
  INV_X1 U8682 ( .A(n8283), .ZN(n8277) );
  OAI222_X1 U8683 ( .A1(n8694), .A2(n6984), .B1(n8696), .B2(n6983), .C1(
        P2_U3152), .C2(n8277), .ZN(P2_U3343) );
  INV_X1 U8684 ( .A(n6985), .ZN(n6987) );
  INV_X1 U8685 ( .A(n8304), .ZN(n8292) );
  OAI222_X1 U8686 ( .A1(n8694), .A2(n6986), .B1(n8696), .B2(n6987), .C1(n8292), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8687 ( .A(n7702), .ZN(n6988) );
  OAI222_X1 U8688 ( .A1(n9522), .A2(n10107), .B1(n6988), .B2(P1_U3084), .C1(
        n9513), .C2(n6987), .ZN(P1_U3337) );
  NAND2_X1 U8689 ( .A1(n6997), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U8690 ( .A1(n6990), .A2(n6989), .ZN(n6993) );
  MUX2_X1 U8691 ( .A(n6991), .B(P2_REG2_REG_11__SCAN_IN), .S(n7107), .Z(n6992)
         );
  NOR2_X1 U8692 ( .A1(n6993), .A2(n6992), .ZN(n7101) );
  AOI21_X1 U8693 ( .B1(n6993), .B2(n6992), .A(n7101), .ZN(n7006) );
  NOR2_X1 U8694 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5292), .ZN(n6994) );
  AOI21_X1 U8695 ( .B1(n9832), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6994), .ZN(
        n7002) );
  INV_X1 U8696 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6995) );
  MUX2_X1 U8697 ( .A(n6995), .B(P2_REG1_REG_11__SCAN_IN), .S(n7107), .Z(n6999)
         );
  AOI21_X1 U8698 ( .B1(n6997), .B2(P2_REG1_REG_10__SCAN_IN), .A(n6996), .ZN(
        n6998) );
  NOR2_X1 U8699 ( .A1(n6998), .A2(n6999), .ZN(n7106) );
  AOI21_X1 U8700 ( .B1(n6999), .B2(n6998), .A(n7106), .ZN(n7000) );
  NAND2_X1 U8701 ( .A1(n9827), .A2(n7000), .ZN(n7001) );
  OAI211_X1 U8702 ( .C1(n9828), .C2(n7003), .A(n7002), .B(n7001), .ZN(n7004)
         );
  INV_X1 U8703 ( .A(n7004), .ZN(n7005) );
  OAI21_X1 U8704 ( .B1(n7006), .B2(n9830), .A(n7005), .ZN(P2_U3256) );
  NAND2_X1 U8705 ( .A1(n7045), .A2(n7932), .ZN(n7904) );
  INV_X1 U8706 ( .A(n7904), .ZN(n9899) );
  INV_X1 U8707 ( .A(n7007), .ZN(n7009) );
  AND2_X1 U8708 ( .A1(n7009), .A2(n7008), .ZN(n7010) );
  NAND2_X1 U8709 ( .A1(n7011), .A2(n7010), .ZN(n7042) );
  NAND3_X1 U8710 ( .A1(n8072), .A2(n7923), .A3(n8069), .ZN(n7373) );
  AND2_X1 U8711 ( .A1(n8547), .A2(n7373), .ZN(n7012) );
  AOI21_X1 U8712 ( .B1(n9838), .B2(n7904), .A(n7013), .ZN(n9895) );
  OAI21_X1 U8713 ( .B1(n10273), .B2(n9845), .A(n9895), .ZN(n7015) );
  INV_X1 U8714 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9548) );
  NOR2_X1 U8715 ( .A1(n8553), .A2(n9548), .ZN(n7014) );
  AOI21_X1 U8716 ( .B1(n8553), .B2(n7015), .A(n7014), .ZN(n7022) );
  INV_X1 U8717 ( .A(n7016), .ZN(n7017) );
  INV_X1 U8718 ( .A(n7042), .ZN(n7019) );
  NAND2_X1 U8719 ( .A1(n7019), .A2(n7018), .ZN(n7525) );
  INV_X1 U8720 ( .A(n7525), .ZN(n7020) );
  OAI21_X1 U8721 ( .B1(n8534), .B2(n7020), .A(n7053), .ZN(n7021) );
  OAI211_X1 U8722 ( .C1(n9899), .C2(n8506), .A(n7022), .B(n7021), .ZN(P2_U3296) );
  NAND2_X1 U8723 ( .A1(n7023), .A2(n9773), .ZN(n7024) );
  INV_X1 U8724 ( .A(n9739), .ZN(n7148) );
  NAND2_X1 U8725 ( .A1(n9138), .A2(n7148), .ZN(n7153) );
  AND2_X1 U8726 ( .A1(n9089), .A2(n7153), .ZN(n7144) );
  NAND2_X1 U8727 ( .A1(n9138), .A2(n9739), .ZN(n7026) );
  INV_X1 U8728 ( .A(n7246), .ZN(n9779) );
  NAND2_X1 U8729 ( .A1(n9779), .A2(n9137), .ZN(n9057) );
  INV_X1 U8730 ( .A(n9137), .ZN(n7027) );
  NAND2_X1 U8731 ( .A1(n7027), .A2(n7246), .ZN(n9090) );
  NAND2_X1 U8732 ( .A1(n9057), .A2(n9090), .ZN(n8932) );
  NAND2_X1 U8733 ( .A1(n9779), .A2(n7027), .ZN(n7028) );
  NAND2_X1 U8734 ( .A1(n7239), .A2(n7028), .ZN(n7029) );
  INV_X1 U8735 ( .A(n9136), .ZN(n7138) );
  OR2_X1 U8736 ( .A1(n7138), .A2(n7219), .ZN(n8941) );
  NAND2_X1 U8737 ( .A1(n7219), .A2(n7138), .ZN(n8940) );
  NAND2_X1 U8738 ( .A1(n8941), .A2(n8940), .ZN(n9061) );
  OAI21_X1 U8739 ( .B1(n7029), .B2(n9061), .A(n7178), .ZN(n7030) );
  INV_X1 U8740 ( .A(n7030), .ZN(n7131) );
  NAND2_X1 U8741 ( .A1(n7151), .A2(n9083), .ZN(n8937) );
  AND2_X1 U8742 ( .A1(n4526), .A2(n9090), .ZN(n9088) );
  NAND2_X1 U8743 ( .A1(n8937), .A2(n9088), .ZN(n7032) );
  NAND2_X1 U8744 ( .A1(n9057), .A2(n7153), .ZN(n7031) );
  NAND2_X1 U8745 ( .A1(n7031), .A2(n9090), .ZN(n8892) );
  NAND2_X1 U8746 ( .A1(n7032), .A2(n8892), .ZN(n7181) );
  XNOR2_X1 U8747 ( .A(n7181), .B(n9061), .ZN(n7033) );
  AOI222_X1 U8748 ( .A1(n9574), .A2(n7033), .B1(n9135), .B2(n9400), .C1(n9137), 
        .C2(n9578), .ZN(n7130) );
  MUX2_X1 U8749 ( .A(n7034), .B(n7130), .S(n9751), .Z(n7039) );
  INV_X1 U8750 ( .A(n7187), .ZN(n7189) );
  AOI211_X1 U8751 ( .C1(n7219), .C2(n7243), .A(n9793), .B(n7189), .ZN(n7128)
         );
  OR2_X1 U8752 ( .A1(n7035), .A2(n9156), .ZN(n7793) );
  INV_X1 U8753 ( .A(n7793), .ZN(n9591) );
  INV_X1 U8754 ( .A(n7219), .ZN(n7036) );
  OAI22_X1 U8755 ( .A1(n9396), .A2(n7036), .B1(n7216), .B2(n9743), .ZN(n7037)
         );
  AOI21_X1 U8756 ( .B1(n7128), .B2(n9591), .A(n7037), .ZN(n7038) );
  OAI211_X1 U8757 ( .C1(n7131), .C2(n9408), .A(n7039), .B(n7038), .ZN(P1_U3284) );
  XNOR2_X1 U8758 ( .A(n7040), .B(n7041), .ZN(n9902) );
  XNOR2_X1 U8759 ( .A(n7054), .B(n9896), .ZN(n7043) );
  NAND2_X1 U8760 ( .A1(n7043), .A2(n9841), .ZN(n9903) );
  OAI22_X1 U8761 ( .A1(n9847), .A2(n9903), .B1(n10120), .B2(n9845), .ZN(n7044)
         );
  AOI21_X1 U8762 ( .B1(n8534), .B2(n7054), .A(n7044), .ZN(n7051) );
  XNOR2_X1 U8763 ( .A(n7045), .B(n7040), .ZN(n7048) );
  OAI22_X1 U8764 ( .A1(n7047), .A2(n9812), .B1(n7046), .B2(n9814), .ZN(n8088)
         );
  AOI21_X1 U8765 ( .B1(n7048), .B2(n9838), .A(n8088), .ZN(n9904) );
  MUX2_X1 U8766 ( .A(n9904), .B(n7049), .S(n9849), .Z(n7050) );
  OAI211_X1 U8767 ( .C1(n9902), .C2(n8506), .A(n7051), .B(n7050), .ZN(P2_U3295) );
  XOR2_X1 U8768 ( .A(n7905), .B(n7052), .Z(n9909) );
  OAI21_X1 U8769 ( .B1(n7054), .B2(n7053), .A(n7057), .ZN(n7055) );
  NAND3_X1 U8770 ( .A1(n7088), .A2(n9841), .A3(n7055), .ZN(n9910) );
  OAI22_X1 U8771 ( .A1(n9847), .A2(n9910), .B1(n10319), .B2(n9845), .ZN(n7056)
         );
  AOI21_X1 U8772 ( .B1(n8534), .B2(n7057), .A(n7056), .ZN(n7063) );
  XNOR2_X1 U8773 ( .A(n7058), .B(n7905), .ZN(n7060) );
  AOI21_X1 U8774 ( .B1(n7060), .B2(n9838), .A(n7059), .ZN(n9911) );
  MUX2_X1 U8775 ( .A(n7061), .B(n9911), .S(n8553), .Z(n7062) );
  OAI211_X1 U8776 ( .C1(n9909), .C2(n8506), .A(n7063), .B(n7062), .ZN(P2_U3294) );
  INV_X1 U8777 ( .A(n8321), .ZN(n8303) );
  INV_X1 U8778 ( .A(n7064), .ZN(n7078) );
  INV_X1 U8779 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7065) );
  OAI222_X1 U8780 ( .A1(P2_U3152), .A2(n8303), .B1(n8696), .B2(n7078), .C1(
        n7065), .C2(n8694), .ZN(P2_U3341) );
  OAI21_X1 U8781 ( .B1(n7068), .B2(n7067), .A(n7066), .ZN(n7076) );
  NAND2_X1 U8782 ( .A1(n9730), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n7069) );
  NAND2_X1 U8783 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3084), .ZN(n7730) );
  OAI211_X1 U8784 ( .C1(n9724), .C2(n7070), .A(n7069), .B(n7730), .ZN(n7075)
         );
  AOI211_X1 U8785 ( .C1(n7073), .C2(n7072), .A(n9690), .B(n7071), .ZN(n7074)
         );
  AOI211_X1 U8786 ( .C1(n9731), .C2(n7076), .A(n7075), .B(n7074), .ZN(n7077)
         );
  INV_X1 U8787 ( .A(n7077), .ZN(P1_U3254) );
  INV_X1 U8788 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7079) );
  INV_X1 U8789 ( .A(n9145), .ZN(n7671) );
  OAI222_X1 U8790 ( .A1(n9522), .A2(n7079), .B1(n7671), .B2(P1_U3084), .C1(
        n9513), .C2(n7078), .ZN(P1_U3336) );
  AOI21_X1 U8791 ( .B1(n7081), .B2(n7080), .A(n4548), .ZN(n7086) );
  AOI22_X1 U8792 ( .A1(n4473), .A2(n9139), .B1(n8811), .B2(n9137), .ZN(n7085)
         );
  NOR2_X1 U8793 ( .A1(n8822), .A2(n9742), .ZN(n7082) );
  AOI211_X1 U8794 ( .C1(n9739), .C2(n8828), .A(n7083), .B(n7082), .ZN(n7084)
         );
  OAI211_X1 U8795 ( .C1(n7086), .C2(n8831), .A(n7085), .B(n7084), .ZN(P1_U3225) );
  XNOR2_X1 U8796 ( .A(n7087), .B(n7095), .ZN(n9922) );
  NAND2_X1 U8797 ( .A1(n7088), .A2(n9917), .ZN(n7089) );
  NAND2_X1 U8798 ( .A1(n7089), .A2(n9841), .ZN(n7090) );
  NOR2_X1 U8799 ( .A1(n9842), .A2(n7090), .ZN(n9916) );
  NAND2_X1 U8800 ( .A1(n8556), .A2(n9916), .ZN(n7092) );
  NAND2_X1 U8801 ( .A1(n9849), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7091) );
  OAI211_X1 U8802 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9845), .A(n7092), .B(
        n7091), .ZN(n7099) );
  OAI21_X1 U8803 ( .B1(n7095), .B2(n7094), .A(n7093), .ZN(n7097) );
  AOI21_X1 U8804 ( .B1(n7097), .B2(n9838), .A(n7096), .ZN(n9920) );
  NOR2_X1 U8805 ( .A1(n9920), .A2(n9849), .ZN(n7098) );
  AOI211_X1 U8806 ( .C1(n8534), .C2(n9917), .A(n7099), .B(n7098), .ZN(n7100)
         );
  OAI21_X1 U8807 ( .B1(n8506), .B2(n9922), .A(n7100), .ZN(P2_U3293) );
  NOR2_X1 U8808 ( .A1(n7107), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7102) );
  NOR2_X1 U8809 ( .A1(n7102), .A2(n7101), .ZN(n7105) );
  MUX2_X1 U8810 ( .A(n7542), .B(P2_REG2_REG_12__SCAN_IN), .S(n7201), .Z(n7103)
         );
  INV_X1 U8811 ( .A(n7103), .ZN(n7104) );
  NAND2_X1 U8812 ( .A1(n7104), .A2(n7105), .ZN(n7196) );
  OAI211_X1 U8813 ( .C1(n7105), .C2(n7104), .A(n9825), .B(n7196), .ZN(n7116)
         );
  MUX2_X1 U8814 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7108), .S(n7201), .Z(n7109)
         );
  OAI21_X1 U8815 ( .B1(n7110), .B2(n7109), .A(n7200), .ZN(n7114) );
  NOR2_X1 U8816 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10257), .ZN(n7113) );
  INV_X1 U8817 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7111) );
  NOR2_X1 U8818 ( .A1(n9537), .A2(n7111), .ZN(n7112) );
  AOI211_X1 U8819 ( .C1(n9827), .C2(n7114), .A(n7113), .B(n7112), .ZN(n7115)
         );
  OAI211_X1 U8820 ( .C1(n9828), .C2(n7117), .A(n7116), .B(n7115), .ZN(P2_U3257) );
  INV_X1 U8821 ( .A(n9743), .ZN(n9583) );
  AOI22_X1 U8822 ( .A1(n9585), .A2(n7119), .B1(n9583), .B2(n7118), .ZN(n7120)
         );
  OAI21_X1 U8823 ( .B1(n9225), .B2(n7121), .A(n7120), .ZN(n7124) );
  MUX2_X1 U8824 ( .A(n7122), .B(P1_REG2_REG_3__SCAN_IN), .S(n9753), .Z(n7123)
         );
  AOI211_X1 U8825 ( .C1(n9592), .C2(n7125), .A(n7124), .B(n7123), .ZN(n7126)
         );
  INV_X1 U8826 ( .A(n7126), .ZN(P1_U3288) );
  INV_X1 U8827 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7133) );
  NAND2_X1 U8828 ( .A1(n7127), .A2(n9490), .ZN(n9788) );
  AOI21_X1 U8829 ( .B1(n9487), .B2(n7219), .A(n7128), .ZN(n7129) );
  OAI211_X1 U8830 ( .C1(n7131), .C2(n9484), .A(n7130), .B(n7129), .ZN(n7164)
         );
  NAND2_X1 U8831 ( .A1(n7164), .A2(n9800), .ZN(n7132) );
  OAI21_X1 U8832 ( .B1(n9800), .B2(n7133), .A(n7132), .ZN(P1_U3475) );
  NAND2_X1 U8833 ( .A1(n7136), .A2(n7135), .ZN(n7137) );
  XNOR2_X1 U8834 ( .A(n7134), .B(n7137), .ZN(n7143) );
  OAI22_X1 U8835 ( .A1(n8824), .A2(n7138), .B1(n8822), .B2(n7244), .ZN(n7139)
         );
  AOI211_X1 U8836 ( .C1(n4473), .C2(n9138), .A(n7140), .B(n7139), .ZN(n7142)
         );
  NAND2_X1 U8837 ( .A1(n8828), .A2(n7246), .ZN(n7141) );
  OAI211_X1 U8838 ( .C1(n7143), .C2(n8831), .A(n7142), .B(n7141), .ZN(P1_U3237) );
  INV_X1 U8839 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7161) );
  NAND2_X1 U8840 ( .A1(n7145), .A2(n7144), .ZN(n7146) );
  AND2_X1 U8841 ( .A1(n5019), .A2(n7146), .ZN(n9736) );
  OAI211_X1 U8842 ( .C1(n7147), .C2(n7148), .A(n7241), .B(n9764), .ZN(n9737)
         );
  NAND2_X1 U8843 ( .A1(n9137), .A2(n9400), .ZN(n9741) );
  OAI211_X1 U8844 ( .C1(n7148), .C2(n9791), .A(n9737), .B(n9741), .ZN(n7159)
         );
  INV_X1 U8845 ( .A(n7149), .ZN(n7150) );
  OR2_X1 U8846 ( .A1(n7151), .A2(n7150), .ZN(n7154) );
  AND2_X1 U8847 ( .A1(n7153), .A2(n9083), .ZN(n9058) );
  AND2_X1 U8848 ( .A1(n9058), .A2(n9089), .ZN(n7152) );
  NAND2_X1 U8849 ( .A1(n7154), .A2(n7152), .ZN(n7155) );
  NAND2_X1 U8850 ( .A1(n7155), .A2(n9089), .ZN(n8933) );
  INV_X1 U8851 ( .A(n7153), .ZN(n8936) );
  NAND3_X1 U8852 ( .A1(n7155), .A2(n9083), .A3(n7154), .ZN(n7156) );
  OAI211_X1 U8853 ( .C1(n8933), .C2(n8936), .A(n7156), .B(n9574), .ZN(n7158)
         );
  NAND2_X1 U8854 ( .A1(n9139), .A2(n9329), .ZN(n7157) );
  NAND2_X1 U8855 ( .A1(n7158), .A2(n7157), .ZN(n9749) );
  AOI211_X1 U8856 ( .C1(n9736), .C2(n9788), .A(n7159), .B(n9749), .ZN(n7162)
         );
  OR2_X1 U8857 ( .A1(n7162), .A2(n9799), .ZN(n7160) );
  OAI21_X1 U8858 ( .B1(n9800), .B2(n7161), .A(n7160), .ZN(P1_U3469) );
  OR2_X1 U8859 ( .A1(n7162), .A2(n9806), .ZN(n7163) );
  OAI21_X1 U8860 ( .B1(n9809), .B2(n6555), .A(n7163), .ZN(P1_U3528) );
  NAND2_X1 U8861 ( .A1(n7164), .A2(n9809), .ZN(n7165) );
  OAI21_X1 U8862 ( .B1(n9809), .B2(n6564), .A(n7165), .ZN(P1_U3530) );
  XOR2_X1 U8863 ( .A(n7167), .B(n7166), .Z(n7175) );
  OR2_X1 U8864 ( .A1(n7261), .A2(n9814), .ZN(n7170) );
  OR2_X1 U8865 ( .A1(n7168), .A2(n9812), .ZN(n7169) );
  NAND2_X1 U8866 ( .A1(n7170), .A2(n7169), .ZN(n7277) );
  AOI21_X1 U8867 ( .B1(n9817), .B2(n7277), .A(n7171), .ZN(n7173) );
  OR2_X1 U8868 ( .A1(n9824), .A2(n7280), .ZN(n7172) );
  OAI211_X1 U8869 ( .C1(n7301), .C2(n9819), .A(n7173), .B(n7172), .ZN(n7174)
         );
  AOI21_X1 U8870 ( .B1(n7175), .B2(n9821), .A(n7174), .ZN(n7176) );
  INV_X1 U8871 ( .A(n7176), .ZN(P2_U3229) );
  INV_X1 U8872 ( .A(n9135), .ZN(n7217) );
  NAND2_X1 U8873 ( .A1(n7436), .A2(n7217), .ZN(n8954) );
  OR2_X1 U8874 ( .A1(n7219), .A2(n9136), .ZN(n7177) );
  INV_X1 U8875 ( .A(n7394), .ZN(n7179) );
  AOI21_X1 U8876 ( .B1(n9063), .B2(n7180), .A(n7179), .ZN(n9789) );
  INV_X1 U8877 ( .A(n9789), .ZN(n7195) );
  INV_X1 U8878 ( .A(n8957), .ZN(n8899) );
  INV_X1 U8879 ( .A(n9063), .ZN(n7182) );
  AOI21_X1 U8880 ( .B1(n7183), .B2(n7182), .A(n7853), .ZN(n7184) );
  OAI21_X1 U8881 ( .B1(n7395), .B2(n8899), .A(n7184), .ZN(n7186) );
  AOI22_X1 U8882 ( .A1(n9329), .A2(n9136), .B1(n9577), .B2(n9400), .ZN(n7185)
         );
  NAND2_X1 U8883 ( .A1(n7186), .A2(n7185), .ZN(n9787) );
  INV_X1 U8884 ( .A(n7436), .ZN(n9784) );
  INV_X1 U8885 ( .A(n7400), .ZN(n7188) );
  OAI21_X1 U8886 ( .B1(n9784), .B2(n7189), .A(n7188), .ZN(n9785) );
  OAI22_X1 U8887 ( .A1(n9751), .A2(n7190), .B1(n7432), .B2(n9743), .ZN(n7191)
         );
  AOI21_X1 U8888 ( .B1(n9585), .B2(n7436), .A(n7191), .ZN(n7192) );
  OAI21_X1 U8889 ( .B1(n9785), .B2(n9225), .A(n7192), .ZN(n7193) );
  AOI21_X1 U8890 ( .B1(n9787), .B2(n9751), .A(n7193), .ZN(n7194) );
  OAI21_X1 U8891 ( .B1(n7195), .B2(n9408), .A(n7194), .ZN(P1_U3283) );
  NAND2_X1 U8892 ( .A1(n7201), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7197) );
  NAND2_X1 U8893 ( .A1(n7197), .A2(n7196), .ZN(n7199) );
  AOI22_X1 U8894 ( .A1(n7335), .A2(n7716), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7331), .ZN(n7198) );
  NOR2_X1 U8895 ( .A1(n7199), .A2(n7198), .ZN(n7330) );
  AOI21_X1 U8896 ( .B1(n7199), .B2(n7198), .A(n7330), .ZN(n7209) );
  AOI22_X1 U8897 ( .A1(n7335), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n5342), .B2(
        n7331), .ZN(n7203) );
  OAI21_X1 U8898 ( .B1(n7203), .B2(n7202), .A(n7334), .ZN(n7204) );
  NAND2_X1 U8899 ( .A1(n7204), .A2(n9827), .ZN(n7208) );
  NOR2_X1 U8900 ( .A1(n7205), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7841) );
  NOR2_X1 U8901 ( .A1(n9828), .A2(n7331), .ZN(n7206) );
  AOI211_X1 U8902 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n9832), .A(n7841), .B(
        n7206), .ZN(n7207) );
  OAI211_X1 U8903 ( .C1(n7209), .C2(n9830), .A(n7208), .B(n7207), .ZN(P2_U3258) );
  INV_X1 U8904 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7211) );
  INV_X1 U8905 ( .A(n7210), .ZN(n7212) );
  INV_X1 U8906 ( .A(n8332), .ZN(n8319) );
  OAI222_X1 U8907 ( .A1(n8694), .A2(n7211), .B1(n8696), .B2(n7212), .C1(
        P2_U3152), .C2(n8319), .ZN(P2_U3340) );
  INV_X1 U8908 ( .A(n9148), .ZN(n9725) );
  OAI222_X1 U8909 ( .A1(n9522), .A2(n10149), .B1(n9513), .B2(n7212), .C1(
        P1_U3084), .C2(n9725), .ZN(P1_U3335) );
  XOR2_X1 U8910 ( .A(n7213), .B(n7214), .Z(n7222) );
  INV_X1 U8911 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7215) );
  NOR2_X1 U8912 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7215), .ZN(n9669) );
  OAI22_X1 U8913 ( .A1(n8824), .A2(n7217), .B1(n8822), .B2(n7216), .ZN(n7218)
         );
  AOI211_X1 U8914 ( .C1(n4473), .C2(n9137), .A(n9669), .B(n7218), .ZN(n7221)
         );
  NAND2_X1 U8915 ( .A1(n8828), .A2(n7219), .ZN(n7220) );
  OAI211_X1 U8916 ( .C1(n7222), .C2(n8831), .A(n7221), .B(n7220), .ZN(P1_U3211) );
  XNOR2_X1 U8917 ( .A(n7223), .B(n7908), .ZN(n7311) );
  INV_X1 U8918 ( .A(n7311), .ZN(n7238) );
  AND2_X1 U8919 ( .A1(n7225), .A2(n7224), .ZN(n7227) );
  XNOR2_X1 U8920 ( .A(n7227), .B(n7226), .ZN(n7231) );
  OR2_X1 U8921 ( .A1(n7345), .A2(n9814), .ZN(n7229) );
  NAND2_X1 U8922 ( .A1(n8270), .A2(n8228), .ZN(n7228) );
  NAND2_X1 U8923 ( .A1(n7229), .A2(n7228), .ZN(n7322) );
  INV_X1 U8924 ( .A(n7322), .ZN(n7230) );
  OAI21_X1 U8925 ( .B1(n7231), .B2(n8527), .A(n7230), .ZN(n7309) );
  INV_X1 U8926 ( .A(n7309), .ZN(n7232) );
  MUX2_X1 U8927 ( .A(n7233), .B(n7232), .S(n8553), .Z(n7237) );
  AOI21_X1 U8928 ( .B1(n7279), .B2(n7312), .A(n9942), .ZN(n7234) );
  AND2_X1 U8929 ( .A1(n7234), .A2(n7256), .ZN(n7310) );
  OAI22_X1 U8930 ( .A1(n9851), .A2(n7325), .B1(n9845), .B2(n7320), .ZN(n7235)
         );
  AOI21_X1 U8931 ( .B1(n8556), .B2(n7310), .A(n7235), .ZN(n7236) );
  OAI211_X1 U8932 ( .C1(n8506), .C2(n7238), .A(n7237), .B(n7236), .ZN(P2_U3290) );
  OAI21_X1 U8933 ( .B1(n7240), .B2(n8932), .A(n7239), .ZN(n9783) );
  NAND2_X1 U8934 ( .A1(n7241), .A2(n7246), .ZN(n7242) );
  NAND2_X1 U8935 ( .A1(n7243), .A2(n7242), .ZN(n9780) );
  INV_X1 U8936 ( .A(n7244), .ZN(n7245) );
  AOI22_X1 U8937 ( .A1(n9585), .A2(n7246), .B1(n7245), .B2(n9583), .ZN(n7247)
         );
  OAI21_X1 U8938 ( .B1(n9780), .B2(n9225), .A(n7247), .ZN(n7252) );
  XNOR2_X1 U8939 ( .A(n8933), .B(n8932), .ZN(n7250) );
  NAND2_X1 U8940 ( .A1(n9783), .A2(n9581), .ZN(n7249) );
  AOI22_X1 U8941 ( .A1(n9348), .A2(n9136), .B1(n9138), .B2(n9329), .ZN(n7248)
         );
  OAI211_X1 U8942 ( .C1(n7853), .C2(n7250), .A(n7249), .B(n7248), .ZN(n9781)
         );
  MUX2_X1 U8943 ( .A(n9781), .B(P1_REG2_REG_6__SCAN_IN), .S(n9753), .Z(n7251)
         );
  AOI211_X1 U8944 ( .C1(n9592), .C2(n9783), .A(n7252), .B(n7251), .ZN(n7253)
         );
  INV_X1 U8945 ( .A(n7253), .ZN(P1_U3285) );
  XOR2_X1 U8946 ( .A(n7254), .B(n7957), .Z(n7288) );
  AOI21_X1 U8947 ( .B1(n7256), .B2(n7255), .A(n9942), .ZN(n7257) );
  NAND2_X1 U8948 ( .A1(n7257), .A2(n7355), .ZN(n7286) );
  INV_X1 U8949 ( .A(n7286), .ZN(n7259) );
  OAI22_X1 U8950 ( .A1(n9851), .A2(n7411), .B1(n7414), .B2(n9845), .ZN(n7258)
         );
  AOI21_X1 U8951 ( .B1(n7259), .B2(n8556), .A(n7258), .ZN(n7267) );
  XNOR2_X1 U8952 ( .A(n7260), .B(n7957), .ZN(n7264) );
  OR2_X1 U8953 ( .A1(n7261), .A2(n9812), .ZN(n7263) );
  OR2_X1 U8954 ( .A1(n7367), .A2(n9814), .ZN(n7262) );
  NAND2_X1 U8955 ( .A1(n7263), .A2(n7262), .ZN(n7410) );
  AOI21_X1 U8956 ( .B1(n7264), .B2(n9838), .A(n7410), .ZN(n7287) );
  MUX2_X1 U8957 ( .A(n7287), .B(n7265), .S(n9849), .Z(n7266) );
  OAI211_X1 U8958 ( .C1(n7288), .C2(n8506), .A(n7267), .B(n7266), .ZN(P2_U3289) );
  NAND2_X1 U8959 ( .A1(n7930), .A2(n7951), .ZN(n7906) );
  NAND2_X1 U8960 ( .A1(n7268), .A2(n9840), .ZN(n7270) );
  NAND2_X1 U8961 ( .A1(n7270), .A2(n7269), .ZN(n7271) );
  XOR2_X1 U8962 ( .A(n7906), .B(n7271), .Z(n7297) );
  INV_X1 U8963 ( .A(n7273), .ZN(n7929) );
  OR2_X1 U8964 ( .A1(n7272), .A2(n7929), .ZN(n7275) );
  NAND2_X1 U8965 ( .A1(n7275), .A2(n7274), .ZN(n7276) );
  XNOR2_X1 U8966 ( .A(n7276), .B(n7906), .ZN(n7278) );
  AOI21_X1 U8967 ( .B1(n7278), .B2(n9838), .A(n7277), .ZN(n7296) );
  INV_X1 U8968 ( .A(n7296), .ZN(n7282) );
  OAI211_X1 U8969 ( .C1(n9843), .C2(n7301), .A(n9841), .B(n7279), .ZN(n7295)
         );
  OAI22_X1 U8970 ( .A1(n7295), .A2(n7923), .B1(n9845), .B2(n7280), .ZN(n7281)
         );
  OAI21_X1 U8971 ( .B1(n7282), .B2(n7281), .A(n8553), .ZN(n7285) );
  AOI22_X1 U8972 ( .A1(n8534), .A2(n7283), .B1(n9849), .B2(
        P2_REG2_REG_5__SCAN_IN), .ZN(n7284) );
  OAI211_X1 U8973 ( .C1(n7297), .C2(n8506), .A(n7285), .B(n7284), .ZN(P2_U3291) );
  OAI211_X1 U8974 ( .C1(n7288), .C2(n9898), .A(n7287), .B(n7286), .ZN(n7293)
         );
  OAI22_X1 U8975 ( .A1(n8634), .A2(n7411), .B1(n9960), .B2(n5186), .ZN(n7289)
         );
  AOI21_X1 U8976 ( .B1(n7293), .B2(n9960), .A(n7289), .ZN(n7290) );
  INV_X1 U8977 ( .A(n7290), .ZN(P2_U3527) );
  INV_X1 U8978 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7291) );
  OAI22_X1 U8979 ( .A1(n8677), .A2(n7411), .B1(n9949), .B2(n7291), .ZN(n7292)
         );
  AOI21_X1 U8980 ( .B1(n7293), .B2(n9949), .A(n7292), .ZN(n7294) );
  INV_X1 U8981 ( .A(n7294), .ZN(P2_U3472) );
  OAI211_X1 U8982 ( .C1(n7297), .C2(n9898), .A(n7296), .B(n7295), .ZN(n7303)
         );
  INV_X1 U8983 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7298) );
  OAI22_X1 U8984 ( .A1(n8634), .A2(n7301), .B1(n9960), .B2(n7298), .ZN(n7299)
         );
  AOI21_X1 U8985 ( .B1(n7303), .B2(n9960), .A(n7299), .ZN(n7300) );
  INV_X1 U8986 ( .A(n7300), .ZN(P2_U3525) );
  OAI22_X1 U8987 ( .A1(n8677), .A2(n7301), .B1(n9949), .B2(n5144), .ZN(n7302)
         );
  AOI21_X1 U8988 ( .B1(n7303), .B2(n9949), .A(n7302), .ZN(n7304) );
  INV_X1 U8989 ( .A(n7304), .ZN(P2_U3466) );
  INV_X1 U8990 ( .A(n7305), .ZN(n7307) );
  OAI222_X1 U8991 ( .A1(n8694), .A2(n7306), .B1(n8696), .B2(n7307), .C1(
        P2_U3152), .C2(n8530), .ZN(P2_U3339) );
  OAI222_X1 U8992 ( .A1(n9522), .A2(n7308), .B1(n9513), .B2(n7307), .C1(
        P1_U3084), .C2(n9745), .ZN(P1_U3334) );
  AOI211_X1 U8993 ( .C1(n7311), .C2(n9946), .A(n7310), .B(n7309), .ZN(n7317)
         );
  INV_X1 U8994 ( .A(n9960), .ZN(n9958) );
  AOI22_X1 U8995 ( .A1(n6508), .A2(n7312), .B1(n9958), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n7313) );
  OAI21_X1 U8996 ( .B1(n7317), .B2(n9958), .A(n7313), .ZN(P2_U3526) );
  INV_X1 U8997 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7314) );
  OAI22_X1 U8998 ( .A1(n8677), .A2(n7325), .B1(n9949), .B2(n7314), .ZN(n7315)
         );
  INV_X1 U8999 ( .A(n7315), .ZN(n7316) );
  OAI21_X1 U9000 ( .B1(n7317), .B2(n9948), .A(n7316), .ZN(P2_U3469) );
  AOI21_X1 U9001 ( .B1(n7319), .B2(n7318), .A(n4550), .ZN(n7329) );
  INV_X1 U9002 ( .A(n7320), .ZN(n7327) );
  INV_X1 U9003 ( .A(n7321), .ZN(n7324) );
  NAND2_X1 U9004 ( .A1(n9817), .A2(n7322), .ZN(n7323) );
  OAI211_X1 U9005 ( .C1(n9819), .C2(n7325), .A(n7324), .B(n7323), .ZN(n7326)
         );
  AOI21_X1 U9006 ( .B1(n7327), .B2(n8231), .A(n7326), .ZN(n7328) );
  OAI21_X1 U9007 ( .B1(n7329), .B2(n8247), .A(n7328), .ZN(P2_U3241) );
  AOI21_X1 U9008 ( .B1(n7331), .B2(n7716), .A(n7330), .ZN(n7333) );
  AOI22_X1 U9009 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7339), .B1(n7592), .B2(
        n7761), .ZN(n7332) );
  NOR2_X1 U9010 ( .A1(n7333), .A2(n7332), .ZN(n7593) );
  AOI21_X1 U9011 ( .B1(n7333), .B2(n7332), .A(n7593), .ZN(n7343) );
  AOI22_X1 U9012 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7592), .B1(n7339), .B2(
        n5367), .ZN(n7337) );
  OAI21_X1 U9013 ( .B1(n7335), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7334), .ZN(
        n7336) );
  OAI21_X1 U9014 ( .B1(n7337), .B2(n7336), .A(n7590), .ZN(n7338) );
  NAND2_X1 U9015 ( .A1(n7338), .A2(n9827), .ZN(n7342) );
  NOR2_X1 U9016 ( .A1(n10260), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8115) );
  NOR2_X1 U9017 ( .A1(n9828), .A2(n7339), .ZN(n7340) );
  AOI211_X1 U9018 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n9832), .A(n8115), .B(
        n7340), .ZN(n7341) );
  OAI211_X1 U9019 ( .C1(n7343), .C2(n9830), .A(n7342), .B(n7341), .ZN(P2_U3259) );
  XNOR2_X1 U9020 ( .A(n7344), .B(n7962), .ZN(n7349) );
  OR2_X1 U9021 ( .A1(n7345), .A2(n9812), .ZN(n7347) );
  OR2_X1 U9022 ( .A1(n7472), .A2(n9814), .ZN(n7346) );
  NAND2_X1 U9023 ( .A1(n7347), .A2(n7346), .ZN(n7496) );
  INV_X1 U9024 ( .A(n7496), .ZN(n7348) );
  OAI21_X1 U9025 ( .B1(n7349), .B2(n8527), .A(n7348), .ZN(n7418) );
  INV_X1 U9026 ( .A(n7418), .ZN(n7362) );
  OR2_X1 U9027 ( .A1(n7254), .A2(n7957), .ZN(n7352) );
  NAND2_X1 U9028 ( .A1(n7352), .A2(n7350), .ZN(n7354) );
  AND2_X1 U9029 ( .A1(n7352), .A2(n7351), .ZN(n7353) );
  AOI21_X1 U9030 ( .B1(n7962), .B2(n7354), .A(n7353), .ZN(n7420) );
  NAND2_X1 U9031 ( .A1(n7420), .A2(n9853), .ZN(n7361) );
  NAND2_X1 U9032 ( .A1(n7355), .A2(n7421), .ZN(n7356) );
  NAND2_X1 U9033 ( .A1(n7356), .A2(n9841), .ZN(n7357) );
  NOR2_X1 U9034 ( .A1(n7374), .A2(n7357), .ZN(n7419) );
  NOR2_X1 U9035 ( .A1(n9851), .A2(n7500), .ZN(n7359) );
  OAI22_X1 U9036 ( .A1(n8553), .A2(n6745), .B1(n7497), .B2(n9845), .ZN(n7358)
         );
  AOI211_X1 U9037 ( .C1(n7419), .C2(n8556), .A(n7359), .B(n7358), .ZN(n7360)
         );
  OAI211_X1 U9038 ( .C1(n9855), .C2(n7362), .A(n7361), .B(n7360), .ZN(P2_U3288) );
  OAI21_X1 U9039 ( .B1(n7364), .B2(n7910), .A(n7363), .ZN(n9936) );
  INV_X1 U9040 ( .A(n8547), .ZN(n9925) );
  NAND2_X1 U9041 ( .A1(n9936), .A2(n9925), .ZN(n7372) );
  INV_X1 U9042 ( .A(n7910), .ZN(n7365) );
  XNOR2_X1 U9043 ( .A(n7366), .B(n7365), .ZN(n7370) );
  OR2_X1 U9044 ( .A1(n7367), .A2(n9812), .ZN(n7369) );
  NAND2_X1 U9045 ( .A1(n8265), .A2(n8218), .ZN(n7368) );
  NAND2_X1 U9046 ( .A1(n7369), .A2(n7368), .ZN(n7551) );
  AOI21_X1 U9047 ( .B1(n7370), .B2(n9838), .A(n7551), .ZN(n7371) );
  AND2_X1 U9048 ( .A1(n7372), .A2(n7371), .ZN(n9938) );
  OR2_X1 U9049 ( .A1(n9855), .A2(n7373), .ZN(n8559) );
  INV_X1 U9050 ( .A(n8559), .ZN(n7380) );
  OAI211_X1 U9051 ( .C1(n7374), .C2(n9933), .A(n7477), .B(n9841), .ZN(n9932)
         );
  OAI22_X1 U9052 ( .A1(n8553), .A2(n7375), .B1(n7554), .B2(n9845), .ZN(n7376)
         );
  AOI21_X1 U9053 ( .B1(n8534), .B2(n7377), .A(n7376), .ZN(n7378) );
  OAI21_X1 U9054 ( .B1(n9932), .B2(n9847), .A(n7378), .ZN(n7379) );
  AOI21_X1 U9055 ( .B1(n9936), .B2(n7380), .A(n7379), .ZN(n7381) );
  OAI21_X1 U9056 ( .B1(n9938), .B2(n9855), .A(n7381), .ZN(P2_U3287) );
  INV_X1 U9057 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7392) );
  OAI21_X1 U9058 ( .B1(n7384), .B2(n7383), .A(n7382), .ZN(n7385) );
  NAND2_X1 U9059 ( .A1(n7385), .A2(n9731), .ZN(n7391) );
  AND2_X1 U9060 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8707) );
  AOI211_X1 U9061 ( .C1(n6091), .C2(n7387), .A(n7386), .B(n9690), .ZN(n7388)
         );
  AOI211_X1 U9062 ( .C1(n9705), .C2(n7389), .A(n8707), .B(n7388), .ZN(n7390)
         );
  OAI211_X1 U9063 ( .C1(n9717), .C2(n7392), .A(n7391), .B(n7390), .ZN(P1_U3255) );
  NAND2_X1 U9064 ( .A1(n7436), .A2(n9135), .ZN(n7393) );
  NAND2_X1 U9065 ( .A1(n7394), .A2(n7393), .ZN(n7455) );
  INV_X1 U9066 ( .A(n9577), .ZN(n7433) );
  OR2_X1 U9067 ( .A1(n7453), .A2(n7433), .ZN(n9570) );
  NAND2_X1 U9068 ( .A1(n7453), .A2(n7433), .ZN(n8955) );
  NAND2_X1 U9069 ( .A1(n9570), .A2(n8955), .ZN(n9065) );
  XNOR2_X1 U9070 ( .A(n7455), .B(n9568), .ZN(n9797) );
  INV_X1 U9071 ( .A(n9797), .ZN(n7406) );
  XNOR2_X1 U9072 ( .A(n9569), .B(n9568), .ZN(n7398) );
  NAND2_X1 U9073 ( .A1(n9797), .A2(n9581), .ZN(n7397) );
  AOI22_X1 U9074 ( .A1(n9348), .A2(n9134), .B1(n9135), .B2(n9578), .ZN(n7396)
         );
  OAI211_X1 U9075 ( .C1(n7853), .C2(n7398), .A(n7397), .B(n7396), .ZN(n9795)
         );
  NAND2_X1 U9076 ( .A1(n9795), .A2(n9751), .ZN(n7405) );
  INV_X1 U9077 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7399) );
  OAI22_X1 U9078 ( .A1(n9751), .A2(n7399), .B1(n7447), .B2(n9743), .ZN(n7403)
         );
  INV_X1 U9079 ( .A(n7453), .ZN(n9792) );
  OR2_X1 U9080 ( .A1(n7400), .A2(n9792), .ZN(n7401) );
  NAND2_X1 U9081 ( .A1(n9586), .A2(n7401), .ZN(n9794) );
  NOR2_X1 U9082 ( .A1(n9794), .A2(n9225), .ZN(n7402) );
  AOI211_X1 U9083 ( .C1(n9585), .C2(n7453), .A(n7403), .B(n7402), .ZN(n7404)
         );
  OAI211_X1 U9084 ( .C1(n7406), .C2(n7661), .A(n7405), .B(n7404), .ZN(P1_U3282) );
  XOR2_X1 U9085 ( .A(n7408), .B(n7407), .Z(n7416) );
  AOI21_X1 U9086 ( .B1(n9817), .B2(n7410), .A(n7409), .ZN(n7413) );
  OR2_X1 U9087 ( .A1(n9819), .A2(n7411), .ZN(n7412) );
  OAI211_X1 U9088 ( .C1(n9824), .C2(n7414), .A(n7413), .B(n7412), .ZN(n7415)
         );
  AOI21_X1 U9089 ( .B1(n7416), .B2(n9821), .A(n7415), .ZN(n7417) );
  INV_X1 U9090 ( .A(n7417), .ZN(P2_U3215) );
  AOI211_X1 U9091 ( .C1(n7420), .C2(n9946), .A(n7419), .B(n7418), .ZN(n7425)
         );
  AOI22_X1 U9092 ( .A1(n6508), .A2(n7421), .B1(n9958), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n7422) );
  OAI21_X1 U9093 ( .B1(n7425), .B2(n9958), .A(n7422), .ZN(P2_U3528) );
  OAI22_X1 U9094 ( .A1(n8677), .A2(n7500), .B1(n9949), .B2(n5211), .ZN(n7423)
         );
  INV_X1 U9095 ( .A(n7423), .ZN(n7424) );
  OAI21_X1 U9096 ( .B1(n7425), .B2(n9948), .A(n7424), .ZN(P2_U3475) );
  INV_X1 U9097 ( .A(n7426), .ZN(n7440) );
  OAI222_X1 U9098 ( .A1(n9513), .A2(n7440), .B1(n4672), .B2(P1_U3084), .C1(
        n7427), .C2(n9522), .ZN(P1_U3333) );
  NAND2_X1 U9099 ( .A1(n7429), .A2(n7428), .ZN(n7430) );
  XOR2_X1 U9100 ( .A(n7431), .B(n7430), .Z(n7439) );
  NAND2_X1 U9101 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9688) );
  INV_X1 U9102 ( .A(n9688), .ZN(n7435) );
  OAI22_X1 U9103 ( .A1(n8824), .A2(n7433), .B1(n8822), .B2(n7432), .ZN(n7434)
         );
  AOI211_X1 U9104 ( .C1(n4473), .C2(n9136), .A(n7435), .B(n7434), .ZN(n7438)
         );
  NAND2_X1 U9105 ( .A1(n8828), .A2(n7436), .ZN(n7437) );
  OAI211_X1 U9106 ( .C1(n7439), .C2(n8831), .A(n7438), .B(n7437), .ZN(P1_U3219) );
  OAI222_X1 U9107 ( .A1(n8694), .A2(n7441), .B1(n8696), .B2(n7440), .C1(n8072), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  INV_X1 U9108 ( .A(n8828), .ZN(n8758) );
  OAI21_X1 U9109 ( .B1(n7444), .B2(n7442), .A(n7443), .ZN(n7445) );
  NAND2_X1 U9110 ( .A1(n7445), .A2(n8808), .ZN(n7450) );
  NOR2_X1 U9111 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7446), .ZN(n9695) );
  INV_X1 U9112 ( .A(n9134), .ZN(n7456) );
  OAI22_X1 U9113 ( .A1(n8824), .A2(n7456), .B1(n8822), .B2(n7447), .ZN(n7448)
         );
  AOI211_X1 U9114 ( .C1(n4473), .C2(n9135), .A(n9695), .B(n7448), .ZN(n7449)
         );
  OAI211_X1 U9115 ( .C1(n9792), .C2(n8758), .A(n7450), .B(n7449), .ZN(P1_U3229) );
  INV_X1 U9116 ( .A(n7451), .ZN(n7463) );
  OAI222_X1 U9117 ( .A1(n9513), .A2(n7463), .B1(n9082), .B2(P1_U3084), .C1(
        n7452), .C2(n9522), .ZN(P1_U3332) );
  INV_X1 U9118 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7460) );
  AND2_X1 U9119 ( .A1(n7453), .A2(n9577), .ZN(n7454) );
  OR2_X1 U9120 ( .A1(n9587), .A2(n7456), .ZN(n8949) );
  NAND2_X1 U9121 ( .A1(n9587), .A2(n7456), .ZN(n8959) );
  NAND2_X1 U9122 ( .A1(n8949), .A2(n8959), .ZN(n9572) );
  XNOR2_X1 U9123 ( .A(n7574), .B(n9576), .ZN(n9051) );
  XNOR2_X1 U9124 ( .A(n7567), .B(n9051), .ZN(n7511) );
  NAND2_X1 U9125 ( .A1(n8949), .A2(n9570), .ZN(n8963) );
  NAND2_X1 U9126 ( .A1(n8959), .A2(n8955), .ZN(n8952) );
  NAND2_X1 U9127 ( .A1(n8952), .A2(n8949), .ZN(n8877) );
  XNOR2_X1 U9128 ( .A(n7575), .B(n9051), .ZN(n7457) );
  AOI222_X1 U9129 ( .A1(n9574), .A2(n7457), .B1(n9133), .B2(n9400), .C1(n9134), 
        .C2(n9329), .ZN(n7506) );
  AOI21_X1 U9130 ( .B1(n7574), .B2(n9588), .A(n7568), .ZN(n7509) );
  AOI22_X1 U9131 ( .A1(n7509), .A2(n9764), .B1(n9487), .B2(n7574), .ZN(n7458)
         );
  OAI211_X1 U9132 ( .C1(n7511), .C2(n9484), .A(n7506), .B(n7458), .ZN(n7461)
         );
  NAND2_X1 U9133 ( .A1(n7461), .A2(n9800), .ZN(n7459) );
  OAI21_X1 U9134 ( .B1(n9800), .B2(n7460), .A(n7459), .ZN(P1_U3487) );
  NAND2_X1 U9135 ( .A1(n7461), .A2(n9809), .ZN(n7462) );
  OAI21_X1 U9136 ( .B1(n9809), .B2(n6022), .A(n7462), .ZN(P1_U3534) );
  OAI222_X1 U9137 ( .A1(n8694), .A2(n7464), .B1(n8696), .B2(n7463), .C1(n7937), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NAND2_X1 U9138 ( .A1(n7465), .A2(n7470), .ZN(n7466) );
  NAND2_X1 U9139 ( .A1(n7467), .A2(n7466), .ZN(n7607) );
  NAND2_X1 U9140 ( .A1(n7469), .A2(n7468), .ZN(n7471) );
  XNOR2_X1 U9141 ( .A(n7471), .B(n6443), .ZN(n7475) );
  OR2_X1 U9142 ( .A1(n7535), .A2(n9814), .ZN(n7474) );
  OR2_X1 U9143 ( .A1(n7472), .A2(n9812), .ZN(n7473) );
  NAND2_X1 U9144 ( .A1(n7474), .A2(n7473), .ZN(n7616) );
  AOI21_X1 U9145 ( .B1(n7475), .B2(n9838), .A(n7616), .ZN(n7606) );
  OR2_X1 U9146 ( .A1(n7606), .A2(n9855), .ZN(n7483) );
  OAI22_X1 U9147 ( .A1(n8553), .A2(n7476), .B1(n7620), .B2(n9845), .ZN(n7480)
         );
  AOI21_X1 U9148 ( .B1(n7477), .B2(n7481), .A(n9942), .ZN(n7478) );
  NAND2_X1 U9149 ( .A1(n7478), .A2(n7518), .ZN(n7605) );
  NOR2_X1 U9150 ( .A1(n7605), .A2(n9847), .ZN(n7479) );
  AOI211_X1 U9151 ( .C1(n8534), .C2(n7481), .A(n7480), .B(n7479), .ZN(n7482)
         );
  OAI211_X1 U9152 ( .C1(n7607), .C2(n8506), .A(n7483), .B(n7482), .ZN(P2_U3286) );
  XNOR2_X1 U9153 ( .A(n7485), .B(n7484), .ZN(n7486) );
  XNOR2_X1 U9154 ( .A(n7487), .B(n7486), .ZN(n7492) );
  INV_X1 U9155 ( .A(n9576), .ZN(n7573) );
  OAI22_X1 U9156 ( .A1(n8824), .A2(n7573), .B1(n8822), .B2(n9582), .ZN(n7488)
         );
  AOI211_X1 U9157 ( .C1(n4473), .C2(n9577), .A(n7489), .B(n7488), .ZN(n7491)
         );
  NAND2_X1 U9158 ( .A1(n8828), .A2(n9587), .ZN(n7490) );
  OAI211_X1 U9159 ( .C1(n7492), .C2(n8831), .A(n7491), .B(n7490), .ZN(P1_U3215) );
  XOR2_X1 U9160 ( .A(n7494), .B(n7493), .Z(n7502) );
  AOI21_X1 U9161 ( .B1(n9817), .B2(n7496), .A(n7495), .ZN(n7499) );
  OR2_X1 U9162 ( .A1(n9824), .A2(n7497), .ZN(n7498) );
  OAI211_X1 U9163 ( .C1(n7500), .C2(n9819), .A(n7499), .B(n7498), .ZN(n7501)
         );
  AOI21_X1 U9164 ( .B1(n7502), .B2(n9821), .A(n7501), .ZN(n7503) );
  INV_X1 U9165 ( .A(n7503), .ZN(P2_U3223) );
  INV_X1 U9166 ( .A(n7562), .ZN(n7504) );
  AOI22_X1 U9167 ( .A1(n9753), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7504), .B2(
        n9583), .ZN(n7505) );
  OAI21_X1 U9168 ( .B1(n4589), .B2(n9396), .A(n7505), .ZN(n7508) );
  NOR2_X1 U9169 ( .A1(n7506), .A2(n9753), .ZN(n7507) );
  AOI211_X1 U9170 ( .C1(n7509), .C2(n9406), .A(n7508), .B(n7507), .ZN(n7510)
         );
  OAI21_X1 U9171 ( .B1(n9408), .B2(n7511), .A(n7510), .ZN(P1_U3280) );
  XNOR2_X1 U9172 ( .A(n7512), .B(n4985), .ZN(n9947) );
  INV_X1 U9173 ( .A(n9947), .ZN(n7528) );
  NAND2_X1 U9174 ( .A1(n7513), .A2(n7971), .ZN(n7515) );
  XNOR2_X1 U9175 ( .A(n7515), .B(n7514), .ZN(n7517) );
  OAI21_X1 U9176 ( .B1(n7517), .B2(n8527), .A(n7516), .ZN(n9944) );
  INV_X1 U9177 ( .A(n7518), .ZN(n7520) );
  INV_X1 U9178 ( .A(n7519), .ZN(n7541) );
  OAI21_X1 U9179 ( .B1(n9941), .B2(n7520), .A(n7541), .ZN(n9943) );
  OAI22_X1 U9180 ( .A1(n8553), .A2(n6991), .B1(n7521), .B2(n9845), .ZN(n7522)
         );
  AOI21_X1 U9181 ( .B1(n8534), .B2(n7523), .A(n7522), .ZN(n7524) );
  OAI21_X1 U9182 ( .B1(n9943), .B2(n7525), .A(n7524), .ZN(n7526) );
  AOI21_X1 U9183 ( .B1(n9944), .B2(n8553), .A(n7526), .ZN(n7527) );
  OAI21_X1 U9184 ( .B1(n7528), .B2(n8506), .A(n7527), .ZN(P2_U3285) );
  INV_X1 U9185 ( .A(n7529), .ZN(n7532) );
  OAI222_X1 U9186 ( .A1(n8694), .A2(n7531), .B1(n8696), .B2(n7532), .C1(
        P2_U3152), .C2(n7530), .ZN(P2_U3336) );
  OAI222_X1 U9187 ( .A1(n9522), .A2(n10122), .B1(n9513), .B2(n7532), .C1(
        P1_U3084), .C2(n9042), .ZN(P1_U3331) );
  NAND2_X1 U9188 ( .A1(n7533), .A2(n7972), .ZN(n7534) );
  XNOR2_X1 U9189 ( .A(n7534), .B(n7913), .ZN(n7539) );
  OR2_X1 U9190 ( .A1(n7753), .A2(n9814), .ZN(n7537) );
  OR2_X1 U9191 ( .A1(n7535), .A2(n9812), .ZN(n7536) );
  NAND2_X1 U9192 ( .A1(n7537), .A2(n7536), .ZN(n7772) );
  INV_X1 U9193 ( .A(n7772), .ZN(n7538) );
  OAI21_X1 U9194 ( .B1(n7539), .B2(n8527), .A(n7538), .ZN(n7662) );
  INV_X1 U9195 ( .A(n7662), .ZN(n7547) );
  XNOR2_X1 U9196 ( .A(n7540), .B(n7913), .ZN(n7664) );
  NAND2_X1 U9197 ( .A1(n7664), .A2(n9853), .ZN(n7546) );
  AOI211_X1 U9198 ( .C1(n7771), .C2(n7541), .A(n9942), .B(n7717), .ZN(n7663)
         );
  NOR2_X1 U9199 ( .A1(n9851), .A2(n7669), .ZN(n7544) );
  OAI22_X1 U9200 ( .A1(n8553), .A2(n7542), .B1(n7775), .B2(n9845), .ZN(n7543)
         );
  AOI211_X1 U9201 ( .C1(n7663), .C2(n8556), .A(n7544), .B(n7543), .ZN(n7545)
         );
  OAI211_X1 U9202 ( .C1(n9849), .C2(n7547), .A(n7546), .B(n7545), .ZN(P2_U3284) );
  OAI21_X1 U9203 ( .B1(n7550), .B2(n7549), .A(n7548), .ZN(n7557) );
  NOR2_X1 U9204 ( .A1(n9819), .A2(n9933), .ZN(n7556) );
  NAND2_X1 U9205 ( .A1(n9817), .A2(n7551), .ZN(n7553) );
  OAI211_X1 U9206 ( .C1(n9824), .C2(n7554), .A(n7553), .B(n7552), .ZN(n7555)
         );
  AOI211_X1 U9207 ( .C1(n7557), .C2(n9821), .A(n7556), .B(n7555), .ZN(n7558)
         );
  INV_X1 U9208 ( .A(n7558), .ZN(P2_U3233) );
  XNOR2_X1 U9209 ( .A(n7560), .B(n7559), .ZN(n7566) );
  INV_X1 U9210 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7561) );
  NOR2_X1 U9211 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7561), .ZN(n9703) );
  INV_X1 U9212 ( .A(n9133), .ZN(n7732) );
  OAI22_X1 U9213 ( .A1(n8824), .A2(n7732), .B1(n8822), .B2(n7562), .ZN(n7563)
         );
  AOI211_X1 U9214 ( .C1(n4473), .C2(n9134), .A(n9703), .B(n7563), .ZN(n7565)
         );
  NAND2_X1 U9215 ( .A1(n7574), .A2(n8828), .ZN(n7564) );
  OAI211_X1 U9216 ( .C1(n7566), .C2(n8831), .A(n7565), .B(n7564), .ZN(P1_U3234) );
  NAND2_X1 U9217 ( .A1(n7745), .A2(n7732), .ZN(n8967) );
  NAND2_X1 U9218 ( .A1(n8968), .A2(n8967), .ZN(n9069) );
  XNOR2_X1 U9219 ( .A(n7624), .B(n9069), .ZN(n7583) );
  INV_X1 U9220 ( .A(n7568), .ZN(n7569) );
  INV_X1 U9221 ( .A(n7745), .ZN(n7572) );
  AOI211_X1 U9222 ( .C1(n7745), .C2(n7569), .A(n9793), .B(n7653), .ZN(n7580)
         );
  INV_X1 U9223 ( .A(n7741), .ZN(n7570) );
  AOI22_X1 U9224 ( .A1(n9753), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7570), .B2(
        n9583), .ZN(n7571) );
  OAI21_X1 U9225 ( .B1(n7572), .B2(n9396), .A(n7571), .ZN(n7578) );
  AND2_X1 U9226 ( .A1(n7574), .A2(n7573), .ZN(n8876) );
  OR2_X1 U9227 ( .A1(n7574), .A2(n7573), .ZN(n8894) );
  OAI21_X1 U9228 ( .B1(n7575), .B2(n8876), .A(n8894), .ZN(n7630) );
  XNOR2_X1 U9229 ( .A(n7630), .B(n9069), .ZN(n7576) );
  AOI222_X1 U9230 ( .A1(n9574), .A2(n7576), .B1(n9132), .B2(n9400), .C1(n9576), 
        .C2(n9329), .ZN(n7582) );
  NOR2_X1 U9231 ( .A1(n7582), .A2(n9753), .ZN(n7577) );
  AOI211_X1 U9232 ( .C1(n7580), .C2(n9591), .A(n7578), .B(n7577), .ZN(n7579)
         );
  OAI21_X1 U9233 ( .B1(n9408), .B2(n7583), .A(n7579), .ZN(P1_U3279) );
  AOI21_X1 U9234 ( .B1(n9487), .B2(n7745), .A(n7580), .ZN(n7581) );
  OAI211_X1 U9235 ( .C1(n7583), .C2(n9484), .A(n7582), .B(n7581), .ZN(n7585)
         );
  NAND2_X1 U9236 ( .A1(n7585), .A2(n9800), .ZN(n7584) );
  OAI21_X1 U9237 ( .B1(n9800), .B2(n6047), .A(n7584), .ZN(P1_U3490) );
  NAND2_X1 U9238 ( .A1(n7585), .A2(n9809), .ZN(n7586) );
  OAI21_X1 U9239 ( .B1(n9809), .B2(n6566), .A(n7586), .ZN(P1_U3535) );
  INV_X1 U9240 ( .A(n7602), .ZN(n7589) );
  OR2_X1 U9241 ( .A1(n7587), .A2(P1_U3084), .ZN(n9129) );
  NAND2_X1 U9242 ( .A1(n9511), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7588) );
  OAI211_X1 U9243 ( .C1(n7589), .C2(n9513), .A(n9129), .B(n7588), .ZN(P1_U3330) );
  INV_X1 U9244 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7870) );
  AOI211_X1 U9245 ( .C1(n7591), .C2(n7870), .A(n8278), .B(n9554), .ZN(n7601)
         );
  NOR2_X1 U9246 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7592), .ZN(n7594) );
  NOR2_X1 U9247 ( .A1(n7594), .A2(n7593), .ZN(n8282) );
  XNOR2_X1 U9248 ( .A(n8282), .B(n8283), .ZN(n7595) );
  NOR2_X1 U9249 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7595), .ZN(n8284) );
  AOI21_X1 U9250 ( .B1(n7595), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8284), .ZN(
        n7596) );
  NOR2_X1 U9251 ( .A1(n7596), .A2(n9830), .ZN(n7600) );
  AND2_X1 U9252 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7597) );
  AOI21_X1 U9253 ( .B1(n9832), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7597), .ZN(
        n7598) );
  OAI21_X1 U9254 ( .B1(n9828), .B2(n8277), .A(n7598), .ZN(n7599) );
  OR3_X1 U9255 ( .A1(n7601), .A2(n7600), .A3(n7599), .ZN(P2_U3260) );
  NAND2_X1 U9256 ( .A1(n7602), .A2(n8690), .ZN(n7603) );
  OAI211_X1 U9257 ( .C1(n7604), .C2(n8694), .A(n7603), .B(n8082), .ZN(P2_U3335) );
  OAI211_X1 U9258 ( .C1(n7607), .C2(n9898), .A(n7606), .B(n7605), .ZN(n7610)
         );
  MUX2_X1 U9259 ( .A(n7610), .B(P2_REG1_REG_10__SCAN_IN), .S(n9958), .Z(n7608)
         );
  INV_X1 U9260 ( .A(n7608), .ZN(n7609) );
  OAI21_X1 U9261 ( .B1(n7617), .B2(n8634), .A(n7609), .ZN(P2_U3530) );
  MUX2_X1 U9262 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n7610), .S(n9949), .Z(n7611)
         );
  INV_X1 U9263 ( .A(n7611), .ZN(n7612) );
  OAI21_X1 U9264 ( .B1(n7617), .B2(n8677), .A(n7612), .ZN(P2_U3481) );
  XOR2_X1 U9265 ( .A(n7614), .B(n7613), .Z(n7622) );
  AOI21_X1 U9266 ( .B1(n9817), .B2(n7616), .A(n7615), .ZN(n7619) );
  OR2_X1 U9267 ( .A1(n9819), .A2(n7617), .ZN(n7618) );
  OAI211_X1 U9268 ( .C1(n9824), .C2(n7620), .A(n7619), .B(n7618), .ZN(n7621)
         );
  AOI21_X1 U9269 ( .B1(n7622), .B2(n9821), .A(n7621), .ZN(n7623) );
  INV_X1 U9270 ( .A(n7623), .ZN(P2_U3219) );
  NAND2_X1 U9271 ( .A1(n7624), .A2(n9069), .ZN(n7626) );
  NAND2_X1 U9272 ( .A1(n7745), .A2(n9133), .ZN(n7625) );
  AND2_X1 U9273 ( .A1(n9486), .A2(n9132), .ZN(n7627) );
  OR2_X1 U9274 ( .A1(n9486), .A2(n9132), .ZN(n7628) );
  INV_X1 U9275 ( .A(n9131), .ZN(n8874) );
  XNOR2_X1 U9276 ( .A(n8875), .B(n8874), .ZN(n7784) );
  XNOR2_X1 U9277 ( .A(n7780), .B(n7784), .ZN(n9617) );
  INV_X1 U9278 ( .A(n9617), .ZN(n7640) );
  INV_X1 U9279 ( .A(n8968), .ZN(n7629) );
  INV_X1 U9280 ( .A(n9132), .ZN(n7742) );
  OR2_X1 U9281 ( .A1(n9486), .A2(n7742), .ZN(n8948) );
  NAND2_X1 U9282 ( .A1(n9486), .A2(n7742), .ZN(n8973) );
  INV_X1 U9283 ( .A(n7784), .ZN(n9070) );
  XNOR2_X1 U9284 ( .A(n7785), .B(n9070), .ZN(n7631) );
  NAND2_X1 U9285 ( .A1(n7631), .A2(n9574), .ZN(n7633) );
  AOI22_X1 U9286 ( .A1(n9130), .A2(n9400), .B1(n9132), .B2(n9578), .ZN(n7632)
         );
  NAND2_X1 U9287 ( .A1(n7633), .A2(n7632), .ZN(n9616) );
  INV_X1 U9288 ( .A(n9486), .ZN(n7656) );
  INV_X1 U9289 ( .A(n7655), .ZN(n7634) );
  OAI211_X1 U9290 ( .C1(n7634), .C2(n9614), .A(n9764), .B(n4546), .ZN(n9613)
         );
  INV_X1 U9291 ( .A(n7635), .ZN(n8704) );
  OAI22_X1 U9292 ( .A1(n9751), .A2(n6091), .B1(n8704), .B2(n9743), .ZN(n7636)
         );
  AOI21_X1 U9293 ( .B1(n8875), .B2(n9585), .A(n7636), .ZN(n7637) );
  OAI21_X1 U9294 ( .B1(n9613), .B2(n7793), .A(n7637), .ZN(n7638) );
  AOI21_X1 U9295 ( .B1(n9616), .B2(n9751), .A(n7638), .ZN(n7639) );
  OAI21_X1 U9296 ( .B1(n7640), .B2(n9408), .A(n7639), .ZN(P1_U3277) );
  INV_X1 U9297 ( .A(n7641), .ZN(n7693) );
  INV_X1 U9298 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10109) );
  OAI222_X1 U9299 ( .A1(n9513), .A2(n7693), .B1(P1_U3084), .B2(n7642), .C1(
        n10109), .C2(n9522), .ZN(P1_U3329) );
  XNOR2_X1 U9300 ( .A(n7643), .B(n9072), .ZN(n7644) );
  INV_X1 U9301 ( .A(n7644), .ZN(n9491) );
  NAND2_X1 U9302 ( .A1(n7644), .A2(n9581), .ZN(n7652) );
  OAI21_X1 U9303 ( .B1(n9072), .B2(n7646), .A(n7645), .ZN(n7650) );
  NAND2_X1 U9304 ( .A1(n9131), .A2(n9400), .ZN(n7648) );
  NAND2_X1 U9305 ( .A1(n9133), .A2(n9578), .ZN(n7647) );
  NAND2_X1 U9306 ( .A1(n7648), .A2(n7647), .ZN(n7649) );
  AOI21_X1 U9307 ( .B1(n7650), .B2(n9574), .A(n7649), .ZN(n7651) );
  NAND2_X1 U9308 ( .A1(n7652), .A2(n7651), .ZN(n9493) );
  NAND2_X1 U9309 ( .A1(n9493), .A2(n9751), .ZN(n7660) );
  OR2_X1 U9310 ( .A1(n7653), .A2(n7656), .ZN(n7654) );
  AND2_X1 U9311 ( .A1(n7655), .A2(n7654), .ZN(n9488) );
  NOR2_X1 U9312 ( .A1(n7656), .A2(n9396), .ZN(n7658) );
  OAI22_X1 U9313 ( .A1(n9751), .A2(n6542), .B1(n7728), .B2(n9743), .ZN(n7657)
         );
  AOI211_X1 U9314 ( .C1(n9488), .C2(n9406), .A(n7658), .B(n7657), .ZN(n7659)
         );
  OAI211_X1 U9315 ( .C1(n9491), .C2(n7661), .A(n7660), .B(n7659), .ZN(P1_U3278) );
  INV_X1 U9316 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7665) );
  AOI211_X1 U9317 ( .C1(n7664), .C2(n9946), .A(n7663), .B(n7662), .ZN(n7667)
         );
  MUX2_X1 U9318 ( .A(n7665), .B(n7667), .S(n9949), .Z(n7666) );
  OAI21_X1 U9319 ( .B1(n7669), .B2(n8677), .A(n7666), .ZN(P2_U3487) );
  MUX2_X1 U9320 ( .A(n7108), .B(n7667), .S(n9960), .Z(n7668) );
  OAI21_X1 U9321 ( .B1(n7669), .B2(n8634), .A(n7668), .ZN(P2_U3532) );
  AND2_X1 U9322 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8755) );
  INV_X1 U9323 ( .A(n8755), .ZN(n7670) );
  OAI21_X1 U9324 ( .B1(n9724), .B2(n7671), .A(n7670), .ZN(n7681) );
  NOR2_X1 U9325 ( .A1(n7682), .A2(n7672), .ZN(n7674) );
  NOR2_X1 U9326 ( .A1(n7674), .A2(n7673), .ZN(n7700) );
  INV_X1 U9327 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7675) );
  OR2_X1 U9328 ( .A1(n7702), .A2(n7675), .ZN(n7677) );
  NAND2_X1 U9329 ( .A1(n7702), .A2(n7675), .ZN(n7676) );
  AND2_X1 U9330 ( .A1(n7677), .A2(n7676), .ZN(n7701) );
  NOR2_X1 U9331 ( .A1(n7700), .A2(n7701), .ZN(n7699) );
  AOI21_X1 U9332 ( .B1(n7702), .B2(P1_REG1_REG_16__SCAN_IN), .A(n7699), .ZN(
        n7679) );
  XNOR2_X1 U9333 ( .A(n9145), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7678) );
  NOR2_X1 U9334 ( .A1(n7679), .A2(n7678), .ZN(n9142) );
  AOI211_X1 U9335 ( .C1(n7679), .C2(n7678), .A(n9673), .B(n9142), .ZN(n7680)
         );
  AOI211_X1 U9336 ( .C1(n9730), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n7681), .B(
        n7680), .ZN(n7691) );
  NOR2_X1 U9337 ( .A1(n7683), .A2(n7682), .ZN(n7685) );
  NOR2_X1 U9338 ( .A1(n7685), .A2(n7684), .ZN(n7698) );
  XNOR2_X1 U9339 ( .A(n7702), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U9340 ( .A1(n7702), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7686) );
  NAND2_X1 U9341 ( .A1(n7695), .A2(n7686), .ZN(n7689) );
  INV_X1 U9342 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7687) );
  XNOR2_X1 U9343 ( .A(n9145), .B(n7687), .ZN(n7688) );
  NAND2_X1 U9344 ( .A1(n7689), .A2(n7688), .ZN(n9147) );
  OAI211_X1 U9345 ( .C1(n7689), .C2(n7688), .A(n9147), .B(n9718), .ZN(n7690)
         );
  NAND2_X1 U9346 ( .A1(n7691), .A2(n7690), .ZN(P1_U3258) );
  OAI222_X1 U9347 ( .A1(n7694), .A2(P2_U3152), .B1(n8696), .B2(n7693), .C1(
        n7692), .C2(n8694), .ZN(P2_U3334) );
  INV_X1 U9348 ( .A(n7695), .ZN(n7696) );
  AOI211_X1 U9349 ( .C1(n7698), .C2(n7697), .A(n9690), .B(n7696), .ZN(n7707)
         );
  AOI211_X1 U9350 ( .C1(n7701), .C2(n7700), .A(n9673), .B(n7699), .ZN(n7706)
         );
  INV_X1 U9351 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7704) );
  AND2_X1 U9352 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8747) );
  AOI21_X1 U9353 ( .B1(n9705), .B2(n7702), .A(n8747), .ZN(n7703) );
  OAI21_X1 U9354 ( .B1(n9717), .B2(n7704), .A(n7703), .ZN(n7705) );
  OR3_X1 U9355 ( .A1(n7707), .A2(n7706), .A3(n7705), .ZN(P1_U3257) );
  XNOR2_X1 U9356 ( .A(n7708), .B(n7977), .ZN(n7712) );
  OR2_X1 U9357 ( .A1(n7823), .A2(n9814), .ZN(n7711) );
  OR2_X1 U9358 ( .A1(n7709), .A2(n9812), .ZN(n7710) );
  NAND2_X1 U9359 ( .A1(n7711), .A2(n7710), .ZN(n7842) );
  AOI21_X1 U9360 ( .B1(n7712), .B2(n9838), .A(n7842), .ZN(n7798) );
  INV_X1 U9361 ( .A(n7713), .ZN(n7714) );
  AOI21_X1 U9362 ( .B1(n7977), .B2(n7715), .A(n7714), .ZN(n7800) );
  NAND2_X1 U9363 ( .A1(n7800), .A2(n9853), .ZN(n7722) );
  OAI22_X1 U9364 ( .A1(n8553), .A2(n7716), .B1(n7839), .B2(n9845), .ZN(n7719)
         );
  OAI211_X1 U9365 ( .C1(n7717), .C2(n7979), .A(n9841), .B(n7760), .ZN(n7797)
         );
  NOR2_X1 U9366 ( .A1(n7797), .A2(n9847), .ZN(n7718) );
  AOI211_X1 U9367 ( .C1(n8534), .C2(n7720), .A(n7719), .B(n7718), .ZN(n7721)
         );
  OAI211_X1 U9368 ( .C1(n9855), .C2(n7798), .A(n7722), .B(n7721), .ZN(P2_U3283) );
  INV_X1 U9369 ( .A(n7723), .ZN(n7725) );
  NAND2_X1 U9370 ( .A1(n7725), .A2(n7724), .ZN(n7726) );
  XNOR2_X1 U9371 ( .A(n7727), .B(n7726), .ZN(n7735) );
  INV_X1 U9372 ( .A(n4473), .ZN(n8800) );
  INV_X1 U9373 ( .A(n7728), .ZN(n7729) );
  AOI22_X1 U9374 ( .A1(n8811), .A2(n9131), .B1(n7729), .B2(n8810), .ZN(n7731)
         );
  OAI211_X1 U9375 ( .C1(n8800), .C2(n7732), .A(n7731), .B(n7730), .ZN(n7733)
         );
  AOI21_X1 U9376 ( .B1(n9486), .B2(n8828), .A(n7733), .ZN(n7734) );
  OAI21_X1 U9377 ( .B1(n7735), .B2(n8831), .A(n7734), .ZN(P1_U3232) );
  INV_X1 U9378 ( .A(n7737), .ZN(n7738) );
  AOI21_X1 U9379 ( .B1(n7739), .B2(n7736), .A(n7738), .ZN(n7748) );
  INV_X1 U9380 ( .A(n7740), .ZN(n7744) );
  OAI22_X1 U9381 ( .A1(n8824), .A2(n7742), .B1(n8822), .B2(n7741), .ZN(n7743)
         );
  AOI211_X1 U9382 ( .C1(n4473), .C2(n9576), .A(n7744), .B(n7743), .ZN(n7747)
         );
  NAND2_X1 U9383 ( .A1(n7745), .A2(n8828), .ZN(n7746) );
  OAI211_X1 U9384 ( .C1(n7748), .C2(n8831), .A(n7747), .B(n7746), .ZN(P1_U3222) );
  NAND2_X1 U9385 ( .A1(n7750), .A2(n7751), .ZN(n7752) );
  NAND3_X1 U9386 ( .A1(n7749), .A2(n9838), .A3(n7752), .ZN(n7757) );
  OR2_X1 U9387 ( .A1(n8170), .A2(n9814), .ZN(n7755) );
  OR2_X1 U9388 ( .A1(n7753), .A2(n9812), .ZN(n7754) );
  NAND2_X1 U9389 ( .A1(n7755), .A2(n7754), .ZN(n8116) );
  INV_X1 U9390 ( .A(n8116), .ZN(n7756) );
  NAND2_X1 U9391 ( .A1(n7757), .A2(n7756), .ZN(n7805) );
  INV_X1 U9392 ( .A(n7805), .ZN(n7766) );
  XNOR2_X1 U9393 ( .A(n7758), .B(n7989), .ZN(n7807) );
  NAND2_X1 U9394 ( .A1(n7807), .A2(n9853), .ZN(n7765) );
  INV_X1 U9395 ( .A(n7829), .ZN(n7759) );
  AOI211_X1 U9396 ( .C1(n8120), .C2(n7760), .A(n9942), .B(n7759), .ZN(n7806)
         );
  INV_X1 U9397 ( .A(n8120), .ZN(n7812) );
  NOR2_X1 U9398 ( .A1(n7812), .A2(n9851), .ZN(n7763) );
  OAI22_X1 U9399 ( .A1(n8553), .A2(n7761), .B1(n8118), .B2(n9845), .ZN(n7762)
         );
  AOI211_X1 U9400 ( .C1(n7806), .C2(n8556), .A(n7763), .B(n7762), .ZN(n7764)
         );
  OAI211_X1 U9401 ( .C1(n9849), .C2(n7766), .A(n7765), .B(n7764), .ZN(P2_U3282) );
  NAND2_X1 U9402 ( .A1(n7768), .A2(n7767), .ZN(n7769) );
  XNOR2_X1 U9403 ( .A(n7770), .B(n7769), .ZN(n7777) );
  NAND2_X1 U9404 ( .A1(n8244), .A2(n7771), .ZN(n7774) );
  AOI22_X1 U9405 ( .A1(n9817), .A2(n7772), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n7773) );
  OAI211_X1 U9406 ( .C1(n9824), .C2(n7775), .A(n7774), .B(n7773), .ZN(n7776)
         );
  AOI21_X1 U9407 ( .B1(n7777), .B2(n9821), .A(n7776), .ZN(n7778) );
  INV_X1 U9408 ( .A(n7778), .ZN(P2_U3226) );
  NOR2_X1 U9409 ( .A1(n8875), .A2(n9131), .ZN(n7779) );
  OR2_X1 U9410 ( .A1(n9606), .A2(n9130), .ZN(n7781) );
  NAND2_X1 U9411 ( .A1(n7849), .A2(n7781), .ZN(n7783) );
  NAND2_X1 U9412 ( .A1(n9606), .A2(n9130), .ZN(n7782) );
  NAND2_X1 U9413 ( .A1(n7783), .A2(n7782), .ZN(n9172) );
  INV_X1 U9414 ( .A(n9402), .ZN(n8823) );
  OR2_X1 U9415 ( .A1(n9173), .A2(n8823), .ZN(n8931) );
  NAND2_X1 U9416 ( .A1(n9173), .A2(n8823), .ZN(n9193) );
  NAND2_X1 U9417 ( .A1(n8931), .A2(n9193), .ZN(n9171) );
  XNOR2_X1 U9418 ( .A(n9172), .B(n8989), .ZN(n9605) );
  INV_X1 U9419 ( .A(n9605), .ZN(n7796) );
  OR2_X1 U9420 ( .A1(n8875), .A2(n8874), .ZN(n8980) );
  INV_X1 U9421 ( .A(n9130), .ZN(n8705) );
  OR2_X1 U9422 ( .A1(n9606), .A2(n8705), .ZN(n8987) );
  NAND2_X1 U9423 ( .A1(n9606), .A2(n8705), .ZN(n8986) );
  NAND2_X1 U9424 ( .A1(n8987), .A2(n8986), .ZN(n7848) );
  NAND3_X1 U9425 ( .A1(n7845), .A2(n8986), .A3(n9171), .ZN(n7786) );
  NAND2_X1 U9426 ( .A1(n9194), .A2(n7786), .ZN(n7787) );
  NAND2_X1 U9427 ( .A1(n7787), .A2(n9574), .ZN(n7789) );
  AOI22_X1 U9428 ( .A1(n9376), .A2(n9400), .B1(n9329), .B2(n9130), .ZN(n7788)
         );
  NAND2_X1 U9429 ( .A1(n7789), .A2(n7788), .ZN(n9604) );
  INV_X1 U9430 ( .A(n9173), .ZN(n9602) );
  OAI211_X1 U9431 ( .C1(n9602), .C2(n7854), .A(n4545), .B(n9764), .ZN(n9601)
         );
  INV_X1 U9432 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7790) );
  OAI22_X1 U9433 ( .A1(n9751), .A2(n7790), .B1(n8745), .B2(n9743), .ZN(n7791)
         );
  AOI21_X1 U9434 ( .B1(n9173), .B2(n9585), .A(n7791), .ZN(n7792) );
  OAI21_X1 U9435 ( .B1(n9601), .B2(n7793), .A(n7792), .ZN(n7794) );
  AOI21_X1 U9436 ( .B1(n9604), .B2(n9751), .A(n7794), .ZN(n7795) );
  OAI21_X1 U9437 ( .B1(n7796), .B2(n9408), .A(n7795), .ZN(P1_U3275) );
  NAND2_X1 U9438 ( .A1(n7798), .A2(n7797), .ZN(n7799) );
  AOI21_X1 U9439 ( .B1(n7800), .B2(n9946), .A(n7799), .ZN(n7802) );
  MUX2_X1 U9440 ( .A(n5342), .B(n7802), .S(n9960), .Z(n7801) );
  OAI21_X1 U9441 ( .B1(n7979), .B2(n8634), .A(n7801), .ZN(P2_U3533) );
  INV_X1 U9442 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7803) );
  MUX2_X1 U9443 ( .A(n7803), .B(n7802), .S(n9949), .Z(n7804) );
  OAI21_X1 U9444 ( .B1(n7979), .B2(n8677), .A(n7804), .ZN(P2_U3490) );
  AOI211_X1 U9445 ( .C1(n7807), .C2(n9946), .A(n7806), .B(n7805), .ZN(n7809)
         );
  MUX2_X1 U9446 ( .A(n5367), .B(n7809), .S(n9960), .Z(n7808) );
  OAI21_X1 U9447 ( .B1(n7812), .B2(n8634), .A(n7808), .ZN(P2_U3534) );
  INV_X1 U9448 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7810) );
  MUX2_X1 U9449 ( .A(n7810), .B(n7809), .S(n9949), .Z(n7811) );
  OAI21_X1 U9450 ( .B1(n7812), .B2(n8677), .A(n7811), .ZN(P2_U3493) );
  INV_X1 U9451 ( .A(n7813), .ZN(n7815) );
  OAI222_X1 U9452 ( .A1(n9522), .A2(n10301), .B1(n9513), .B2(n7815), .C1(n6336), .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U9453 ( .A1(n8694), .A2(n7816), .B1(n8696), .B2(n7815), .C1(n7814), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  INV_X1 U9454 ( .A(n7817), .ZN(n7863) );
  OAI222_X1 U9455 ( .A1(n9513), .A2(n7863), .B1(P1_U3084), .B2(n7818), .C1(
        n10124), .C2(n9522), .ZN(P1_U3327) );
  OAI21_X1 U9456 ( .B1(n7820), .B2(n7903), .A(n7819), .ZN(n7867) );
  INV_X1 U9457 ( .A(n7867), .ZN(n7835) );
  XNOR2_X1 U9458 ( .A(n7821), .B(n7903), .ZN(n7822) );
  NAND2_X1 U9459 ( .A1(n7822), .A2(n9838), .ZN(n7828) );
  OR2_X1 U9460 ( .A1(n7823), .A2(n9812), .ZN(n7826) );
  OR2_X1 U9461 ( .A1(n7824), .A2(n9814), .ZN(n7825) );
  NAND2_X1 U9462 ( .A1(n7826), .A2(n7825), .ZN(n8240) );
  INV_X1 U9463 ( .A(n8240), .ZN(n7827) );
  NAND2_X1 U9464 ( .A1(n7828), .A2(n7827), .ZN(n7865) );
  AOI211_X1 U9465 ( .C1(n8245), .C2(n7829), .A(n9942), .B(n8548), .ZN(n7866)
         );
  NAND2_X1 U9466 ( .A1(n7866), .A2(n8556), .ZN(n7832) );
  INV_X1 U9467 ( .A(n8242), .ZN(n7830) );
  INV_X1 U9468 ( .A(n9845), .ZN(n8483) );
  AOI22_X1 U9469 ( .A1(n9849), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7830), .B2(
        n8483), .ZN(n7831) );
  OAI211_X1 U9470 ( .C1(n4703), .C2(n9851), .A(n7832), .B(n7831), .ZN(n7833)
         );
  AOI21_X1 U9471 ( .B1(n7865), .B2(n8553), .A(n7833), .ZN(n7834) );
  OAI21_X1 U9472 ( .B1(n7835), .B2(n8506), .A(n7834), .ZN(P2_U3281) );
  OAI211_X1 U9473 ( .C1(n7838), .C2(n7837), .A(n7836), .B(n9821), .ZN(n7844)
         );
  NOR2_X1 U9474 ( .A1(n9824), .A2(n7839), .ZN(n7840) );
  AOI211_X1 U9475 ( .C1(n9817), .C2(n7842), .A(n7841), .B(n7840), .ZN(n7843)
         );
  OAI211_X1 U9476 ( .C1(n7979), .C2(n9819), .A(n7844), .B(n7843), .ZN(P2_U3236) );
  INV_X1 U9477 ( .A(n7845), .ZN(n7846) );
  AOI21_X1 U9478 ( .B1(n7848), .B2(n7847), .A(n7846), .ZN(n7852) );
  INV_X1 U9479 ( .A(n7848), .ZN(n9073) );
  XNOR2_X1 U9480 ( .A(n7849), .B(n9073), .ZN(n9611) );
  NAND2_X1 U9481 ( .A1(n9611), .A2(n9581), .ZN(n7851) );
  AOI22_X1 U9482 ( .A1(n9402), .A2(n9400), .B1(n9329), .B2(n9131), .ZN(n7850)
         );
  OAI211_X1 U9483 ( .C1(n7853), .C2(n7852), .A(n7851), .B(n7850), .ZN(n9609)
         );
  INV_X1 U9484 ( .A(n9609), .ZN(n7861) );
  AND2_X1 U9485 ( .A1(n4546), .A2(n9606), .ZN(n7855) );
  OR2_X1 U9486 ( .A1(n7855), .A2(n7854), .ZN(n9608) );
  AOI22_X1 U9487 ( .A1(n9753), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7856), .B2(
        n9583), .ZN(n7858) );
  NAND2_X1 U9488 ( .A1(n9606), .A2(n9585), .ZN(n7857) );
  OAI211_X1 U9489 ( .C1(n9608), .C2(n9225), .A(n7858), .B(n7857), .ZN(n7859)
         );
  AOI21_X1 U9490 ( .B1(n9611), .B2(n9592), .A(n7859), .ZN(n7860) );
  OAI21_X1 U9491 ( .B1(n7861), .B2(n9753), .A(n7860), .ZN(P1_U3276) );
  OAI222_X1 U9492 ( .A1(n7864), .A2(P2_U3152), .B1(n8696), .B2(n7863), .C1(
        n7862), .C2(n8694), .ZN(P2_U3332) );
  AOI211_X1 U9493 ( .C1(n7867), .C2(n9946), .A(n7866), .B(n7865), .ZN(n7869)
         );
  MUX2_X1 U9494 ( .A(n5414), .B(n7869), .S(n9949), .Z(n7868) );
  OAI21_X1 U9495 ( .B1(n4703), .B2(n8677), .A(n7868), .ZN(P2_U3496) );
  MUX2_X1 U9496 ( .A(n7870), .B(n7869), .S(n9960), .Z(n7871) );
  OAI21_X1 U9497 ( .B1(n4703), .B2(n8634), .A(n7871), .ZN(P2_U3535) );
  INV_X1 U9498 ( .A(n7874), .ZN(n7875) );
  NAND2_X1 U9499 ( .A1(n7875), .A2(n10172), .ZN(n7876) );
  INV_X1 U9500 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8685) );
  INV_X1 U9501 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10146) );
  MUX2_X1 U9502 ( .A(n8685), .B(n10146), .S(n6469), .Z(n7884) );
  INV_X1 U9503 ( .A(n8841), .ZN(n8686) );
  OAI222_X1 U9504 ( .A1(n9513), .A2(n8686), .B1(n5785), .B2(P1_U3084), .C1(
        n10146), .C2(n9522), .ZN(P1_U3323) );
  INV_X1 U9505 ( .A(n8052), .ZN(n7878) );
  INV_X1 U9506 ( .A(n7896), .ZN(n7897) );
  NAND2_X1 U9507 ( .A1(n8841), .A2(n7890), .ZN(n7881) );
  OR2_X1 U9508 ( .A1(n4476), .A2(n8685), .ZN(n7880) );
  INV_X1 U9509 ( .A(n8642), .ZN(n7895) );
  INV_X1 U9510 ( .A(n8249), .ZN(n7894) );
  INV_X1 U9511 ( .A(n7883), .ZN(n7886) );
  INV_X1 U9512 ( .A(n7884), .ZN(n7885) );
  NAND2_X1 U9513 ( .A1(n7886), .A2(n7885), .ZN(n7887) );
  MUX2_X1 U9514 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6469), .Z(n7888) );
  XNOR2_X1 U9515 ( .A(n7888), .B(SI_31_), .ZN(n7889) );
  NAND2_X1 U9516 ( .A1(n8833), .A2(n7890), .ZN(n7893) );
  INV_X1 U9517 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7891) );
  OR2_X1 U9518 ( .A1(n5199), .A2(n7891), .ZN(n7892) );
  INV_X1 U9519 ( .A(n8347), .ZN(n7898) );
  OR2_X1 U9520 ( .A1(n8560), .A2(n7898), .ZN(n8060) );
  NAND2_X1 U9521 ( .A1(n7895), .A2(n7894), .ZN(n8055) );
  NAND2_X1 U9522 ( .A1(n8060), .A2(n8055), .ZN(n8058) );
  XNOR2_X1 U9523 ( .A(n7899), .B(n8530), .ZN(n8077) );
  NAND2_X1 U9524 ( .A1(n7901), .A2(n7900), .ZN(n8076) );
  INV_X1 U9525 ( .A(n7902), .ZN(n8061) );
  NAND2_X1 U9526 ( .A1(n8061), .A2(n8056), .ZN(n8057) );
  INV_X1 U9527 ( .A(n8417), .ZN(n7918) );
  INV_X1 U9528 ( .A(n8469), .ZN(n8461) );
  NAND2_X1 U9529 ( .A1(n8007), .A2(n8012), .ZN(n8511) );
  INV_X1 U9530 ( .A(n7903), .ZN(n7994) );
  NOR4_X1 U9531 ( .A1(n9840), .A2(n7905), .A3(n7904), .A4(n7040), .ZN(n7909)
         );
  NOR3_X1 U9532 ( .A1(n7944), .A2(n7906), .A3(n8072), .ZN(n7907) );
  NAND4_X1 U9533 ( .A1(n7909), .A2(n7957), .A3(n7908), .A4(n7907), .ZN(n7911)
         );
  NOR4_X1 U9534 ( .A1(n7911), .A2(n6443), .A3(n7910), .A4(n6439), .ZN(n7912)
         );
  AND4_X1 U9535 ( .A1(n7977), .A2(n7913), .A3(n4985), .A4(n7912), .ZN(n7914)
         );
  NAND4_X1 U9536 ( .A1(n8542), .A2(n7994), .A3(n7989), .A4(n7914), .ZN(n7915)
         );
  NOR4_X1 U9537 ( .A1(n8496), .A2(n8532), .A3(n8511), .A4(n7915), .ZN(n7916)
         );
  NAND4_X1 U9538 ( .A1(n8450), .A2(n4786), .A3(n8461), .A4(n7916), .ZN(n7917)
         );
  NOR4_X1 U9539 ( .A1(n8393), .A2(n7918), .A3(n8435), .A4(n7917), .ZN(n7920)
         );
  INV_X1 U9540 ( .A(n8368), .ZN(n7919) );
  NAND4_X1 U9541 ( .A1(n8051), .A2(n7920), .A3(n8405), .A4(n7919), .ZN(n7921)
         );
  XNOR2_X1 U9542 ( .A(n7922), .B(n7923), .ZN(n8068) );
  NOR2_X1 U9543 ( .A1(n8252), .A2(n8059), .ZN(n8045) );
  INV_X1 U9544 ( .A(n7924), .ZN(n7928) );
  INV_X1 U9545 ( .A(n7950), .ZN(n7925) );
  INV_X1 U9546 ( .A(n7952), .ZN(n7927) );
  OAI21_X1 U9547 ( .B1(n7929), .B2(n7928), .A(n7927), .ZN(n7931) );
  NAND3_X1 U9548 ( .A1(n7931), .A2(n7958), .A3(n7930), .ZN(n7947) );
  NAND2_X1 U9549 ( .A1(n7933), .A2(n7932), .ZN(n7936) );
  NAND3_X1 U9550 ( .A1(n7936), .A2(n7938), .A3(n7934), .ZN(n7935) );
  AND2_X1 U9551 ( .A1(n7935), .A2(n7940), .ZN(n7943) );
  OAI21_X1 U9552 ( .B1(n7937), .B2(n7936), .A(n7058), .ZN(n7941) );
  INV_X1 U9553 ( .A(n7938), .ZN(n7939) );
  AOI21_X1 U9554 ( .B1(n7941), .B2(n7940), .A(n7939), .ZN(n7942) );
  MUX2_X1 U9555 ( .A(n7943), .B(n7942), .S(n8059), .Z(n7945) );
  NOR3_X1 U9556 ( .A1(n7945), .A2(n7944), .A3(n7952), .ZN(n7946) );
  AOI21_X1 U9557 ( .B1(n8059), .B2(n7947), .A(n7946), .ZN(n7956) );
  INV_X1 U9558 ( .A(n7948), .ZN(n7955) );
  AOI22_X1 U9559 ( .A1(n7952), .A2(n7951), .B1(n7950), .B2(n7949), .ZN(n7953)
         );
  NOR2_X1 U9560 ( .A1(n7953), .A2(n7955), .ZN(n7954) );
  MUX2_X1 U9561 ( .A(n7960), .B(n7959), .S(n8059), .Z(n7961) );
  MUX2_X1 U9562 ( .A(n7964), .B(n7963), .S(n8059), .Z(n7965) );
  INV_X1 U9563 ( .A(n7970), .ZN(n7968) );
  OAI21_X1 U9564 ( .B1(n7968), .B2(n4765), .A(n7967), .ZN(n7975) );
  INV_X1 U9565 ( .A(n7971), .ZN(n7973) );
  MUX2_X1 U9566 ( .A(n7975), .B(n7974), .S(n8059), .Z(n7980) );
  OAI21_X1 U9567 ( .B1(n7978), .B2(n8059), .A(n7977), .ZN(n7988) );
  NAND3_X1 U9568 ( .A1(n7979), .A2(n4722), .A3(n8262), .ZN(n7987) );
  INV_X1 U9569 ( .A(n7980), .ZN(n7985) );
  NAND2_X1 U9570 ( .A1(n7982), .A2(n7981), .ZN(n7984) );
  OAI21_X1 U9571 ( .B1(n4722), .B2(n7990), .A(n7989), .ZN(n7995) );
  MUX2_X1 U9572 ( .A(n7992), .B(n7991), .S(n8059), .Z(n7993) );
  MUX2_X1 U9573 ( .A(n7997), .B(n7996), .S(n8059), .Z(n7998) );
  MUX2_X1 U9574 ( .A(n8000), .B(n7999), .S(n8059), .Z(n8001) );
  NOR2_X1 U9575 ( .A1(n8673), .A2(n8259), .ZN(n8004) );
  NAND2_X1 U9576 ( .A1(n8007), .A2(n8002), .ZN(n8003) );
  MUX2_X1 U9577 ( .A(n8004), .B(n8003), .S(n8059), .Z(n8005) );
  INV_X1 U9578 ( .A(n8013), .ZN(n8009) );
  INV_X1 U9579 ( .A(n8015), .ZN(n8008) );
  AOI211_X1 U9580 ( .C1(n8009), .C2(n8012), .A(n4785), .B(n8008), .ZN(n8011)
         );
  INV_X1 U9581 ( .A(n8018), .ZN(n8010) );
  NOR2_X1 U9582 ( .A1(n8011), .A2(n8010), .ZN(n8022) );
  NAND2_X1 U9583 ( .A1(n8013), .A2(n8012), .ZN(n8016) );
  INV_X1 U9584 ( .A(n8014), .ZN(n8023) );
  INV_X1 U9585 ( .A(n8019), .ZN(n8021) );
  AOI22_X1 U9586 ( .A1(n8019), .A2(n8018), .B1(n4722), .B2(n8017), .ZN(n8020)
         );
  AOI21_X1 U9587 ( .B1(n8022), .B2(n8021), .A(n8020), .ZN(n8032) );
  AOI21_X1 U9588 ( .B1(n8027), .B2(n4536), .A(n8026), .ZN(n8029) );
  OAI211_X1 U9589 ( .C1(n8029), .C2(n8435), .A(n8417), .B(n8028), .ZN(n8030)
         );
  AND3_X1 U9590 ( .A1(n8030), .A2(n8405), .A3(n8035), .ZN(n8039) );
  INV_X1 U9591 ( .A(n8393), .ZN(n8388) );
  OAI211_X1 U9592 ( .C1(n8653), .C2(n8253), .A(n8037), .B(n8388), .ZN(n8038)
         );
  MUX2_X1 U9593 ( .A(n8039), .B(n8038), .S(n8059), .Z(n8043) );
  AOI21_X1 U9594 ( .B1(n8042), .B2(n8040), .A(n8059), .ZN(n8041) );
  AOI21_X1 U9595 ( .B1(n8043), .B2(n8042), .A(n8041), .ZN(n8044) );
  INV_X1 U9596 ( .A(n8227), .ZN(n8251) );
  NOR2_X1 U9597 ( .A1(n4707), .A2(n8251), .ZN(n8046) );
  MUX2_X1 U9598 ( .A(n8047), .B(n8046), .S(n8059), .Z(n8048) );
  NAND3_X1 U9599 ( .A1(n8364), .A2(n8250), .A3(n8059), .ZN(n8050) );
  NAND3_X1 U9600 ( .A1(n8569), .A2(n8105), .A3(n4722), .ZN(n8049) );
  MUX2_X1 U9601 ( .A(n8053), .B(n8052), .S(n8059), .Z(n8054) );
  MUX2_X1 U9602 ( .A(n8058), .B(n8057), .S(n8059), .Z(n8063) );
  MUX2_X1 U9603 ( .A(n8061), .B(n8060), .S(n8059), .Z(n8062) );
  OAI21_X1 U9604 ( .B1(n8064), .B2(n8063), .A(n8062), .ZN(n8073) );
  INV_X1 U9605 ( .A(n8065), .ZN(n8066) );
  OAI21_X1 U9606 ( .B1(n8069), .B2(n8068), .A(n8067), .ZN(n8075) );
  INV_X1 U9607 ( .A(n8070), .ZN(n8071) );
  NAND3_X1 U9608 ( .A1(n8073), .A2(n8072), .A3(n8071), .ZN(n8074) );
  AOI22_X1 U9609 ( .A1(n8077), .A2(n8076), .B1(n8075), .B2(n8074), .ZN(n8083)
         );
  NOR3_X1 U9610 ( .A1(n8078), .A2(n9812), .A3(n6496), .ZN(n8081) );
  OAI21_X1 U9611 ( .B1(n8082), .B2(n8079), .A(P2_B_REG_SCAN_IN), .ZN(n8080) );
  OAI21_X1 U9612 ( .B1(n4554), .B2(n8085), .A(n8084), .ZN(n8086) );
  NAND2_X1 U9613 ( .A1(n8086), .A2(n9821), .ZN(n8090) );
  AOI22_X1 U9614 ( .A1(n9817), .A2(n8088), .B1(n8087), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n8089) );
  OAI211_X1 U9615 ( .C1(n6422), .C2(n9819), .A(n8090), .B(n8089), .ZN(P2_U3224) );
  INV_X1 U9616 ( .A(n8851), .ZN(n8688) );
  INV_X1 U9617 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8091) );
  OAI222_X1 U9618 ( .A1(n9513), .A2(n8688), .B1(n8092), .B2(P1_U3084), .C1(
        n8091), .C2(n9522), .ZN(P1_U3324) );
  NAND2_X1 U9619 ( .A1(n8093), .A2(n9853), .ZN(n8101) );
  INV_X1 U9620 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8095) );
  OAI22_X1 U9621 ( .A1(n8553), .A2(n8095), .B1(n8094), .B2(n9845), .ZN(n8098)
         );
  NOR2_X1 U9622 ( .A1(n8096), .A2(n9847), .ZN(n8097) );
  AOI211_X1 U9623 ( .C1(n8534), .C2(n8099), .A(n8098), .B(n8097), .ZN(n8100)
         );
  OAI211_X1 U9624 ( .C1(n8102), .C2(n9849), .A(n8101), .B(n8100), .ZN(P2_U3267) );
  XNOR2_X1 U9625 ( .A(n8104), .B(n8103), .ZN(n8110) );
  INV_X1 U9626 ( .A(n8378), .ZN(n8107) );
  OAI22_X1 U9627 ( .A1(n8105), .A2(n9814), .B1(n8157), .B2(n9812), .ZN(n8373)
         );
  AOI22_X1 U9628 ( .A1(n8373), .A2(n9817), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8106) );
  OAI21_X1 U9629 ( .B1(n8107), .B2(n9824), .A(n8106), .ZN(n8108) );
  AOI21_X1 U9630 ( .B1(n8377), .B2(n8244), .A(n8108), .ZN(n8109) );
  OAI21_X1 U9631 ( .B1(n8110), .B2(n8247), .A(n8109), .ZN(P2_U3216) );
  INV_X1 U9632 ( .A(n8111), .ZN(n8112) );
  AOI21_X1 U9633 ( .B1(n8114), .B2(n8113), .A(n8112), .ZN(n8122) );
  AOI21_X1 U9634 ( .B1(n9817), .B2(n8116), .A(n8115), .ZN(n8117) );
  OAI21_X1 U9635 ( .B1(n8118), .B2(n9824), .A(n8117), .ZN(n8119) );
  AOI21_X1 U9636 ( .B1(n8120), .B2(n8244), .A(n8119), .ZN(n8121) );
  OAI21_X1 U9637 ( .B1(n8122), .B2(n8247), .A(n8121), .ZN(P2_U3217) );
  INV_X1 U9638 ( .A(n8441), .ZN(n8125) );
  OAI22_X1 U9639 ( .A1(n8123), .A2(n9814), .B1(n8147), .B2(n9812), .ZN(n8437)
         );
  AOI22_X1 U9640 ( .A1(n8437), .A2(n9817), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8124) );
  OAI21_X1 U9641 ( .B1(n8125), .B2(n9824), .A(n8124), .ZN(n8130) );
  INV_X1 U9642 ( .A(n8126), .ZN(n8128) );
  NOR2_X1 U9643 ( .A1(n8128), .A2(n8127), .ZN(n8187) );
  AOI211_X1 U9644 ( .C1(n8128), .C2(n8127), .A(n8247), .B(n8187), .ZN(n8129)
         );
  AOI211_X1 U9645 ( .C1(n8442), .C2(n8244), .A(n8130), .B(n8129), .ZN(n8131)
         );
  INV_X1 U9646 ( .A(n8131), .ZN(P2_U3218) );
  INV_X1 U9647 ( .A(n8132), .ZN(n8133) );
  AOI21_X1 U9648 ( .B1(n8135), .B2(n8134), .A(n8133), .ZN(n8141) );
  OR2_X1 U9649 ( .A1(n8146), .A2(n9814), .ZN(n8137) );
  NAND2_X1 U9650 ( .A1(n8258), .A2(n8228), .ZN(n8136) );
  NAND2_X1 U9651 ( .A1(n8137), .A2(n8136), .ZN(n8498) );
  AOI22_X1 U9652 ( .A1(n9817), .A2(n8498), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8138) );
  OAI21_X1 U9653 ( .B1(n8494), .B2(n9824), .A(n8138), .ZN(n8139) );
  AOI21_X1 U9654 ( .B1(n8614), .B2(n8244), .A(n8139), .ZN(n8140) );
  OAI21_X1 U9655 ( .B1(n8141), .B2(n8247), .A(n8140), .ZN(P2_U3221) );
  OAI211_X1 U9656 ( .C1(n8144), .C2(n8143), .A(n8142), .B(n9821), .ZN(n8151)
         );
  INV_X1 U9657 ( .A(n8145), .ZN(n8466) );
  OAI22_X1 U9658 ( .A1(n8147), .A2(n9814), .B1(n8146), .B2(n9812), .ZN(n8473)
         );
  INV_X1 U9659 ( .A(n8473), .ZN(n8148) );
  OAI22_X1 U9660 ( .A1(n8148), .A2(n8233), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10176), .ZN(n8149) );
  AOI21_X1 U9661 ( .B1(n8466), .B2(n8231), .A(n8149), .ZN(n8150) );
  OAI211_X1 U9662 ( .C1(n8468), .C2(n9819), .A(n8151), .B(n8150), .ZN(P2_U3225) );
  INV_X1 U9663 ( .A(n8152), .ZN(n8154) );
  NOR2_X1 U9664 ( .A1(n8154), .A2(n8153), .ZN(n8155) );
  XNOR2_X1 U9665 ( .A(n8156), .B(n8155), .ZN(n8163) );
  OR2_X1 U9666 ( .A1(n8157), .A2(n9814), .ZN(n8159) );
  NAND2_X1 U9667 ( .A1(n4999), .A2(n8228), .ZN(n8158) );
  NAND2_X1 U9668 ( .A1(n8159), .A2(n8158), .ZN(n8402) );
  AOI22_X1 U9669 ( .A1(n8402), .A2(n9817), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8160) );
  OAI21_X1 U9670 ( .B1(n8407), .B2(n9824), .A(n8160), .ZN(n8161) );
  AOI21_X1 U9671 ( .B1(n8410), .B2(n8244), .A(n8161), .ZN(n8162) );
  OAI21_X1 U9672 ( .B1(n8163), .B2(n8247), .A(n8162), .ZN(P2_U3227) );
  XNOR2_X1 U9673 ( .A(n8164), .B(n8165), .ZN(n8238) );
  NOR2_X1 U9674 ( .A1(n8238), .A2(n8239), .ZN(n8237) );
  AOI21_X1 U9675 ( .B1(n8164), .B2(n8165), .A(n8237), .ZN(n8169) );
  XNOR2_X1 U9676 ( .A(n8167), .B(n8166), .ZN(n8168) );
  XNOR2_X1 U9677 ( .A(n8169), .B(n8168), .ZN(n8176) );
  OAI22_X1 U9678 ( .A1(n8170), .A2(n9812), .B1(n8217), .B2(n9814), .ZN(n8544)
         );
  NAND2_X1 U9679 ( .A1(n9817), .A2(n8544), .ZN(n8173) );
  NOR2_X1 U9680 ( .A1(n8171), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8289) );
  INV_X1 U9681 ( .A(n8289), .ZN(n8172) );
  OAI211_X1 U9682 ( .C1(n9824), .C2(n8551), .A(n8173), .B(n8172), .ZN(n8174)
         );
  AOI21_X1 U9683 ( .B1(n8550), .B2(n8244), .A(n8174), .ZN(n8175) );
  OAI21_X1 U9684 ( .B1(n8176), .B2(n8247), .A(n8175), .ZN(P2_U3228) );
  AOI21_X1 U9685 ( .B1(n8178), .B2(n8177), .A(n8247), .ZN(n8180) );
  NAND2_X1 U9686 ( .A1(n8180), .A2(n8179), .ZN(n8185) );
  INV_X1 U9687 ( .A(n8524), .ZN(n8183) );
  AOI22_X1 U9688 ( .A1(n8260), .A2(n8228), .B1(n8218), .B2(n8258), .ZN(n8526)
         );
  OAI22_X1 U9689 ( .A1(n8526), .A2(n8233), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8181), .ZN(n8182) );
  AOI21_X1 U9690 ( .B1(n8183), .B2(n8231), .A(n8182), .ZN(n8184) );
  OAI211_X1 U9691 ( .C1(n8673), .C2(n9819), .A(n8185), .B(n8184), .ZN(P2_U3230) );
  NOR2_X1 U9692 ( .A1(n8187), .A2(n8186), .ZN(n8191) );
  XNOR2_X1 U9693 ( .A(n8189), .B(n8188), .ZN(n8190) );
  XNOR2_X1 U9694 ( .A(n8191), .B(n8190), .ZN(n8197) );
  NAND2_X1 U9695 ( .A1(n8253), .A2(n8218), .ZN(n8193) );
  NAND2_X1 U9696 ( .A1(n8254), .A2(n8228), .ZN(n8192) );
  NAND2_X1 U9697 ( .A1(n8193), .A2(n8192), .ZN(n8419) );
  AOI22_X1 U9698 ( .A1(n8419), .A2(n9817), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8194) );
  OAI21_X1 U9699 ( .B1(n8424), .B2(n9824), .A(n8194), .ZN(n8195) );
  AOI21_X1 U9700 ( .B1(n8590), .B2(n8244), .A(n8195), .ZN(n8196) );
  OAI21_X1 U9701 ( .B1(n8197), .B2(n8247), .A(n8196), .ZN(P2_U3231) );
  OAI211_X1 U9702 ( .C1(n4547), .C2(n8199), .A(n8198), .B(n9821), .ZN(n8204)
         );
  OAI22_X1 U9703 ( .A1(n8207), .A2(n9814), .B1(n8200), .B2(n9812), .ZN(n8481)
         );
  AOI22_X1 U9704 ( .A1(n9817), .A2(n8481), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8201) );
  OAI21_X1 U9705 ( .B1(n8478), .B2(n9824), .A(n8201), .ZN(n8202) );
  AOI21_X1 U9706 ( .B1(n8487), .B2(n8244), .A(n8202), .ZN(n8203) );
  NAND2_X1 U9707 ( .A1(n8204), .A2(n8203), .ZN(P2_U3235) );
  XOR2_X1 U9708 ( .A(n8206), .B(n8205), .Z(n8213) );
  INV_X1 U9709 ( .A(n8455), .ZN(n8210) );
  OAI22_X1 U9710 ( .A1(n8208), .A2(n9814), .B1(n8207), .B2(n9812), .ZN(n8451)
         );
  AOI22_X1 U9711 ( .A1(n8451), .A2(n9817), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8209) );
  OAI21_X1 U9712 ( .B1(n8210), .B2(n9824), .A(n8209), .ZN(n8211) );
  AOI21_X1 U9713 ( .B1(n8600), .B2(n8244), .A(n8211), .ZN(n8212) );
  OAI21_X1 U9714 ( .B1(n8213), .B2(n8247), .A(n8212), .ZN(P2_U3237) );
  OAI211_X1 U9715 ( .C1(n8216), .C2(n8215), .A(n8214), .B(n9821), .ZN(n8224)
         );
  INV_X1 U9716 ( .A(n8515), .ZN(n8222) );
  OR2_X1 U9717 ( .A1(n8217), .A2(n9812), .ZN(n8220) );
  NAND2_X1 U9718 ( .A1(n8257), .A2(n8218), .ZN(n8219) );
  AND2_X1 U9719 ( .A1(n8220), .A2(n8219), .ZN(n8509) );
  OAI22_X1 U9720 ( .A1(n8509), .A2(n8233), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8317), .ZN(n8221) );
  AOI21_X1 U9721 ( .B1(n8222), .B2(n8231), .A(n8221), .ZN(n8223) );
  OAI211_X1 U9722 ( .C1(n8669), .C2(n9819), .A(n8224), .B(n8223), .ZN(P2_U3240) );
  XNOR2_X1 U9723 ( .A(n8226), .B(n8225), .ZN(n8236) );
  OR2_X1 U9724 ( .A1(n8227), .A2(n9814), .ZN(n8230) );
  NAND2_X1 U9725 ( .A1(n8253), .A2(n8228), .ZN(n8229) );
  AND2_X1 U9726 ( .A1(n8230), .A2(n8229), .ZN(n8390) );
  AOI22_X1 U9727 ( .A1(n8231), .A2(n8386), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8232) );
  OAI21_X1 U9728 ( .B1(n8390), .B2(n8233), .A(n8232), .ZN(n8234) );
  AOI21_X1 U9729 ( .B1(n8577), .B2(n8244), .A(n8234), .ZN(n8235) );
  OAI21_X1 U9730 ( .B1(n8236), .B2(n8247), .A(n8235), .ZN(P2_U3242) );
  AOI21_X1 U9731 ( .B1(n8239), .B2(n8238), .A(n8237), .ZN(n8248) );
  AOI22_X1 U9732 ( .A1(n9817), .A2(n8240), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n8241) );
  OAI21_X1 U9733 ( .B1(n8242), .B2(n9824), .A(n8241), .ZN(n8243) );
  AOI21_X1 U9734 ( .B1(n8245), .B2(n8244), .A(n8243), .ZN(n8246) );
  OAI21_X1 U9735 ( .B1(n8248), .B2(n8247), .A(n8246), .ZN(P2_U3243) );
  MUX2_X1 U9736 ( .A(n8249), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8275), .Z(
        P2_U3582) );
  MUX2_X1 U9737 ( .A(n8250), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8275), .Z(
        P2_U3580) );
  MUX2_X1 U9738 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8251), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9739 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8252), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U9740 ( .A(n8253), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8275), .Z(
        P2_U3577) );
  MUX2_X1 U9741 ( .A(n4999), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8275), .Z(
        P2_U3576) );
  MUX2_X1 U9742 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8254), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9743 ( .A(n8255), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8275), .Z(
        P2_U3573) );
  MUX2_X1 U9744 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8256), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9745 ( .A(n8257), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8275), .Z(
        P2_U3571) );
  MUX2_X1 U9746 ( .A(n8258), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8275), .Z(
        P2_U3570) );
  MUX2_X1 U9747 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8259), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9748 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8260), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9749 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8261), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9750 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8262), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9751 ( .A(n8263), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8275), .Z(
        P2_U3564) );
  MUX2_X1 U9752 ( .A(n8264), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8275), .Z(
        P2_U3563) );
  MUX2_X1 U9753 ( .A(n8265), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8275), .Z(
        P2_U3562) );
  MUX2_X1 U9754 ( .A(n8266), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8275), .Z(
        P2_U3561) );
  MUX2_X1 U9755 ( .A(n8267), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8275), .Z(
        P2_U3560) );
  MUX2_X1 U9756 ( .A(n8268), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8275), .Z(
        P2_U3559) );
  MUX2_X1 U9757 ( .A(n8269), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8275), .Z(
        P2_U3558) );
  MUX2_X1 U9758 ( .A(n8270), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8275), .Z(
        P2_U3557) );
  MUX2_X1 U9759 ( .A(n8271), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8275), .Z(
        P2_U3556) );
  MUX2_X1 U9760 ( .A(n8272), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8275), .Z(
        P2_U3555) );
  MUX2_X1 U9761 ( .A(n8273), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8275), .Z(
        P2_U3554) );
  MUX2_X1 U9762 ( .A(n8274), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8275), .Z(
        P2_U3553) );
  MUX2_X1 U9763 ( .A(n6475), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8275), .Z(
        P2_U3552) );
  NOR2_X1 U9764 ( .A1(n8277), .A2(n8276), .ZN(n8279) );
  NOR2_X1 U9765 ( .A1(n8279), .A2(n8278), .ZN(n8281) );
  XNOR2_X1 U9766 ( .A(n8304), .B(n8632), .ZN(n8280) );
  NAND2_X1 U9767 ( .A1(n8280), .A2(n8281), .ZN(n8305) );
  OAI21_X1 U9768 ( .B1(n8281), .B2(n8280), .A(n8305), .ZN(n8294) );
  NOR2_X1 U9769 ( .A1(n8283), .A2(n8282), .ZN(n8285) );
  NOR2_X1 U9770 ( .A1(n8285), .A2(n8284), .ZN(n8288) );
  NAND2_X1 U9771 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8304), .ZN(n8297) );
  INV_X1 U9772 ( .A(n8297), .ZN(n8286) );
  AOI21_X1 U9773 ( .B1(n8552), .B2(n8292), .A(n8286), .ZN(n8287) );
  NAND2_X1 U9774 ( .A1(n8287), .A2(n8288), .ZN(n8296) );
  OAI211_X1 U9775 ( .C1(n8288), .C2(n8287), .A(n9825), .B(n8296), .ZN(n8291)
         );
  AOI21_X1 U9776 ( .B1(n9832), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8289), .ZN(
        n8290) );
  OAI211_X1 U9777 ( .C1(n9828), .C2(n8292), .A(n8291), .B(n8290), .ZN(n8293)
         );
  AOI21_X1 U9778 ( .B1(n8294), .B2(n9827), .A(n8293), .ZN(n8295) );
  INV_X1 U9779 ( .A(n8295), .ZN(P2_U3261) );
  NAND2_X1 U9780 ( .A1(n8297), .A2(n8296), .ZN(n8301) );
  INV_X1 U9781 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8299) );
  NAND2_X1 U9782 ( .A1(n8321), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8315) );
  INV_X1 U9783 ( .A(n8315), .ZN(n8298) );
  AOI21_X1 U9784 ( .B1(n8299), .B2(n8303), .A(n8298), .ZN(n8300) );
  NAND2_X1 U9785 ( .A1(n8300), .A2(n8301), .ZN(n8314) );
  OAI211_X1 U9786 ( .C1(n8301), .C2(n8300), .A(n9825), .B(n8314), .ZN(n8313)
         );
  NOR2_X1 U9787 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8181), .ZN(n8302) );
  AOI21_X1 U9788 ( .B1(n9832), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8302), .ZN(
        n8312) );
  OR2_X1 U9789 ( .A1(n9828), .A2(n8303), .ZN(n8311) );
  XNOR2_X1 U9790 ( .A(n8321), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8308) );
  OR2_X1 U9791 ( .A1(n8304), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U9792 ( .A1(n8306), .A2(n8305), .ZN(n8307) );
  NOR2_X1 U9793 ( .A1(n8308), .A2(n8307), .ZN(n8320) );
  AOI21_X1 U9794 ( .B1(n8308), .B2(n8307), .A(n8320), .ZN(n8309) );
  NAND2_X1 U9795 ( .A1(n9827), .A2(n8309), .ZN(n8310) );
  NAND4_X1 U9796 ( .A1(n8313), .A2(n8312), .A3(n8311), .A4(n8310), .ZN(
        P2_U3262) );
  NAND2_X1 U9797 ( .A1(n8315), .A2(n8314), .ZN(n8331) );
  XOR2_X1 U9798 ( .A(n8332), .B(n8331), .Z(n8316) );
  NAND2_X1 U9799 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8316), .ZN(n8334) );
  OAI211_X1 U9800 ( .C1(n8316), .C2(P2_REG2_REG_18__SCAN_IN), .A(n9825), .B(
        n8334), .ZN(n8328) );
  NOR2_X1 U9801 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8317), .ZN(n8318) );
  AOI21_X1 U9802 ( .B1(n9832), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8318), .ZN(
        n8327) );
  OR2_X1 U9803 ( .A1(n9828), .A2(n8319), .ZN(n8326) );
  XNOR2_X1 U9804 ( .A(n8332), .B(n8621), .ZN(n8323) );
  OAI21_X1 U9805 ( .B1(n8323), .B2(n8322), .A(n8329), .ZN(n8324) );
  NAND2_X1 U9806 ( .A1(n9827), .A2(n8324), .ZN(n8325) );
  NAND4_X1 U9807 ( .A1(n8328), .A2(n8327), .A3(n8326), .A4(n8325), .ZN(
        P2_U3263) );
  INV_X1 U9808 ( .A(n8339), .ZN(n8337) );
  NAND2_X1 U9809 ( .A1(n8332), .A2(n8331), .ZN(n8333) );
  NAND2_X1 U9810 ( .A1(n8334), .A2(n8333), .ZN(n8335) );
  XOR2_X1 U9811 ( .A(n8335), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8338) );
  OAI21_X1 U9812 ( .B1(n8338), .B2(n9830), .A(n9828), .ZN(n8336) );
  AOI21_X1 U9813 ( .B1(n8337), .B2(n9827), .A(n8336), .ZN(n8341) );
  AOI22_X1 U9814 ( .A1(n8339), .A2(n9827), .B1(n9825), .B2(n8338), .ZN(n8340)
         );
  MUX2_X1 U9815 ( .A(n8341), .B(n8340), .S(n8530), .Z(n8343) );
  NAND2_X1 U9816 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8342) );
  OAI211_X1 U9817 ( .C1(n9537), .C2(n4856), .A(n8343), .B(n8342), .ZN(P2_U3264) );
  INV_X1 U9818 ( .A(n8344), .ZN(n8351) );
  NAND2_X1 U9819 ( .A1(n8642), .A2(n8351), .ZN(n8350) );
  NOR2_X1 U9820 ( .A1(n8553), .A2(n8345), .ZN(n8348) );
  NAND2_X1 U9821 ( .A1(n8347), .A2(n8346), .ZN(n8563) );
  NOR2_X1 U9822 ( .A1(n9849), .A2(n8563), .ZN(n8353) );
  AOI211_X1 U9823 ( .C1(n8560), .C2(n8534), .A(n8348), .B(n8353), .ZN(n8349)
         );
  OAI21_X1 U9824 ( .B1(n8561), .B2(n9847), .A(n8349), .ZN(P2_U3265) );
  OAI211_X1 U9825 ( .C1(n8642), .C2(n8351), .A(n9841), .B(n8350), .ZN(n8564)
         );
  NOR2_X1 U9826 ( .A1(n8642), .A2(n9851), .ZN(n8352) );
  AOI211_X1 U9827 ( .C1(n9849), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8353), .B(
        n8352), .ZN(n8354) );
  OAI21_X1 U9828 ( .B1(n9847), .B2(n8564), .A(n8354), .ZN(P2_U3266) );
  XOR2_X1 U9829 ( .A(n8356), .B(n8355), .Z(n8571) );
  OAI21_X1 U9830 ( .B1(n4517), .B2(n4774), .A(n9838), .ZN(n8359) );
  OAI21_X1 U9831 ( .B1(n8359), .B2(n8358), .A(n8357), .ZN(n8567) );
  AOI211_X1 U9832 ( .C1(n8569), .C2(n4709), .A(n9942), .B(n8360), .ZN(n8568)
         );
  NAND2_X1 U9833 ( .A1(n8568), .A2(n8556), .ZN(n8363) );
  AOI22_X1 U9834 ( .A1(n8361), .A2(n8483), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9849), .ZN(n8362) );
  OAI211_X1 U9835 ( .C1(n8364), .C2(n9851), .A(n8363), .B(n8362), .ZN(n8365)
         );
  AOI21_X1 U9836 ( .B1(n8567), .B2(n8553), .A(n8365), .ZN(n8366) );
  OAI21_X1 U9837 ( .B1(n8571), .B2(n8506), .A(n8366), .ZN(P2_U3268) );
  XNOR2_X1 U9838 ( .A(n8367), .B(n8368), .ZN(n8574) );
  INV_X1 U9839 ( .A(n8574), .ZN(n8383) );
  NAND2_X1 U9840 ( .A1(n8369), .A2(n8368), .ZN(n8370) );
  NAND2_X1 U9841 ( .A1(n8370), .A2(n9838), .ZN(n8371) );
  OR2_X1 U9842 ( .A1(n8372), .A2(n8371), .ZN(n8375) );
  INV_X1 U9843 ( .A(n8373), .ZN(n8374) );
  NAND2_X1 U9844 ( .A1(n8375), .A2(n8374), .ZN(n8572) );
  AOI211_X1 U9845 ( .C1(n8377), .C2(n8384), .A(n9942), .B(n8376), .ZN(n8573)
         );
  NAND2_X1 U9846 ( .A1(n8573), .A2(n8556), .ZN(n8380) );
  AOI22_X1 U9847 ( .A1(n8378), .A2(n8483), .B1(n9849), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8379) );
  OAI211_X1 U9848 ( .C1(n4707), .C2(n9851), .A(n8380), .B(n8379), .ZN(n8381)
         );
  AOI21_X1 U9849 ( .B1(n8572), .B2(n8553), .A(n8381), .ZN(n8382) );
  OAI21_X1 U9850 ( .B1(n8383), .B2(n8506), .A(n8382), .ZN(P2_U3269) );
  INV_X1 U9851 ( .A(n8384), .ZN(n8385) );
  AOI211_X1 U9852 ( .C1(n8577), .C2(n8398), .A(n9942), .B(n8385), .ZN(n8579)
         );
  INV_X1 U9853 ( .A(n8386), .ZN(n8387) );
  NOR2_X1 U9854 ( .A1(n8387), .A2(n9845), .ZN(n8392) );
  XNOR2_X1 U9855 ( .A(n8389), .B(n8388), .ZN(n8391) );
  OAI21_X1 U9856 ( .B1(n8391), .B2(n8527), .A(n8390), .ZN(n8578) );
  AOI211_X1 U9857 ( .C1(n8579), .C2(n8530), .A(n8392), .B(n8578), .ZN(n8397)
         );
  XNOR2_X1 U9858 ( .A(n8394), .B(n8393), .ZN(n8580) );
  NAND2_X1 U9859 ( .A1(n8580), .A2(n9853), .ZN(n8396) );
  AOI22_X1 U9860 ( .A1(n8577), .A2(n8534), .B1(n9849), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8395) );
  OAI211_X1 U9861 ( .C1(n9855), .C2(n8397), .A(n8396), .B(n8395), .ZN(P2_U3270) );
  INV_X1 U9862 ( .A(n8423), .ZN(n8400) );
  INV_X1 U9863 ( .A(n8398), .ZN(n8399) );
  AOI211_X1 U9864 ( .C1(n8410), .C2(n8400), .A(n9942), .B(n8399), .ZN(n8584)
         );
  XNOR2_X1 U9865 ( .A(n8401), .B(n8405), .ZN(n8404) );
  INV_X1 U9866 ( .A(n8402), .ZN(n8403) );
  OAI21_X1 U9867 ( .B1(n8404), .B2(n8527), .A(n8403), .ZN(n8583) );
  AOI21_X1 U9868 ( .B1(n8584), .B2(n8530), .A(n8583), .ZN(n8413) );
  XNOR2_X1 U9869 ( .A(n8406), .B(n8405), .ZN(n8585) );
  NAND2_X1 U9870 ( .A1(n8585), .A2(n9853), .ZN(n8412) );
  INV_X1 U9871 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8408) );
  OAI22_X1 U9872 ( .A1(n8553), .A2(n8408), .B1(n8407), .B2(n9845), .ZN(n8409)
         );
  AOI21_X1 U9873 ( .B1(n8410), .B2(n8534), .A(n8409), .ZN(n8411) );
  OAI211_X1 U9874 ( .C1(n9855), .C2(n8413), .A(n8412), .B(n8411), .ZN(P2_U3271) );
  AOI21_X1 U9875 ( .B1(n8417), .B2(n8415), .A(n8414), .ZN(n8592) );
  OAI211_X1 U9876 ( .C1(n8418), .C2(n8417), .A(n8416), .B(n9838), .ZN(n8421)
         );
  INV_X1 U9877 ( .A(n8419), .ZN(n8420) );
  NAND2_X1 U9878 ( .A1(n8421), .A2(n8420), .ZN(n8588) );
  INV_X1 U9879 ( .A(n8422), .ZN(n8440) );
  AOI211_X1 U9880 ( .C1(n8590), .C2(n8440), .A(n9942), .B(n8423), .ZN(n8589)
         );
  NAND2_X1 U9881 ( .A1(n8589), .A2(n8556), .ZN(n8427) );
  INV_X1 U9882 ( .A(n8424), .ZN(n8425) );
  AOI22_X1 U9883 ( .A1(n9849), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8425), .B2(
        n8483), .ZN(n8426) );
  OAI211_X1 U9884 ( .C1(n8428), .C2(n9851), .A(n8427), .B(n8426), .ZN(n8429)
         );
  AOI21_X1 U9885 ( .B1(n8588), .B2(n8553), .A(n8429), .ZN(n8430) );
  OAI21_X1 U9886 ( .B1(n8592), .B2(n8506), .A(n8430), .ZN(P2_U3272) );
  OAI21_X1 U9887 ( .B1(n8432), .B2(n8435), .A(n8431), .ZN(n8595) );
  NAND2_X1 U9888 ( .A1(n8433), .A2(n8434), .ZN(n8436) );
  XNOR2_X1 U9889 ( .A(n8436), .B(n8435), .ZN(n8438) );
  AOI21_X1 U9890 ( .B1(n8438), .B2(n9838), .A(n8437), .ZN(n8594) );
  INV_X1 U9891 ( .A(n8594), .ZN(n8446) );
  INV_X1 U9892 ( .A(n8439), .ZN(n8454) );
  OAI211_X1 U9893 ( .C1(n8658), .C2(n8454), .A(n8440), .B(n9841), .ZN(n8593)
         );
  AOI22_X1 U9894 ( .A1(n9849), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8441), .B2(
        n8483), .ZN(n8444) );
  NAND2_X1 U9895 ( .A1(n8442), .A2(n8534), .ZN(n8443) );
  OAI211_X1 U9896 ( .C1(n8593), .C2(n9847), .A(n8444), .B(n8443), .ZN(n8445)
         );
  AOI21_X1 U9897 ( .B1(n8446), .B2(n8553), .A(n8445), .ZN(n8447) );
  OAI21_X1 U9898 ( .B1(n8595), .B2(n8506), .A(n8447), .ZN(P2_U3273) );
  XNOR2_X1 U9899 ( .A(n8448), .B(n8450), .ZN(n8602) );
  OAI211_X1 U9900 ( .C1(n8450), .C2(n8449), .A(n8433), .B(n9838), .ZN(n8453)
         );
  INV_X1 U9901 ( .A(n8451), .ZN(n8452) );
  NAND2_X1 U9902 ( .A1(n8453), .A2(n8452), .ZN(n8598) );
  AOI211_X1 U9903 ( .C1(n8600), .C2(n8463), .A(n9942), .B(n8454), .ZN(n8599)
         );
  NAND2_X1 U9904 ( .A1(n8599), .A2(n8556), .ZN(n8457) );
  AOI22_X1 U9905 ( .A1(n9849), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8455), .B2(
        n8483), .ZN(n8456) );
  OAI211_X1 U9906 ( .C1(n8458), .C2(n9851), .A(n8457), .B(n8456), .ZN(n8459)
         );
  AOI21_X1 U9907 ( .B1(n8598), .B2(n8553), .A(n8459), .ZN(n8460) );
  OAI21_X1 U9908 ( .B1(n8602), .B2(n8506), .A(n8460), .ZN(P2_U3274) );
  XNOR2_X1 U9909 ( .A(n8462), .B(n8461), .ZN(n8607) );
  INV_X1 U9910 ( .A(n8486), .ZN(n8465) );
  INV_X1 U9911 ( .A(n8463), .ZN(n8464) );
  AOI211_X1 U9912 ( .C1(n8604), .C2(n8465), .A(n9942), .B(n8464), .ZN(n8603)
         );
  AOI22_X1 U9913 ( .A1(n9849), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8466), .B2(
        n8483), .ZN(n8467) );
  OAI21_X1 U9914 ( .B1(n8468), .B2(n9851), .A(n8467), .ZN(n8476) );
  OAI21_X1 U9915 ( .B1(n4489), .B2(n8470), .A(n8469), .ZN(n8472) );
  AOI21_X1 U9916 ( .B1(n8472), .B2(n8471), .A(n8527), .ZN(n8474) );
  NOR2_X1 U9917 ( .A1(n8474), .A2(n8473), .ZN(n8606) );
  NOR2_X1 U9918 ( .A1(n8606), .A2(n9849), .ZN(n8475) );
  AOI211_X1 U9919 ( .C1(n8603), .C2(n8556), .A(n8476), .B(n8475), .ZN(n8477)
         );
  OAI21_X1 U9920 ( .B1(n8607), .B2(n8506), .A(n8477), .ZN(P2_U3275) );
  INV_X1 U9921 ( .A(n8478), .ZN(n8484) );
  AOI211_X1 U9922 ( .C1(n8480), .C2(n8479), .A(n8527), .B(n4489), .ZN(n8482)
         );
  OR2_X1 U9923 ( .A1(n8482), .A2(n8481), .ZN(n8608) );
  AOI21_X1 U9924 ( .B1(n8484), .B2(n8483), .A(n8608), .ZN(n8492) );
  XNOR2_X1 U9925 ( .A(n8485), .B(n4786), .ZN(n8610) );
  NAND2_X1 U9926 ( .A1(n8610), .A2(n9853), .ZN(n8491) );
  AOI211_X1 U9927 ( .C1(n8487), .C2(n8500), .A(n9942), .B(n8486), .ZN(n8609)
         );
  INV_X1 U9928 ( .A(n8487), .ZN(n8664) );
  OAI22_X1 U9929 ( .A1(n8664), .A2(n9851), .B1(n8488), .B2(n8553), .ZN(n8489)
         );
  AOI21_X1 U9930 ( .B1(n8609), .B2(n8556), .A(n8489), .ZN(n8490) );
  OAI211_X1 U9931 ( .C1(n9855), .C2(n8492), .A(n8491), .B(n8490), .ZN(P2_U3276) );
  XNOR2_X1 U9932 ( .A(n8493), .B(n8496), .ZN(n8617) );
  OAI22_X1 U9933 ( .A1(n8553), .A2(n8495), .B1(n8494), .B2(n9845), .ZN(n8504)
         );
  XNOR2_X1 U9934 ( .A(n8497), .B(n8496), .ZN(n8499) );
  AOI21_X1 U9935 ( .B1(n8499), .B2(n9838), .A(n8498), .ZN(n8616) );
  INV_X1 U9936 ( .A(n8500), .ZN(n8501) );
  AOI211_X1 U9937 ( .C1(n8614), .C2(n8513), .A(n9942), .B(n8501), .ZN(n8613)
         );
  NAND2_X1 U9938 ( .A1(n8613), .A2(n8530), .ZN(n8502) );
  AOI21_X1 U9939 ( .B1(n8616), .B2(n8502), .A(n9849), .ZN(n8503) );
  AOI211_X1 U9940 ( .C1(n8534), .C2(n8614), .A(n8504), .B(n8503), .ZN(n8505)
         );
  OAI21_X1 U9941 ( .B1(n8617), .B2(n8506), .A(n8505), .ZN(P2_U3277) );
  XNOR2_X1 U9942 ( .A(n8507), .B(n8511), .ZN(n8508) );
  NAND2_X1 U9943 ( .A1(n8508), .A2(n9838), .ZN(n8510) );
  NAND2_X1 U9944 ( .A1(n8510), .A2(n8509), .ZN(n8618) );
  INV_X1 U9945 ( .A(n8618), .ZN(n8521) );
  XNOR2_X1 U9946 ( .A(n8512), .B(n8511), .ZN(n8620) );
  NAND2_X1 U9947 ( .A1(n8620), .A2(n9853), .ZN(n8520) );
  AOI211_X1 U9948 ( .C1(n8514), .C2(n8523), .A(n9942), .B(n4699), .ZN(n8619)
         );
  NOR2_X1 U9949 ( .A1(n8669), .A2(n9851), .ZN(n8518) );
  OAI22_X1 U9950 ( .A1(n8553), .A2(n8516), .B1(n8515), .B2(n9845), .ZN(n8517)
         );
  AOI211_X1 U9951 ( .C1(n8619), .C2(n8556), .A(n8518), .B(n8517), .ZN(n8519)
         );
  OAI211_X1 U9952 ( .C1(n9849), .C2(n8521), .A(n8520), .B(n8519), .ZN(P2_U3278) );
  OR2_X1 U9953 ( .A1(n8549), .A2(n8673), .ZN(n8522) );
  AND3_X1 U9954 ( .A1(n8523), .A2(n8522), .A3(n9841), .ZN(n8624) );
  NOR2_X1 U9955 ( .A1(n9845), .A2(n8524), .ZN(n8529) );
  XNOR2_X1 U9956 ( .A(n8525), .B(n8532), .ZN(n8528) );
  OAI21_X1 U9957 ( .B1(n8528), .B2(n8527), .A(n8526), .ZN(n8623) );
  AOI211_X1 U9958 ( .C1(n8624), .C2(n8530), .A(n8529), .B(n8623), .ZN(n8538)
         );
  OAI21_X1 U9959 ( .B1(n8533), .B2(n8532), .A(n8531), .ZN(n8625) );
  NAND2_X1 U9960 ( .A1(n8625), .A2(n9853), .ZN(n8537) );
  AOI22_X1 U9961 ( .A1(n8535), .A2(n8534), .B1(P2_REG2_REG_17__SCAN_IN), .B2(
        n9849), .ZN(n8536) );
  OAI211_X1 U9962 ( .C1(n9855), .C2(n8538), .A(n8537), .B(n8536), .ZN(P2_U3279) );
  AND2_X1 U9963 ( .A1(n8539), .A2(n8542), .ZN(n8540) );
  XNOR2_X1 U9964 ( .A(n8543), .B(n8542), .ZN(n8545) );
  AOI21_X1 U9965 ( .B1(n8545), .B2(n9838), .A(n8544), .ZN(n8546) );
  OAI21_X1 U9966 ( .B1(n8628), .B2(n8547), .A(n8546), .ZN(n8629) );
  NAND2_X1 U9967 ( .A1(n8629), .A2(n8553), .ZN(n8558) );
  AOI211_X1 U9968 ( .C1(n8550), .C2(n4705), .A(n9942), .B(n8549), .ZN(n8630)
         );
  NOR2_X1 U9969 ( .A1(n8678), .A2(n9851), .ZN(n8555) );
  OAI22_X1 U9970 ( .A1(n8553), .A2(n8552), .B1(n8551), .B2(n9845), .ZN(n8554)
         );
  AOI211_X1 U9971 ( .C1(n8630), .C2(n8556), .A(n8555), .B(n8554), .ZN(n8557)
         );
  OAI211_X1 U9972 ( .C1(n8628), .C2(n8559), .A(n8558), .B(n8557), .ZN(P2_U3280) );
  INV_X1 U9973 ( .A(n8560), .ZN(n8638) );
  INV_X1 U9974 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8565) );
  AND2_X1 U9975 ( .A1(n8564), .A2(n8563), .ZN(n8639) );
  MUX2_X1 U9976 ( .A(n8565), .B(n8639), .S(n9960), .Z(n8566) );
  OAI21_X1 U9977 ( .B1(n8642), .B2(n8634), .A(n8566), .ZN(P2_U3550) );
  AOI211_X1 U9978 ( .C1(n9918), .C2(n8569), .A(n8568), .B(n8567), .ZN(n8570)
         );
  OAI21_X1 U9979 ( .B1(n8571), .B2(n9898), .A(n8570), .ZN(n8643) );
  MUX2_X1 U9980 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8643), .S(n9960), .Z(
        P2_U3548) );
  INV_X1 U9981 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8575) );
  AOI211_X1 U9982 ( .C1(n8574), .C2(n9946), .A(n8573), .B(n8572), .ZN(n8644)
         );
  MUX2_X1 U9983 ( .A(n8575), .B(n8644), .S(n9960), .Z(n8576) );
  OAI21_X1 U9984 ( .B1(n4707), .B2(n8634), .A(n8576), .ZN(P2_U3547) );
  INV_X1 U9985 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8581) );
  AOI211_X1 U9986 ( .C1(n8580), .C2(n9946), .A(n8579), .B(n8578), .ZN(n8647)
         );
  MUX2_X1 U9987 ( .A(n8581), .B(n8647), .S(n9960), .Z(n8582) );
  OAI21_X1 U9988 ( .B1(n6456), .B2(n8634), .A(n8582), .ZN(P2_U3546) );
  INV_X1 U9989 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8586) );
  AOI211_X1 U9990 ( .C1(n8585), .C2(n9946), .A(n8584), .B(n8583), .ZN(n8650)
         );
  MUX2_X1 U9991 ( .A(n8586), .B(n8650), .S(n9960), .Z(n8587) );
  OAI21_X1 U9992 ( .B1(n8653), .B2(n8634), .A(n8587), .ZN(P2_U3545) );
  AOI211_X1 U9993 ( .C1(n9918), .C2(n8590), .A(n8589), .B(n8588), .ZN(n8591)
         );
  OAI21_X1 U9994 ( .B1(n8592), .B2(n9898), .A(n8591), .ZN(n8654) );
  MUX2_X1 U9995 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8654), .S(n9960), .Z(
        P2_U3544) );
  OAI211_X1 U9996 ( .C1(n8595), .C2(n9898), .A(n8594), .B(n8593), .ZN(n8655)
         );
  MUX2_X1 U9997 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8655), .S(n9960), .Z(n8596)
         );
  INV_X1 U9998 ( .A(n8596), .ZN(n8597) );
  OAI21_X1 U9999 ( .B1(n8658), .B2(n8634), .A(n8597), .ZN(P2_U3543) );
  AOI211_X1 U10000 ( .C1(n9918), .C2(n8600), .A(n8599), .B(n8598), .ZN(n8601)
         );
  OAI21_X1 U10001 ( .B1(n8602), .B2(n9898), .A(n8601), .ZN(n8659) );
  MUX2_X1 U10002 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8659), .S(n9960), .Z(
        P2_U3542) );
  AOI21_X1 U10003 ( .B1(n9918), .B2(n8604), .A(n8603), .ZN(n8605) );
  OAI211_X1 U10004 ( .C1(n8607), .C2(n9898), .A(n8606), .B(n8605), .ZN(n8660)
         );
  MUX2_X1 U10005 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8660), .S(n9960), .Z(
        P2_U3541) );
  INV_X1 U10006 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8611) );
  AOI211_X1 U10007 ( .C1(n8610), .C2(n9946), .A(n8609), .B(n8608), .ZN(n8661)
         );
  MUX2_X1 U10008 ( .A(n8611), .B(n8661), .S(n9960), .Z(n8612) );
  OAI21_X1 U10009 ( .B1(n8664), .B2(n8634), .A(n8612), .ZN(P2_U3540) );
  AOI21_X1 U10010 ( .B1(n9918), .B2(n8614), .A(n8613), .ZN(n8615) );
  OAI211_X1 U10011 ( .C1(n8617), .C2(n9898), .A(n8616), .B(n8615), .ZN(n8665)
         );
  MUX2_X1 U10012 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8665), .S(n9960), .Z(
        P2_U3539) );
  AOI211_X1 U10013 ( .C1(n8620), .C2(n9946), .A(n8619), .B(n8618), .ZN(n8666)
         );
  MUX2_X1 U10014 ( .A(n8621), .B(n8666), .S(n9960), .Z(n8622) );
  OAI21_X1 U10015 ( .B1(n8669), .B2(n8634), .A(n8622), .ZN(P2_U3538) );
  INV_X1 U10016 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8626) );
  AOI211_X1 U10017 ( .C1(n8625), .C2(n9946), .A(n8624), .B(n8623), .ZN(n8670)
         );
  MUX2_X1 U10018 ( .A(n8626), .B(n8670), .S(n9960), .Z(n8627) );
  OAI21_X1 U10019 ( .B1(n8673), .B2(n8634), .A(n8627), .ZN(P2_U3537) );
  INV_X1 U10020 ( .A(n8628), .ZN(n8631) );
  INV_X1 U10021 ( .A(n9921), .ZN(n9935) );
  AOI211_X1 U10022 ( .C1(n8631), .C2(n9935), .A(n8630), .B(n8629), .ZN(n8674)
         );
  MUX2_X1 U10023 ( .A(n8632), .B(n8674), .S(n9960), .Z(n8633) );
  OAI21_X1 U10024 ( .B1(n8678), .B2(n8634), .A(n8633), .ZN(P2_U3536) );
  INV_X1 U10025 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8636) );
  MUX2_X1 U10026 ( .A(n8636), .B(n8635), .S(n9949), .Z(n8637) );
  OAI21_X1 U10027 ( .B1(n8638), .B2(n8677), .A(n8637), .ZN(P2_U3519) );
  MUX2_X1 U10028 ( .A(n8640), .B(n8639), .S(n9949), .Z(n8641) );
  OAI21_X1 U10029 ( .B1(n8642), .B2(n8677), .A(n8641), .ZN(P2_U3518) );
  MUX2_X1 U10030 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8643), .S(n9949), .Z(
        P2_U3516) );
  MUX2_X1 U10031 ( .A(n8645), .B(n8644), .S(n9949), .Z(n8646) );
  OAI21_X1 U10032 ( .B1(n4707), .B2(n8677), .A(n8646), .ZN(P2_U3515) );
  MUX2_X1 U10033 ( .A(n8648), .B(n8647), .S(n9949), .Z(n8649) );
  OAI21_X1 U10034 ( .B1(n6456), .B2(n8677), .A(n8649), .ZN(P2_U3514) );
  MUX2_X1 U10035 ( .A(n8651), .B(n8650), .S(n9949), .Z(n8652) );
  OAI21_X1 U10036 ( .B1(n8653), .B2(n8677), .A(n8652), .ZN(P2_U3513) );
  MUX2_X1 U10037 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8654), .S(n9949), .Z(
        P2_U3512) );
  MUX2_X1 U10038 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8655), .S(n9949), .Z(n8656) );
  INV_X1 U10039 ( .A(n8656), .ZN(n8657) );
  OAI21_X1 U10040 ( .B1(n8658), .B2(n8677), .A(n8657), .ZN(P2_U3511) );
  MUX2_X1 U10041 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8659), .S(n9949), .Z(
        P2_U3510) );
  MUX2_X1 U10042 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8660), .S(n9949), .Z(
        P2_U3509) );
  MUX2_X1 U10043 ( .A(n8662), .B(n8661), .S(n9949), .Z(n8663) );
  OAI21_X1 U10044 ( .B1(n8664), .B2(n8677), .A(n8663), .ZN(P2_U3508) );
  MUX2_X1 U10045 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8665), .S(n9949), .Z(
        P2_U3507) );
  INV_X1 U10046 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8667) );
  MUX2_X1 U10047 ( .A(n8667), .B(n8666), .S(n9949), .Z(n8668) );
  OAI21_X1 U10048 ( .B1(n8669), .B2(n8677), .A(n8668), .ZN(P2_U3505) );
  MUX2_X1 U10049 ( .A(n8671), .B(n8670), .S(n9949), .Z(n8672) );
  OAI21_X1 U10050 ( .B1(n8673), .B2(n8677), .A(n8672), .ZN(P2_U3502) );
  INV_X1 U10051 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8675) );
  MUX2_X1 U10052 ( .A(n8675), .B(n8674), .S(n9949), .Z(n8676) );
  OAI21_X1 U10053 ( .B1(n8678), .B2(n8677), .A(n8676), .ZN(P2_U3499) );
  INV_X1 U10054 ( .A(n8833), .ZN(n9514) );
  INV_X1 U10055 ( .A(n8679), .ZN(n8681) );
  NOR4_X1 U10056 ( .A1(n8681), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8680), .A4(
        P2_U3152), .ZN(n8682) );
  AOI21_X1 U10057 ( .B1(n8683), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8682), .ZN(
        n8684) );
  OAI21_X1 U10058 ( .B1(n9514), .B2(n8696), .A(n8684), .ZN(P2_U3327) );
  OAI222_X1 U10059 ( .A1(n5046), .A2(P2_U3152), .B1(n8696), .B2(n8686), .C1(
        n8685), .C2(n8694), .ZN(P2_U3328) );
  OAI222_X1 U10060 ( .A1(P2_U3152), .A2(n8689), .B1(n8696), .B2(n8688), .C1(
        n8687), .C2(n8694), .ZN(P2_U3329) );
  NAND2_X1 U10061 ( .A1(n9515), .A2(n8690), .ZN(n8692) );
  OAI211_X1 U10062 ( .C1(n8694), .C2(n8693), .A(n8692), .B(n8691), .ZN(
        P2_U3330) );
  INV_X1 U10063 ( .A(n9519), .ZN(n8695) );
  OAI222_X1 U10064 ( .A1(n8694), .A2(n8697), .B1(n8696), .B2(n8695), .C1(n6496), .C2(P2_U3152), .ZN(P2_U3331) );
  MUX2_X1 U10065 ( .A(n8698), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10066 ( .A1(n8700), .A2(n8699), .ZN(n8702) );
  XNOR2_X1 U10067 ( .A(n8702), .B(n8701), .ZN(n8703) );
  NAND2_X1 U10068 ( .A1(n8703), .A2(n8808), .ZN(n8709) );
  OAI22_X1 U10069 ( .A1(n8824), .A2(n8705), .B1(n8822), .B2(n8704), .ZN(n8706)
         );
  AOI211_X1 U10070 ( .C1(n4473), .C2(n9132), .A(n8707), .B(n8706), .ZN(n8708)
         );
  OAI211_X1 U10071 ( .C1(n9614), .C2(n8758), .A(n8709), .B(n8708), .ZN(
        P1_U3213) );
  NAND2_X1 U10072 ( .A1(n4927), .A2(n8711), .ZN(n8713) );
  XNOR2_X1 U10073 ( .A(n8713), .B(n8712), .ZN(n8718) );
  INV_X1 U10074 ( .A(n9303), .ZN(n9187) );
  INV_X1 U10075 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8714) );
  OAI22_X1 U10076 ( .A1(n8824), .A2(n9187), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8714), .ZN(n8716) );
  INV_X1 U10077 ( .A(n9330), .ZN(n9182) );
  OAI22_X1 U10078 ( .A1(n8800), .A2(n9182), .B1(n8822), .B2(n9298), .ZN(n8715)
         );
  AOI211_X1 U10079 ( .C1(n9447), .C2(n8828), .A(n8716), .B(n8715), .ZN(n8717)
         );
  OAI21_X1 U10080 ( .B1(n8718), .B2(n8831), .A(n8717), .ZN(P1_U3214) );
  INV_X1 U10081 ( .A(n9468), .ZN(n9360) );
  OAI21_X1 U10082 ( .B1(n8720), .B2(n4543), .A(n8719), .ZN(n8721) );
  NAND2_X1 U10083 ( .A1(n8721), .A2(n8808), .ZN(n8724) );
  AND2_X1 U10084 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9158) );
  INV_X1 U10085 ( .A(n9401), .ZN(n8864) );
  OAI22_X1 U10086 ( .A1(n8800), .A2(n8864), .B1(n8822), .B2(n9357), .ZN(n8722)
         );
  AOI211_X1 U10087 ( .C1(n8811), .C2(n9367), .A(n9158), .B(n8722), .ZN(n8723)
         );
  OAI211_X1 U10088 ( .C1(n9360), .C2(n8758), .A(n8724), .B(n8723), .ZN(
        P1_U3217) );
  XOR2_X1 U10089 ( .A(n8726), .B(n8725), .Z(n8731) );
  INV_X1 U10090 ( .A(n9367), .ZN(n8865) );
  INV_X1 U10091 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8727) );
  OAI22_X1 U10092 ( .A1(n8800), .A2(n8865), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8727), .ZN(n8729) );
  OAI22_X1 U10093 ( .A1(n8824), .A2(n9182), .B1(n8822), .B2(n9323), .ZN(n8728)
         );
  AOI211_X1 U10094 ( .C1(n9458), .C2(n8828), .A(n8729), .B(n8728), .ZN(n8730)
         );
  OAI21_X1 U10095 ( .B1(n8731), .B2(n8831), .A(n8730), .ZN(P1_U3221) );
  AOI21_X1 U10096 ( .B1(n8734), .B2(n8733), .A(n8732), .ZN(n8735) );
  OR2_X1 U10097 ( .A1(n8735), .A2(n8831), .ZN(n8740) );
  AOI22_X1 U10098 ( .A1(n8811), .A2(n9277), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8739) );
  INV_X1 U10099 ( .A(n8736), .ZN(n9273) );
  AOI22_X1 U10100 ( .A1(n4473), .A2(n9303), .B1(n9273), .B2(n8810), .ZN(n8738)
         );
  NAND2_X1 U10101 ( .A1(n9437), .A2(n8828), .ZN(n8737) );
  NAND4_X1 U10102 ( .A1(n8740), .A2(n8739), .A3(n8738), .A4(n8737), .ZN(
        P1_U3223) );
  INV_X1 U10103 ( .A(n8741), .ZN(n8742) );
  AOI21_X1 U10104 ( .B1(n8744), .B2(n8743), .A(n8742), .ZN(n8750) );
  INV_X1 U10105 ( .A(n9376), .ZN(n8872) );
  OAI22_X1 U10106 ( .A1(n8824), .A2(n8872), .B1(n8822), .B2(n8745), .ZN(n8746)
         );
  AOI211_X1 U10107 ( .C1(n4473), .C2(n9130), .A(n8747), .B(n8746), .ZN(n8749)
         );
  NAND2_X1 U10108 ( .A1(n9173), .A2(n8828), .ZN(n8748) );
  OAI211_X1 U10109 ( .C1(n8750), .C2(n8831), .A(n8749), .B(n8748), .ZN(
        P1_U3224) );
  INV_X1 U10110 ( .A(n9480), .ZN(n9397) );
  XNOR2_X1 U10111 ( .A(n8752), .B(n8751), .ZN(n8753) );
  NAND2_X1 U10112 ( .A1(n8753), .A2(n8808), .ZN(n8757) );
  OAI22_X1 U10113 ( .A1(n8824), .A2(n8864), .B1(n8822), .B2(n9393), .ZN(n8754)
         );
  AOI211_X1 U10114 ( .C1(n4473), .C2(n9402), .A(n8755), .B(n8754), .ZN(n8756)
         );
  OAI211_X1 U10115 ( .C1(n9397), .C2(n8758), .A(n8757), .B(n8756), .ZN(
        P1_U3226) );
  AOI21_X1 U10116 ( .B1(n8760), .B2(n8759), .A(n4515), .ZN(n8765) );
  INV_X1 U10117 ( .A(n9286), .ZN(n8911) );
  OAI22_X1 U10118 ( .A1(n8824), .A2(n8911), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8761), .ZN(n8763) );
  INV_X1 U10119 ( .A(n9316), .ZN(n9183) );
  OAI22_X1 U10120 ( .A1(n8800), .A2(n9183), .B1(n8822), .B2(n9289), .ZN(n8762)
         );
  AOI211_X1 U10121 ( .C1(n9442), .C2(n8828), .A(n8763), .B(n8762), .ZN(n8764)
         );
  OAI21_X1 U10122 ( .B1(n8765), .B2(n8831), .A(n8764), .ZN(P1_U3227) );
  NAND2_X1 U10123 ( .A1(n8767), .A2(n8766), .ZN(n8768) );
  XNOR2_X1 U10124 ( .A(n8769), .B(n8768), .ZN(n8774) );
  INV_X1 U10125 ( .A(n9349), .ZN(n8861) );
  OAI22_X1 U10126 ( .A1(n8824), .A2(n8861), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8770), .ZN(n8772) );
  INV_X1 U10127 ( .A(n9375), .ZN(n8866) );
  OAI22_X1 U10128 ( .A1(n8800), .A2(n8866), .B1(n8822), .B2(n9342), .ZN(n8771)
         );
  AOI211_X1 U10129 ( .C1(n9464), .C2(n8828), .A(n8772), .B(n8771), .ZN(n8773)
         );
  OAI21_X1 U10130 ( .B1(n8774), .B2(n8831), .A(n8773), .ZN(P1_U3231) );
  INV_X1 U10131 ( .A(n8778), .ZN(n8781) );
  AOI21_X1 U10132 ( .B1(n8778), .B2(n8776), .A(n8777), .ZN(n8779) );
  NOR2_X1 U10133 ( .A1(n8779), .A2(n8831), .ZN(n8780) );
  OAI21_X1 U10134 ( .B1(n8781), .B2(n8775), .A(n8780), .ZN(n8787) );
  NOR2_X1 U10135 ( .A1(n8782), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8783) );
  AOI21_X1 U10136 ( .B1(n8811), .B2(n9316), .A(n8783), .ZN(n8786) );
  AOI22_X1 U10137 ( .A1(n4473), .A2(n9349), .B1(n9310), .B2(n8810), .ZN(n8785)
         );
  NAND2_X1 U10138 ( .A1(n9451), .A2(n8828), .ZN(n8784) );
  NAND4_X1 U10139 ( .A1(n8787), .A2(n8786), .A3(n8785), .A4(n8784), .ZN(
        P1_U3233) );
  OAI21_X1 U10140 ( .B1(n8790), .B2(n8788), .A(n8789), .ZN(n8791) );
  NAND2_X1 U10141 ( .A1(n8791), .A2(n8808), .ZN(n8796) );
  AOI22_X1 U10142 ( .A1(n8793), .A2(n8828), .B1(n8792), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n8795) );
  NAND3_X1 U10143 ( .A1(n8796), .A2(n8795), .A3(n8794), .ZN(P1_U3235) );
  NAND2_X1 U10144 ( .A1(n4523), .A2(n8797), .ZN(n8798) );
  XOR2_X1 U10145 ( .A(n8799), .B(n8798), .Z(n8804) );
  NAND2_X1 U10146 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9722) );
  OAI21_X1 U10147 ( .B1(n8824), .B2(n8866), .A(n9722), .ZN(n8802) );
  OAI22_X1 U10148 ( .A1(n8800), .A2(n8872), .B1(n8822), .B2(n9380), .ZN(n8801)
         );
  AOI211_X1 U10149 ( .C1(n9475), .C2(n8828), .A(n8802), .B(n8801), .ZN(n8803)
         );
  OAI21_X1 U10150 ( .B1(n8804), .B2(n8831), .A(n8803), .ZN(P1_U3236) );
  OAI21_X1 U10151 ( .B1(n8732), .B2(n8806), .A(n8805), .ZN(n8807) );
  NAND3_X1 U10152 ( .A1(n4529), .A2(n8808), .A3(n8807), .ZN(n8815) );
  AOI22_X1 U10153 ( .A1(n4473), .A2(n9286), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8814) );
  INV_X1 U10154 ( .A(n8809), .ZN(n9258) );
  AOI22_X1 U10155 ( .A1(n8811), .A2(n9265), .B1(n9258), .B2(n8810), .ZN(n8813)
         );
  NAND2_X1 U10156 ( .A1(n9432), .A2(n8828), .ZN(n8812) );
  NAND4_X1 U10157 ( .A1(n8815), .A2(n8814), .A3(n8813), .A4(n8812), .ZN(
        P1_U3238) );
  NAND2_X1 U10158 ( .A1(n8817), .A2(n8816), .ZN(n8818) );
  XOR2_X1 U10159 ( .A(n8819), .B(n8818), .Z(n8832) );
  INV_X1 U10160 ( .A(n8820), .ZN(n8826) );
  OAI22_X1 U10161 ( .A1(n8824), .A2(n8823), .B1(n8822), .B2(n8821), .ZN(n8825)
         );
  AOI211_X1 U10162 ( .C1(n4473), .C2(n9131), .A(n8826), .B(n8825), .ZN(n8830)
         );
  NAND2_X1 U10163 ( .A1(n9606), .A2(n8828), .ZN(n8829) );
  OAI211_X1 U10164 ( .C1(n8832), .C2(n8831), .A(n8830), .B(n8829), .ZN(
        P1_U3239) );
  NAND2_X1 U10165 ( .A1(n8833), .A2(n8850), .ZN(n8835) );
  NAND2_X1 U10166 ( .A1(n5845), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8834) );
  INV_X1 U10167 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8839) );
  NAND2_X1 U10168 ( .A1(n5921), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8838) );
  INV_X1 U10169 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8836) );
  OR2_X1 U10170 ( .A1(n5852), .A2(n8836), .ZN(n8837) );
  OAI211_X1 U10171 ( .C1(n8840), .C2(n8839), .A(n8838), .B(n8837), .ZN(n9164)
         );
  INV_X1 U10172 ( .A(n9164), .ZN(n8916) );
  NAND2_X1 U10173 ( .A1(n8841), .A2(n8850), .ZN(n8843) );
  NAND2_X1 U10174 ( .A1(n4474), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8842) );
  INV_X1 U10175 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8847) );
  NAND2_X1 U10176 ( .A1(n5921), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8846) );
  INV_X1 U10177 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8844) );
  OR2_X1 U10178 ( .A1(n5852), .A2(n8844), .ZN(n8845) );
  OAI211_X1 U10179 ( .C1(n8840), .C2(n8847), .A(n8846), .B(n8845), .ZN(n9215)
         );
  INV_X1 U10180 ( .A(n9215), .ZN(n8849) );
  NAND2_X1 U10181 ( .A1(n9167), .A2(n8849), .ZN(n8848) );
  OR2_X1 U10182 ( .A1(n9167), .A2(n8849), .ZN(n9045) );
  NAND2_X1 U10183 ( .A1(n8851), .A2(n8850), .ZN(n8853) );
  NAND2_X1 U10184 ( .A1(n5845), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8852) );
  INV_X1 U10185 ( .A(n9234), .ZN(n9034) );
  OR2_X1 U10186 ( .A1(n9223), .A2(n9034), .ZN(n8854) );
  INV_X1 U10187 ( .A(n9250), .ZN(n8855) );
  AND2_X1 U10188 ( .A1(n8854), .A2(n9209), .ZN(n8860) );
  NAND2_X1 U10189 ( .A1(n9422), .A2(n8855), .ZN(n9026) );
  INV_X1 U10190 ( .A(n9265), .ZN(n8856) );
  NAND2_X1 U10191 ( .A1(n9426), .A2(n8856), .ZN(n9023) );
  INV_X1 U10192 ( .A(n9277), .ZN(n9014) );
  NAND2_X1 U10193 ( .A1(n9432), .A2(n9014), .ZN(n9207) );
  NAND2_X1 U10194 ( .A1(n9208), .A2(n4638), .ZN(n8857) );
  NAND3_X1 U10195 ( .A1(n9026), .A2(n9023), .A3(n8857), .ZN(n8859) );
  AND2_X1 U10196 ( .A1(n9223), .A2(n9034), .ZN(n8858) );
  AOI21_X1 U10197 ( .B1(n8860), .B2(n8859), .A(n8858), .ZN(n9110) );
  INV_X1 U10198 ( .A(n8860), .ZN(n9108) );
  OR2_X1 U10199 ( .A1(n9442), .A2(n9187), .ZN(n9046) );
  OR2_X1 U10200 ( .A1(n9447), .A2(n9183), .ZN(n9203) );
  NAND2_X1 U10201 ( .A1(n9046), .A2(n9203), .ZN(n9007) );
  NAND2_X1 U10202 ( .A1(n9451), .A2(n9182), .ZN(n9202) );
  NAND2_X1 U10203 ( .A1(n9048), .A2(n9199), .ZN(n8862) );
  NAND2_X1 U10204 ( .A1(n9458), .A2(n8861), .ZN(n9201) );
  AND2_X1 U10205 ( .A1(n8862), .A2(n9201), .ZN(n8863) );
  AND2_X1 U10206 ( .A1(n9202), .A2(n8863), .ZN(n9001) );
  OR2_X1 U10207 ( .A1(n9475), .A2(n8864), .ZN(n9050) );
  OR2_X1 U10208 ( .A1(n9480), .A2(n8872), .ZN(n9372) );
  AND2_X1 U10209 ( .A1(n9050), .A2(n9372), .ZN(n9196) );
  NAND2_X1 U10210 ( .A1(n9468), .A2(n8866), .ZN(n9198) );
  NAND2_X1 U10211 ( .A1(n9475), .A2(n8864), .ZN(n9363) );
  AND2_X1 U10212 ( .A1(n9198), .A2(n9363), .ZN(n8995) );
  INV_X1 U10213 ( .A(n8995), .ZN(n8868) );
  NOR2_X1 U10214 ( .A1(n9464), .A2(n8865), .ZN(n9325) );
  OR2_X1 U10215 ( .A1(n9468), .A2(n8866), .ZN(n9049) );
  INV_X1 U10216 ( .A(n9049), .ZN(n8867) );
  NOR2_X1 U10217 ( .A1(n9325), .A2(n8867), .ZN(n8997) );
  OAI211_X1 U10218 ( .C1(n9196), .C2(n8868), .A(n8997), .B(n9048), .ZN(n8869)
         );
  NAND2_X1 U10219 ( .A1(n9001), .A2(n8869), .ZN(n8870) );
  OR2_X1 U10220 ( .A1(n9451), .A2(n9182), .ZN(n9047) );
  NAND2_X1 U10221 ( .A1(n8870), .A2(n9047), .ZN(n8871) );
  NOR2_X1 U10222 ( .A1(n9007), .A2(n8871), .ZN(n9104) );
  AND2_X1 U10223 ( .A1(n9001), .A2(n9198), .ZN(n9101) );
  AND2_X1 U10224 ( .A1(n9480), .A2(n8872), .ZN(n9195) );
  NOR2_X1 U10225 ( .A1(n9195), .A2(n4644), .ZN(n8873) );
  NAND2_X1 U10226 ( .A1(n8873), .A2(n9363), .ZN(n8905) );
  NAND2_X1 U10227 ( .A1(n8875), .A2(n8874), .ZN(n8977) );
  NAND2_X1 U10228 ( .A1(n8977), .A2(n8973), .ZN(n8961) );
  INV_X1 U10229 ( .A(n8961), .ZN(n8879) );
  INV_X1 U10230 ( .A(n8876), .ZN(n8966) );
  AND3_X1 U10231 ( .A1(n8967), .A2(n8966), .A3(n8877), .ZN(n8878) );
  NAND3_X1 U10232 ( .A1(n8986), .A2(n8879), .A3(n8878), .ZN(n8901) );
  NAND2_X1 U10233 ( .A1(n8954), .A2(n8940), .ZN(n8880) );
  OR3_X1 U10234 ( .A1(n8905), .A2(n8901), .A3(n8880), .ZN(n9099) );
  INV_X1 U10235 ( .A(n8881), .ZN(n8883) );
  NAND3_X1 U10236 ( .A1(n8883), .A2(n4673), .A3(n8882), .ZN(n8884) );
  NAND2_X1 U10237 ( .A1(n8885), .A2(n8884), .ZN(n8887) );
  OAI21_X1 U10238 ( .B1(n8888), .B2(n8887), .A(n8886), .ZN(n8889) );
  NAND2_X1 U10239 ( .A1(n8889), .A2(n9087), .ZN(n8891) );
  NAND3_X1 U10240 ( .A1(n8891), .A2(n9083), .A3(n8890), .ZN(n8893) );
  NAND2_X1 U10241 ( .A1(n8892), .A2(n8941), .ZN(n9084) );
  AOI21_X1 U10242 ( .B1(n8893), .B2(n9088), .A(n9084), .ZN(n8906) );
  NAND2_X1 U10243 ( .A1(n8968), .A2(n8894), .ZN(n8895) );
  NAND2_X1 U10244 ( .A1(n8895), .A2(n8967), .ZN(n8896) );
  NAND2_X1 U10245 ( .A1(n8948), .A2(n8896), .ZN(n8974) );
  INV_X1 U10246 ( .A(n8974), .ZN(n8897) );
  OAI21_X1 U10247 ( .B1(n8961), .B2(n8897), .A(n8980), .ZN(n8898) );
  NAND2_X1 U10248 ( .A1(n8898), .A2(n8986), .ZN(n8903) );
  NOR2_X1 U10249 ( .A1(n8963), .A2(n8899), .ZN(n8900) );
  OR2_X1 U10250 ( .A1(n8901), .A2(n8900), .ZN(n8902) );
  AND4_X1 U10251 ( .A1(n8931), .A2(n8987), .A3(n8903), .A4(n8902), .ZN(n8904)
         );
  OR2_X1 U10252 ( .A1(n8905), .A2(n8904), .ZN(n9097) );
  OAI21_X1 U10253 ( .B1(n9099), .B2(n8906), .A(n9097), .ZN(n8907) );
  NAND2_X1 U10254 ( .A1(n9101), .A2(n8907), .ZN(n8910) );
  NAND2_X1 U10255 ( .A1(n9442), .A2(n9187), .ZN(n9204) );
  NAND2_X1 U10256 ( .A1(n9447), .A2(n9183), .ZN(n8908) );
  NAND2_X1 U10257 ( .A1(n9204), .A2(n8908), .ZN(n9006) );
  NAND2_X1 U10258 ( .A1(n9006), .A2(n9046), .ZN(n8909) );
  NAND2_X1 U10259 ( .A1(n9205), .A2(n8909), .ZN(n9102) );
  AOI21_X1 U10260 ( .B1(n9104), .B2(n8910), .A(n9102), .ZN(n8913) );
  OR2_X1 U10261 ( .A1(n9432), .A2(n9014), .ZN(n8912) );
  AND2_X1 U10262 ( .A1(n8912), .A2(n9261), .ZN(n9206) );
  INV_X1 U10263 ( .A(n9206), .ZN(n9106) );
  OR4_X1 U10264 ( .A1(n9108), .A2(n4560), .A3(n8913), .A4(n9106), .ZN(n8914)
         );
  NAND2_X1 U10265 ( .A1(n9110), .A2(n8914), .ZN(n8915) );
  AND2_X1 U10266 ( .A1(n9045), .A2(n8915), .ZN(n8917) );
  NAND2_X1 U10267 ( .A1(n8919), .A2(n8916), .ZN(n9044) );
  OAI21_X1 U10268 ( .B1(n9081), .B2(n8917), .A(n9044), .ZN(n8918) );
  XNOR2_X1 U10269 ( .A(n8918), .B(n9156), .ZN(n9123) );
  NAND2_X1 U10270 ( .A1(n9045), .A2(n9164), .ZN(n8920) );
  NAND2_X1 U10271 ( .A1(n8920), .A2(n8919), .ZN(n9113) );
  NAND2_X1 U10272 ( .A1(n9164), .A2(n9215), .ZN(n8921) );
  NAND2_X1 U10273 ( .A1(n9167), .A2(n8921), .ZN(n9111) );
  NAND2_X1 U10274 ( .A1(n9432), .A2(n9261), .ZN(n8922) );
  NAND2_X1 U10275 ( .A1(n9023), .A2(n8922), .ZN(n8925) );
  NAND2_X1 U10276 ( .A1(n9205), .A2(n9277), .ZN(n8923) );
  NAND2_X1 U10277 ( .A1(n9208), .A2(n8923), .ZN(n8924) );
  MUX2_X1 U10278 ( .A(n8925), .B(n8924), .S(n9030), .Z(n9012) );
  NAND2_X1 U10279 ( .A1(n9007), .A2(n9204), .ZN(n8926) );
  NAND2_X1 U10280 ( .A1(n9261), .A2(n8926), .ZN(n8927) );
  MUX2_X1 U10281 ( .A(n9102), .B(n8927), .S(n9030), .Z(n8928) );
  INV_X1 U10282 ( .A(n8928), .ZN(n9010) );
  INV_X1 U10283 ( .A(n9195), .ZN(n8930) );
  AND2_X1 U10284 ( .A1(n9363), .A2(n8930), .ZN(n8929) );
  INV_X1 U10285 ( .A(n9030), .ZN(n9032) );
  MUX2_X1 U10286 ( .A(n9196), .B(n8929), .S(n9032), .Z(n8994) );
  MUX2_X1 U10287 ( .A(n8931), .B(n9193), .S(n9030), .Z(n8992) );
  AOI21_X1 U10288 ( .B1(n8933), .B2(n9032), .A(n8932), .ZN(n8939) );
  INV_X1 U10289 ( .A(n8939), .ZN(n8935) );
  AND2_X1 U10290 ( .A1(n8941), .A2(n9057), .ZN(n9093) );
  INV_X1 U10291 ( .A(n8940), .ZN(n8934) );
  AOI21_X1 U10292 ( .B1(n8935), .B2(n9093), .A(n8934), .ZN(n8946) );
  AOI21_X1 U10293 ( .B1(n8937), .B2(n4526), .A(n8936), .ZN(n8938) );
  NAND2_X1 U10294 ( .A1(n8939), .A2(n8938), .ZN(n8944) );
  AND2_X1 U10295 ( .A1(n8940), .A2(n9090), .ZN(n8943) );
  INV_X1 U10296 ( .A(n8941), .ZN(n8942) );
  AOI21_X1 U10297 ( .B1(n8944), .B2(n8943), .A(n8942), .ZN(n8945) );
  MUX2_X1 U10298 ( .A(n8946), .B(n8945), .S(n9030), .Z(n8958) );
  NAND2_X1 U10299 ( .A1(n9570), .A2(n8957), .ZN(n8947) );
  AOI21_X1 U10300 ( .B1(n8958), .B2(n8954), .A(n8947), .ZN(n8953) );
  NAND2_X1 U10301 ( .A1(n8980), .A2(n8948), .ZN(n8965) );
  NAND4_X1 U10302 ( .A1(n8968), .A2(n9032), .A3(n8949), .A4(n9051), .ZN(n8950)
         );
  NOR2_X1 U10303 ( .A1(n8965), .A2(n8950), .ZN(n8951) );
  OAI21_X1 U10304 ( .B1(n8953), .B2(n8952), .A(n8951), .ZN(n8984) );
  NAND2_X1 U10305 ( .A1(n8955), .A2(n8954), .ZN(n8956) );
  AOI21_X1 U10306 ( .B1(n8958), .B2(n8957), .A(n8956), .ZN(n8964) );
  NAND4_X1 U10307 ( .A1(n8967), .A2(n8959), .A3(n9030), .A4(n9051), .ZN(n8960)
         );
  NOR2_X1 U10308 ( .A1(n8961), .A2(n8960), .ZN(n8962) );
  OAI21_X1 U10309 ( .B1(n8964), .B2(n8963), .A(n8962), .ZN(n8983) );
  INV_X1 U10310 ( .A(n8965), .ZN(n8972) );
  NAND2_X1 U10311 ( .A1(n8967), .A2(n8966), .ZN(n8969) );
  NAND2_X1 U10312 ( .A1(n8969), .A2(n8968), .ZN(n8970) );
  AOI21_X1 U10313 ( .B1(n8973), .B2(n8970), .A(n9030), .ZN(n8971) );
  NAND2_X1 U10314 ( .A1(n8972), .A2(n8971), .ZN(n8979) );
  NAND3_X1 U10315 ( .A1(n8974), .A2(n8973), .A3(n9030), .ZN(n8975) );
  NAND2_X1 U10316 ( .A1(n8975), .A2(n8977), .ZN(n8976) );
  OAI21_X1 U10317 ( .B1(n9032), .B2(n8977), .A(n8976), .ZN(n8978) );
  OAI211_X1 U10318 ( .C1(n9032), .C2(n8980), .A(n8979), .B(n8978), .ZN(n8981)
         );
  INV_X1 U10319 ( .A(n8981), .ZN(n8982) );
  NAND3_X1 U10320 ( .A1(n8984), .A2(n8983), .A3(n8982), .ZN(n8985) );
  NAND2_X1 U10321 ( .A1(n8985), .A2(n9073), .ZN(n8990) );
  MUX2_X1 U10322 ( .A(n8987), .B(n8986), .S(n9032), .Z(n8988) );
  NAND3_X1 U10323 ( .A1(n8990), .A2(n8989), .A3(n8988), .ZN(n8991) );
  NAND3_X1 U10324 ( .A1(n9398), .A2(n8992), .A3(n8991), .ZN(n8993) );
  NAND2_X1 U10325 ( .A1(n8994), .A2(n8993), .ZN(n8996) );
  INV_X1 U10326 ( .A(n9325), .ZN(n8998) );
  NAND2_X1 U10327 ( .A1(n8999), .A2(n9201), .ZN(n9000) );
  INV_X1 U10328 ( .A(n9048), .ZN(n9002) );
  OAI21_X1 U10329 ( .B1(n9003), .B2(n9002), .A(n9001), .ZN(n9004) );
  NAND2_X1 U10330 ( .A1(n9004), .A2(n9047), .ZN(n9005) );
  NOR2_X1 U10331 ( .A1(n9007), .A2(n9006), .ZN(n9008) );
  NAND2_X1 U10332 ( .A1(n9012), .A2(n9011), .ZN(n9022) );
  INV_X1 U10333 ( .A(n9189), .ZN(n9020) );
  NOR2_X1 U10334 ( .A1(n9205), .A2(n9277), .ZN(n9013) );
  NOR2_X1 U10335 ( .A1(n9013), .A2(n9432), .ZN(n9017) );
  NAND2_X1 U10336 ( .A1(n9261), .A2(n9014), .ZN(n9015) );
  NAND2_X1 U10337 ( .A1(n9207), .A2(n9015), .ZN(n9016) );
  MUX2_X1 U10338 ( .A(n9017), .B(n9016), .S(n9032), .Z(n9018) );
  OAI21_X1 U10339 ( .B1(n9020), .B2(n9019), .A(n9018), .ZN(n9021) );
  NAND2_X1 U10340 ( .A1(n9022), .A2(n9021), .ZN(n9025) );
  MUX2_X1 U10341 ( .A(n9023), .B(n9208), .S(n9032), .Z(n9024) );
  NAND3_X1 U10342 ( .A1(n9025), .A2(n9233), .A3(n9024), .ZN(n9028) );
  MUX2_X1 U10343 ( .A(n9026), .B(n9209), .S(n9030), .Z(n9027) );
  AND2_X1 U10344 ( .A1(n9028), .A2(n9027), .ZN(n9033) );
  NAND3_X1 U10345 ( .A1(n9113), .A2(n9033), .A3(n9223), .ZN(n9029) );
  AND2_X1 U10346 ( .A1(n9234), .A2(n9030), .ZN(n9031) );
  AOI21_X1 U10347 ( .B1(n9223), .B2(n9032), .A(n9031), .ZN(n9037) );
  INV_X1 U10348 ( .A(n9033), .ZN(n9035) );
  INV_X1 U10349 ( .A(n9223), .ZN(n9415) );
  NAND3_X1 U10350 ( .A1(n9035), .A2(n9415), .A3(n9034), .ZN(n9036) );
  NAND4_X1 U10351 ( .A1(n9113), .A2(n9037), .A3(n9111), .A4(n9036), .ZN(n9038)
         );
  NAND2_X1 U10352 ( .A1(n9039), .A2(n4673), .ZN(n9041) );
  OR3_X1 U10353 ( .A1(n9043), .A2(n9040), .A3(n9041), .ZN(n9121) );
  INV_X1 U10354 ( .A(n9041), .ZN(n9115) );
  NAND3_X1 U10355 ( .A1(n9043), .A2(n9115), .A3(n9042), .ZN(n9120) );
  XNOR2_X1 U10356 ( .A(n9223), .B(n9234), .ZN(n9211) );
  NAND2_X1 U10357 ( .A1(n9048), .A2(n9201), .ZN(n9334) );
  INV_X1 U10358 ( .A(n9051), .ZN(n9068) );
  INV_X1 U10359 ( .A(n9052), .ZN(n9055) );
  NAND4_X1 U10360 ( .A1(n9056), .A2(n9055), .A3(n9054), .A4(n9053), .ZN(n9060)
         );
  INV_X1 U10361 ( .A(n9057), .ZN(n9059) );
  INV_X1 U10362 ( .A(n9058), .ZN(n9091) );
  NOR3_X1 U10363 ( .A1(n9060), .A2(n9059), .A3(n9091), .ZN(n9064) );
  INV_X1 U10364 ( .A(n9061), .ZN(n9062) );
  NAND4_X1 U10365 ( .A1(n9064), .A2(n9088), .A3(n9063), .A4(n9062), .ZN(n9066)
         );
  OR3_X1 U10366 ( .A1(n9066), .A2(n9572), .A3(n9065), .ZN(n9067) );
  NOR3_X1 U10367 ( .A1(n9069), .A2(n9068), .A3(n9067), .ZN(n9071) );
  NAND4_X1 U10368 ( .A1(n9073), .A2(n9072), .A3(n9071), .A4(n9070), .ZN(n9074)
         );
  NOR2_X1 U10369 ( .A1(n9171), .A2(n9074), .ZN(n9075) );
  NAND4_X1 U10370 ( .A1(n9361), .A2(n9398), .A3(n9385), .A4(n9075), .ZN(n9076)
         );
  NOR3_X1 U10371 ( .A1(n9334), .A2(n9347), .A3(n9076), .ZN(n9077) );
  XNOR2_X1 U10372 ( .A(n9447), .B(n9183), .ZN(n9293) );
  AND4_X1 U10373 ( .A1(n9285), .A2(n9315), .A3(n9077), .A4(n4647), .ZN(n9079)
         );
  NAND2_X1 U10374 ( .A1(n9432), .A2(n9277), .ZN(n9188) );
  INV_X1 U10375 ( .A(n9188), .ZN(n9078) );
  AND4_X1 U10376 ( .A1(n9248), .A2(n9276), .A3(n9079), .A4(n9264), .ZN(n9080)
         );
  INV_X1 U10377 ( .A(n9208), .ZN(n9107) );
  INV_X1 U10378 ( .A(n9083), .ZN(n9085) );
  OR3_X1 U10379 ( .A1(n9086), .A2(n9085), .A3(n9084), .ZN(n9096) );
  NAND2_X1 U10380 ( .A1(n9088), .A2(n9087), .ZN(n9094) );
  NAND3_X1 U10381 ( .A1(n9091), .A2(n9090), .A3(n9089), .ZN(n9092) );
  NAND3_X1 U10382 ( .A1(n9094), .A2(n9093), .A3(n9092), .ZN(n9095) );
  NAND2_X1 U10383 ( .A1(n9096), .A2(n9095), .ZN(n9098) );
  OAI21_X1 U10384 ( .B1(n9099), .B2(n9098), .A(n9097), .ZN(n9100) );
  NAND2_X1 U10385 ( .A1(n9101), .A2(n9100), .ZN(n9103) );
  AOI21_X1 U10386 ( .B1(n9104), .B2(n9103), .A(n9102), .ZN(n9105) );
  OR4_X1 U10387 ( .A1(n9108), .A2(n9107), .A3(n9106), .A4(n9105), .ZN(n9109)
         );
  NAND3_X1 U10388 ( .A1(n9111), .A2(n9110), .A3(n9109), .ZN(n9112) );
  NAND2_X1 U10389 ( .A1(n9113), .A2(n9112), .ZN(n9114) );
  NAND2_X1 U10390 ( .A1(n9115), .A2(n9114), .ZN(n9116) );
  MUX2_X1 U10391 ( .A(n9118), .B(n9117), .S(n9745), .Z(n9119) );
  NAND3_X1 U10392 ( .A1(n9125), .A2(n9124), .A3(n9162), .ZN(n9126) );
  OAI21_X1 U10393 ( .B1(n9127), .B2(n9129), .A(P1_B_REG_SCAN_IN), .ZN(n9128)
         );
  CLKBUF_X1 U10394 ( .A(P1_U4006), .Z(n9631) );
  MUX2_X1 U10395 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9164), .S(n9631), .Z(
        P1_U3586) );
  MUX2_X1 U10396 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9215), .S(n9631), .Z(
        P1_U3585) );
  MUX2_X1 U10397 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9234), .S(n9631), .Z(
        P1_U3584) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9250), .S(n9631), .Z(
        P1_U3583) );
  MUX2_X1 U10399 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9265), .S(n9631), .Z(
        P1_U3582) );
  MUX2_X1 U10400 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9277), .S(n9631), .Z(
        P1_U3581) );
  MUX2_X1 U10401 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9286), .S(n9631), .Z(
        P1_U3580) );
  MUX2_X1 U10402 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9303), .S(n9631), .Z(
        P1_U3579) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9316), .S(n9631), .Z(
        P1_U3578) );
  MUX2_X1 U10404 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9330), .S(n9631), .Z(
        P1_U3577) );
  MUX2_X1 U10405 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9349), .S(n9631), .Z(
        P1_U3576) );
  MUX2_X1 U10406 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9367), .S(n9631), .Z(
        P1_U3575) );
  MUX2_X1 U10407 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9375), .S(n9631), .Z(
        P1_U3574) );
  MUX2_X1 U10408 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9401), .S(n9631), .Z(
        P1_U3573) );
  MUX2_X1 U10409 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9376), .S(n9631), .Z(
        P1_U3572) );
  MUX2_X1 U10410 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9402), .S(n9631), .Z(
        P1_U3571) );
  MUX2_X1 U10411 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9130), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10412 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9131), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10413 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9132), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10414 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9133), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10415 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9576), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10416 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9134), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10417 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9577), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10418 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9135), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10419 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9136), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10420 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9137), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10421 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9138), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10422 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9139), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10423 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9140), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10424 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9141), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10425 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6776), .S(n9631), .Z(
        P1_U3555) );
  AOI21_X1 U10426 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9145), .A(n9142), .ZN(
        n9728) );
  XNOR2_X1 U10427 ( .A(n9148), .B(n9143), .ZN(n9729) );
  NAND2_X1 U10428 ( .A1(n9728), .A2(n9729), .ZN(n9727) );
  OAI21_X1 U10429 ( .B1(n9148), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9727), .ZN(
        n9144) );
  XNOR2_X1 U10430 ( .A(n9144), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9153) );
  NAND2_X1 U10431 ( .A1(n9145), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U10432 ( .A1(n9147), .A2(n9146), .ZN(n9721) );
  NAND2_X1 U10433 ( .A1(n9148), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9150) );
  OR2_X1 U10434 ( .A1(n9148), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9149) );
  AND2_X1 U10435 ( .A1(n9150), .A2(n9149), .ZN(n9720) );
  NAND2_X1 U10436 ( .A1(n9721), .A2(n9720), .ZN(n9719) );
  NAND2_X1 U10437 ( .A1(n9719), .A2(n9150), .ZN(n9151) );
  XNOR2_X1 U10438 ( .A(n9151), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9155) );
  INV_X1 U10439 ( .A(n9155), .ZN(n9152) );
  OAI21_X1 U10440 ( .B1(n9153), .B2(n9673), .A(n9724), .ZN(n9154) );
  AOI21_X1 U10441 ( .B1(n9155), .B2(n9718), .A(n9154), .ZN(n9157) );
  INV_X1 U10442 ( .A(n9158), .ZN(n9159) );
  OAI211_X1 U10443 ( .C1(n9161), .C2(n9717), .A(n9160), .B(n9159), .ZN(
        P1_U3260) );
  INV_X1 U10444 ( .A(n9426), .ZN(n9247) );
  INV_X1 U10445 ( .A(n9447), .ZN(n9301) );
  NOR2_X1 U10446 ( .A1(n9378), .A2(n9468), .ZN(n9356) );
  INV_X1 U10447 ( .A(n9464), .ZN(n9345) );
  NAND2_X1 U10448 ( .A1(n9356), .A2(n9345), .ZN(n9339) );
  NAND2_X1 U10449 ( .A1(n9247), .A2(n9256), .ZN(n9242) );
  NAND2_X1 U10450 ( .A1(n9162), .A2(P1_B_REG_SCAN_IN), .ZN(n9163) );
  AND2_X1 U10451 ( .A1(n9348), .A2(n9163), .ZN(n9214) );
  NAND2_X1 U10452 ( .A1(n9164), .A2(n9214), .ZN(n9411) );
  NOR2_X1 U10453 ( .A1(n9753), .A2(n9411), .ZN(n9168) );
  AOI21_X1 U10454 ( .B1(n9753), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9168), .ZN(
        n9166) );
  NAND2_X1 U10455 ( .A1(n8919), .A2(n9585), .ZN(n9165) );
  OAI211_X1 U10456 ( .C1(n9409), .C2(n9225), .A(n9166), .B(n9165), .ZN(
        P1_U3261) );
  INV_X1 U10457 ( .A(n9167), .ZN(n9413) );
  NAND2_X1 U10458 ( .A1(n9167), .A2(n9219), .ZN(n9410) );
  NAND3_X1 U10459 ( .A1(n4588), .A2(n9406), .A3(n9410), .ZN(n9170) );
  AOI21_X1 U10460 ( .B1(n9753), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9168), .ZN(
        n9169) );
  OAI211_X1 U10461 ( .C1(n9413), .C2(n9396), .A(n9170), .B(n9169), .ZN(
        P1_U3262) );
  INV_X1 U10462 ( .A(n9442), .ZN(n9186) );
  NAND2_X1 U10463 ( .A1(n9172), .A2(n9171), .ZN(n9175) );
  NAND2_X1 U10464 ( .A1(n9173), .A2(n9402), .ZN(n9174) );
  AND2_X1 U10465 ( .A1(n9480), .A2(n9376), .ZN(n9176) );
  OR2_X1 U10466 ( .A1(n9480), .A2(n9376), .ZN(n9177) );
  NAND2_X1 U10467 ( .A1(n9475), .A2(n9401), .ZN(n9178) );
  NAND2_X1 U10468 ( .A1(n9474), .A2(n9178), .ZN(n9355) );
  OR2_X1 U10469 ( .A1(n9468), .A2(n9375), .ZN(n9180) );
  AND2_X1 U10470 ( .A1(n9468), .A2(n9375), .ZN(n9179) );
  AOI21_X2 U10471 ( .B1(n9355), .B2(n9180), .A(n9179), .ZN(n9338) );
  NAND2_X1 U10472 ( .A1(n9464), .A2(n9367), .ZN(n9181) );
  INV_X1 U10473 ( .A(n9451), .ZN(n9312) );
  INV_X1 U10474 ( .A(n9294), .ZN(n9185) );
  NOR2_X1 U10475 ( .A1(n9229), .A2(n9190), .ZN(n9192) );
  INV_X1 U10476 ( .A(n9211), .ZN(n9191) );
  XNOR2_X1 U10477 ( .A(n9192), .B(n9191), .ZN(n9414) );
  INV_X1 U10478 ( .A(n9414), .ZN(n9228) );
  NAND2_X1 U10479 ( .A1(n9197), .A2(n9361), .ZN(n9366) );
  NAND2_X1 U10480 ( .A1(n9366), .A2(n9198), .ZN(n9346) );
  NOR2_X1 U10481 ( .A1(n9334), .A2(n9325), .ZN(n9200) );
  NAND2_X1 U10482 ( .A1(n9324), .A2(n9200), .ZN(n9327) );
  NAND2_X1 U10483 ( .A1(n9327), .A2(n9201), .ZN(n9314) );
  AND2_X2 U10484 ( .A1(n9283), .A2(n9204), .ZN(n9275) );
  INV_X1 U10485 ( .A(n9209), .ZN(n9210) );
  AOI21_X1 U10486 ( .B1(n9232), .B2(n9233), .A(n9210), .ZN(n9212) );
  XNOR2_X1 U10487 ( .A(n9212), .B(n9211), .ZN(n9213) );
  NAND2_X1 U10488 ( .A1(n9213), .A2(n9574), .ZN(n9217) );
  AOI22_X1 U10489 ( .A1(n9329), .A2(n9250), .B1(n9215), .B2(n9214), .ZN(n9216)
         );
  NAND2_X1 U10490 ( .A1(n9217), .A2(n9216), .ZN(n9418) );
  NAND2_X1 U10491 ( .A1(n9223), .A2(n9235), .ZN(n9218) );
  NAND2_X1 U10492 ( .A1(n9219), .A2(n9218), .ZN(n9416) );
  INV_X1 U10493 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9221) );
  OAI22_X1 U10494 ( .A1(n9751), .A2(n9221), .B1(n9220), .B2(n9743), .ZN(n9222)
         );
  AOI21_X1 U10495 ( .B1(n9223), .B2(n9585), .A(n9222), .ZN(n9224) );
  OAI21_X1 U10496 ( .B1(n9416), .B2(n9225), .A(n9224), .ZN(n9226) );
  AOI21_X1 U10497 ( .B1(n9418), .B2(n9751), .A(n9226), .ZN(n9227) );
  OAI21_X1 U10498 ( .B1(n9228), .B2(n9408), .A(n9227), .ZN(P1_U3355) );
  AOI21_X1 U10499 ( .B1(n9233), .B2(n9230), .A(n9229), .ZN(n9231) );
  INV_X1 U10500 ( .A(n9231), .ZN(n9425) );
  AOI22_X1 U10501 ( .A1(n9422), .A2(n9585), .B1(n9753), .B2(
        P1_REG2_REG_28__SCAN_IN), .ZN(n9240) );
  AOI211_X1 U10502 ( .C1(n9422), .C2(n9242), .A(n9793), .B(n4897), .ZN(n9421)
         );
  NAND2_X1 U10503 ( .A1(n9421), .A2(n9745), .ZN(n9236) );
  OAI211_X1 U10504 ( .C1(n9743), .C2(n9237), .A(n9424), .B(n9236), .ZN(n9238)
         );
  NAND2_X1 U10505 ( .A1(n9238), .A2(n9751), .ZN(n9239) );
  OAI211_X1 U10506 ( .C1(n9425), .C2(n9408), .A(n9240), .B(n9239), .ZN(
        P1_U3263) );
  XNOR2_X1 U10507 ( .A(n9241), .B(n4560), .ZN(n9430) );
  INV_X1 U10508 ( .A(n9256), .ZN(n9244) );
  INV_X1 U10509 ( .A(n9242), .ZN(n9243) );
  AOI21_X1 U10510 ( .B1(n9426), .B2(n9244), .A(n9243), .ZN(n9427) );
  AOI22_X1 U10511 ( .A1(n9753), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9245), .B2(
        n9583), .ZN(n9246) );
  OAI21_X1 U10512 ( .B1(n9247), .B2(n9396), .A(n9246), .ZN(n9253) );
  XNOR2_X1 U10513 ( .A(n9249), .B(n9248), .ZN(n9251) );
  AOI222_X1 U10514 ( .A1(n9574), .A2(n9251), .B1(n9250), .B2(n9400), .C1(n9277), .C2(n9329), .ZN(n9429) );
  NOR2_X1 U10515 ( .A1(n9429), .A2(n9753), .ZN(n9252) );
  AOI211_X1 U10516 ( .C1(n9406), .C2(n9427), .A(n9253), .B(n9252), .ZN(n9254)
         );
  OAI21_X1 U10517 ( .B1(n9430), .B2(n9408), .A(n9254), .ZN(P1_U3264) );
  XNOR2_X1 U10518 ( .A(n9255), .B(n9264), .ZN(n9435) );
  AOI211_X1 U10519 ( .C1(n9432), .C2(n9271), .A(n9793), .B(n9256), .ZN(n9431)
         );
  INV_X1 U10520 ( .A(n9257), .ZN(n9353) );
  INV_X1 U10521 ( .A(n9432), .ZN(n9260) );
  AOI22_X1 U10522 ( .A1(n9753), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9258), .B2(
        n9583), .ZN(n9259) );
  OAI21_X1 U10523 ( .B1(n9260), .B2(n9396), .A(n9259), .ZN(n9268) );
  NAND2_X1 U10524 ( .A1(n9262), .A2(n9261), .ZN(n9263) );
  XOR2_X1 U10525 ( .A(n9264), .B(n9263), .Z(n9266) );
  AOI222_X1 U10526 ( .A1(n9574), .A2(n9266), .B1(n9265), .B2(n9348), .C1(n9286), .C2(n9329), .ZN(n9434) );
  NOR2_X1 U10527 ( .A1(n9434), .A2(n9753), .ZN(n9267) );
  AOI211_X1 U10528 ( .C1(n9431), .C2(n9353), .A(n9268), .B(n9267), .ZN(n9269)
         );
  OAI21_X1 U10529 ( .B1(n9435), .B2(n9408), .A(n9269), .ZN(P1_U3265) );
  XOR2_X1 U10530 ( .A(n9276), .B(n9270), .Z(n9440) );
  INV_X1 U10531 ( .A(n9271), .ZN(n9272) );
  AOI211_X1 U10532 ( .C1(n9437), .C2(n4595), .A(n9793), .B(n9272), .ZN(n9436)
         );
  AOI22_X1 U10533 ( .A1(n9753), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9273), .B2(
        n9583), .ZN(n9274) );
  OAI21_X1 U10534 ( .B1(n4898), .B2(n9396), .A(n9274), .ZN(n9280) );
  XOR2_X1 U10535 ( .A(n9276), .B(n9275), .Z(n9278) );
  AOI222_X1 U10536 ( .A1(n9574), .A2(n9278), .B1(n9277), .B2(n9348), .C1(n9303), .C2(n9329), .ZN(n9439) );
  NOR2_X1 U10537 ( .A1(n9439), .A2(n9753), .ZN(n9279) );
  AOI211_X1 U10538 ( .C1(n9436), .C2(n9353), .A(n9280), .B(n9279), .ZN(n9281)
         );
  OAI21_X1 U10539 ( .B1(n9440), .B2(n9408), .A(n9281), .ZN(P1_U3266) );
  XOR2_X1 U10540 ( .A(n9282), .B(n9285), .Z(n9445) );
  AOI22_X1 U10541 ( .A1(n9442), .A2(n9585), .B1(n9753), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9292) );
  OAI21_X1 U10542 ( .B1(n9285), .B2(n9284), .A(n9283), .ZN(n9287) );
  AOI222_X1 U10543 ( .A1(n9574), .A2(n9287), .B1(n9286), .B2(n9348), .C1(n9316), .C2(n9329), .ZN(n9444) );
  AOI211_X1 U10544 ( .C1(n9442), .C2(n9295), .A(n9793), .B(n4899), .ZN(n9441)
         );
  NAND2_X1 U10545 ( .A1(n9441), .A2(n9745), .ZN(n9288) );
  OAI211_X1 U10546 ( .C1(n9743), .C2(n9289), .A(n9444), .B(n9288), .ZN(n9290)
         );
  NAND2_X1 U10547 ( .A1(n9290), .A2(n9751), .ZN(n9291) );
  OAI211_X1 U10548 ( .C1(n9445), .C2(n9408), .A(n9292), .B(n9291), .ZN(
        P1_U3267) );
  XNOR2_X1 U10549 ( .A(n9294), .B(n9293), .ZN(n9450) );
  INV_X1 U10550 ( .A(n9309), .ZN(n9297) );
  INV_X1 U10551 ( .A(n9295), .ZN(n9296) );
  AOI211_X1 U10552 ( .C1(n9447), .C2(n9297), .A(n9793), .B(n9296), .ZN(n9446)
         );
  INV_X1 U10553 ( .A(n9298), .ZN(n9299) );
  AOI22_X1 U10554 ( .A1(n9753), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9299), .B2(
        n9583), .ZN(n9300) );
  OAI21_X1 U10555 ( .B1(n9301), .B2(n9396), .A(n9300), .ZN(n9306) );
  XNOR2_X1 U10556 ( .A(n9302), .B(n4647), .ZN(n9304) );
  AOI222_X1 U10557 ( .A1(n9574), .A2(n9304), .B1(n9330), .B2(n9578), .C1(n9303), .C2(n9400), .ZN(n9449) );
  NOR2_X1 U10558 ( .A1(n9449), .A2(n9753), .ZN(n9305) );
  AOI211_X1 U10559 ( .C1(n9446), .C2(n9353), .A(n9306), .B(n9305), .ZN(n9307)
         );
  OAI21_X1 U10560 ( .B1(n9450), .B2(n9408), .A(n9307), .ZN(P1_U3268) );
  XNOR2_X1 U10561 ( .A(n9308), .B(n9315), .ZN(n9455) );
  AOI21_X1 U10562 ( .B1(n9451), .B2(n9321), .A(n9309), .ZN(n9452) );
  AOI22_X1 U10563 ( .A1(n9753), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9310), .B2(
        n9583), .ZN(n9311) );
  OAI21_X1 U10564 ( .B1(n9312), .B2(n9396), .A(n9311), .ZN(n9319) );
  OAI21_X1 U10565 ( .B1(n9315), .B2(n9314), .A(n9313), .ZN(n9317) );
  AOI222_X1 U10566 ( .A1(n9574), .A2(n9317), .B1(n9349), .B2(n9578), .C1(n9316), .C2(n9348), .ZN(n9454) );
  NOR2_X1 U10567 ( .A1(n9454), .A2(n9753), .ZN(n9318) );
  AOI211_X1 U10568 ( .C1(n9452), .C2(n9406), .A(n9319), .B(n9318), .ZN(n9320)
         );
  OAI21_X1 U10569 ( .B1(n9455), .B2(n9408), .A(n9320), .ZN(P1_U3269) );
  INV_X1 U10570 ( .A(n9321), .ZN(n9322) );
  AOI211_X1 U10571 ( .C1(n9458), .C2(n9339), .A(n9793), .B(n9322), .ZN(n9457)
         );
  NOR2_X1 U10572 ( .A1(n9743), .A2(n9323), .ZN(n9333) );
  INV_X1 U10573 ( .A(n9324), .ZN(n9326) );
  OAI21_X1 U10574 ( .B1(n9326), .B2(n9325), .A(n9334), .ZN(n9328) );
  NAND2_X1 U10575 ( .A1(n9328), .A2(n9327), .ZN(n9331) );
  AOI222_X1 U10576 ( .A1(n9574), .A2(n9331), .B1(n9330), .B2(n9400), .C1(n9367), .C2(n9329), .ZN(n9460) );
  INV_X1 U10577 ( .A(n9460), .ZN(n9332) );
  AOI211_X1 U10578 ( .C1(n9457), .C2(n9745), .A(n9333), .B(n9332), .ZN(n9337)
         );
  AOI22_X1 U10579 ( .A1(n9458), .A2(n9585), .B1(n9753), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9336) );
  INV_X1 U10580 ( .A(n9408), .ZN(n9387) );
  OR2_X1 U10581 ( .A1(n4544), .A2(n9334), .ZN(n9456) );
  NAND3_X1 U10582 ( .A1(n4945), .A2(n9387), .A3(n9456), .ZN(n9335) );
  OAI211_X1 U10583 ( .C1(n9337), .C2(n9753), .A(n9336), .B(n9335), .ZN(
        P1_U3270) );
  XOR2_X1 U10584 ( .A(n9347), .B(n9338), .Z(n9467) );
  INV_X1 U10585 ( .A(n9356), .ZN(n9341) );
  INV_X1 U10586 ( .A(n9339), .ZN(n9340) );
  AOI211_X1 U10587 ( .C1(n9464), .C2(n9341), .A(n9793), .B(n9340), .ZN(n9463)
         );
  INV_X1 U10588 ( .A(n9342), .ZN(n9343) );
  AOI22_X1 U10589 ( .A1(n9753), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9343), .B2(
        n9583), .ZN(n9344) );
  OAI21_X1 U10590 ( .B1(n9345), .B2(n9396), .A(n9344), .ZN(n9352) );
  XOR2_X1 U10591 ( .A(n9347), .B(n9346), .Z(n9350) );
  AOI222_X1 U10592 ( .A1(n9574), .A2(n9350), .B1(n9375), .B2(n9578), .C1(n9349), .C2(n9348), .ZN(n9466) );
  NOR2_X1 U10593 ( .A1(n9466), .A2(n9753), .ZN(n9351) );
  AOI211_X1 U10594 ( .C1(n9463), .C2(n9353), .A(n9352), .B(n9351), .ZN(n9354)
         );
  OAI21_X1 U10595 ( .B1(n9408), .B2(n9467), .A(n9354), .ZN(P1_U3271) );
  XOR2_X1 U10596 ( .A(n9361), .B(n9355), .Z(n9472) );
  AOI21_X1 U10597 ( .B1(n9468), .B2(n9378), .A(n9356), .ZN(n9469) );
  INV_X1 U10598 ( .A(n9357), .ZN(n9358) );
  AOI22_X1 U10599 ( .A1(n9753), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9358), .B2(
        n9583), .ZN(n9359) );
  OAI21_X1 U10600 ( .B1(n9360), .B2(n9396), .A(n9359), .ZN(n9370) );
  INV_X1 U10601 ( .A(n9361), .ZN(n9362) );
  NAND3_X1 U10602 ( .A1(n9364), .A2(n9363), .A3(n9362), .ZN(n9365) );
  NAND2_X1 U10603 ( .A1(n9366), .A2(n9365), .ZN(n9368) );
  AOI222_X1 U10604 ( .A1(n9574), .A2(n9368), .B1(n9401), .B2(n9578), .C1(n9367), .C2(n9348), .ZN(n9471) );
  NOR2_X1 U10605 ( .A1(n9471), .A2(n9753), .ZN(n9369) );
  AOI211_X1 U10606 ( .C1(n9469), .C2(n9406), .A(n9370), .B(n9369), .ZN(n9371)
         );
  OAI21_X1 U10607 ( .B1(n9408), .B2(n9472), .A(n9371), .ZN(P1_U3272) );
  NAND2_X1 U10608 ( .A1(n9373), .A2(n9372), .ZN(n9374) );
  XOR2_X1 U10609 ( .A(n9385), .B(n9374), .Z(n9377) );
  AOI222_X1 U10610 ( .A1(n9574), .A2(n9377), .B1(n9376), .B2(n9578), .C1(n9375), .C2(n9400), .ZN(n9478) );
  INV_X1 U10611 ( .A(n9378), .ZN(n9379) );
  AOI21_X1 U10612 ( .B1(n9475), .B2(n9391), .A(n9379), .ZN(n9476) );
  INV_X1 U10613 ( .A(n9475), .ZN(n9383) );
  INV_X1 U10614 ( .A(n9380), .ZN(n9381) );
  AOI22_X1 U10615 ( .A1(n9753), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9381), .B2(
        n9583), .ZN(n9382) );
  OAI21_X1 U10616 ( .B1(n9383), .B2(n9396), .A(n9382), .ZN(n9384) );
  AOI21_X1 U10617 ( .B1(n9476), .B2(n9406), .A(n9384), .ZN(n9389) );
  NAND2_X1 U10618 ( .A1(n9386), .A2(n9385), .ZN(n9473) );
  NAND3_X1 U10619 ( .A1(n9474), .A2(n9473), .A3(n9387), .ZN(n9388) );
  OAI211_X1 U10620 ( .C1(n9478), .C2(n9753), .A(n9389), .B(n9388), .ZN(
        P1_U3273) );
  XOR2_X1 U10621 ( .A(n9398), .B(n9390), .Z(n9485) );
  INV_X1 U10622 ( .A(n9391), .ZN(n9392) );
  AOI21_X1 U10623 ( .B1(n9480), .B2(n4545), .A(n9392), .ZN(n9481) );
  INV_X1 U10624 ( .A(n9393), .ZN(n9394) );
  AOI22_X1 U10625 ( .A1(n9753), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9394), .B2(
        n9583), .ZN(n9395) );
  OAI21_X1 U10626 ( .B1(n9397), .B2(n9396), .A(n9395), .ZN(n9405) );
  XNOR2_X1 U10627 ( .A(n9399), .B(n9398), .ZN(n9403) );
  AOI222_X1 U10628 ( .A1(n9574), .A2(n9403), .B1(n9402), .B2(n9578), .C1(n9401), .C2(n9400), .ZN(n9483) );
  NOR2_X1 U10629 ( .A1(n9483), .A2(n9753), .ZN(n9404) );
  AOI211_X1 U10630 ( .C1(n9481), .C2(n9406), .A(n9405), .B(n9404), .ZN(n9407)
         );
  OAI21_X1 U10631 ( .B1(n9408), .B2(n9485), .A(n9407), .ZN(P1_U3274) );
  MUX2_X1 U10632 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9494), .S(n9809), .Z(
        P1_U3554) );
  NAND3_X1 U10633 ( .A1(n4588), .A2(n9764), .A3(n9410), .ZN(n9412) );
  OAI211_X1 U10634 ( .C1(n9413), .C2(n9791), .A(n9412), .B(n9411), .ZN(n9495)
         );
  MUX2_X1 U10635 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9495), .S(n9809), .Z(
        P1_U3553) );
  NAND2_X1 U10636 ( .A1(n9414), .A2(n9788), .ZN(n9420) );
  OAI22_X1 U10637 ( .A1(n9416), .A2(n9793), .B1(n9415), .B2(n9791), .ZN(n9417)
         );
  NAND2_X1 U10638 ( .A1(n9420), .A2(n9419), .ZN(n9496) );
  MUX2_X1 U10639 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9496), .S(n9809), .Z(
        P1_U3552) );
  AOI21_X1 U10640 ( .B1(n9487), .B2(n9422), .A(n9421), .ZN(n9423) );
  OAI211_X1 U10641 ( .C1(n9425), .C2(n9484), .A(n9424), .B(n9423), .ZN(n9497)
         );
  MUX2_X1 U10642 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9497), .S(n9809), .Z(
        P1_U3551) );
  AOI22_X1 U10643 ( .A1(n9427), .A2(n9764), .B1(n9487), .B2(n9426), .ZN(n9428)
         );
  OAI211_X1 U10644 ( .C1(n9430), .C2(n9484), .A(n9429), .B(n9428), .ZN(n9498)
         );
  MUX2_X1 U10645 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9498), .S(n9809), .Z(
        P1_U3550) );
  AOI21_X1 U10646 ( .B1(n9487), .B2(n9432), .A(n9431), .ZN(n9433) );
  OAI211_X1 U10647 ( .C1(n9435), .C2(n9484), .A(n9434), .B(n9433), .ZN(n9499)
         );
  MUX2_X1 U10648 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9499), .S(n9809), .Z(
        P1_U3549) );
  AOI21_X1 U10649 ( .B1(n9487), .B2(n9437), .A(n9436), .ZN(n9438) );
  OAI211_X1 U10650 ( .C1(n9440), .C2(n9484), .A(n9439), .B(n9438), .ZN(n9500)
         );
  MUX2_X1 U10651 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9500), .S(n9809), .Z(
        P1_U3548) );
  AOI21_X1 U10652 ( .B1(n9487), .B2(n9442), .A(n9441), .ZN(n9443) );
  OAI211_X1 U10653 ( .C1(n9445), .C2(n9484), .A(n9444), .B(n9443), .ZN(n9501)
         );
  MUX2_X1 U10654 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9501), .S(n9809), .Z(
        P1_U3547) );
  AOI21_X1 U10655 ( .B1(n9487), .B2(n9447), .A(n9446), .ZN(n9448) );
  OAI211_X1 U10656 ( .C1(n9450), .C2(n9484), .A(n9449), .B(n9448), .ZN(n9502)
         );
  MUX2_X1 U10657 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9502), .S(n9809), .Z(
        P1_U3546) );
  AOI22_X1 U10658 ( .A1(n9452), .A2(n9764), .B1(n9487), .B2(n9451), .ZN(n9453)
         );
  OAI211_X1 U10659 ( .C1(n9455), .C2(n9484), .A(n9454), .B(n9453), .ZN(n9503)
         );
  MUX2_X1 U10660 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9503), .S(n9809), .Z(
        P1_U3545) );
  NAND2_X1 U10661 ( .A1(n9456), .A2(n9788), .ZN(n9462) );
  AOI21_X1 U10662 ( .B1(n9487), .B2(n9458), .A(n9457), .ZN(n9459) );
  OAI211_X1 U10663 ( .C1(n9462), .C2(n9461), .A(n9460), .B(n9459), .ZN(n9504)
         );
  MUX2_X1 U10664 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9504), .S(n9809), .Z(
        P1_U3544) );
  AOI21_X1 U10665 ( .B1(n9487), .B2(n9464), .A(n9463), .ZN(n9465) );
  OAI211_X1 U10666 ( .C1(n9467), .C2(n9484), .A(n9466), .B(n9465), .ZN(n9505)
         );
  MUX2_X1 U10667 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9505), .S(n9809), .Z(
        P1_U3543) );
  AOI22_X1 U10668 ( .A1(n9469), .A2(n9764), .B1(n9487), .B2(n9468), .ZN(n9470)
         );
  OAI211_X1 U10669 ( .C1(n9472), .C2(n9484), .A(n9471), .B(n9470), .ZN(n9506)
         );
  MUX2_X1 U10670 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9506), .S(n9809), .Z(
        P1_U3542) );
  NAND3_X1 U10671 ( .A1(n9474), .A2(n9788), .A3(n9473), .ZN(n9479) );
  AOI22_X1 U10672 ( .A1(n9476), .A2(n9764), .B1(n9487), .B2(n9475), .ZN(n9477)
         );
  NAND3_X1 U10673 ( .A1(n9479), .A2(n9478), .A3(n9477), .ZN(n9507) );
  MUX2_X1 U10674 ( .A(n9507), .B(P1_REG1_REG_18__SCAN_IN), .S(n9806), .Z(
        P1_U3541) );
  AOI22_X1 U10675 ( .A1(n9481), .A2(n9764), .B1(n9487), .B2(n9480), .ZN(n9482)
         );
  OAI211_X1 U10676 ( .C1(n9485), .C2(n9484), .A(n9483), .B(n9482), .ZN(n9508)
         );
  MUX2_X1 U10677 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9508), .S(n9809), .Z(
        P1_U3540) );
  AOI22_X1 U10678 ( .A1(n9488), .A2(n9764), .B1(n9487), .B2(n9486), .ZN(n9489)
         );
  OAI21_X1 U10679 ( .B1(n9491), .B2(n9490), .A(n9489), .ZN(n9492) );
  MUX2_X1 U10680 ( .A(n9509), .B(P1_REG1_REG_13__SCAN_IN), .S(n9806), .Z(
        P1_U3536) );
  MUX2_X1 U10681 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9494), .S(n9800), .Z(
        P1_U3522) );
  MUX2_X1 U10682 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9495), .S(n9800), .Z(
        P1_U3521) );
  MUX2_X1 U10683 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9496), .S(n9800), .Z(
        P1_U3520) );
  MUX2_X1 U10684 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9497), .S(n9800), .Z(
        P1_U3519) );
  MUX2_X1 U10685 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9498), .S(n9800), .Z(
        P1_U3518) );
  MUX2_X1 U10686 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9499), .S(n9800), .Z(
        P1_U3517) );
  MUX2_X1 U10687 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9500), .S(n9800), .Z(
        P1_U3516) );
  MUX2_X1 U10688 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9501), .S(n9800), .Z(
        P1_U3515) );
  MUX2_X1 U10689 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9502), .S(n9800), .Z(
        P1_U3514) );
  MUX2_X1 U10690 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9503), .S(n9800), .Z(
        P1_U3513) );
  MUX2_X1 U10691 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9504), .S(n9800), .Z(
        P1_U3512) );
  MUX2_X1 U10692 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9505), .S(n9800), .Z(
        P1_U3511) );
  MUX2_X1 U10693 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9506), .S(n9800), .Z(
        P1_U3510) );
  MUX2_X1 U10694 ( .A(n9507), .B(P1_REG0_REG_18__SCAN_IN), .S(n9799), .Z(
        P1_U3508) );
  MUX2_X1 U10695 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9508), .S(n9800), .Z(
        P1_U3505) );
  MUX2_X1 U10696 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9509), .S(n9800), .Z(
        P1_U3493) );
  NOR4_X1 U10697 ( .A1(n5778), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n5754), .ZN(n9510) );
  AOI21_X1 U10698 ( .B1(n9511), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9510), .ZN(
        n9512) );
  OAI21_X1 U10699 ( .B1(n9514), .B2(n9513), .A(n9512), .ZN(P1_U3322) );
  INV_X1 U10700 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10173) );
  NAND2_X1 U10701 ( .A1(n9515), .A2(n9518), .ZN(n9517) );
  OAI211_X1 U10702 ( .C1(n9522), .C2(n10173), .A(n9517), .B(n9516), .ZN(
        P1_U3325) );
  NAND2_X1 U10703 ( .A1(n9519), .A2(n9518), .ZN(n9521) );
  OAI211_X1 U10704 ( .C1(n9522), .C2(n10244), .A(n9521), .B(n9520), .ZN(
        P1_U3326) );
  MUX2_X1 U10705 ( .A(n9523), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U10706 ( .A1(n9724), .A2(n9524), .ZN(n9525) );
  AOI211_X1 U10707 ( .C1(n9730), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9526), .B(
        n9525), .ZN(n9536) );
  NAND2_X1 U10708 ( .A1(n9528), .A2(n9527), .ZN(n9529) );
  NAND3_X1 U10709 ( .A1(n9718), .A2(n9530), .A3(n9529), .ZN(n9535) );
  OAI211_X1 U10710 ( .C1(n9533), .C2(n9532), .A(n9731), .B(n9531), .ZN(n9534)
         );
  NAND3_X1 U10711 ( .A1(n9536), .A2(n9535), .A3(n9534), .ZN(P1_U3244) );
  INV_X1 U10712 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9964) );
  OAI22_X1 U10713 ( .A1(n9537), .A2(n9964), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10120), .ZN(n9538) );
  INV_X1 U10714 ( .A(n9538), .ZN(n9545) );
  INV_X1 U10715 ( .A(n9539), .ZN(n9543) );
  NAND2_X1 U10716 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9540) );
  NAND2_X1 U10717 ( .A1(n9541), .A2(n9540), .ZN(n9542) );
  NAND3_X1 U10718 ( .A1(n9827), .A2(n9543), .A3(n9542), .ZN(n9544) );
  OAI211_X1 U10719 ( .C1(n9828), .C2(n9546), .A(n9545), .B(n9544), .ZN(n9547)
         );
  INV_X1 U10720 ( .A(n9547), .ZN(n9553) );
  NOR2_X1 U10721 ( .A1(n9835), .A2(n9548), .ZN(n9551) );
  OAI211_X1 U10722 ( .C1(n9551), .C2(n9550), .A(n9825), .B(n9549), .ZN(n9552)
         );
  NAND2_X1 U10723 ( .A1(n9553), .A2(n9552), .ZN(P2_U3246) );
  AOI22_X1 U10724 ( .A1(n9832), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9566) );
  INV_X1 U10725 ( .A(n9828), .ZN(n9560) );
  AOI211_X1 U10726 ( .C1(n9557), .C2(n9556), .A(n9555), .B(n9554), .ZN(n9558)
         );
  AOI21_X1 U10727 ( .B1(n9560), .B2(n9559), .A(n9558), .ZN(n9565) );
  OAI211_X1 U10728 ( .C1(n9563), .C2(n9562), .A(n9825), .B(n9561), .ZN(n9564)
         );
  NAND3_X1 U10729 ( .A1(n9566), .A2(n9565), .A3(n9564), .ZN(P2_U3247) );
  XNOR2_X1 U10730 ( .A(n9567), .B(n9572), .ZN(n9599) );
  NAND2_X1 U10731 ( .A1(n9569), .A2(n9568), .ZN(n9571) );
  NAND2_X1 U10732 ( .A1(n9571), .A2(n9570), .ZN(n9573) );
  XNOR2_X1 U10733 ( .A(n9573), .B(n9572), .ZN(n9575) );
  NAND2_X1 U10734 ( .A1(n9575), .A2(n9574), .ZN(n9580) );
  AOI22_X1 U10735 ( .A1(n9578), .A2(n9577), .B1(n9576), .B2(n9400), .ZN(n9579)
         );
  NAND2_X1 U10736 ( .A1(n9580), .A2(n9579), .ZN(n9598) );
  AOI21_X1 U10737 ( .B1(n9599), .B2(n9581), .A(n9598), .ZN(n9595) );
  INV_X1 U10738 ( .A(n9582), .ZN(n9584) );
  AOI222_X1 U10739 ( .A1(n9587), .A2(n9585), .B1(n9584), .B2(n9583), .C1(
        P1_REG2_REG_10__SCAN_IN), .C2(n9753), .ZN(n9594) );
  INV_X1 U10740 ( .A(n9586), .ZN(n9589) );
  OAI211_X1 U10741 ( .C1(n9589), .C2(n4893), .A(n9764), .B(n9588), .ZN(n9596)
         );
  INV_X1 U10742 ( .A(n9596), .ZN(n9590) );
  AOI22_X1 U10743 ( .A1(n9599), .A2(n9592), .B1(n9591), .B2(n9590), .ZN(n9593)
         );
  OAI211_X1 U10744 ( .C1(n9753), .C2(n9595), .A(n9594), .B(n9593), .ZN(
        P1_U3281) );
  OAI21_X1 U10745 ( .B1(n4893), .B2(n9791), .A(n9596), .ZN(n9597) );
  AOI211_X1 U10746 ( .C1(n9599), .C2(n9788), .A(n9598), .B(n9597), .ZN(n9600)
         );
  AOI22_X1 U10747 ( .A1(n9800), .A2(n9600), .B1(n6005), .B2(n9799), .ZN(
        P1_U3484) );
  AOI22_X1 U10748 ( .A1(n9809), .A2(n9600), .B1(n6552), .B2(n9806), .ZN(
        P1_U3533) );
  OAI21_X1 U10749 ( .B1(n9602), .B2(n9791), .A(n9601), .ZN(n9603) );
  AOI211_X1 U10750 ( .C1(n9605), .C2(n9788), .A(n9604), .B(n9603), .ZN(n9619)
         );
  AOI22_X1 U10751 ( .A1(n9809), .A2(n9619), .B1(n7675), .B2(n9806), .ZN(
        P1_U3539) );
  INV_X1 U10752 ( .A(n9606), .ZN(n9607) );
  OAI22_X1 U10753 ( .A1(n9608), .A2(n9793), .B1(n9607), .B2(n9791), .ZN(n9610)
         );
  AOI211_X1 U10754 ( .C1(n9798), .C2(n9611), .A(n9610), .B(n9609), .ZN(n9621)
         );
  AOI22_X1 U10755 ( .A1(n9809), .A2(n9621), .B1(n9612), .B2(n9806), .ZN(
        P1_U3538) );
  OAI21_X1 U10756 ( .B1(n9614), .B2(n9791), .A(n9613), .ZN(n9615) );
  AOI211_X1 U10757 ( .C1(n9617), .C2(n9788), .A(n9616), .B(n9615), .ZN(n9622)
         );
  AOI22_X1 U10758 ( .A1(n9809), .A2(n9622), .B1(n6551), .B2(n9806), .ZN(
        P1_U3537) );
  INV_X1 U10759 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9618) );
  AOI22_X1 U10760 ( .A1(n9800), .A2(n9619), .B1(n9618), .B2(n9799), .ZN(
        P1_U3502) );
  INV_X1 U10761 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9620) );
  AOI22_X1 U10762 ( .A1(n9800), .A2(n9621), .B1(n9620), .B2(n9799), .ZN(
        P1_U3499) );
  AOI22_X1 U10763 ( .A1(n9800), .A2(n9622), .B1(n6092), .B2(n9799), .ZN(
        P1_U3496) );
  INV_X1 U10764 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10283) );
  XOR2_X1 U10765 ( .A(n10283), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XOR2_X1 U10766 ( .A(n4858), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  OAI22_X1 U10767 ( .A1(n9724), .A2(n9624), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9623), .ZN(n9625) );
  AOI21_X1 U10768 ( .B1(n9730), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n9625), .ZN(
        n9644) );
  MUX2_X1 U10769 ( .A(n9628), .B(n9627), .S(n9626), .Z(n9633) );
  NAND2_X1 U10770 ( .A1(n9629), .A2(n10275), .ZN(n9630) );
  OAI211_X1 U10771 ( .C1(n9633), .C2(n9632), .A(n9631), .B(n9630), .ZN(n9658)
         );
  NAND2_X1 U10772 ( .A1(n9635), .A2(n9634), .ZN(n9636) );
  NAND3_X1 U10773 ( .A1(n9731), .A2(n9637), .A3(n9636), .ZN(n9643) );
  AOI211_X1 U10774 ( .C1(n9640), .C2(n9639), .A(n9638), .B(n9690), .ZN(n9641)
         );
  INV_X1 U10775 ( .A(n9641), .ZN(n9642) );
  NAND4_X1 U10776 ( .A1(n9644), .A2(n9658), .A3(n9643), .A4(n9642), .ZN(
        P1_U3243) );
  INV_X1 U10777 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9660) );
  AOI21_X1 U10778 ( .B1(n9647), .B2(n9646), .A(n9645), .ZN(n9656) );
  AOI21_X1 U10779 ( .B1(n9650), .B2(n9649), .A(n9648), .ZN(n9651) );
  NOR2_X1 U10780 ( .A1(n9690), .A2(n9651), .ZN(n9652) );
  AOI211_X1 U10781 ( .C1(n9705), .C2(n9654), .A(n9653), .B(n9652), .ZN(n9655)
         );
  OAI21_X1 U10782 ( .B1(n9656), .B2(n9673), .A(n9655), .ZN(n9657) );
  INV_X1 U10783 ( .A(n9657), .ZN(n9659) );
  OAI211_X1 U10784 ( .C1(n9660), .C2(n9717), .A(n9659), .B(n9658), .ZN(
        P1_U3245) );
  INV_X1 U10785 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9677) );
  AOI21_X1 U10786 ( .B1(n9663), .B2(n9662), .A(n9661), .ZN(n9674) );
  AOI21_X1 U10787 ( .B1(n9666), .B2(n9665), .A(n9664), .ZN(n9667) );
  OR2_X1 U10788 ( .A1(n9667), .A2(n9690), .ZN(n9672) );
  INV_X1 U10789 ( .A(n9668), .ZN(n9670) );
  AOI21_X1 U10790 ( .B1(n9705), .B2(n9670), .A(n9669), .ZN(n9671) );
  OAI211_X1 U10791 ( .C1(n9674), .C2(n9673), .A(n9672), .B(n9671), .ZN(n9675)
         );
  INV_X1 U10792 ( .A(n9675), .ZN(n9676) );
  OAI21_X1 U10793 ( .B1(n9717), .B2(n9677), .A(n9676), .ZN(P1_U3248) );
  NAND3_X1 U10794 ( .A1(n9731), .A2(P1_REG1_REG_8__SCAN_IN), .A3(n9683), .ZN(
        n9679) );
  NAND3_X1 U10795 ( .A1(n9718), .A2(P1_REG2_REG_8__SCAN_IN), .A3(n9685), .ZN(
        n9678) );
  NAND3_X1 U10796 ( .A1(n9679), .A2(n9724), .A3(n9678), .ZN(n9680) );
  AOI22_X1 U10797 ( .A1(n9681), .A2(n9680), .B1(n9730), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n9689) );
  OAI211_X1 U10798 ( .C1(n9683), .C2(n9682), .A(n9731), .B(n9698), .ZN(n9687)
         );
  OAI211_X1 U10799 ( .C1(n9685), .C2(n9684), .A(n9718), .B(n9693), .ZN(n9686)
         );
  NAND4_X1 U10800 ( .A1(n9689), .A2(n9688), .A3(n9687), .A4(n9686), .ZN(
        P1_U3249) );
  AOI211_X1 U10801 ( .C1(n9693), .C2(n9692), .A(n9691), .B(n9690), .ZN(n9694)
         );
  AOI211_X1 U10802 ( .C1(n9705), .C2(n9696), .A(n9695), .B(n9694), .ZN(n9702)
         );
  OAI21_X1 U10803 ( .B1(n9699), .B2(n9698), .A(n9697), .ZN(n9700) );
  AOI22_X1 U10804 ( .A1(n9700), .A2(n9731), .B1(n9730), .B2(
        P1_ADDR_REG_9__SCAN_IN), .ZN(n9701) );
  NAND2_X1 U10805 ( .A1(n9702), .A2(n9701), .ZN(P1_U3250) );
  INV_X1 U10806 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9716) );
  AOI21_X1 U10807 ( .B1(n9705), .B2(n9704), .A(n9703), .ZN(n9715) );
  OAI21_X1 U10808 ( .B1(n9708), .B2(n9707), .A(n9706), .ZN(n9713) );
  OAI21_X1 U10809 ( .B1(n9711), .B2(n9710), .A(n9709), .ZN(n9712) );
  AOI22_X1 U10810 ( .A1(n9713), .A2(n9718), .B1(n9731), .B2(n9712), .ZN(n9714)
         );
  OAI211_X1 U10811 ( .C1(n9717), .C2(n9716), .A(n9715), .B(n9714), .ZN(
        P1_U3252) );
  OAI211_X1 U10812 ( .C1(n9721), .C2(n9720), .A(n9719), .B(n9718), .ZN(n9723)
         );
  OAI211_X1 U10813 ( .C1(n9725), .C2(n9724), .A(n9723), .B(n9722), .ZN(n9726)
         );
  INV_X1 U10814 ( .A(n9726), .ZN(n9734) );
  OAI21_X1 U10815 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n9732) );
  AOI22_X1 U10816 ( .A1(n9732), .A2(n9731), .B1(n9730), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9733) );
  NAND2_X1 U10817 ( .A1(n9734), .A2(n9733), .ZN(P1_U3259) );
  NAND2_X1 U10818 ( .A1(n9736), .A2(n9735), .ZN(n9748) );
  INV_X1 U10819 ( .A(n9737), .ZN(n9746) );
  NAND2_X1 U10820 ( .A1(n9739), .A2(n9738), .ZN(n9740) );
  OAI211_X1 U10821 ( .C1(n9743), .C2(n9742), .A(n9741), .B(n9740), .ZN(n9744)
         );
  AOI21_X1 U10822 ( .B1(n9746), .B2(n9745), .A(n9744), .ZN(n9747) );
  NAND2_X1 U10823 ( .A1(n9748), .A2(n9747), .ZN(n9750) );
  NOR2_X1 U10824 ( .A1(n9750), .A2(n9749), .ZN(n9752) );
  AOI22_X1 U10825 ( .A1(n9753), .A2(n5887), .B1(n9752), .B2(n9751), .ZN(
        P1_U3286) );
  AND2_X1 U10826 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9757), .ZN(P1_U3292) );
  AND2_X1 U10827 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9757), .ZN(P1_U3293) );
  AND2_X1 U10828 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9757), .ZN(P1_U3294) );
  AND2_X1 U10829 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9757), .ZN(P1_U3295) );
  AND2_X1 U10830 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9757), .ZN(P1_U3296) );
  AND2_X1 U10831 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9757), .ZN(P1_U3297) );
  AND2_X1 U10832 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9757), .ZN(P1_U3298) );
  AND2_X1 U10833 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9757), .ZN(P1_U3299) );
  AND2_X1 U10834 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9757), .ZN(P1_U3300) );
  AND2_X1 U10835 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9757), .ZN(P1_U3301) );
  AND2_X1 U10836 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9757), .ZN(P1_U3302) );
  AND2_X1 U10837 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9757), .ZN(P1_U3303) );
  AND2_X1 U10838 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9757), .ZN(P1_U3304) );
  AND2_X1 U10839 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9757), .ZN(P1_U3305) );
  AND2_X1 U10840 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9757), .ZN(P1_U3306) );
  AND2_X1 U10841 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9757), .ZN(P1_U3307) );
  AND2_X1 U10842 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9757), .ZN(P1_U3308) );
  AND2_X1 U10843 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9757), .ZN(P1_U3309) );
  AND2_X1 U10844 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9757), .ZN(P1_U3310) );
  AND2_X1 U10845 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9757), .ZN(P1_U3311) );
  AND2_X1 U10846 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9757), .ZN(P1_U3312) );
  AND2_X1 U10847 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9757), .ZN(P1_U3313) );
  AND2_X1 U10848 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9757), .ZN(P1_U3314) );
  AND2_X1 U10849 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9757), .ZN(P1_U3315) );
  AND2_X1 U10850 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9757), .ZN(P1_U3316) );
  AND2_X1 U10851 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9757), .ZN(P1_U3317) );
  AND2_X1 U10852 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9757), .ZN(P1_U3318) );
  INV_X1 U10853 ( .A(n9757), .ZN(n9756) );
  INV_X1 U10854 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10245) );
  NOR2_X1 U10855 ( .A1(n9756), .A2(n10245), .ZN(P1_U3319) );
  INV_X1 U10856 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10082) );
  NOR2_X1 U10857 ( .A1(n9756), .A2(n10082), .ZN(P1_U3320) );
  AND2_X1 U10858 ( .A1(n9757), .A2(P1_D_REG_2__SCAN_IN), .ZN(P1_U3321) );
  INV_X1 U10859 ( .A(n9758), .ZN(n9762) );
  OAI21_X1 U10860 ( .B1(n4675), .B2(n9791), .A(n9759), .ZN(n9761) );
  AOI211_X1 U10861 ( .C1(n9798), .C2(n9762), .A(n9761), .B(n9760), .ZN(n9801)
         );
  AOI22_X1 U10862 ( .A1(n9800), .A2(n9801), .B1(n5814), .B2(n9799), .ZN(
        P1_U3457) );
  INV_X1 U10863 ( .A(n9763), .ZN(n9771) );
  NAND2_X1 U10864 ( .A1(n9765), .A2(n9764), .ZN(n9768) );
  OAI22_X1 U10865 ( .A1(n9768), .A2(n9767), .B1(n9766), .B2(n9791), .ZN(n9770)
         );
  AOI211_X1 U10866 ( .C1(n9798), .C2(n9771), .A(n9770), .B(n9769), .ZN(n9802)
         );
  INV_X1 U10867 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9772) );
  AOI22_X1 U10868 ( .A1(n9800), .A2(n9802), .B1(n9772), .B2(n9799), .ZN(
        P1_U3460) );
  OAI22_X1 U10869 ( .A1(n9774), .A2(n9793), .B1(n9773), .B2(n9791), .ZN(n9776)
         );
  AOI211_X1 U10870 ( .C1(n9798), .C2(n9777), .A(n9776), .B(n9775), .ZN(n9803)
         );
  INV_X1 U10871 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9778) );
  AOI22_X1 U10872 ( .A1(n9800), .A2(n9803), .B1(n9778), .B2(n9799), .ZN(
        P1_U3466) );
  OAI22_X1 U10873 ( .A1(n9780), .A2(n9793), .B1(n9779), .B2(n9791), .ZN(n9782)
         );
  AOI211_X1 U10874 ( .C1(n9798), .C2(n9783), .A(n9782), .B(n9781), .ZN(n9804)
         );
  AOI22_X1 U10875 ( .A1(n9800), .A2(n9804), .B1(n5923), .B2(n9799), .ZN(
        P1_U3472) );
  OAI22_X1 U10876 ( .A1(n9785), .A2(n9793), .B1(n9784), .B2(n9791), .ZN(n9786)
         );
  AOI211_X1 U10877 ( .C1(n9789), .C2(n9788), .A(n9787), .B(n9786), .ZN(n9805)
         );
  INV_X1 U10878 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9790) );
  AOI22_X1 U10879 ( .A1(n9800), .A2(n9805), .B1(n9790), .B2(n9799), .ZN(
        P1_U3478) );
  OAI22_X1 U10880 ( .A1(n9794), .A2(n9793), .B1(n9792), .B2(n9791), .ZN(n9796)
         );
  AOI211_X1 U10881 ( .C1(n9798), .C2(n9797), .A(n9796), .B(n9795), .ZN(n9808)
         );
  AOI22_X1 U10882 ( .A1(n9800), .A2(n9808), .B1(n5984), .B2(n9799), .ZN(
        P1_U3481) );
  AOI22_X1 U10883 ( .A1(n9809), .A2(n9801), .B1(n5813), .B2(n9806), .ZN(
        P1_U3524) );
  AOI22_X1 U10884 ( .A1(n9809), .A2(n9802), .B1(n6558), .B2(n9806), .ZN(
        P1_U3525) );
  AOI22_X1 U10885 ( .A1(n9809), .A2(n9803), .B1(n5870), .B2(n9806), .ZN(
        P1_U3527) );
  AOI22_X1 U10886 ( .A1(n9809), .A2(n9804), .B1(n5922), .B2(n9806), .ZN(
        P1_U3529) );
  AOI22_X1 U10887 ( .A1(n9809), .A2(n9805), .B1(n6554), .B2(n9806), .ZN(
        P1_U3531) );
  INV_X1 U10888 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9807) );
  AOI22_X1 U10889 ( .A1(n9809), .A2(n9808), .B1(n9807), .B2(n9806), .ZN(
        P1_U3532) );
  OAI21_X1 U10890 ( .B1(n4487), .B2(n9811), .A(n9810), .ZN(n9822) );
  OAI22_X1 U10891 ( .A1(n9815), .A2(n9814), .B1(n9813), .B2(n9812), .ZN(n9837)
         );
  AOI21_X1 U10892 ( .B1(n9817), .B2(n9837), .A(n9816), .ZN(n9818) );
  OAI21_X1 U10893 ( .B1(n9929), .B2(n9819), .A(n9818), .ZN(n9820) );
  AOI21_X1 U10894 ( .B1(n9822), .B2(n9821), .A(n9820), .ZN(n9823) );
  OAI21_X1 U10895 ( .B1(n9824), .B2(n9846), .A(n9823), .ZN(P2_U3232) );
  AOI22_X1 U10896 ( .A1(n9825), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9827), .ZN(n9836) );
  NAND2_X1 U10897 ( .A1(n9827), .A2(n9826), .ZN(n9829) );
  OAI211_X1 U10898 ( .C1(n9830), .C2(P2_REG2_REG_0__SCAN_IN), .A(n9829), .B(
        n9828), .ZN(n9831) );
  INV_X1 U10899 ( .A(n9831), .ZN(n9834) );
  AOI22_X1 U10900 ( .A1(n9832), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9833) );
  OAI221_X1 U10901 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9836), .C1(n9835), .C2(
        n9834), .A(n9833), .ZN(P2_U3245) );
  XOR2_X1 U10902 ( .A(n9840), .B(n7272), .Z(n9839) );
  AOI21_X1 U10903 ( .B1(n9839), .B2(n9838), .A(n9837), .ZN(n9928) );
  XNOR2_X1 U10904 ( .A(n7268), .B(n9840), .ZN(n9931) );
  OAI21_X1 U10905 ( .B1(n9842), .B2(n9929), .A(n9841), .ZN(n9844) );
  OR2_X1 U10906 ( .A1(n9844), .A2(n9843), .ZN(n9927) );
  OAI22_X1 U10907 ( .A1(n9927), .A2(n9847), .B1(n9846), .B2(n9845), .ZN(n9848)
         );
  AOI21_X1 U10908 ( .B1(n9849), .B2(P2_REG2_REG_4__SCAN_IN), .A(n9848), .ZN(
        n9850) );
  OAI21_X1 U10909 ( .B1(n9929), .B2(n9851), .A(n9850), .ZN(n9852) );
  AOI21_X1 U10910 ( .B1(n9853), .B2(n9931), .A(n9852), .ZN(n9854) );
  OAI21_X1 U10911 ( .B1(n9855), .B2(n9928), .A(n9854), .ZN(P2_U3292) );
  INV_X1 U10912 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9858) );
  NOR2_X1 U10913 ( .A1(n9893), .A2(n9858), .ZN(P2_U3297) );
  INV_X1 U10914 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9859) );
  NOR2_X1 U10915 ( .A1(n9893), .A2(n9859), .ZN(P2_U3298) );
  INV_X1 U10916 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9860) );
  NOR2_X1 U10917 ( .A1(n9893), .A2(n9860), .ZN(P2_U3299) );
  INV_X1 U10918 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9861) );
  NOR2_X1 U10919 ( .A1(n9893), .A2(n9861), .ZN(P2_U3300) );
  INV_X1 U10920 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9862) );
  NOR2_X1 U10921 ( .A1(n9872), .A2(n9862), .ZN(P2_U3301) );
  INV_X1 U10922 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9863) );
  NOR2_X1 U10923 ( .A1(n9872), .A2(n9863), .ZN(P2_U3302) );
  INV_X1 U10924 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9864) );
  NOR2_X1 U10925 ( .A1(n9872), .A2(n9864), .ZN(P2_U3303) );
  INV_X1 U10926 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n9865) );
  NOR2_X1 U10927 ( .A1(n9872), .A2(n9865), .ZN(P2_U3304) );
  INV_X1 U10928 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9866) );
  NOR2_X1 U10929 ( .A1(n9872), .A2(n9866), .ZN(P2_U3305) );
  INV_X1 U10930 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9867) );
  NOR2_X1 U10931 ( .A1(n9872), .A2(n9867), .ZN(P2_U3306) );
  INV_X1 U10932 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9868) );
  NOR2_X1 U10933 ( .A1(n9872), .A2(n9868), .ZN(P2_U3307) );
  INV_X1 U10934 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9869) );
  NOR2_X1 U10935 ( .A1(n9872), .A2(n9869), .ZN(P2_U3308) );
  INV_X1 U10936 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9870) );
  NOR2_X1 U10937 ( .A1(n9872), .A2(n9870), .ZN(P2_U3309) );
  INV_X1 U10938 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9871) );
  NOR2_X1 U10939 ( .A1(n9872), .A2(n9871), .ZN(P2_U3310) );
  INV_X1 U10940 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9873) );
  NOR2_X1 U10941 ( .A1(n9893), .A2(n9873), .ZN(P2_U3311) );
  INV_X1 U10942 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9874) );
  NOR2_X1 U10943 ( .A1(n9893), .A2(n9874), .ZN(P2_U3312) );
  INV_X1 U10944 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n9875) );
  NOR2_X1 U10945 ( .A1(n9893), .A2(n9875), .ZN(P2_U3313) );
  INV_X1 U10946 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9876) );
  NOR2_X1 U10947 ( .A1(n9893), .A2(n9876), .ZN(P2_U3314) );
  INV_X1 U10948 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9877) );
  NOR2_X1 U10949 ( .A1(n9893), .A2(n9877), .ZN(P2_U3315) );
  INV_X1 U10950 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9878) );
  NOR2_X1 U10951 ( .A1(n9893), .A2(n9878), .ZN(P2_U3316) );
  INV_X1 U10952 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9879) );
  NOR2_X1 U10953 ( .A1(n9893), .A2(n9879), .ZN(P2_U3317) );
  INV_X1 U10954 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9880) );
  NOR2_X1 U10955 ( .A1(n9893), .A2(n9880), .ZN(P2_U3318) );
  INV_X1 U10956 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9881) );
  NOR2_X1 U10957 ( .A1(n9893), .A2(n9881), .ZN(P2_U3319) );
  INV_X1 U10958 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9882) );
  NOR2_X1 U10959 ( .A1(n9893), .A2(n9882), .ZN(P2_U3320) );
  INV_X1 U10960 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9883) );
  NOR2_X1 U10961 ( .A1(n9893), .A2(n9883), .ZN(P2_U3321) );
  INV_X1 U10962 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9884) );
  NOR2_X1 U10963 ( .A1(n9893), .A2(n9884), .ZN(P2_U3322) );
  NOR2_X1 U10964 ( .A1(n9893), .A2(n9885), .ZN(P2_U3323) );
  NOR2_X1 U10965 ( .A1(n9893), .A2(n9886), .ZN(P2_U3324) );
  NOR2_X1 U10966 ( .A1(n9893), .A2(n9887), .ZN(P2_U3325) );
  NOR2_X1 U10967 ( .A1(n9893), .A2(n9888), .ZN(P2_U3326) );
  OAI22_X1 U10968 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9893), .B1(n9892), .B2(
        n9889), .ZN(n9890) );
  INV_X1 U10969 ( .A(n9890), .ZN(P2_U3437) );
  OAI22_X1 U10970 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n9893), .B1(n9892), .B2(
        n9891), .ZN(n9894) );
  INV_X1 U10971 ( .A(n9894), .ZN(P2_U3438) );
  INV_X1 U10972 ( .A(n9895), .ZN(n9901) );
  OAI22_X1 U10973 ( .A1(n9899), .A2(n9898), .B1(n9897), .B2(n9896), .ZN(n9900)
         );
  NOR2_X1 U10974 ( .A1(n9901), .A2(n9900), .ZN(n9950) );
  AOI22_X1 U10975 ( .A1(n9949), .A2(n9950), .B1(n5074), .B2(n9948), .ZN(
        P2_U3451) );
  INV_X1 U10976 ( .A(n9902), .ZN(n9907) );
  OAI21_X1 U10977 ( .B1(n6422), .B2(n9940), .A(n9903), .ZN(n9906) );
  INV_X1 U10978 ( .A(n9904), .ZN(n9905) );
  AOI211_X1 U10979 ( .C1(n9946), .C2(n9907), .A(n9906), .B(n9905), .ZN(n9951)
         );
  INV_X1 U10980 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9908) );
  AOI22_X1 U10981 ( .A1(n9949), .A2(n9951), .B1(n9908), .B2(n9948), .ZN(
        P2_U3454) );
  INV_X1 U10982 ( .A(n9909), .ZN(n9914) );
  OAI211_X1 U10983 ( .C1(n9912), .C2(n9940), .A(n9911), .B(n9910), .ZN(n9913)
         );
  AOI21_X1 U10984 ( .B1(n9914), .B2(n9946), .A(n9913), .ZN(n9953) );
  INV_X1 U10985 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9915) );
  AOI22_X1 U10986 ( .A1(n9949), .A2(n9953), .B1(n9915), .B2(n9948), .ZN(
        P2_U3457) );
  INV_X1 U10987 ( .A(n9922), .ZN(n9924) );
  AOI21_X1 U10988 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(n9919) );
  OAI211_X1 U10989 ( .C1(n9922), .C2(n9921), .A(n9920), .B(n9919), .ZN(n9923)
         );
  AOI21_X1 U10990 ( .B1(n9925), .B2(n9924), .A(n9923), .ZN(n9954) );
  INV_X1 U10991 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9926) );
  AOI22_X1 U10992 ( .A1(n9949), .A2(n9954), .B1(n9926), .B2(n9948), .ZN(
        P2_U3460) );
  OAI211_X1 U10993 ( .C1(n9929), .C2(n9940), .A(n9928), .B(n9927), .ZN(n9930)
         );
  AOI21_X1 U10994 ( .B1(n9946), .B2(n9931), .A(n9930), .ZN(n9956) );
  AOI22_X1 U10995 ( .A1(n9949), .A2(n9956), .B1(n5122), .B2(n9948), .ZN(
        P2_U3463) );
  OAI21_X1 U10996 ( .B1(n9933), .B2(n9940), .A(n9932), .ZN(n9934) );
  AOI21_X1 U10997 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(n9937) );
  AND2_X1 U10998 ( .A1(n9938), .A2(n9937), .ZN(n9957) );
  INV_X1 U10999 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9939) );
  AOI22_X1 U11000 ( .A1(n9949), .A2(n9957), .B1(n9939), .B2(n9948), .ZN(
        P2_U3478) );
  OAI22_X1 U11001 ( .A1(n9943), .A2(n9942), .B1(n9941), .B2(n9940), .ZN(n9945)
         );
  AOI211_X1 U11002 ( .C1(n9947), .C2(n9946), .A(n9945), .B(n9944), .ZN(n9959)
         );
  AOI22_X1 U11003 ( .A1(n9949), .A2(n9959), .B1(n5295), .B2(n9948), .ZN(
        P2_U3484) );
  AOI22_X1 U11004 ( .A1(n9960), .A2(n9950), .B1(n9826), .B2(n9958), .ZN(
        P2_U3520) );
  AOI22_X1 U11005 ( .A1(n9960), .A2(n9951), .B1(n6683), .B2(n9958), .ZN(
        P2_U3521) );
  INV_X1 U11006 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9952) );
  AOI22_X1 U11007 ( .A1(n9960), .A2(n9953), .B1(n9952), .B2(n9958), .ZN(
        P2_U3522) );
  AOI22_X1 U11008 ( .A1(n9960), .A2(n9954), .B1(n5104), .B2(n9958), .ZN(
        P2_U3523) );
  INV_X1 U11009 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U11010 ( .A1(n9960), .A2(n9956), .B1(n9955), .B2(n9958), .ZN(
        P2_U3524) );
  AOI22_X1 U11011 ( .A1(n9960), .A2(n9957), .B1(n6790), .B2(n9958), .ZN(
        P2_U3529) );
  AOI22_X1 U11012 ( .A1(n9960), .A2(n9959), .B1(n6995), .B2(n9958), .ZN(
        P2_U3531) );
  NAND3_X1 U11013 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9963) );
  AND2_X1 U11014 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n9961) );
  NOR2_X1 U11015 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9961), .ZN(n9962) );
  INV_X1 U11016 ( .A(n9962), .ZN(n9979) );
  NAND2_X1 U11017 ( .A1(n9964), .A2(n9963), .ZN(n9978) );
  OAI222_X1 U11018 ( .A1(n9964), .A2(n9963), .B1(n9964), .B2(n9979), .C1(n9962), .C2(n9978), .ZN(ADD_1071_U5) );
  XOR2_X1 U11019 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  NOR2_X1 U11020 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n9965) );
  AOI21_X1 U11021 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9965), .ZN(n9984) );
  NOR2_X1 U11022 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n9966) );
  AOI21_X1 U11023 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9966), .ZN(n9987) );
  NOR2_X1 U11024 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n9967) );
  AOI21_X1 U11025 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9967), .ZN(n9990) );
  NOR2_X1 U11026 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9968) );
  AOI21_X1 U11027 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9968), .ZN(n9993) );
  NOR2_X1 U11028 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9969) );
  AOI21_X1 U11029 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9969), .ZN(n9996) );
  NOR2_X1 U11030 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9970) );
  AOI21_X1 U11031 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9970), .ZN(n9999) );
  NOR2_X1 U11032 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9971) );
  AOI21_X1 U11033 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9971), .ZN(n10002) );
  NOR2_X1 U11034 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9972) );
  AOI21_X1 U11035 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9972), .ZN(n10005) );
  NOR2_X1 U11036 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(P2_ADDR_REG_9__SCAN_IN), 
        .ZN(n9973) );
  AOI21_X1 U11037 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n9973), .ZN(n10386) );
  NOR2_X1 U11038 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(P2_ADDR_REG_8__SCAN_IN), 
        .ZN(n9974) );
  AOI21_X1 U11039 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n9974), .ZN(n10401) );
  NOR2_X1 U11040 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n9975) );
  AOI21_X1 U11041 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n9975), .ZN(n10389) );
  NOR2_X1 U11042 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n9976) );
  AOI21_X1 U11043 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n9976), .ZN(n10404) );
  NOR2_X1 U11044 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n9977) );
  AOI21_X1 U11045 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n9977), .ZN(n10395) );
  NAND2_X1 U11046 ( .A1(n9979), .A2(n9978), .ZN(n10392) );
  NAND2_X1 U11047 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9980) );
  OAI21_X1 U11048 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n9980), .ZN(n10391) );
  NOR2_X1 U11049 ( .A1(n10392), .A2(n10391), .ZN(n10390) );
  AOI21_X1 U11050 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10390), .ZN(n10407) );
  NAND2_X1 U11051 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9981) );
  OAI21_X1 U11052 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n9981), .ZN(n10406) );
  NOR2_X1 U11053 ( .A1(n10407), .A2(n10406), .ZN(n10405) );
  AOI21_X1 U11054 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10405), .ZN(n10410) );
  NOR2_X1 U11055 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9982) );
  AOI21_X1 U11056 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n9982), .ZN(n10409) );
  NAND2_X1 U11057 ( .A1(n10410), .A2(n10409), .ZN(n10408) );
  OAI21_X1 U11058 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10408), .ZN(n10394) );
  NAND2_X1 U11059 ( .A1(n10395), .A2(n10394), .ZN(n10393) );
  OAI21_X1 U11060 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10393), .ZN(n10403) );
  NAND2_X1 U11061 ( .A1(n10404), .A2(n10403), .ZN(n10402) );
  OAI21_X1 U11062 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10402), .ZN(n10388) );
  NAND2_X1 U11063 ( .A1(n10389), .A2(n10388), .ZN(n10387) );
  OAI21_X1 U11064 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10387), .ZN(n10400) );
  NAND2_X1 U11065 ( .A1(n10401), .A2(n10400), .ZN(n10399) );
  OAI21_X1 U11066 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10399), .ZN(n10385) );
  NAND2_X1 U11067 ( .A1(n10386), .A2(n10385), .ZN(n10384) );
  OAI21_X1 U11068 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10384), .ZN(n10004) );
  NAND2_X1 U11069 ( .A1(n10005), .A2(n10004), .ZN(n10003) );
  OAI21_X1 U11070 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10003), .ZN(n10001) );
  NAND2_X1 U11071 ( .A1(n10002), .A2(n10001), .ZN(n10000) );
  OAI21_X1 U11072 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10000), .ZN(n9998) );
  NAND2_X1 U11073 ( .A1(n9999), .A2(n9998), .ZN(n9997) );
  OAI21_X1 U11074 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9997), .ZN(n9995) );
  NAND2_X1 U11075 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  OAI21_X1 U11076 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9994), .ZN(n9992) );
  NAND2_X1 U11077 ( .A1(n9993), .A2(n9992), .ZN(n9991) );
  OAI21_X1 U11078 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9991), .ZN(n9989) );
  NAND2_X1 U11079 ( .A1(n9990), .A2(n9989), .ZN(n9988) );
  OAI21_X1 U11080 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9988), .ZN(n9986) );
  NAND2_X1 U11081 ( .A1(n9987), .A2(n9986), .ZN(n9985) );
  OAI21_X1 U11082 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9985), .ZN(n9983) );
  NAND2_X1 U11083 ( .A1(n9984), .A2(n9983), .ZN(n10007) );
  OAI21_X1 U11084 ( .B1(n9984), .B2(n9983), .A(n10007), .ZN(ADD_1071_U56) );
  OAI21_X1 U11085 ( .B1(n9987), .B2(n9986), .A(n9985), .ZN(ADD_1071_U57) );
  OAI21_X1 U11086 ( .B1(n9990), .B2(n9989), .A(n9988), .ZN(ADD_1071_U58) );
  OAI21_X1 U11087 ( .B1(n9993), .B2(n9992), .A(n9991), .ZN(ADD_1071_U59) );
  OAI21_X1 U11088 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(ADD_1071_U60) );
  OAI21_X1 U11089 ( .B1(n9999), .B2(n9998), .A(n9997), .ZN(ADD_1071_U61) );
  OAI21_X1 U11090 ( .B1(n10002), .B2(n10001), .A(n10000), .ZN(ADD_1071_U62) );
  OAI21_X1 U11091 ( .B1(n10005), .B2(n10004), .A(n10003), .ZN(ADD_1071_U63) );
  NOR2_X1 U11092 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(P2_ADDR_REG_18__SCAN_IN), 
        .ZN(n10006) );
  AOI21_X1 U11093 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10006), .ZN(n10398) );
  OAI21_X1 U11094 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10007), .ZN(n10397) );
  NAND2_X1 U11095 ( .A1(n10398), .A2(n10397), .ZN(n10396) );
  OAI21_X1 U11096 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n10396), .ZN(n10383) );
  XNOR2_X1 U11097 ( .A(n6342), .B(keyinput_g123), .ZN(n10014) );
  AOI22_X1 U11098 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(
        SI_18_), .B2(keyinput_g14), .ZN(n10008) );
  OAI221_X1 U11099 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        SI_18_), .C2(keyinput_g14), .A(n10008), .ZN(n10013) );
  AOI22_X1 U11100 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        SI_17_), .B2(keyinput_g15), .ZN(n10009) );
  OAI221_X1 U11101 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        SI_17_), .C2(keyinput_g15), .A(n10009), .ZN(n10012) );
  AOI22_X1 U11102 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_g58), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n10010) );
  OAI221_X1 U11103 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n10010), .ZN(n10011)
         );
  NOR4_X1 U11104 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10042) );
  AOI22_X1 U11105 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(
        SI_20_), .B2(keyinput_g12), .ZN(n10015) );
  OAI221_X1 U11106 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .C1(
        SI_20_), .C2(keyinput_g12), .A(n10015), .ZN(n10022) );
  AOI22_X1 U11107 ( .A1(SI_4_), .A2(keyinput_g28), .B1(P1_IR_REG_1__SCAN_IN), 
        .B2(keyinput_g92), .ZN(n10016) );
  OAI221_X1 U11108 ( .B1(SI_4_), .B2(keyinput_g28), .C1(P1_IR_REG_1__SCAN_IN), 
        .C2(keyinput_g92), .A(n10016), .ZN(n10021) );
  AOI22_X1 U11109 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_g120), .B1(SI_15_), .B2(keyinput_g17), .ZN(n10017) );
  OAI221_X1 U11110 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_g120), .C1(
        SI_15_), .C2(keyinput_g17), .A(n10017), .ZN(n10020) );
  AOI22_X1 U11111 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        P1_IR_REG_8__SCAN_IN), .B2(keyinput_g99), .ZN(n10018) );
  OAI221_X1 U11112 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_g99), .A(n10018), .ZN(n10019) );
  NOR4_X1 U11113 ( .A1(n10022), .A2(n10021), .A3(n10020), .A4(n10019), .ZN(
        n10041) );
  AOI22_X1 U11114 ( .A1(SI_16_), .A2(keyinput_g16), .B1(P1_D_REG_4__SCAN_IN), 
        .B2(keyinput_g127), .ZN(n10023) );
  OAI221_X1 U11115 ( .B1(SI_16_), .B2(keyinput_g16), .C1(P1_D_REG_4__SCAN_IN), 
        .C2(keyinput_g127), .A(n10023), .ZN(n10030) );
  AOI22_X1 U11116 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_g55), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput_g93), .ZN(n10024) );
  OAI221_X1 U11117 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .C1(
        P1_IR_REG_2__SCAN_IN), .C2(keyinput_g93), .A(n10024), .ZN(n10029) );
  AOI22_X1 U11118 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput_g75), .B1(
        P1_IR_REG_24__SCAN_IN), .B2(keyinput_g115), .ZN(n10025) );
  OAI221_X1 U11119 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .C1(
        P1_IR_REG_24__SCAN_IN), .C2(keyinput_g115), .A(n10025), .ZN(n10028) );
  AOI22_X1 U11120 ( .A1(SI_31_), .A2(keyinput_g1), .B1(SI_10_), .B2(
        keyinput_g22), .ZN(n10026) );
  OAI221_X1 U11121 ( .B1(SI_31_), .B2(keyinput_g1), .C1(SI_10_), .C2(
        keyinput_g22), .A(n10026), .ZN(n10027) );
  NOR4_X1 U11122 ( .A1(n10030), .A2(n10029), .A3(n10028), .A4(n10027), .ZN(
        n10040) );
  AOI22_X1 U11123 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .ZN(n10031) );
  OAI221_X1 U11124 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P2_DATAO_REG_10__SCAN_IN), .C2(keyinput_g86), .A(n10031), .ZN(n10038)
         );
  AOI22_X1 U11125 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_g121), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .ZN(n10032) );
  OAI221_X1 U11126 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_g121), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput_g84), .A(n10032), .ZN(n10037)
         );
  AOI22_X1 U11127 ( .A1(SI_2_), .A2(keyinput_g30), .B1(P1_IR_REG_27__SCAN_IN), 
        .B2(keyinput_g118), .ZN(n10033) );
  OAI221_X1 U11128 ( .B1(SI_2_), .B2(keyinput_g30), .C1(P1_IR_REG_27__SCAN_IN), 
        .C2(keyinput_g118), .A(n10033), .ZN(n10036) );
  AOI22_X1 U11129 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_g95), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_g107), .ZN(n10034) );
  OAI221_X1 U11130 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_g95), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_g107), .A(n10034), .ZN(n10035) );
  NOR4_X1 U11131 ( .A1(n10038), .A2(n10037), .A3(n10036), .A4(n10035), .ZN(
        n10039) );
  NAND4_X1 U11132 ( .A1(n10042), .A2(n10041), .A3(n10040), .A4(n10039), .ZN(
        n10190) );
  AOI22_X1 U11133 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_g94), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_g101), .ZN(n10043) );
  OAI221_X1 U11134 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_g94), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_g101), .A(n10043), .ZN(n10050) );
  AOI22_X1 U11135 ( .A1(SI_21_), .A2(keyinput_g11), .B1(SI_23_), .B2(
        keyinput_g9), .ZN(n10044) );
  OAI221_X1 U11136 ( .B1(SI_21_), .B2(keyinput_g11), .C1(SI_23_), .C2(
        keyinput_g9), .A(n10044), .ZN(n10049) );
  AOI22_X1 U11137 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(keyinput_g76), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_g73), .ZN(n10045) );
  OAI221_X1 U11138 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .C1(
        P2_DATAO_REG_23__SCAN_IN), .C2(keyinput_g73), .A(n10045), .ZN(n10048)
         );
  AOI22_X1 U11139 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_g34), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput_g102), .ZN(n10046) );
  OAI221_X1 U11140 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_g102), .A(n10046), .ZN(n10047) );
  NOR4_X1 U11141 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        n10080) );
  AOI22_X1 U11142 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(keyinput_g90), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .ZN(n10051) );
  OAI221_X1 U11143 ( .B1(P2_DATAO_REG_6__SCAN_IN), .B2(keyinput_g90), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput_g88), .A(n10051), .ZN(n10058)
         );
  AOI22_X1 U11144 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_g67), .B1(
        SI_3_), .B2(keyinput_g29), .ZN(n10052) );
  OAI221_X1 U11145 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_g67), .C1(
        SI_3_), .C2(keyinput_g29), .A(n10052), .ZN(n10057) );
  AOI22_X1 U11146 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput_g82), .B1(
        SI_22_), .B2(keyinput_g10), .ZN(n10053) );
  OAI221_X1 U11147 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .C1(
        SI_22_), .C2(keyinput_g10), .A(n10053), .ZN(n10056) );
  AOI22_X1 U11148 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_g77), .ZN(n10054) );
  OAI221_X1 U11149 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput_g77), .A(n10054), .ZN(n10055)
         );
  NOR4_X1 U11150 ( .A1(n10058), .A2(n10057), .A3(n10056), .A4(n10055), .ZN(
        n10079) );
  AOI22_X1 U11151 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_g96), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput_g106), .ZN(n10059) );
  OAI221_X1 U11152 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_g96), .C1(
        P1_IR_REG_15__SCAN_IN), .C2(keyinput_g106), .A(n10059), .ZN(n10066) );
  AOI22_X1 U11153 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_g53), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput_g125), .ZN(n10060) );
  OAI221_X1 U11154 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_g53), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput_g125), .A(n10060), .ZN(n10065) );
  AOI22_X1 U11155 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n10061) );
  OAI221_X1 U11156 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n10061), .ZN(n10064)
         );
  AOI22_X1 U11157 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput_g104), .ZN(n10062) );
  OAI221_X1 U11158 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput_g104), .A(n10062), .ZN(n10063) );
  NOR4_X1 U11159 ( .A1(n10066), .A2(n10065), .A3(n10064), .A4(n10063), .ZN(
        n10078) );
  AOI22_X1 U11160 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .ZN(n10067) );
  OAI221_X1 U11161 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        P2_DATAO_REG_9__SCAN_IN), .C2(keyinput_g87), .A(n10067), .ZN(n10076)
         );
  AOI22_X1 U11162 ( .A1(SI_9_), .A2(keyinput_g23), .B1(SI_24_), .B2(
        keyinput_g8), .ZN(n10068) );
  OAI221_X1 U11163 ( .B1(SI_9_), .B2(keyinput_g23), .C1(SI_24_), .C2(
        keyinput_g8), .A(n10068), .ZN(n10075) );
  AOI22_X1 U11164 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_g41), .B1(
        P1_IR_REG_26__SCAN_IN), .B2(keyinput_g117), .ZN(n10069) );
  OAI221_X1 U11165 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .C1(
        P1_IR_REG_26__SCAN_IN), .C2(keyinput_g117), .A(n10069), .ZN(n10074) );
  AOI22_X1 U11166 ( .A1(n10072), .A2(keyinput_g114), .B1(keyinput_g13), .B2(
        n10071), .ZN(n10070) );
  OAI221_X1 U11167 ( .B1(n10072), .B2(keyinput_g114), .C1(n10071), .C2(
        keyinput_g13), .A(n10070), .ZN(n10073) );
  NOR4_X1 U11168 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(
        n10077) );
  NAND4_X1 U11169 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n10189) );
  AOI22_X1 U11170 ( .A1(n10083), .A2(keyinput_g65), .B1(n10082), .B2(
        keyinput_g126), .ZN(n10081) );
  OAI221_X1 U11171 ( .B1(n10083), .B2(keyinput_g65), .C1(n10082), .C2(
        keyinput_g126), .A(n10081), .ZN(n10092) );
  INV_X1 U11172 ( .A(SI_6_), .ZN(n10085) );
  AOI22_X1 U11173 ( .A1(n5142), .A2(keyinput_g49), .B1(n10085), .B2(
        keyinput_g26), .ZN(n10084) );
  OAI221_X1 U11174 ( .B1(n5142), .B2(keyinput_g49), .C1(n10085), .C2(
        keyinput_g26), .A(n10084), .ZN(n10091) );
  XNOR2_X1 U11175 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_g91), .ZN(n10089) );
  XNOR2_X1 U11176 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_g111), .ZN(n10088)
         );
  XNOR2_X1 U11177 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g97), .ZN(n10087) );
  XNOR2_X1 U11178 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_g51), .ZN(n10086)
         );
  NAND4_X1 U11179 ( .A1(n10089), .A2(n10088), .A3(n10087), .A4(n10086), .ZN(
        n10090) );
  NOR3_X1 U11180 ( .A1(n10092), .A2(n10091), .A3(n10090), .ZN(n10135) );
  AOI22_X1 U11181 ( .A1(n10244), .A2(keyinput_g69), .B1(n6354), .B2(
        keyinput_g124), .ZN(n10093) );
  OAI221_X1 U11182 ( .B1(n10244), .B2(keyinput_g69), .C1(n6354), .C2(
        keyinput_g124), .A(n10093), .ZN(n10104) );
  AOI22_X1 U11183 ( .A1(n10095), .A2(keyinput_g6), .B1(keyinput_g43), .B2(
        n10318), .ZN(n10094) );
  OAI221_X1 U11184 ( .B1(n10095), .B2(keyinput_g6), .C1(n10318), .C2(
        keyinput_g43), .A(n10094), .ZN(n10103) );
  INV_X1 U11185 ( .A(SI_30_), .ZN(n10098) );
  AOI22_X1 U11186 ( .A1(n10098), .A2(keyinput_g2), .B1(n10097), .B2(
        keyinput_g81), .ZN(n10096) );
  OAI221_X1 U11187 ( .B1(n10098), .B2(keyinput_g2), .C1(n10097), .C2(
        keyinput_g81), .A(n10096), .ZN(n10102) );
  XOR2_X1 U11188 ( .A(n5183), .B(keyinput_g35), .Z(n10100) );
  XNOR2_X1 U11189 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_g112), .ZN(n10099)
         );
  NAND2_X1 U11190 ( .A1(n10100), .A2(n10099), .ZN(n10101) );
  NOR4_X1 U11191 ( .A1(n10104), .A2(n10103), .A3(n10102), .A4(n10101), .ZN(
        n10134) );
  AOI22_X1 U11192 ( .A1(n10107), .A2(keyinput_g80), .B1(n10106), .B2(
        keyinput_g5), .ZN(n10105) );
  OAI221_X1 U11193 ( .B1(n10107), .B2(keyinput_g80), .C1(n10106), .C2(
        keyinput_g5), .A(n10105), .ZN(n10118) );
  AOI22_X1 U11194 ( .A1(n10110), .A2(keyinput_g7), .B1(keyinput_g72), .B2(
        n10109), .ZN(n10108) );
  OAI221_X1 U11195 ( .B1(n10110), .B2(keyinput_g7), .C1(n10109), .C2(
        keyinput_g72), .A(n10108), .ZN(n10117) );
  AOI22_X1 U11196 ( .A1(n10113), .A2(keyinput_g18), .B1(keyinput_g39), .B2(
        n10112), .ZN(n10111) );
  OAI221_X1 U11197 ( .B1(n10113), .B2(keyinput_g18), .C1(n10112), .C2(
        keyinput_g39), .A(n10111), .ZN(n10116) );
  AOI22_X1 U11198 ( .A1(n10234), .A2(keyinput_g100), .B1(keyinput_g33), .B2(
        n4858), .ZN(n10114) );
  OAI221_X1 U11199 ( .B1(n10234), .B2(keyinput_g100), .C1(n4858), .C2(
        keyinput_g33), .A(n10114), .ZN(n10115) );
  NOR4_X1 U11200 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10133) );
  AOI22_X1 U11201 ( .A1(n10120), .A2(keyinput_g44), .B1(n5603), .B2(
        keyinput_g47), .ZN(n10119) );
  OAI221_X1 U11202 ( .B1(n10120), .B2(keyinput_g44), .C1(n5603), .C2(
        keyinput_g47), .A(n10119), .ZN(n10131) );
  AOI22_X1 U11203 ( .A1(n10301), .A2(keyinput_g71), .B1(keyinput_g74), .B2(
        n10122), .ZN(n10121) );
  OAI221_X1 U11204 ( .B1(n10301), .B2(keyinput_g71), .C1(n10122), .C2(
        keyinput_g74), .A(n10121), .ZN(n10130) );
  AOI22_X1 U11205 ( .A1(n10125), .A2(keyinput_g21), .B1(n10124), .B2(
        keyinput_g70), .ZN(n10123) );
  OAI221_X1 U11206 ( .B1(n10125), .B2(keyinput_g21), .C1(n10124), .C2(
        keyinput_g70), .A(n10123), .ZN(n10129) );
  XNOR2_X1 U11207 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_g108), .ZN(n10127)
         );
  XNOR2_X1 U11208 ( .A(SI_0_), .B(keyinput_g32), .ZN(n10126) );
  NAND2_X1 U11209 ( .A1(n10127), .A2(n10126), .ZN(n10128) );
  NOR4_X1 U11210 ( .A1(n10131), .A2(n10130), .A3(n10129), .A4(n10128), .ZN(
        n10132) );
  NAND4_X1 U11211 ( .A1(n10135), .A2(n10134), .A3(n10133), .A4(n10132), .ZN(
        n10188) );
  INV_X1 U11212 ( .A(SI_13_), .ZN(n10303) );
  AOI22_X1 U11213 ( .A1(n10288), .A2(keyinput_g62), .B1(n10303), .B2(
        keyinput_g19), .ZN(n10136) );
  OAI221_X1 U11214 ( .B1(n10288), .B2(keyinput_g62), .C1(n10303), .C2(
        keyinput_g19), .A(n10136), .ZN(n10144) );
  XOR2_X1 U11215 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_g119), .Z(n10143) );
  XNOR2_X1 U11216 ( .A(keyinput_g40), .B(n10300), .ZN(n10142) );
  XNOR2_X1 U11217 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_g79), .ZN(n10140) );
  XNOR2_X1 U11218 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_g110), .ZN(n10139)
         );
  XNOR2_X1 U11219 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_g89), .ZN(n10138)
         );
  XNOR2_X1 U11220 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_g109), .ZN(n10137)
         );
  NAND4_X1 U11221 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n10141) );
  NOR4_X1 U11222 ( .A1(n10144), .A2(n10143), .A3(n10142), .A4(n10141), .ZN(
        n10186) );
  AOI22_X1 U11223 ( .A1(n10146), .A2(keyinput_g66), .B1(n8181), .B2(
        keyinput_g50), .ZN(n10145) );
  OAI221_X1 U11224 ( .B1(n10146), .B2(keyinput_g66), .C1(n8181), .C2(
        keyinput_g50), .A(n10145), .ZN(n10156) );
  AOI22_X1 U11225 ( .A1(n10149), .A2(keyinput_g78), .B1(keyinput_g64), .B2(
        n10148), .ZN(n10147) );
  OAI221_X1 U11226 ( .B1(n10149), .B2(keyinput_g78), .C1(n10148), .C2(
        keyinput_g64), .A(n10147), .ZN(n10155) );
  XOR2_X1 U11227 ( .A(n5577), .B(keyinput_g38), .Z(n10153) );
  XNOR2_X1 U11228 ( .A(SI_8_), .B(keyinput_g24), .ZN(n10152) );
  XNOR2_X1 U11229 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_g103), .ZN(n10151)
         );
  XNOR2_X1 U11230 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10150) );
  NAND4_X1 U11231 ( .A1(n10153), .A2(n10152), .A3(n10151), .A4(n10150), .ZN(
        n10154) );
  NOR3_X1 U11232 ( .A1(n10156), .A2(n10155), .A3(n10154), .ZN(n10185) );
  AOI22_X1 U11233 ( .A1(n10159), .A2(keyinput_g20), .B1(keyinput_g85), .B2(
        n10158), .ZN(n10157) );
  OAI221_X1 U11234 ( .B1(n10159), .B2(keyinput_g20), .C1(n10158), .C2(
        keyinput_g85), .A(n10157), .ZN(n10168) );
  AOI22_X1 U11235 ( .A1(n10161), .A2(keyinput_g27), .B1(keyinput_g59), .B2(
        n10319), .ZN(n10160) );
  OAI221_X1 U11236 ( .B1(n10161), .B2(keyinput_g27), .C1(n10319), .C2(
        keyinput_g59), .A(n10160), .ZN(n10167) );
  XNOR2_X1 U11237 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g98), .ZN(n10165) );
  XNOR2_X1 U11238 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_g116), .ZN(n10164)
         );
  XNOR2_X1 U11239 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_g122), .ZN(n10163)
         );
  XNOR2_X1 U11240 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_g61), .ZN(n10162)
         );
  NAND4_X1 U11241 ( .A1(n10165), .A2(n10164), .A3(n10163), .A4(n10162), .ZN(
        n10166) );
  NOR3_X1 U11242 ( .A1(n10168), .A2(n10167), .A3(n10166), .ZN(n10184) );
  AOI22_X1 U11243 ( .A1(n6465), .A2(keyinput_g4), .B1(keyinput_g52), .B2(
        n10170), .ZN(n10169) );
  OAI221_X1 U11244 ( .B1(n6465), .B2(keyinput_g4), .C1(n10170), .C2(
        keyinput_g52), .A(n10169), .ZN(n10182) );
  AOI22_X1 U11245 ( .A1(n10173), .A2(keyinput_g68), .B1(keyinput_g3), .B2(
        n10172), .ZN(n10171) );
  OAI221_X1 U11246 ( .B1(n10173), .B2(keyinput_g68), .C1(n10172), .C2(
        keyinput_g3), .A(n10171), .ZN(n10181) );
  AOI22_X1 U11247 ( .A1(n10176), .A2(keyinput_g45), .B1(n10175), .B2(
        keyinput_g25), .ZN(n10174) );
  OAI221_X1 U11248 ( .B1(n10176), .B2(keyinput_g45), .C1(n10175), .C2(
        keyinput_g25), .A(n10174), .ZN(n10180) );
  XNOR2_X1 U11249 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_g113), .ZN(n10178)
         );
  XNOR2_X1 U11250 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_g83), .ZN(n10177) );
  NAND2_X1 U11251 ( .A1(n10178), .A2(n10177), .ZN(n10179) );
  NOR4_X1 U11252 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10183) );
  NAND4_X1 U11253 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n10187) );
  NOR4_X1 U11254 ( .A1(n10190), .A2(n10189), .A3(n10188), .A4(n10187), .ZN(
        n10377) );
  OAI22_X1 U11255 ( .A1(SI_10_), .A2(keyinput_f22), .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .ZN(n10191) );
  AOI221_X1 U11256 ( .B1(SI_10_), .B2(keyinput_f22), .C1(keyinput_f35), .C2(
        P2_REG3_REG_7__SCAN_IN), .A(n10191), .ZN(n10198) );
  OAI22_X1 U11257 ( .A1(SI_26_), .A2(keyinput_f6), .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n10192) );
  AOI221_X1 U11258 ( .B1(SI_26_), .B2(keyinput_f6), .C1(keyinput_f39), .C2(
        P2_REG3_REG_10__SCAN_IN), .A(n10192), .ZN(n10197) );
  OAI22_X1 U11259 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_f125), .B1(SI_15_), 
        .B2(keyinput_f17), .ZN(n10193) );
  AOI221_X1 U11260 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_f125), .C1(
        keyinput_f17), .C2(SI_15_), .A(n10193), .ZN(n10196) );
  OAI22_X1 U11261 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_f124), .B1(
        keyinput_f65), .B2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10194) );
  AOI221_X1 U11262 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_f124), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput_f65), .A(n10194), .ZN(n10195)
         );
  NAND4_X1 U11263 ( .A1(n10198), .A2(n10197), .A3(n10196), .A4(n10195), .ZN(
        n10336) );
  AOI22_X1 U11264 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput_f109), .ZN(n10199) );
  OAI221_X1 U11265 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput_f109), .A(n10199), .ZN(n10206) );
  AOI22_X1 U11266 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_f85), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput_f106), .ZN(n10200) );
  OAI221_X1 U11267 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_f85), .C1(
        P1_IR_REG_15__SCAN_IN), .C2(keyinput_f106), .A(n10200), .ZN(n10205) );
  AOI22_X1 U11268 ( .A1(SI_28_), .A2(keyinput_f4), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_f73), .ZN(n10201) );
  OAI221_X1 U11269 ( .B1(SI_28_), .B2(keyinput_f4), .C1(
        P2_DATAO_REG_23__SCAN_IN), .C2(keyinput_f73), .A(n10201), .ZN(n10204)
         );
  AOI22_X1 U11270 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_f87), .B1(
        SI_25_), .B2(keyinput_f7), .ZN(n10202) );
  OAI221_X1 U11271 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .C1(
        SI_25_), .C2(keyinput_f7), .A(n10202), .ZN(n10203) );
  NOR4_X1 U11272 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10224) );
  AOI22_X1 U11273 ( .A1(SI_7_), .A2(keyinput_f25), .B1(P1_IR_REG_20__SCAN_IN), 
        .B2(keyinput_f111), .ZN(n10207) );
  OAI221_X1 U11274 ( .B1(SI_7_), .B2(keyinput_f25), .C1(P1_IR_REG_20__SCAN_IN), 
        .C2(keyinput_f111), .A(n10207), .ZN(n10214) );
  AOI22_X1 U11275 ( .A1(SI_14_), .A2(keyinput_f18), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_f79), .ZN(n10208) );
  OAI221_X1 U11276 ( .B1(SI_14_), .B2(keyinput_f18), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput_f79), .A(n10208), .ZN(n10213)
         );
  AOI22_X1 U11277 ( .A1(SI_31_), .A2(keyinput_f1), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_f77), .ZN(n10209) );
  OAI221_X1 U11278 ( .B1(SI_31_), .B2(keyinput_f1), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput_f77), .A(n10209), .ZN(n10212)
         );
  AOI22_X1 U11279 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_f66), .B1(
        SI_0_), .B2(keyinput_f32), .ZN(n10210) );
  OAI221_X1 U11280 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .C1(
        SI_0_), .C2(keyinput_f32), .A(n10210), .ZN(n10211) );
  NOR4_X1 U11281 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10223) );
  OAI22_X1 U11282 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f104), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_f96), .ZN(n10215) );
  AOI221_X1 U11283 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f104), .C1(
        keyinput_f96), .C2(P1_IR_REG_5__SCAN_IN), .A(n10215), .ZN(n10221) );
  OAI22_X1 U11284 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_f112), .B1(
        keyinput_f26), .B2(SI_6_), .ZN(n10216) );
  AOI221_X1 U11285 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_f112), .C1(SI_6_), .C2(keyinput_f26), .A(n10216), .ZN(n10220) );
  OAI22_X1 U11286 ( .A1(SI_11_), .A2(keyinput_f21), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_f86), .ZN(n10217) );
  AOI221_X1 U11287 ( .B1(SI_11_), .B2(keyinput_f21), .C1(keyinput_f86), .C2(
        P2_DATAO_REG_10__SCAN_IN), .A(n10217), .ZN(n10219) );
  XNOR2_X1 U11288 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_f122), .ZN(n10218)
         );
  AND4_X1 U11289 ( .A1(n10221), .A2(n10220), .A3(n10219), .A4(n10218), .ZN(
        n10222) );
  NAND3_X1 U11290 ( .A1(n10224), .A2(n10223), .A3(n10222), .ZN(n10335) );
  AOI22_X1 U11291 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_f89), .ZN(n10225) );
  OAI221_X1 U11292 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput_f89), .A(n10225), .ZN(n10232)
         );
  AOI22_X1 U11293 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_f72), .ZN(n10226) );
  OAI221_X1 U11294 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput_f72), .A(n10226), .ZN(n10231)
         );
  AOI22_X1 U11295 ( .A1(SI_29_), .A2(keyinput_f3), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_f75), .ZN(n10227) );
  OAI221_X1 U11296 ( .B1(SI_29_), .B2(keyinput_f3), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n10227), .ZN(n10230)
         );
  AOI22_X1 U11297 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_f63), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n10228) );
  OAI221_X1 U11298 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n10228), .ZN(n10229)
         );
  NOR4_X1 U11299 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(n10229), .ZN(
        n10271) );
  AOI22_X1 U11300 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_f50), .B1(
        n10234), .B2(keyinput_f100), .ZN(n10233) );
  OAI221_X1 U11301 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .C1(
        n10234), .C2(keyinput_f100), .A(n10233), .ZN(n10242) );
  AOI22_X1 U11302 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_f52), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .ZN(n10235) );
  OAI221_X1 U11303 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_f80), .A(n10235), .ZN(n10241)
         );
  XNOR2_X1 U11304 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_f48), .ZN(n10239)
         );
  XNOR2_X1 U11305 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_f103), .ZN(n10238)
         );
  XNOR2_X1 U11306 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_f119), .ZN(n10237)
         );
  XNOR2_X1 U11307 ( .A(SI_8_), .B(keyinput_f24), .ZN(n10236) );
  NAND4_X1 U11308 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10240) );
  NOR3_X1 U11309 ( .A1(n10242), .A2(n10241), .A3(n10240), .ZN(n10270) );
  AOI22_X1 U11310 ( .A1(n10245), .A2(keyinput_f127), .B1(keyinput_f69), .B2(
        n10244), .ZN(n10243) );
  OAI221_X1 U11311 ( .B1(n10245), .B2(keyinput_f127), .C1(n10244), .C2(
        keyinput_f69), .A(n10243), .ZN(n10253) );
  XOR2_X1 U11312 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_f117), .Z(n10252) );
  XNOR2_X1 U11313 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_f120), .ZN(n10249)
         );
  XNOR2_X1 U11314 ( .A(SI_17_), .B(keyinput_f15), .ZN(n10248) );
  XNOR2_X1 U11315 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_f60), .ZN(n10247)
         );
  XNOR2_X1 U11316 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_f93), .ZN(n10246) );
  NAND4_X1 U11317 ( .A1(n10249), .A2(n10248), .A3(n10247), .A4(n10246), .ZN(
        n10251) );
  XNOR2_X1 U11318 ( .A(keyinput_f123), .B(n6342), .ZN(n10250) );
  NOR4_X1 U11319 ( .A1(n10253), .A2(n10252), .A3(n10251), .A4(n10250), .ZN(
        n10269) );
  AOI22_X1 U11320 ( .A1(n4858), .A2(keyinput_f33), .B1(keyinput_f36), .B2(
        n10255), .ZN(n10254) );
  OAI221_X1 U11321 ( .B1(n4858), .B2(keyinput_f33), .C1(n10255), .C2(
        keyinput_f36), .A(n10254), .ZN(n10267) );
  INV_X1 U11322 ( .A(SI_21_), .ZN(n10258) );
  AOI22_X1 U11323 ( .A1(n10258), .A2(keyinput_f11), .B1(keyinput_f46), .B2(
        n10257), .ZN(n10256) );
  OAI221_X1 U11324 ( .B1(n10258), .B2(keyinput_f11), .C1(n10257), .C2(
        keyinput_f46), .A(n10256), .ZN(n10266) );
  AOI22_X1 U11325 ( .A1(n10261), .A2(keyinput_f10), .B1(keyinput_f37), .B2(
        n10260), .ZN(n10259) );
  OAI221_X1 U11326 ( .B1(n10261), .B2(keyinput_f10), .C1(n10260), .C2(
        keyinput_f37), .A(n10259), .ZN(n10265) );
  XNOR2_X1 U11327 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_f110), .ZN(n10263)
         );
  XNOR2_X1 U11328 ( .A(SI_19_), .B(keyinput_f13), .ZN(n10262) );
  NAND2_X1 U11329 ( .A1(n10263), .A2(n10262), .ZN(n10264) );
  NOR4_X1 U11330 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10268) );
  NAND4_X1 U11331 ( .A1(n10271), .A2(n10270), .A3(n10269), .A4(n10268), .ZN(
        n10334) );
  AOI22_X1 U11332 ( .A1(n10274), .A2(keyinput_f8), .B1(keyinput_f54), .B2(
        n10273), .ZN(n10272) );
  OAI221_X1 U11333 ( .B1(n10274), .B2(keyinput_f8), .C1(n10273), .C2(
        keyinput_f54), .A(n10272), .ZN(n10278) );
  XOR2_X1 U11334 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_f68), .Z(n10277)
         );
  XNOR2_X1 U11335 ( .A(n10275), .B(keyinput_f91), .ZN(n10276) );
  NOR3_X1 U11336 ( .A1(n10278), .A2(n10277), .A3(n10276), .ZN(n10282) );
  XNOR2_X1 U11337 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_f107), .ZN(n10281)
         );
  XNOR2_X1 U11338 ( .A(SI_9_), .B(keyinput_f23), .ZN(n10280) );
  XNOR2_X1 U11339 ( .A(SI_1_), .B(keyinput_f31), .ZN(n10279) );
  NAND4_X1 U11340 ( .A1(n10282), .A2(n10281), .A3(n10280), .A4(n10279), .ZN(
        n10285) );
  XNOR2_X1 U11341 ( .A(n10283), .B(keyinput_f0), .ZN(n10284) );
  NOR2_X1 U11342 ( .A1(n10285), .A2(n10284), .ZN(n10332) );
  AOI22_X1 U11343 ( .A1(n10288), .A2(keyinput_f62), .B1(n10287), .B2(
        keyinput_f9), .ZN(n10286) );
  OAI221_X1 U11344 ( .B1(n10288), .B2(keyinput_f62), .C1(n10287), .C2(
        keyinput_f9), .A(n10286), .ZN(n10298) );
  XNOR2_X1 U11345 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_f98), .ZN(n10292) );
  XNOR2_X1 U11346 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_f88), .ZN(n10291)
         );
  XNOR2_X1 U11347 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_f115), .ZN(n10290)
         );
  XNOR2_X1 U11348 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_f74), .ZN(n10289) );
  NAND4_X1 U11349 ( .A1(n10292), .A2(n10291), .A3(n10290), .A4(n10289), .ZN(
        n10297) );
  XNOR2_X1 U11350 ( .A(n10293), .B(keyinput_f116), .ZN(n10296) );
  XNOR2_X1 U11351 ( .A(n10294), .B(keyinput_f108), .ZN(n10295) );
  NOR4_X1 U11352 ( .A1(n10298), .A2(n10297), .A3(n10296), .A4(n10295), .ZN(
        n10331) );
  AOI22_X1 U11353 ( .A1(n10301), .A2(keyinput_f71), .B1(keyinput_f40), .B2(
        n10300), .ZN(n10299) );
  OAI221_X1 U11354 ( .B1(n10301), .B2(keyinput_f71), .C1(n10300), .C2(
        keyinput_f40), .A(n10299), .ZN(n10313) );
  AOI22_X1 U11355 ( .A1(n10304), .A2(keyinput_f41), .B1(n10303), .B2(
        keyinput_f19), .ZN(n10302) );
  OAI221_X1 U11356 ( .B1(n10304), .B2(keyinput_f41), .C1(n10303), .C2(
        keyinput_f19), .A(n10302), .ZN(n10312) );
  AOI22_X1 U11357 ( .A1(n10307), .A2(keyinput_f28), .B1(n10306), .B2(
        keyinput_f12), .ZN(n10305) );
  OAI221_X1 U11358 ( .B1(n10307), .B2(keyinput_f28), .C1(n10306), .C2(
        keyinput_f12), .A(n10305), .ZN(n10311) );
  XNOR2_X1 U11359 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_f92), .ZN(n10309) );
  XNOR2_X1 U11360 ( .A(SI_5_), .B(keyinput_f27), .ZN(n10308) );
  NAND2_X1 U11361 ( .A1(n10309), .A2(n10308), .ZN(n10310) );
  NOR4_X1 U11362 ( .A1(n10313), .A2(n10312), .A3(n10311), .A4(n10310), .ZN(
        n10330) );
  AOI22_X1 U11363 ( .A1(n10316), .A2(keyinput_f82), .B1(keyinput_f51), .B2(
        n10315), .ZN(n10314) );
  OAI221_X1 U11364 ( .B1(n10316), .B2(keyinput_f82), .C1(n10315), .C2(
        keyinput_f51), .A(n10314), .ZN(n10328) );
  AOI22_X1 U11365 ( .A1(n10319), .A2(keyinput_f59), .B1(n10318), .B2(
        keyinput_f43), .ZN(n10317) );
  OAI221_X1 U11366 ( .B1(n10319), .B2(keyinput_f59), .C1(n10318), .C2(
        keyinput_f43), .A(n10317), .ZN(n10327) );
  AOI22_X1 U11367 ( .A1(n10321), .A2(keyinput_f83), .B1(keyinput_f42), .B2(
        n5655), .ZN(n10320) );
  OAI221_X1 U11368 ( .B1(n10321), .B2(keyinput_f83), .C1(n5655), .C2(
        keyinput_f42), .A(n10320), .ZN(n10326) );
  AOI22_X1 U11369 ( .A1(n10324), .A2(keyinput_f29), .B1(n10323), .B2(
        keyinput_f16), .ZN(n10322) );
  OAI221_X1 U11370 ( .B1(n10324), .B2(keyinput_f29), .C1(n10323), .C2(
        keyinput_f16), .A(n10322), .ZN(n10325) );
  NOR4_X1 U11371 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10329) );
  NAND4_X1 U11372 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10333) );
  NOR4_X1 U11373 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n10375) );
  OAI22_X1 U11374 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_f102), .B1(
        keyinput_f5), .B2(SI_27_), .ZN(n10337) );
  AOI221_X1 U11375 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_f102), .C1(
        SI_27_), .C2(keyinput_f5), .A(n10337), .ZN(n10344) );
  OAI22_X1 U11376 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_f113), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .ZN(n10338) );
  AOI221_X1 U11377 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_f113), .C1(
        keyinput_f56), .C2(P2_REG3_REG_13__SCAN_IN), .A(n10338), .ZN(n10343)
         );
  OAI22_X1 U11378 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(keyinput_f76), .B1(
        P1_IR_REG_30__SCAN_IN), .B2(keyinput_f121), .ZN(n10339) );
  AOI221_X1 U11379 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_f76), .C1(
        keyinput_f121), .C2(P1_IR_REG_30__SCAN_IN), .A(n10339), .ZN(n10342) );
  OAI22_X1 U11380 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_f99), .B1(
        keyinput_f57), .B2(P2_REG3_REG_22__SCAN_IN), .ZN(n10340) );
  AOI221_X1 U11381 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_f99), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n10340), .ZN(n10341)
         );
  NAND4_X1 U11382 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10372) );
  OAI22_X1 U11383 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        keyinput_f67), .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n10345) );
  AOI221_X1 U11384 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput_f67), .A(n10345), .ZN(n10352)
         );
  OAI22_X1 U11385 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput_f70), .B1(
        SI_12_), .B2(keyinput_f20), .ZN(n10346) );
  AOI221_X1 U11386 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_f70), .C1(
        keyinput_f20), .C2(SI_12_), .A(n10346), .ZN(n10351) );
  OAI22_X1 U11387 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_f126), .B1(
        keyinput_f49), .B2(P2_REG3_REG_5__SCAN_IN), .ZN(n10347) );
  AOI221_X1 U11388 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_f126), .C1(
        P2_REG3_REG_5__SCAN_IN), .C2(keyinput_f49), .A(n10347), .ZN(n10350) );
  OAI22_X1 U11389 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_f95), .B1(
        keyinput_f38), .B2(P2_REG3_REG_23__SCAN_IN), .ZN(n10348) );
  AOI221_X1 U11390 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_f95), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n10348), .ZN(n10349)
         );
  NAND4_X1 U11391 ( .A1(n10352), .A2(n10351), .A3(n10350), .A4(n10349), .ZN(
        n10371) );
  OAI22_X1 U11392 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput_f64), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n10353) );
  AOI221_X1 U11393 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput_f64), .C1(
        keyinput_f58), .C2(P2_REG3_REG_11__SCAN_IN), .A(n10353), .ZN(n10360)
         );
  OAI22_X1 U11394 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput_f78), .B1(
        keyinput_f90), .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n10354) );
  AOI221_X1 U11395 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_f78), .C1(
        P2_DATAO_REG_6__SCAN_IN), .C2(keyinput_f90), .A(n10354), .ZN(n10359)
         );
  OAI22_X1 U11396 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_f97), .B1(
        P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n10355) );
  AOI221_X1 U11397 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_f97), .C1(
        keyinput_f45), .C2(P2_REG3_REG_21__SCAN_IN), .A(n10355), .ZN(n10358)
         );
  OAI22_X1 U11398 ( .A1(SI_18_), .A2(keyinput_f14), .B1(keyinput_f84), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n10356) );
  AOI221_X1 U11399 ( .B1(SI_18_), .B2(keyinput_f14), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput_f84), .A(n10356), .ZN(n10357)
         );
  NAND4_X1 U11400 ( .A1(n10360), .A2(n10359), .A3(n10358), .A4(n10357), .ZN(
        n10370) );
  OAI22_X1 U11401 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_f114), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_f101), .ZN(n10361) );
  AOI221_X1 U11402 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_f114), .C1(
        keyinput_f101), .C2(P1_IR_REG_10__SCAN_IN), .A(n10361), .ZN(n10368) );
  OAI22_X1 U11403 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput_f81), .B1(
        SI_30_), .B2(keyinput_f2), .ZN(n10362) );
  AOI221_X1 U11404 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_f81), .C1(
        keyinput_f2), .C2(SI_30_), .A(n10362), .ZN(n10367) );
  OAI22_X1 U11405 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput_f118), .B1(
        keyinput_f30), .B2(SI_2_), .ZN(n10363) );
  AOI221_X1 U11406 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput_f118), .C1(SI_2_), .C2(keyinput_f30), .A(n10363), .ZN(n10366) );
  OAI22_X1 U11407 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_f94), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .ZN(n10364) );
  AOI221_X1 U11408 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_f94), .C1(
        keyinput_f34), .C2(P2_STATE_REG_SCAN_IN), .A(n10364), .ZN(n10365) );
  NAND4_X1 U11409 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10369) );
  NOR4_X1 U11410 ( .A1(n10372), .A2(n10371), .A3(n10370), .A4(n10369), .ZN(
        n10374) );
  NOR2_X1 U11411 ( .A1(n10379), .A2(keyinput_f105), .ZN(n10373) );
  AOI221_X1 U11412 ( .B1(n10375), .B2(n10374), .C1(keyinput_f105), .C2(n10379), 
        .A(n10373), .ZN(n10376) );
  AOI211_X1 U11413 ( .C1(keyinput_g105), .C2(n10379), .A(n10377), .B(n10376), 
        .ZN(n10378) );
  OAI21_X1 U11414 ( .B1(n10379), .B2(keyinput_g105), .A(n10378), .ZN(n10381)
         );
  XNOR2_X1 U11415 ( .A(n4856), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n10380) );
  XNOR2_X1 U11416 ( .A(n10381), .B(n10380), .ZN(n10382) );
  XNOR2_X1 U11417 ( .A(n10383), .B(n10382), .ZN(ADD_1071_U4) );
  OAI21_X1 U11418 ( .B1(n10386), .B2(n10385), .A(n10384), .ZN(ADD_1071_U47) );
  OAI21_X1 U11419 ( .B1(n10389), .B2(n10388), .A(n10387), .ZN(ADD_1071_U49) );
  AOI21_X1 U11420 ( .B1(n10392), .B2(n10391), .A(n10390), .ZN(ADD_1071_U54) );
  OAI21_X1 U11421 ( .B1(n10395), .B2(n10394), .A(n10393), .ZN(ADD_1071_U51) );
  OAI21_X1 U11422 ( .B1(n10398), .B2(n10397), .A(n10396), .ZN(ADD_1071_U55) );
  OAI21_X1 U11423 ( .B1(n10401), .B2(n10400), .A(n10399), .ZN(ADD_1071_U48) );
  OAI21_X1 U11424 ( .B1(n10404), .B2(n10403), .A(n10402), .ZN(ADD_1071_U50) );
  AOI21_X1 U11425 ( .B1(n10407), .B2(n10406), .A(n10405), .ZN(ADD_1071_U53) );
  OAI21_X1 U11426 ( .B1(n10410), .B2(n10409), .A(n10408), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4987 ( .A(n5163), .Z(n5658) );
  AND2_X1 U8029 ( .A1(n7991), .A2(n7992), .ZN(n7989) );
endmodule

