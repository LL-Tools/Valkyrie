

module b17_C_AntiSAT_k_128_7 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21259;

  AOI21_X1 U11096 ( .B1(n14669), .B2(n14668), .A(n14316), .ZN(n15060) );
  INV_X1 U11097 ( .A(n18935), .ZN(n18330) );
  INV_X1 U11098 ( .A(n17144), .ZN(n9942) );
  BUF_X1 U11099 ( .A(n10703), .Z(n10736) );
  OR2_X1 U11100 ( .A1(n11170), .A2(n13303), .ZN(n12105) );
  AND2_X1 U11101 ( .A1(n10408), .A2(n10389), .ZN(n10542) );
  AND2_X1 U11102 ( .A1(n10407), .A2(n10390), .ZN(n10540) );
  CLKBUF_X2 U11103 ( .A(n12249), .Z(n14205) );
  INV_X2 U11104 ( .A(n11086), .ZN(n11236) );
  INV_X4 U11105 ( .A(n12237), .ZN(n17406) );
  INV_X1 U11106 ( .A(n12367), .ZN(n17438) );
  INV_X1 U11107 ( .A(n14411), .ZN(n10604) );
  CLKBUF_X2 U11108 ( .A(n11061), .Z(n11791) );
  NAND2_X1 U11109 ( .A1(n10337), .A2(n10336), .ZN(n10344) );
  CLKBUF_X2 U11110 ( .A(n12225), .Z(n9658) );
  AND2_X1 U11111 ( .A1(n14440), .A2(n10419), .ZN(n14431) );
  INV_X1 U11112 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16267) );
  CLKBUF_X2 U11113 ( .A(n9672), .Z(n11215) );
  CLKBUF_X2 U11114 ( .A(n9662), .Z(n9686) );
  CLKBUF_X2 U11115 ( .A(n9666), .Z(n11861) );
  CLKBUF_X2 U11116 ( .A(n11220), .Z(n9690) );
  BUF_X2 U11117 ( .A(n19535), .Z(n9676) );
  INV_X1 U11119 ( .A(n11170), .ZN(n13310) );
  INV_X2 U11120 ( .A(n11168), .ZN(n20446) );
  NAND2_X1 U11121 ( .A1(n11016), .A2(n11015), .ZN(n11168) );
  NOR2_X2 U11122 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10418) );
  AND2_X1 U11123 ( .A1(n11009), .A2(n13570), .ZN(n11061) );
  AND2_X1 U11124 ( .A1(n11007), .A2(n9806), .ZN(n11220) );
  AND3_X2 U11126 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13219) );
  INV_X2 U11127 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11302) );
  CLKBUF_X1 U11128 ( .A(n21027), .Z(n9652) );
  NOR2_X1 U11129 ( .A1(n20982), .A2(n21059), .ZN(n21027) );
  INV_X1 U11132 ( .A(n14412), .ZN(n10607) );
  INV_X1 U11133 ( .A(n14417), .ZN(n10605) );
  CLKBUF_X2 U11134 ( .A(n11118), .Z(n11839) );
  INV_X1 U11135 ( .A(n20438), .ZN(n9954) );
  AND2_X1 U11136 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13570) );
  AND2_X1 U11137 ( .A1(n14440), .A2(n10418), .ZN(n14421) );
  INV_X1 U11138 ( .A(n10164), .ZN(n14404) );
  AND2_X1 U11139 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10431) );
  AND2_X1 U11140 ( .A1(n10038), .A2(n13642), .ZN(n11164) );
  NAND2_X1 U11141 ( .A1(n11164), .A2(n11113), .ZN(n11169) );
  AND2_X1 U11142 ( .A1(n20438), .A2(n20442), .ZN(n11172) );
  NAND2_X1 U11143 ( .A1(n11129), .A2(n11128), .ZN(n13303) );
  CLKBUF_X2 U11144 ( .A(n10310), .Z(n9663) );
  CLKBUF_X2 U11145 ( .A(n12537), .Z(n9657) );
  MUX2_X1 U11146 ( .A(n17801), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .S(
        n18038), .Z(n12301) );
  CLKBUF_X2 U11149 ( .A(n10695), .Z(n12963) );
  NOR2_X1 U11150 ( .A1(n15674), .A2(n15667), .ZN(n15658) );
  XNOR2_X1 U11152 ( .A(n14298), .B(n14297), .ZN(n19333) );
  NAND2_X1 U11153 ( .A1(n10823), .A2(n19286), .ZN(n10862) );
  AND2_X1 U11154 ( .A1(n9888), .A2(n18140), .ZN(n17773) );
  INV_X1 U11155 ( .A(n17933), .ZN(n18038) );
  INV_X1 U11157 ( .A(n20308), .ZN(n20335) );
  NAND4_X2 U11158 ( .A1(n11112), .A2(n11111), .A3(n11110), .A4(n11109), .ZN(
        n11165) );
  INV_X2 U11159 ( .A(n13637), .ZN(n11968) );
  INV_X1 U11160 ( .A(n20393), .ZN(n20407) );
  NOR2_X1 U11162 ( .A1(n16165), .A2(n15521), .ZN(n15520) );
  INV_X1 U11163 ( .A(n18125), .ZN(n18079) );
  INV_X1 U11164 ( .A(n18937), .ZN(n18921) );
  INV_X2 U11165 ( .A(n20339), .ZN(n20330) );
  INV_X1 U11166 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20963) );
  OR2_X1 U11167 ( .A1(n12179), .A2(n12181), .ZN(n9653) );
  AND2_X2 U11168 ( .A1(n9806), .A2(n13569), .ZN(n9654) );
  NAND2_X2 U11169 ( .A1(n11009), .A2(n11006), .ZN(n11885) );
  NOR3_X2 U11170 ( .A1(n17078), .A2(n17451), .A3(n17452), .ZN(n17418) );
  BUF_X1 U11171 ( .A(n14257), .Z(n9655) );
  OAI21_X2 U11172 ( .B1(n10370), .B2(n16575), .A(n10357), .ZN(n10363) );
  AND2_X1 U11173 ( .A1(n13303), .A2(n13637), .ZN(n13202) );
  AND2_X1 U11174 ( .A1(n9675), .A2(n20041), .ZN(n12537) );
  XNOR2_X2 U11175 ( .A(n10862), .B(n10824), .ZN(n14068) );
  XNOR2_X2 U11176 ( .A(n14522), .B(n10185), .ZN(n15544) );
  NAND2_X2 U11177 ( .A1(n15550), .A2(n14506), .ZN(n14522) );
  XNOR2_X2 U11178 ( .A(n9952), .B(n11232), .ZN(n11320) );
  OAI22_X2 U11179 ( .A1(n13223), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n13669), 
        .B2(n11334), .ZN(n11230) );
  NOR2_X1 U11180 ( .A1(n12177), .A2(n17176), .ZN(n12225) );
  NOR2_X2 U11182 ( .A1(n17900), .A2(n18038), .ZN(n17819) );
  OR2_X1 U11183 ( .A1(n15014), .A2(n15015), .ZN(n15118) );
  NAND2_X1 U11184 ( .A1(n14217), .A2(n9980), .ZN(n15197) );
  NAND2_X1 U11185 ( .A1(n14214), .A2(n14213), .ZN(n14217) );
  NAND2_X1 U11186 ( .A1(n10861), .A2(n10860), .ZN(n14067) );
  NAND2_X1 U11187 ( .A1(n17773), .A2(n17755), .ZN(n12305) );
  INV_X1 U11188 ( .A(n15011), .ZN(n15135) );
  NAND2_X1 U11189 ( .A1(n13476), .A2(n13477), .ZN(n13621) );
  NAND2_X1 U11190 ( .A1(n11312), .A2(n11311), .ZN(n13103) );
  NAND2_X1 U11191 ( .A1(n13647), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13656) );
  AND2_X1 U11192 ( .A1(n12818), .A2(n15501), .ZN(n15676) );
  BUF_X1 U11193 ( .A(n10547), .Z(n19752) );
  NAND2_X1 U11194 ( .A1(n11269), .A2(n14091), .ZN(n11295) );
  CLKBUF_X2 U11195 ( .A(n10380), .Z(n13689) );
  NAND2_X1 U11196 ( .A1(n11287), .A2(n11288), .ZN(n11290) );
  NOR2_X1 U11197 ( .A1(n12425), .A2(n12424), .ZN(n18917) );
  NAND2_X2 U11198 ( .A1(n12009), .A2(n12942), .ZN(n12008) );
  AND2_X1 U11200 ( .A1(n10309), .A2(n13047), .ZN(n10310) );
  NAND2_X1 U11201 ( .A1(n10297), .A2(n9675), .ZN(n10695) );
  INV_X2 U11202 ( .A(n13107), .ZN(n12033) );
  OR2_X1 U11204 ( .A1(n13637), .A2(n11170), .ZN(n14094) );
  BUF_X1 U11205 ( .A(n10296), .Z(n19539) );
  INV_X1 U11206 ( .A(n10307), .ZN(n9661) );
  AND4_X1 U11207 ( .A1(n11077), .A2(n11076), .A3(n11075), .A4(n11074), .ZN(
        n11090) );
  AND3_X1 U11208 ( .A1(n11127), .A2(n11126), .A3(n9746), .ZN(n11128) );
  INV_X1 U11209 ( .A(n14416), .ZN(n10606) );
  BUF_X2 U11210 ( .A(n9654), .Z(n9698) );
  BUF_X2 U11211 ( .A(n11069), .Z(n11270) );
  AND2_X2 U11212 ( .A1(n14593), .A2(n10261), .ZN(n10468) );
  BUF_X1 U11213 ( .A(n10211), .Z(n9696) );
  INV_X2 U11214 ( .A(n11885), .ZN(n9662) );
  INV_X1 U11215 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19072) );
  NAND2_X1 U11216 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17176) );
  NOR2_X2 U11217 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13810) );
  INV_X2 U11218 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13581) );
  INV_X2 U11219 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10996) );
  AOI21_X1 U11220 ( .B1(n14663), .B2(n16529), .A(n14662), .ZN(n14664) );
  XNOR2_X1 U11221 ( .A(n14313), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14663) );
  OAI21_X1 U11222 ( .B1(n15047), .B2(n20422), .A(n15046), .ZN(n15048) );
  XNOR2_X1 U11223 ( .A(n12145), .B(n12144), .ZN(n15026) );
  NAND2_X1 U11224 ( .A1(n14679), .A2(n10030), .ZN(n12141) );
  OR2_X1 U11225 ( .A1(n16030), .A2(n15772), .ZN(n15788) );
  AND2_X2 U11226 ( .A1(n14770), .A2(n14769), .ZN(n14757) );
  NOR2_X1 U11227 ( .A1(n10092), .A2(n10093), .ZN(n15700) );
  AND2_X1 U11228 ( .A1(n16032), .A2(n16031), .ZN(n16492) );
  OAI21_X1 U11229 ( .B1(n10092), .B2(n9713), .A(n10981), .ZN(n10987) );
  AOI21_X1 U11230 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(n16319) );
  NAND2_X1 U11231 ( .A1(n9921), .A2(n9920), .ZN(n10092) );
  NAND2_X1 U11232 ( .A1(n15745), .A2(n15947), .ZN(n9921) );
  NOR2_X1 U11233 ( .A1(n16121), .A2(n16128), .ZN(n16120) );
  NOR2_X1 U11234 ( .A1(n14830), .A2(n14831), .ZN(n14829) );
  NOR2_X1 U11235 ( .A1(n15967), .A2(n10959), .ZN(n15745) );
  NAND2_X1 U11236 ( .A1(n11555), .A2(n11554), .ZN(n14830) );
  NOR2_X1 U11237 ( .A1(n15544), .A2(n15543), .ZN(n15542) );
  AOI21_X1 U11238 ( .B1(n16659), .B2(n18367), .A(n9790), .ZN(n16209) );
  AOI211_X1 U11239 ( .C1(n15525), .C2(n19505), .A(n14312), .B(n14311), .ZN(
        n14315) );
  XNOR2_X1 U11240 ( .A(n9904), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16659) );
  NAND2_X1 U11241 ( .A1(n14661), .A2(n14660), .ZN(n14662) );
  XNOR2_X1 U11242 ( .A(n14282), .B(n14281), .ZN(n15888) );
  NOR2_X1 U11243 ( .A1(n12305), .A2(n10143), .ZN(n16634) );
  NAND2_X1 U11244 ( .A1(n9983), .A2(n9981), .ZN(n14503) );
  NOR2_X1 U11245 ( .A1(n9744), .A2(n15135), .ZN(n9978) );
  OAI211_X1 U11246 ( .C1(n16343), .C2(n9963), .A(n14003), .B(n9815), .ZN(n9814) );
  OR2_X1 U11247 ( .A1(n9963), .A2(n16342), .ZN(n9815) );
  AOI211_X1 U11248 ( .C1(n15432), .C2(n19317), .A(n15431), .B(n15430), .ZN(
        n15433) );
  AND2_X1 U11249 ( .A1(n10181), .A2(n14216), .ZN(n9980) );
  NOR2_X1 U11250 ( .A1(n15568), .A2(n15567), .ZN(n15566) );
  NOR2_X1 U11251 ( .A1(n9979), .A2(n9977), .ZN(n9976) );
  INV_X1 U11252 ( .A(n15135), .ZN(n16312) );
  AND2_X1 U11253 ( .A1(n9739), .A2(n10664), .ZN(n9816) );
  AND2_X1 U11254 ( .A1(n17800), .A2(n10191), .ZN(n12303) );
  NAND2_X1 U11255 ( .A1(n10662), .A2(n10661), .ZN(n10664) );
  XNOR2_X1 U11256 ( .A(n13994), .B(n16409), .ZN(n16342) );
  OR2_X1 U11257 ( .A1(n14609), .A2(n14608), .ZN(n16447) );
  NAND2_X1 U11259 ( .A1(n13993), .A2(n13992), .ZN(n13994) );
  NAND2_X1 U11260 ( .A1(n9812), .A2(n9811), .ZN(n14093) );
  NAND2_X1 U11261 ( .A1(n10625), .A2(n10624), .ZN(n10638) );
  NOR2_X1 U11262 ( .A1(n13911), .A2(n13914), .ZN(n14127) );
  NAND2_X1 U11263 ( .A1(n10630), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10636) );
  AND2_X1 U11264 ( .A1(n10030), .A2(n10028), .ZN(n10027) );
  NAND2_X1 U11265 ( .A1(n17815), .A2(n17814), .ZN(n17813) );
  NAND2_X1 U11266 ( .A1(n13103), .A2(n13102), .ZN(n13426) );
  NOR2_X1 U11267 ( .A1(n19961), .A2(n19760), .ZN(n19745) );
  NAND2_X1 U11268 ( .A1(n11391), .A2(n11354), .ZN(n13626) );
  XNOR2_X1 U11269 ( .A(n10844), .B(n10851), .ZN(n10859) );
  AND2_X1 U11270 ( .A1(n15657), .A2(n15999), .ZN(n16001) );
  OR2_X1 U11271 ( .A1(n20263), .A2(n20280), .ZN(n20270) );
  NOR2_X1 U11272 ( .A1(n17806), .A2(n18272), .ZN(n18170) );
  NOR2_X1 U11273 ( .A1(n17517), .A2(n17649), .ZN(n17512) );
  NAND2_X1 U11274 ( .A1(n13656), .A2(n13655), .ZN(n13666) );
  NOR2_X2 U11275 ( .A1(n10960), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10969) );
  NAND2_X1 U11276 ( .A1(n10623), .A2(n10622), .ZN(n10631) );
  AND2_X1 U11277 ( .A1(n10587), .A2(n9858), .ZN(n9857) );
  OR2_X1 U11278 ( .A1(n10603), .A2(n10602), .ZN(n10623) );
  OR2_X1 U11279 ( .A1(n10570), .A2(n10569), .ZN(n10587) );
  XNOR2_X1 U11280 ( .A(n13653), .B(n13646), .ZN(n13647) );
  NAND2_X1 U11281 ( .A1(n15676), .A2(n15675), .ZN(n15674) );
  AND4_X1 U11282 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        n10414) );
  INV_X2 U11283 ( .A(n16264), .ZN(n13741) );
  NOR2_X2 U11284 ( .A1(n18129), .A2(n17605), .ZN(n18039) );
  AOI21_X1 U11285 ( .B1(n18050), .B2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n9891), .ZN(n9890) );
  OAI22_X1 U11286 ( .A1(n10552), .A2(n10396), .B1(n10551), .B2(n13145), .ZN(
        n10397) );
  CLKBUF_X1 U11287 ( .A(n10552), .Z(n19600) );
  NOR2_X1 U11288 ( .A1(n16125), .A2(n10106), .ZN(n12818) );
  XNOR2_X1 U11289 ( .A(n11295), .B(n11293), .ZN(n11307) );
  OR2_X1 U11290 ( .A1(n11295), .A2(n11294), .ZN(n11296) );
  NAND2_X1 U11291 ( .A1(n15520), .A2(n13724), .ZN(n16125) );
  NAND2_X2 U11292 ( .A1(n20356), .A2(n11165), .ZN(n14890) );
  NOR2_X2 U11293 ( .A1(n16828), .A2(n16794), .ZN(n18115) );
  INV_X2 U11294 ( .A(n13114), .ZN(n13366) );
  OAI21_X2 U11295 ( .B1(n13937), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11291), 
        .ZN(n11292) );
  NAND2_X1 U11296 ( .A1(n9970), .A2(n11318), .ZN(n13302) );
  AND2_X1 U11297 ( .A1(n13237), .A2(n13158), .ZN(n9991) );
  NOR2_X1 U11298 ( .A1(n13181), .A2(n13243), .ZN(n13276) );
  INV_X1 U11299 ( .A(n12289), .ZN(n9892) );
  NAND2_X1 U11300 ( .A1(n11204), .A2(n11203), .ZN(n11328) );
  AND2_X1 U11301 ( .A1(n13173), .A2(n13172), .ZN(n13237) );
  AND2_X1 U11302 ( .A1(n13268), .A2(n12943), .ZN(n21047) );
  OR2_X1 U11303 ( .A1(n13045), .A2(n13044), .ZN(n13159) );
  NAND2_X1 U11304 ( .A1(n16564), .A2(n9769), .ZN(n16165) );
  XNOR2_X1 U11305 ( .A(n12287), .B(n12288), .ZN(n18051) );
  AND3_X1 U11306 ( .A1(n9901), .A2(n9753), .A3(n9900), .ZN(n12287) );
  NAND2_X1 U11307 ( .A1(n9803), .A2(n19112), .ZN(n18303) );
  NAND2_X1 U11308 ( .A1(n9803), .A2(n16193), .ZN(n18912) );
  NAND2_X1 U11309 ( .A1(n12950), .A2(n12949), .ZN(n13155) );
  BUF_X1 U11310 ( .A(n10404), .Z(n13845) );
  INV_X1 U11311 ( .A(n13737), .ZN(n12043) );
  OR2_X1 U11312 ( .A1(n18071), .A2(n9903), .ZN(n9900) );
  AND2_X1 U11313 ( .A1(n10392), .A2(n19314), .ZN(n10389) );
  AND2_X1 U11314 ( .A1(n19314), .A2(n10379), .ZN(n10390) );
  NOR3_X1 U11315 ( .A1(n17487), .A2(n17486), .A3(n17485), .ZN(n17577) );
  AND2_X1 U11316 ( .A1(n12007), .A2(n12006), .ZN(n13285) );
  AND2_X2 U11317 ( .A1(n10393), .A2(n10376), .ZN(n19314) );
  NAND2_X1 U11318 ( .A1(n11333), .A2(n11332), .ZN(n20552) );
  AND2_X1 U11319 ( .A1(n10718), .A2(n10713), .ZN(n10124) );
  AND2_X1 U11320 ( .A1(n9843), .A2(n12811), .ZN(n19199) );
  NAND2_X1 U11321 ( .A1(n12566), .A2(n12565), .ZN(n14074) );
  NAND2_X1 U11322 ( .A1(n10043), .A2(n10042), .ZN(n9828) );
  OR2_X1 U11323 ( .A1(n13681), .A2(n10095), .ZN(n12566) );
  XNOR2_X1 U11324 ( .A(n10378), .B(n10377), .ZN(n10392) );
  NOR2_X1 U11325 ( .A1(n13469), .A2(n13468), .ZN(n13471) );
  NOR3_X1 U11326 ( .A1(n18988), .A2(n14254), .A3(n16786), .ZN(n16271) );
  AND2_X1 U11327 ( .A1(n10717), .A2(n10716), .ZN(n13182) );
  OAI21_X1 U11328 ( .B1(n18918), .B2(n14250), .A(n18917), .ZN(n18935) );
  INV_X1 U11329 ( .A(n10351), .ZN(n10378) );
  AND2_X1 U11330 ( .A1(n10722), .A2(n10721), .ZN(n13243) );
  AND2_X1 U11331 ( .A1(n10730), .A2(n10729), .ZN(n13256) );
  XNOR2_X1 U11332 ( .A(n10710), .B(n10712), .ZN(n10708) );
  INV_X2 U11333 ( .A(n17482), .ZN(n17470) );
  NAND2_X1 U11334 ( .A1(n9735), .A2(n12530), .ZN(n10967) );
  INV_X2 U11335 ( .A(n17751), .ZN(n17745) );
  NAND2_X1 U11336 ( .A1(n10343), .A2(n10342), .ZN(n10375) );
  NOR2_X1 U11337 ( .A1(n18094), .A2(n12278), .ZN(n18089) );
  NOR2_X1 U11338 ( .A1(n18096), .A2(n18095), .ZN(n18094) );
  NAND2_X1 U11339 ( .A1(n10355), .A2(n10354), .ZN(n10377) );
  AOI21_X1 U11340 ( .B1(n13716), .B2(n10195), .A(n12555), .ZN(n12558) );
  AOI21_X1 U11341 ( .B1(n10366), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10369), .ZN(n10710) );
  XNOR2_X1 U11342 ( .A(n10149), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18096) );
  CLKBUF_X1 U11343 ( .A(n10365), .Z(n10366) );
  NOR2_X1 U11344 ( .A1(n12424), .A2(n12418), .ZN(n14249) );
  XNOR2_X1 U11345 ( .A(n12486), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14658) );
  NOR2_X1 U11346 ( .A1(n17706), .A2(n14253), .ZN(n12422) );
  XNOR2_X1 U11347 ( .A(n12552), .B(n12545), .ZN(n13712) );
  AOI21_X1 U11348 ( .B1(n10341), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10340), 
        .ZN(n10342) );
  NAND2_X1 U11349 ( .A1(n9895), .A2(n9745), .ZN(n10149) );
  AND2_X1 U11350 ( .A1(n16792), .A2(n12421), .ZN(n14253) );
  AOI211_X1 U11351 ( .C1(n12414), .C2(n18475), .A(n12413), .B(n12412), .ZN(
        n14257) );
  AND2_X1 U11352 ( .A1(n13003), .A2(n13001), .ZN(n12552) );
  AND2_X1 U11353 ( .A1(n10353), .A2(n10352), .ZN(n10355) );
  OAI21_X1 U11354 ( .B1(n12740), .B2(n12540), .A(n12539), .ZN(n13003) );
  NAND2_X1 U11355 ( .A1(n12423), .A2(n12417), .ZN(n14255) );
  NOR2_X1 U11356 ( .A1(n17613), .A2(n12281), .ZN(n12260) );
  AND2_X1 U11357 ( .A1(n10314), .A2(n10313), .ZN(n13066) );
  NOR2_X1 U11358 ( .A1(n10308), .A2(n10301), .ZN(n12998) );
  AND2_X1 U11359 ( .A1(n12840), .A2(n10299), .ZN(n13011) );
  OR2_X1 U11360 ( .A1(n12408), .A2(n9794), .ZN(n12418) );
  NAND2_X1 U11361 ( .A1(n10695), .A2(n10298), .ZN(n12840) );
  NAND2_X1 U11362 ( .A1(n11335), .A2(n11334), .ZN(n11990) );
  NAND2_X1 U11363 ( .A1(n10327), .A2(n13056), .ZN(n12987) );
  NOR2_X1 U11364 ( .A1(n10308), .A2(n10695), .ZN(n13047) );
  NOR2_X1 U11365 ( .A1(n18123), .A2(n18117), .ZN(n18116) );
  AND3_X1 U11366 ( .A1(n9752), .A2(n10332), .A3(n10303), .ZN(n10327) );
  INV_X1 U11367 ( .A(n14094), .ZN(n16235) );
  XNOR2_X1 U11368 ( .A(n17634), .B(n19073), .ZN(n18117) );
  NOR2_X1 U11369 ( .A1(n12146), .A2(n20457), .ZN(n11134) );
  NOR2_X1 U11370 ( .A1(n18503), .A2(n16194), .ZN(n18936) );
  NOR2_X1 U11371 ( .A1(n18518), .A2(n18491), .ZN(n12423) );
  INV_X1 U11372 ( .A(n11130), .ZN(n11113) );
  INV_X1 U11373 ( .A(n17642), .ZN(n18475) );
  INV_X4 U11374 ( .A(n13056), .ZN(n10297) );
  INV_X1 U11375 ( .A(n18503), .ZN(n17495) );
  NAND3_X2 U11376 ( .A1(n9727), .A2(n10168), .A3(n12224), .ZN(n17634) );
  INV_X1 U11377 ( .A(n10321), .ZN(n12989) );
  NAND3_X1 U11378 ( .A1(n12272), .A2(n12271), .A3(n10169), .ZN(n18124) );
  CLKBUF_X1 U11379 ( .A(n10302), .Z(n13078) );
  INV_X2 U11380 ( .A(U212), .ZN(n16725) );
  NAND4_X2 U11381 ( .A1(n11036), .A2(n11035), .A3(n11034), .A4(n11033), .ZN(
        n13642) );
  AND4_X1 U11382 ( .A1(n11143), .A2(n11142), .A3(n11141), .A4(n11140), .ZN(
        n11155) );
  AND2_X2 U11383 ( .A1(n11051), .A2(n11050), .ZN(n11170) );
  NAND2_X1 U11384 ( .A1(n10242), .A2(n10241), .ZN(n10296) );
  AND4_X1 U11385 ( .A1(n11122), .A2(n11121), .A3(n11120), .A4(n11119), .ZN(
        n11129) );
  NAND2_X1 U11386 ( .A1(n10267), .A2(n10266), .ZN(n10307) );
  NAND2_X1 U11387 ( .A1(n9867), .A2(n9865), .ZN(n10321) );
  NAND2_X1 U11388 ( .A1(n9729), .A2(n10259), .ZN(n10267) );
  AND4_X1 U11389 ( .A1(n11073), .A2(n11072), .A3(n11071), .A4(n11070), .ZN(
        n11091) );
  NAND2_X1 U11390 ( .A1(n10283), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10291) );
  NAND2_X1 U11391 ( .A1(n9743), .A2(n9866), .ZN(n9865) );
  AND4_X1 U11392 ( .A1(n11104), .A2(n11103), .A3(n11102), .A4(n11101), .ZN(
        n11110) );
  AND4_X1 U11393 ( .A1(n11040), .A2(n11039), .A3(n11038), .A4(n11037), .ZN(
        n11051) );
  AND4_X1 U11394 ( .A1(n11024), .A2(n11023), .A3(n11022), .A4(n11021), .ZN(
        n11035) );
  AND4_X1 U11395 ( .A1(n11147), .A2(n11146), .A3(n11145), .A4(n11144), .ZN(
        n11154) );
  AND4_X1 U11396 ( .A1(n11028), .A2(n11027), .A3(n11026), .A4(n11025), .ZN(
        n11034) );
  INV_X2 U11397 ( .A(U214), .ZN(n16743) );
  AND4_X1 U11398 ( .A1(n11066), .A2(n11065), .A3(n11064), .A4(n11063), .ZN(
        n11067) );
  NOR2_X2 U11399 ( .A1(n20419), .A2(n20422), .ZN(n20420) );
  AND4_X1 U11400 ( .A1(n11100), .A2(n11099), .A3(n11098), .A4(n11097), .ZN(
        n11111) );
  AND4_X1 U11401 ( .A1(n11014), .A2(n11013), .A3(n11012), .A4(n11011), .ZN(
        n11015) );
  INV_X4 U11402 ( .A(n9653), .ZN(n9673) );
  INV_X2 U11403 ( .A(n12367), .ZN(n17423) );
  AND2_X2 U11404 ( .A1(n10284), .A2(n10261), .ZN(n14430) );
  AND4_X1 U11405 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11036) );
  AND4_X1 U11406 ( .A1(n11108), .A2(n11107), .A3(n11106), .A4(n11105), .ZN(
        n11109) );
  OAI22_X1 U11407 ( .A1(n17148), .A2(n12220), .B1(n12367), .B2(n12219), .ZN(
        n12221) );
  AND4_X1 U11408 ( .A1(n11139), .A2(n11138), .A3(n11137), .A4(n11136), .ZN(
        n11156) );
  NAND2_X2 U11409 ( .A1(n19121), .A2(n18996), .ZN(n19044) );
  INV_X2 U11410 ( .A(n19002), .ZN(n9664) );
  AND2_X1 U11411 ( .A1(n10258), .A2(n10257), .ZN(n10259) );
  NAND2_X2 U11412 ( .A1(n20163), .A2(n20120), .ZN(n20166) );
  NAND2_X2 U11413 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20163), .ZN(n20162) );
  INV_X1 U11414 ( .A(n17392), .ZN(n17208) );
  NAND2_X1 U11415 ( .A1(n9691), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14416) );
  INV_X2 U11416 ( .A(n11078), .ZN(n11787) );
  BUF_X2 U11417 ( .A(n11221), .Z(n11940) );
  INV_X2 U11418 ( .A(n14264), .ZN(n17196) );
  INV_X1 U11419 ( .A(n12265), .ZN(n12367) );
  CLKBUF_X3 U11420 ( .A(n12266), .Z(n17382) );
  OR2_X2 U11421 ( .A1(n12841), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19277) );
  INV_X2 U11422 ( .A(n16782), .ZN(n16784) );
  BUF_X4 U11423 ( .A(n11062), .Z(n11941) );
  NAND2_X1 U11424 ( .A1(n10416), .A2(n10261), .ZN(n14417) );
  NOR2_X1 U11425 ( .A1(n12180), .A2(n17175), .ZN(n12265) );
  NOR2_X4 U11426 ( .A1(n17175), .A2(n12177), .ZN(n12249) );
  INV_X1 U11427 ( .A(n17440), .ZN(n9665) );
  CLKBUF_X2 U11428 ( .A(n10211), .Z(n14590) );
  AND2_X2 U11429 ( .A1(n10994), .A2(n13574), .ZN(n9678) );
  OR2_X1 U11430 ( .A1(n17176), .A2(n12181), .ZN(n17148) );
  NOR2_X1 U11431 ( .A1(n12178), .A2(n12180), .ZN(n12266) );
  NOR2_X1 U11432 ( .A1(n12177), .A2(n12179), .ZN(n14166) );
  AND2_X2 U11433 ( .A1(n11006), .A2(n11010), .ZN(n9672) );
  OR2_X2 U11434 ( .A1(n13333), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20393) );
  AND2_X1 U11435 ( .A1(n10418), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9679) );
  NAND2_X1 U11436 ( .A1(n12318), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12179) );
  AND2_X2 U11437 ( .A1(n10418), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9680) );
  NAND2_X1 U11438 ( .A1(n19072), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12181) );
  NAND2_X1 U11439 ( .A1(n12318), .A2(n17147), .ZN(n17175) );
  INV_X2 U11440 ( .A(n11123), .ZN(n9666) );
  AND2_X1 U11441 ( .A1(n16215), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10994) );
  AND2_X1 U11442 ( .A1(n13810), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10206) );
  NAND2_X1 U11443 ( .A1(n19072), .A2(n12320), .ZN(n12180) );
  AND2_X2 U11444 ( .A1(n10197), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14442) );
  NOR2_X1 U11445 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10197) );
  INV_X1 U11446 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10339) );
  NAND2_X1 U11447 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14265) );
  INV_X2 U11448 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12318) );
  INV_X1 U11449 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16575) );
  INV_X1 U11450 ( .A(n9665), .ZN(n9689) );
  NOR2_X4 U11451 ( .A1(n17176), .A2(n12180), .ZN(n17440) );
  NAND3_X1 U11452 ( .A1(n9675), .A2(n10300), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n14477) );
  NAND2_X1 U11453 ( .A1(n10300), .A2(n9661), .ZN(n12984) );
  AND2_X1 U11454 ( .A1(n10300), .A2(n10307), .ZN(n10312) );
  OR2_X1 U11455 ( .A1(n15242), .A2(n20325), .ZN(n9667) );
  NAND2_X1 U11456 ( .A1(n9667), .A2(n9869), .ZN(P1_U2810) );
  OR2_X1 U11457 ( .A1(n14830), .A2(n14831), .ZN(n9668) );
  XNOR2_X1 U11458 ( .A(n9872), .B(n9871), .ZN(n15242) );
  NOR2_X1 U11459 ( .A1(n12139), .A2(n9870), .ZN(n9869) );
  NOR2_X1 U11460 ( .A1(n12296), .A2(n12295), .ZN(n17914) );
  NAND2_X1 U11461 ( .A1(n15062), .A2(n15020), .ZN(n9669) );
  CLKBUF_X1 U11462 ( .A(n13299), .Z(n9670) );
  CLKBUF_X1 U11463 ( .A(n13978), .Z(n9671) );
  NAND2_X1 U11464 ( .A1(n15062), .A2(n15020), .ZN(n15022) );
  NOR2_X2 U11465 ( .A1(n17573), .A2(n17671), .ZN(n17568) );
  NOR3_X2 U11467 ( .A1(n12511), .A2(n9839), .A3(n10799), .ZN(n12485) );
  NAND2_X1 U11468 ( .A1(n12008), .A2(n11157), .ZN(n13299) );
  INV_X1 U11469 ( .A(n11215), .ZN(n9674) );
  BUF_X4 U11470 ( .A(n19535), .Z(n9675) );
  NAND2_X2 U11471 ( .A1(n10291), .A2(n10290), .ZN(n19535) );
  NOR2_X2 U11472 ( .A1(n13030), .A2(n13310), .ZN(n11133) );
  OAI21_X2 U11473 ( .B1(n18130), .B2(n18324), .A(n9800), .ZN(n18020) );
  AND2_X1 U11474 ( .A1(n10994), .A2(n13574), .ZN(n9677) );
  AND2_X1 U11475 ( .A1(n10994), .A2(n13574), .ZN(n11213) );
  AND2_X2 U11476 ( .A1(n13581), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11006) );
  NAND2_X2 U11477 ( .A1(n15063), .A2(n15072), .ZN(n15062) );
  INV_X2 U11478 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13840) );
  NAND2_X1 U11479 ( .A1(n15197), .A2(n9751), .ZN(n15010) );
  XNOR2_X1 U11480 ( .A(n11328), .B(n20552), .ZN(n20426) );
  INV_X1 U11481 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n9681) );
  OR2_X1 U11482 ( .A1(n11180), .A2(n11196), .ZN(n11206) );
  AOI21_X2 U11483 ( .B1(n14068), .B2(n14067), .A(n10863), .ZN(n14237) );
  AOI21_X1 U11484 ( .B1(n11197), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11198), .ZN(n11207) );
  INV_X1 U11485 ( .A(n9654), .ZN(n9682) );
  AND2_X2 U11486 ( .A1(n11008), .A2(n11007), .ZN(n11838) );
  CLKBUF_X1 U11487 ( .A(n11838), .Z(n9704) );
  CLKBUF_X1 U11488 ( .A(n11838), .Z(n9703) );
  INV_X2 U11489 ( .A(n14264), .ZN(n9683) );
  OR2_X1 U11490 ( .A1(n12179), .A2(n14265), .ZN(n14264) );
  AND2_X1 U11491 ( .A1(n13661), .A2(n20387), .ZN(n9712) );
  NAND2_X1 U11492 ( .A1(n14093), .A2(n14092), .ZN(n9685) );
  OAI21_X2 U11493 ( .B1(n13627), .B2(n9971), .A(n13660), .ZN(n13661) );
  OAI22_X2 U11494 ( .A1(n9681), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19332) );
  OAI22_X1 U11495 ( .A1(n16267), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14338), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13720) );
  OAI22_X4 U11496 ( .A1(n16267), .A2(n14285), .B1(n14658), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n12811) );
  NAND2_X1 U11497 ( .A1(n20359), .A2(n20358), .ZN(n20361) );
  NAND2_X2 U11498 ( .A1(n11180), .A2(n11176), .ZN(n11197) );
  NAND2_X2 U11499 ( .A1(n11162), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11180) );
  AND2_X4 U11500 ( .A1(n15869), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15850) );
  AND2_X2 U11501 ( .A1(n9818), .A2(n9817), .ZN(n15869) );
  INV_X2 U11502 ( .A(n17209), .ZN(n9687) );
  INV_X1 U11503 ( .A(n17209), .ZN(n9688) );
  XNOR2_X1 U11504 ( .A(n11308), .B(n11292), .ZN(n13630) );
  AND2_X2 U11505 ( .A1(n14757), .A2(n10013), .ZN(n14701) );
  BUF_X4 U11506 ( .A(n10206), .Z(n9691) );
  BUF_X4 U11507 ( .A(n10206), .Z(n9692) );
  AND2_X1 U11508 ( .A1(n11009), .A2(n13570), .ZN(n9693) );
  AND3_X2 U11509 ( .A1(n20450), .A2(n20446), .A3(n10038), .ZN(n13031) );
  NAND2_X1 U11510 ( .A1(n11183), .A2(n11182), .ZN(n9952) );
  NOR2_X2 U11511 ( .A1(n13704), .A2(n13837), .ZN(n13802) );
  NAND2_X2 U11512 ( .A1(n11353), .A2(n11300), .ZN(n13627) );
  NOR2_X1 U11513 ( .A1(n11970), .A2(n20446), .ZN(n11999) );
  BUF_X1 U11514 ( .A(n10211), .Z(n9695) );
  OAI21_X2 U11515 ( .B1(n13626), .B2(n11503), .A(n11364), .ZN(n13467) );
  NAND2_X2 U11516 ( .A1(n11134), .A2(n13031), .ZN(n12149) );
  NAND2_X2 U11517 ( .A1(n11328), .A2(n11208), .ZN(n13223) );
  AND2_X1 U11518 ( .A1(n14679), .A2(n10027), .ZN(n12145) );
  NOR2_X4 U11519 ( .A1(n14691), .A2(n14692), .ZN(n14679) );
  NAND2_X1 U11520 ( .A1(n13219), .A2(n13581), .ZN(n11078) );
  INV_X2 U11521 ( .A(n12155), .ZN(n10038) );
  AND2_X1 U11522 ( .A1(n11009), .A2(n13569), .ZN(n9699) );
  NAND2_X2 U11523 ( .A1(n11133), .A2(n11163), .ZN(n12009) );
  AND2_X1 U11524 ( .A1(n13569), .A2(n11008), .ZN(n9700) );
  NOR2_X2 U11525 ( .A1(n13801), .A2(n10034), .ZN(n14027) );
  INV_X1 U11526 ( .A(n13630), .ZN(n9701) );
  INV_X1 U11527 ( .A(n9701), .ZN(n9702) );
  NAND2_X1 U11528 ( .A1(n10046), .A2(n10045), .ZN(n10359) );
  OR2_X1 U11529 ( .A1(n15412), .A2(n20963), .ZN(n11953) );
  INV_X1 U11530 ( .A(n10196), .ZN(n11928) );
  OAI22_X1 U11531 ( .A1(n14114), .A2(n10546), .B1(n10547), .B2(n14107), .ZN(
        n10387) );
  INV_X1 U11532 ( .A(n11415), .ZN(n9812) );
  NAND2_X1 U11533 ( .A1(n10310), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10048) );
  AOI21_X1 U11534 ( .B1(n10091), .B2(n10089), .A(n10087), .ZN(n10086) );
  INV_X1 U11535 ( .A(n15861), .ZN(n10087) );
  NOR2_X1 U11536 ( .A1(n13944), .A2(n10036), .ZN(n10035) );
  INV_X1 U11537 ( .A(n10176), .ZN(n10036) );
  NOR2_X1 U11538 ( .A1(n11165), .A2(n20966), .ZN(n11359) );
  NOR2_X1 U11539 ( .A1(n15153), .A2(n15001), .ZN(n9810) );
  OR2_X1 U11540 ( .A1(n11430), .A2(n11429), .ZN(n14008) );
  INV_X1 U11541 ( .A(n11032), .ZN(n11033) );
  NAND2_X1 U11542 ( .A1(n10930), .A2(n15583), .ZN(n10951) );
  NAND2_X1 U11543 ( .A1(n10000), .A2(n9999), .ZN(n9998) );
  NAND2_X1 U11544 ( .A1(n10165), .A2(n10000), .ZN(n9997) );
  INV_X1 U11545 ( .A(n15543), .ZN(n9999) );
  NAND2_X1 U11546 ( .A1(n10789), .A2(n15436), .ZN(n10135) );
  NAND2_X1 U11547 ( .A1(n10115), .A2(n10297), .ZN(n10345) );
  NAND2_X1 U11548 ( .A1(n12320), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12177) );
  AND2_X1 U11549 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12279), .ZN(
        n12280) );
  INV_X1 U11550 ( .A(n10076), .ZN(n10075) );
  NAND2_X1 U11551 ( .A1(n20261), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13854) );
  AOI21_X1 U11552 ( .B1(n11928), .B2(n15065), .A(n11875), .ZN(n14680) );
  OR2_X1 U11553 ( .A1(n13285), .A2(n12152), .ZN(n13188) );
  INV_X1 U11554 ( .A(n11902), .ZN(n12143) );
  NAND2_X1 U11555 ( .A1(n13627), .A2(n11306), .ZN(n10012) );
  AOI21_X1 U11556 ( .B1(n11306), .B2(n11503), .A(n10011), .ZN(n10010) );
  INV_X1 U11557 ( .A(n11327), .ZN(n10011) );
  OR2_X1 U11558 ( .A1(n13285), .A2(n20238), .ZN(n13332) );
  INV_X1 U11559 ( .A(n9965), .ZN(n15037) );
  INV_X2 U11560 ( .A(n9656), .ZN(n12472) );
  INV_X1 U11561 ( .A(n11165), .ZN(n20457) );
  OR2_X1 U11562 ( .A1(n20213), .A2(n13081), .ZN(n10698) );
  NAND2_X1 U11563 ( .A1(n12505), .A2(n12811), .ZN(n19183) );
  AND2_X1 U11564 ( .A1(n16590), .A2(n20095), .ZN(n12837) );
  NAND2_X1 U11565 ( .A1(n15700), .A2(n9906), .ZN(n9905) );
  NAND2_X1 U11566 ( .A1(n9756), .A2(n9915), .ZN(n9906) );
  AND2_X1 U11567 ( .A1(n15775), .A2(n9918), .ZN(n9917) );
  AND2_X1 U11568 ( .A1(n9788), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9831) );
  OR2_X1 U11569 ( .A1(n13689), .A2(n13165), .ZN(n13173) );
  NOR2_X1 U11570 ( .A1(n17992), .A2(n17995), .ZN(n17977) );
  INV_X1 U11571 ( .A(n10586), .ZN(n9859) );
  AOI22_X1 U11572 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10542), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10399) );
  AND4_X1 U11573 ( .A1(n10656), .A2(n10655), .A3(n10654), .A4(n10653), .ZN(
        n10658) );
  AND2_X1 U11574 ( .A1(n10201), .A2(n10198), .ZN(n9868) );
  AND2_X1 U11575 ( .A1(n20820), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11973) );
  NOR2_X1 U11576 ( .A1(n11963), .A2(n11964), .ZN(n11962) );
  AND2_X2 U11577 ( .A1(n11302), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11007) );
  AND2_X1 U11578 ( .A1(n12105), .A2(n9877), .ZN(n9875) );
  AND4_X1 U11579 ( .A1(n10321), .A2(n10302), .A3(n10296), .A4(n10305), .ZN(
        n10331) );
  NAND2_X1 U11580 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10047) );
  OR2_X1 U11581 ( .A1(n10584), .A2(n10583), .ZN(n10809) );
  NAND2_X1 U11582 ( .A1(n9663), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U11583 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10061) );
  AOI21_X1 U11584 ( .B1(n10540), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n10443), .ZN(n10451) );
  NAND2_X1 U11585 ( .A1(n10344), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10350) );
  NAND2_X1 U11586 ( .A1(n10331), .A2(n10312), .ZN(n10330) );
  AND2_X1 U11587 ( .A1(n10315), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10309) );
  NAND2_X1 U11588 ( .A1(n10604), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10467) );
  AND2_X1 U11589 ( .A1(n12989), .A2(n10305), .ZN(n10299) );
  AOI21_X1 U11590 ( .B1(n12989), .B2(n12984), .A(n10322), .ZN(n10313) );
  AOI21_X1 U11591 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20182), .A(
        n10675), .ZN(n10679) );
  AND3_X1 U11592 ( .A1(n10237), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10236), .ZN(n10239) );
  AOI22_X1 U11593 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10237) );
  NAND2_X1 U11594 ( .A1(n12408), .A2(n18491), .ZN(n12410) );
  NOR2_X1 U11595 ( .A1(n10019), .A2(n10016), .ZN(n10015) );
  INV_X1 U11596 ( .A(n10017), .ZN(n10016) );
  INV_X1 U11597 ( .A(n14730), .ZN(n10019) );
  NOR2_X1 U11598 ( .A1(n14743), .A2(n10018), .ZN(n10017) );
  INV_X1 U11599 ( .A(n14758), .ZN(n10018) );
  NOR2_X1 U11600 ( .A1(n11694), .A2(n21227), .ZN(n11716) );
  AND2_X1 U11601 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n11670), .ZN(
        n11671) );
  NAND2_X1 U11602 ( .A1(n10022), .A2(n10021), .ZN(n10020) );
  INV_X1 U11603 ( .A(n14783), .ZN(n10021) );
  NOR2_X1 U11604 ( .A1(n10023), .A2(n14796), .ZN(n10022) );
  INV_X1 U11605 ( .A(n10025), .ZN(n10023) );
  XNOR2_X1 U11606 ( .A(n14093), .B(n11440), .ZN(n14006) );
  AOI21_X1 U11607 ( .B1(n9978), .B2(n9976), .A(n9974), .ZN(n9973) );
  INV_X1 U11608 ( .A(n9976), .ZN(n9975) );
  NOR2_X1 U11609 ( .A1(n13736), .A2(n16398), .ZN(n9880) );
  NAND2_X1 U11610 ( .A1(n9812), .A2(n11416), .ZN(n11435) );
  INV_X1 U11611 ( .A(n13662), .ZN(n9960) );
  INV_X1 U11612 ( .A(n13667), .ZN(n9962) );
  AND2_X1 U11613 ( .A1(n13107), .A2(n9656), .ZN(n12112) );
  NAND2_X1 U11614 ( .A1(n13645), .A2(n13644), .ZN(n13653) );
  NOR2_X1 U11615 ( .A1(n9969), .A2(n9971), .ZN(n9968) );
  INV_X1 U11616 ( .A(n11318), .ZN(n9969) );
  AND2_X1 U11617 ( .A1(n11286), .A2(n11285), .ZN(n11293) );
  INV_X1 U11618 ( .A(n13583), .ZN(n16217) );
  OR2_X1 U11619 ( .A1(n10956), .A2(n10954), .ZN(n10960) );
  NAND2_X1 U11620 ( .A1(n10951), .A2(n10967), .ZN(n10932) );
  AND2_X1 U11621 ( .A1(n10911), .A2(n9770), .ZN(n10930) );
  INV_X1 U11622 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n9929) );
  NAND2_X1 U11623 ( .A1(n10907), .A2(n10967), .ZN(n10911) );
  AND2_X1 U11624 ( .A1(n10911), .A2(n10910), .ZN(n10913) );
  AND2_X1 U11625 ( .A1(n10925), .A2(n10923), .ZN(n10916) );
  AND2_X1 U11626 ( .A1(n10888), .A2(n10893), .ZN(n10925) );
  AND2_X1 U11627 ( .A1(n10871), .A2(n13423), .ZN(n10879) );
  NAND2_X1 U11628 ( .A1(n9925), .A2(n10864), .ZN(n9924) );
  INV_X1 U11629 ( .A(n9926), .ZN(n9925) );
  NAND2_X1 U11630 ( .A1(n9663), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10074) );
  NAND2_X1 U11631 ( .A1(n9663), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10070) );
  NAND2_X1 U11632 ( .A1(n9680), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14411) );
  OAI22_X1 U11633 ( .A1(n10370), .A2(n10261), .B1(n20220), .B2(n20182), .ZN(
        n10712) );
  INV_X1 U11634 ( .A(n15454), .ZN(n10103) );
  AOI21_X1 U11635 ( .B1(n9982), .B2(n14479), .A(n9780), .ZN(n9981) );
  AND2_X1 U11636 ( .A1(n12754), .A2(n10105), .ZN(n10104) );
  INV_X1 U11637 ( .A(n15624), .ZN(n10105) );
  INV_X1 U11638 ( .A(n10005), .ZN(n10004) );
  AND2_X1 U11639 ( .A1(n10007), .A2(n10006), .ZN(n10005) );
  INV_X1 U11640 ( .A(n15574), .ZN(n10006) );
  OR2_X1 U11641 ( .A1(n10110), .A2(n10109), .ZN(n10108) );
  INV_X1 U11642 ( .A(n16098), .ZN(n10109) );
  NAND2_X1 U11643 ( .A1(n10111), .A2(n16108), .ZN(n10110) );
  INV_X1 U11644 ( .A(n16124), .ZN(n10111) );
  NOR2_X1 U11645 ( .A1(n9676), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12531) );
  NAND2_X1 U11646 ( .A1(n9663), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10068) );
  NOR2_X1 U11647 ( .A1(n15469), .A2(n10128), .ZN(n10127) );
  NAND2_X1 U11648 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9835) );
  NAND2_X1 U11649 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9836) );
  NAND2_X1 U11650 ( .A1(n9663), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10064) );
  NAND2_X1 U11651 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U11652 ( .A1(n9663), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10060) );
  NAND2_X1 U11653 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10059) );
  INV_X1 U11654 ( .A(n13418), .ZN(n10117) );
  NOR2_X1 U11655 ( .A1(n13256), .A2(n10120), .ZN(n10119) );
  INV_X1 U11656 ( .A(n13528), .ZN(n10120) );
  NAND2_X1 U11657 ( .A1(n9663), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10058) );
  NAND2_X1 U11658 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10057) );
  NAND2_X1 U11659 ( .A1(n9824), .A2(n9828), .ZN(n9823) );
  INV_X1 U11660 ( .A(n10364), .ZN(n9824) );
  NAND2_X1 U11661 ( .A1(n10501), .A2(n10502), .ZN(n10696) );
  NAND2_X1 U11662 ( .A1(n10127), .A2(n15453), .ZN(n10126) );
  OR2_X1 U11663 ( .A1(n15487), .A2(n10869), .ZN(n10953) );
  NAND2_X1 U11664 ( .A1(n9663), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10066) );
  NAND2_X1 U11665 ( .A1(n9663), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U11666 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10051) );
  INV_X1 U11667 ( .A(n10631), .ZN(n10624) );
  INV_X1 U11668 ( .A(n10626), .ZN(n10625) );
  NAND2_X1 U11669 ( .A1(n9663), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10054) );
  NAND2_X1 U11670 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10053) );
  NAND2_X2 U11671 ( .A1(n13004), .A2(n12531), .ZN(n12766) );
  AND2_X1 U11672 ( .A1(n14655), .A2(n10390), .ZN(n10382) );
  NAND2_X1 U11674 ( .A1(n16200), .A2(n12405), .ZN(n12417) );
  INV_X1 U11675 ( .A(n12373), .ZN(n9798) );
  NAND2_X1 U11676 ( .A1(n17933), .A2(n12306), .ZN(n10143) );
  INV_X1 U11677 ( .A(n18106), .ZN(n9895) );
  NAND2_X1 U11678 ( .A1(n18475), .A2(n17597), .ZN(n12408) );
  AOI22_X1 U11679 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18942), .B2(n12318), .ZN(
        n12429) );
  NOR2_X1 U11680 ( .A1(n16822), .A2(n9844), .ZN(n14254) );
  AND2_X1 U11681 ( .A1(n17706), .A2(n16828), .ZN(n9844) );
  INV_X1 U11682 ( .A(n13213), .ZN(n9813) );
  INV_X1 U11683 ( .A(n10031), .ZN(n10029) );
  OR2_X1 U11684 ( .A1(n11851), .A2(n14693), .ZN(n11852) );
  NAND2_X1 U11685 ( .A1(n11803), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11851) );
  OAI21_X1 U11686 ( .B1(n10196), .B2(n15096), .A(n11802), .ZN(n14717) );
  NAND2_X1 U11687 ( .A1(n11716), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11741) );
  AND2_X1 U11688 ( .A1(n11697), .A2(n11696), .ZN(n14769) );
  NAND2_X1 U11689 ( .A1(n10035), .A2(n14028), .ZN(n10034) );
  INV_X1 U11690 ( .A(n11431), .ZN(n11441) );
  AOI21_X1 U11691 ( .B1(n13986), .B2(n11590), .A(n11412), .ZN(n13706) );
  NAND2_X1 U11692 ( .A1(n13668), .A2(n13667), .ZN(n13976) );
  INV_X1 U11693 ( .A(n13426), .ZN(n11326) );
  AND2_X1 U11694 ( .A1(n9708), .A2(n15023), .ZN(n9805) );
  NOR2_X1 U11695 ( .A1(n15135), .A2(n15211), .ZN(n9966) );
  NAND2_X1 U11696 ( .A1(n14881), .A2(n9779), .ZN(n14801) );
  NOR2_X1 U11697 ( .A1(n14800), .A2(n15365), .ZN(n9887) );
  NAND2_X1 U11698 ( .A1(n9728), .A2(n13822), .ZN(n14025) );
  NOR2_X2 U11699 ( .A1(n11968), .A2(n11170), .ZN(n13107) );
  NOR2_X1 U11700 ( .A1(n11005), .A2(n11004), .ZN(n11016) );
  NAND2_X1 U11701 ( .A1(n13298), .A2(n13297), .ZN(n13324) );
  OR2_X1 U11702 ( .A1(n13332), .A2(n13296), .ZN(n13297) );
  INV_X1 U11703 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20786) );
  INV_X1 U11704 ( .A(n13303), .ZN(n20442) );
  NAND2_X1 U11705 ( .A1(n20963), .A2(n20423), .ZN(n20557) );
  INV_X1 U11706 ( .A(n14281), .ZN(n10132) );
  INV_X1 U11707 ( .A(n12828), .ZN(n10133) );
  INV_X1 U11708 ( .A(n10135), .ZN(n10134) );
  INV_X1 U11709 ( .A(n19199), .ZN(n9842) );
  OR2_X1 U11710 ( .A1(n10920), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10907) );
  NAND2_X1 U11711 ( .A1(n10072), .A2(n10071), .ZN(n10782) );
  NAND2_X1 U11712 ( .A1(n13623), .A2(n9996), .ZN(n9995) );
  INV_X1 U11713 ( .A(n13831), .ZN(n9996) );
  NAND2_X1 U11714 ( .A1(n10050), .A2(n10049), .ZN(n10715) );
  INV_X1 U11715 ( .A(n12766), .ZN(n14296) );
  CLKBUF_X2 U11716 ( .A(n12543), .Z(n14295) );
  AND2_X1 U11717 ( .A1(n15443), .A2(n14607), .ZN(n14609) );
  NAND2_X1 U11718 ( .A1(n14582), .A2(n14604), .ZN(n9990) );
  NOR2_X1 U11719 ( .A1(n9987), .A2(n14604), .ZN(n9986) );
  INV_X1 U11720 ( .A(n15526), .ZN(n9987) );
  NOR2_X2 U11721 ( .A1(n9723), .A2(n15444), .ZN(n15443) );
  NOR2_X1 U11722 ( .A1(n15542), .A2(n10165), .ZN(n14545) );
  AND2_X1 U11723 ( .A1(n10307), .A2(n10305), .ZN(n13004) );
  INV_X1 U11724 ( .A(n12977), .ZN(n19416) );
  AND2_X1 U11725 ( .A1(n12485), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12486) );
  NAND2_X1 U11726 ( .A1(n10056), .A2(n10055), .ZN(n10705) );
  AND2_X1 U11727 ( .A1(n15450), .A2(n14277), .ZN(n15702) );
  NAND2_X1 U11728 ( .A1(n9911), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9908) );
  NAND2_X1 U11729 ( .A1(n9913), .A2(n9912), .ZN(n9911) );
  NOR2_X1 U11730 ( .A1(n10948), .A2(n10947), .ZN(n10949) );
  OR2_X1 U11731 ( .A1(n10953), .A2(n15977), .ZN(n15974) );
  INV_X1 U11732 ( .A(n10130), .ZN(n13618) );
  NAND2_X1 U11733 ( .A1(n9754), .A2(n9706), .ZN(n10089) );
  NAND2_X1 U11734 ( .A1(n9755), .A2(n10664), .ZN(n9818) );
  NAND2_X1 U11735 ( .A1(n13276), .A2(n13275), .ZN(n13277) );
  AND2_X1 U11736 ( .A1(n10862), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10863) );
  AND2_X1 U11737 ( .A1(n13065), .A2(n20095), .ZN(n13091) );
  NAND2_X1 U11738 ( .A1(n19314), .A2(n13147), .ZN(n12950) );
  NAND2_X1 U11739 ( .A1(n9991), .A2(n13159), .ZN(n13240) );
  CLKBUF_X1 U11740 ( .A(n13088), .Z(n13809) );
  INV_X1 U11741 ( .A(n19719), .ZN(n19658) );
  INV_X1 U11742 ( .A(n20183), .ZN(n19989) );
  INV_X1 U11743 ( .A(n19898), .ZN(n19886) );
  INV_X1 U11744 ( .A(n19959), .ZN(n19961) );
  AND2_X1 U11745 ( .A1(n20184), .A2(n20193), .ZN(n20174) );
  AND2_X1 U11746 ( .A1(n20225), .A2(n20200), .ZN(n16266) );
  AND2_X1 U11747 ( .A1(n10681), .A2(n12974), .ZN(n16590) );
  NOR2_X1 U11748 ( .A1(n16865), .A2(n17144), .ZN(n16855) );
  OR2_X1 U11749 ( .A1(n16855), .A2(n16856), .ZN(n9931) );
  NOR2_X1 U11750 ( .A1(n16866), .A2(n17759), .ZN(n16865) );
  AND2_X1 U11751 ( .A1(n9944), .A2(n9943), .ZN(n9940) );
  OR2_X1 U11752 ( .A1(n17144), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9944) );
  NAND2_X1 U11753 ( .A1(n9940), .A2(n16959), .ZN(n9941) );
  NOR2_X1 U11754 ( .A1(n18909), .A2(n17641), .ZN(n19122) );
  AOI22_X1 U11755 ( .A1(n14259), .A2(n18907), .B1(n14134), .B2(n14133), .ZN(
        n16269) );
  NAND2_X1 U11756 ( .A1(n12263), .A2(n12262), .ZN(n12264) );
  NAND2_X1 U11757 ( .A1(n12191), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12262) );
  OAI21_X1 U11758 ( .B1(n17148), .B2(n9899), .A(n9897), .ZN(n9896) );
  INV_X1 U11759 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n9899) );
  AOI21_X1 U11760 ( .B1(n12335), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(n9898), .ZN(n9897) );
  NOR2_X1 U11761 ( .A1(n9721), .A2(n18478), .ZN(n9898) );
  NOR2_X1 U11762 ( .A1(n18967), .A2(n16786), .ZN(n17705) );
  AND2_X1 U11763 ( .A1(n12458), .A2(n9946), .ZN(n16660) );
  NOR2_X1 U11764 ( .A1(n9947), .A2(n16862), .ZN(n9946) );
  INV_X1 U11765 ( .A(n9948), .ZN(n9947) );
  NOR2_X1 U11766 ( .A1(n17794), .A2(n17795), .ZN(n12458) );
  INV_X1 U11767 ( .A(n17813), .ZN(n17801) );
  NOR2_X1 U11768 ( .A1(n17863), .A2(n17838), .ZN(n16819) );
  NOR2_X1 U11769 ( .A1(n17919), .A2(n12456), .ZN(n17903) );
  NAND2_X1 U11770 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12456) );
  NOR2_X1 U11771 ( .A1(n17946), .A2(n17947), .ZN(n17916) );
  NAND2_X1 U11772 ( .A1(n18029), .A2(n9734), .ZN(n17992) );
  NOR2_X1 U11773 ( .A1(n12305), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16627) );
  NAND2_X1 U11774 ( .A1(n10146), .A2(n12306), .ZN(n10144) );
  NOR2_X1 U11775 ( .A1(n18038), .A2(n16628), .ZN(n10146) );
  NAND2_X1 U11776 ( .A1(n9718), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10145) );
  INV_X1 U11777 ( .A(n16634), .ZN(n10142) );
  NOR2_X1 U11778 ( .A1(n12289), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10150) );
  OR2_X1 U11779 ( .A1(n18059), .A2(n18072), .ZN(n9903) );
  NAND2_X1 U11780 ( .A1(n12284), .A2(n9902), .ZN(n9901) );
  INV_X1 U11781 ( .A(n18059), .ZN(n9902) );
  OR2_X1 U11782 ( .A1(n18071), .A2(n18072), .ZN(n10138) );
  OR2_X1 U11783 ( .A1(n16453), .A2(n10973), .ZN(n10985) );
  OR2_X1 U11784 ( .A1(n10984), .A2(n15937), .ZN(n15731) );
  NAND2_X1 U11785 ( .A1(n10094), .A2(n15732), .ZN(n10093) );
  INV_X1 U11786 ( .A(n15727), .ZN(n10094) );
  NAND2_X1 U11787 ( .A1(n10964), .A2(n10963), .ZN(n9920) );
  NOR2_X2 U11788 ( .A1(n12128), .A2(n12119), .ZN(n20334) );
  AND2_X1 U11789 ( .A1(n14988), .A2(n14329), .ZN(n14959) );
  INV_X1 U11790 ( .A(n14988), .ZN(n14991) );
  INV_X1 U11791 ( .A(n13268), .ZN(n13267) );
  INV_X1 U11792 ( .A(n12471), .ZN(n9871) );
  INV_X1 U11793 ( .A(n12118), .ZN(n9872) );
  AND2_X1 U11794 ( .A1(n19480), .A2(n12777), .ZN(n19319) );
  INV_X1 U11795 ( .A(n20184), .ZN(n19520) );
  INV_X1 U11796 ( .A(n20193), .ZN(n19657) );
  INV_X1 U11797 ( .A(n15572), .ZN(n15592) );
  AND2_X1 U11798 ( .A1(n19371), .A2(n13004), .ZN(n19338) );
  AND2_X1 U11799 ( .A1(n19414), .A2(n19413), .ZN(n19456) );
  NAND2_X1 U11800 ( .A1(n12847), .A2(n10791), .ZN(n16541) );
  INV_X1 U11801 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20182) );
  AND2_X1 U11802 ( .A1(n16597), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16616) );
  INV_X1 U11803 ( .A(n17190), .ZN(n17177) );
  NOR2_X1 U11804 ( .A1(n17597), .A2(n17303), .ZN(n17291) );
  NAND2_X1 U11805 ( .A1(n17579), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n17573) );
  CLKBUF_X1 U11806 ( .A(n14442), .Z(n14589) );
  AOI22_X1 U11807 ( .A1(n10562), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10561), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10411) );
  NAND2_X1 U11808 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10045) );
  AOI21_X1 U11809 ( .B1(n10318), .B2(n19545), .A(n13056), .ZN(n10316) );
  AND2_X1 U11810 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10216) );
  OAI21_X1 U11811 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n12320), .A(
        n12323), .ZN(n12324) );
  OR2_X1 U11812 ( .A1(n12322), .A2(n12321), .ZN(n12323) );
  NAND2_X1 U11813 ( .A1(n11959), .A2(n11958), .ZN(n11986) );
  AOI22_X1 U11814 ( .A1(n11986), .A2(n11985), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20787), .ZN(n11963) );
  AND2_X1 U11815 ( .A1(n11167), .A2(n11186), .ZN(n12148) );
  INV_X1 U11816 ( .A(n15143), .ZN(n9974) );
  OR2_X1 U11817 ( .A1(n11406), .A2(n11405), .ZN(n13997) );
  OR2_X1 U11818 ( .A1(n11170), .A2(n20963), .ZN(n11970) );
  NAND2_X1 U11819 ( .A1(n12148), .A2(n20446), .ZN(n13193) );
  OR2_X1 U11820 ( .A1(n11246), .A2(n11245), .ZN(n14010) );
  NAND2_X1 U11821 ( .A1(n10009), .A2(n9656), .ZN(n13204) );
  INV_X1 U11822 ( .A(n12148), .ZN(n10009) );
  NAND2_X1 U11823 ( .A1(n11092), .A2(n20438), .ZN(n11093) );
  NAND2_X1 U11824 ( .A1(n11168), .A2(n11165), .ZN(n11130) );
  OR2_X1 U11825 ( .A1(n9927), .A2(n10846), .ZN(n9926) );
  INV_X1 U11826 ( .A(n10820), .ZN(n9927) );
  NOR2_X1 U11827 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14440) );
  INV_X1 U11828 ( .A(n13807), .ZN(n14595) );
  INV_X1 U11829 ( .A(n14544), .ZN(n10000) );
  INV_X1 U11830 ( .A(n10178), .ZN(n9982) );
  AND2_X1 U11831 ( .A1(n10254), .A2(n10253), .ZN(n10256) );
  AOI21_X1 U11832 ( .B1(n9692), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A(n10260), .ZN(n10265) );
  OR2_X1 U11833 ( .A1(n10621), .A2(n10620), .ZN(n10811) );
  NOR2_X1 U11834 ( .A1(n9859), .A2(n12533), .ZN(n9858) );
  OAI211_X1 U11835 ( .C1(n19993), .C2(n12597), .A(n10456), .B(n10455), .ZN(
        n10457) );
  AND4_X1 U11836 ( .A1(n10644), .A2(n10643), .A3(n10642), .A4(n10641), .ZN(
        n10660) );
  OR2_X1 U11837 ( .A1(n10310), .A2(n10044), .ZN(n10340) );
  NOR2_X1 U11838 ( .A1(n20220), .A2(n20208), .ZN(n10044) );
  OAI21_X1 U11839 ( .B1(n10295), .B2(n13078), .A(n10294), .ZN(n13012) );
  NAND2_X1 U11840 ( .A1(n10293), .A2(n13078), .ZN(n10294) );
  NAND2_X1 U11841 ( .A1(n19545), .A2(n10296), .ZN(n10308) );
  NAND2_X1 U11842 ( .A1(n13263), .A2(n10386), .ZN(n10547) );
  NAND2_X1 U11843 ( .A1(n10416), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10271) );
  AND4_X1 U11844 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(n10261), .ZN(
        n10233) );
  NAND2_X1 U11845 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10231) );
  NAND2_X1 U11846 ( .A1(n9868), .A2(n9737), .ZN(n9867) );
  AND2_X1 U11847 ( .A1(n10205), .A2(n10203), .ZN(n9866) );
  INV_X1 U11848 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10153) );
  NAND2_X1 U11849 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n9797) );
  AOI21_X1 U11850 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18942), .A(
        n12319), .ZN(n12321) );
  NOR2_X1 U11851 ( .A1(n12429), .A2(n12326), .ZN(n12319) );
  AND2_X1 U11852 ( .A1(n11924), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11925) );
  NAND2_X1 U11853 ( .A1(n10032), .A2(n14680), .ZN(n10031) );
  INV_X1 U11854 ( .A(n14669), .ZN(n10032) );
  NOR2_X1 U11855 ( .A1(n11776), .A2(n14721), .ZN(n11803) );
  NOR2_X1 U11856 ( .A1(n10026), .A2(n14813), .ZN(n10025) );
  INV_X1 U11857 ( .A(n14956), .ZN(n10026) );
  NAND2_X1 U11858 ( .A1(n11498), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11504) );
  AND2_X1 U11859 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n11441), .ZN(
        n11442) );
  NAND2_X1 U11860 ( .A1(n12109), .A2(n9883), .ZN(n9882) );
  NOR2_X1 U11861 ( .A1(n9884), .A2(n14704), .ZN(n9883) );
  INV_X1 U11862 ( .A(n14688), .ZN(n9884) );
  NOR2_X1 U11863 ( .A1(n9685), .A2(n15009), .ZN(n9977) );
  INV_X1 U11864 ( .A(n12112), .ZN(n12106) );
  NOR2_X1 U11865 ( .A1(n14025), .A2(n14024), .ZN(n14023) );
  INV_X1 U11866 ( .A(n13995), .ZN(n9963) );
  AND2_X1 U11867 ( .A1(n11437), .A2(n11416), .ZN(n9811) );
  INV_X1 U11868 ( .A(n11436), .ZN(n11437) );
  OR2_X1 U11869 ( .A1(n11349), .A2(n11348), .ZN(n13988) );
  INV_X1 U11870 ( .A(n12105), .ZN(n12053) );
  NAND2_X1 U11871 ( .A1(n12472), .A2(n9742), .ZN(n9876) );
  NAND2_X1 U11872 ( .A1(n9875), .A2(n12472), .ZN(n9874) );
  AND2_X1 U11873 ( .A1(n12024), .A2(n9774), .ZN(n9873) );
  OR2_X1 U11874 ( .A1(n11259), .A2(n11258), .ZN(n13641) );
  NAND2_X1 U11875 ( .A1(n11320), .A2(n20963), .ZN(n11313) );
  NAND2_X1 U11876 ( .A1(n20446), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11334) );
  NAND2_X1 U11877 ( .A1(n11170), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11335) );
  OR2_X1 U11878 ( .A1(n13194), .A2(n13853), .ZN(n13224) );
  NAND2_X1 U11879 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11046) );
  INV_X1 U11880 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20787) );
  INV_X1 U11881 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20722) );
  AND2_X1 U11882 ( .A1(n11999), .A2(n14005), .ZN(n11998) );
  AOI221_X1 U11883 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n11961), 
        .C1(n16422), .C2(n11961), .A(n11960), .ZN(n12015) );
  OR2_X1 U11884 ( .A1(n10675), .A2(n10674), .ZN(n12967) );
  AND3_X1 U11885 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10679), .A3(
        n13026), .ZN(n12972) );
  NAND2_X1 U11886 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9839) );
  NAND2_X1 U11887 ( .A1(n10969), .A2(n15553), .ZN(n10971) );
  NAND2_X1 U11888 ( .A1(n10967), .A2(n9732), .ZN(n10970) );
  NAND2_X1 U11889 ( .A1(n10911), .A2(n9781), .ZN(n10901) );
  NAND2_X1 U11890 ( .A1(n10879), .A2(n9930), .ZN(n10891) );
  AND2_X1 U11891 ( .A1(n21083), .A2(n10704), .ZN(n9930) );
  NAND2_X1 U11892 ( .A1(n10891), .A2(n10967), .ZN(n10888) );
  NOR2_X1 U11893 ( .A1(n10847), .A2(n9926), .ZN(n10866) );
  NAND2_X1 U11894 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10073) );
  NAND2_X1 U11895 ( .A1(n9663), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10072) );
  NAND2_X1 U11896 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10071) );
  NAND2_X1 U11897 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U11898 ( .A1(n14590), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14412) );
  NAND2_X1 U11899 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10049) );
  NAND2_X1 U11900 ( .A1(n10048), .A2(n10047), .ZN(n10367) );
  AND2_X1 U11901 ( .A1(n15486), .A2(n15471), .ZN(n12754) );
  AND2_X1 U11902 ( .A1(n15585), .A2(n15580), .ZN(n10007) );
  NOR2_X1 U11903 ( .A1(n10102), .A2(n12591), .ZN(n10101) );
  INV_X1 U11904 ( .A(n16563), .ZN(n10102) );
  NAND2_X1 U11905 ( .A1(n10318), .A2(n10317), .ZN(n12999) );
  INV_X1 U11906 ( .A(n13072), .ZN(n10317) );
  NAND2_X1 U11907 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10067) );
  NAND2_X1 U11908 ( .A1(n10062), .A2(n10061), .ZN(n10749) );
  NAND2_X1 U11909 ( .A1(n9663), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10056) );
  NAND2_X1 U11910 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10055) );
  NOR2_X1 U11911 ( .A1(n19262), .A2(n9838), .ZN(n9837) );
  INV_X1 U11912 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n9838) );
  NOR2_X1 U11913 ( .A1(n15882), .A2(n14612), .ZN(n10163) );
  AND2_X1 U11914 ( .A1(n10958), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10959) );
  AND2_X1 U11915 ( .A1(n10933), .A2(n15824), .ZN(n9918) );
  AOI21_X1 U11916 ( .B1(n9862), .B2(n10083), .A(n9766), .ZN(n9861) );
  INV_X1 U11917 ( .A(n9733), .ZN(n9862) );
  INV_X1 U11918 ( .A(n10083), .ZN(n9863) );
  OR2_X1 U11919 ( .A1(n19188), .A2(n10869), .ZN(n10941) );
  AND2_X1 U11920 ( .A1(n15811), .A2(n15813), .ZN(n15771) );
  OR2_X1 U11921 ( .A1(n10108), .A2(n10107), .ZN(n10106) );
  INV_X1 U11922 ( .A(n12819), .ZN(n10107) );
  INV_X1 U11923 ( .A(n10736), .ZN(n12788) );
  AOI21_X1 U11924 ( .B1(n10086), .B2(n10088), .A(n10084), .ZN(n10083) );
  INV_X1 U11925 ( .A(n15860), .ZN(n10084) );
  INV_X1 U11926 ( .A(n10089), .ZN(n10088) );
  INV_X1 U11927 ( .A(n16516), .ZN(n9819) );
  NAND2_X1 U11928 ( .A1(n10519), .A2(n10518), .ZN(n10533) );
  NAND2_X1 U11929 ( .A1(n10508), .A2(n10507), .ZN(n10538) );
  NAND2_X1 U11930 ( .A1(n10373), .A2(n10378), .ZN(n9826) );
  NAND2_X1 U11931 ( .A1(n10041), .A2(n10356), .ZN(n9827) );
  INV_X1 U11932 ( .A(n10363), .ZN(n10043) );
  INV_X1 U11933 ( .A(n10362), .ZN(n10042) );
  AND2_X1 U11934 ( .A1(n10812), .A2(n13235), .ZN(n10831) );
  NOR2_X1 U11935 ( .A1(n10473), .A2(n10112), .ZN(n12540) );
  NAND2_X1 U11936 ( .A1(n10696), .A2(n9916), .ZN(n12554) );
  NOR2_X1 U11937 ( .A1(n14477), .A2(n13145), .ZN(n13153) );
  INV_X1 U11938 ( .A(n10284), .ZN(n13807) );
  INV_X1 U11939 ( .A(n10308), .ZN(n13073) );
  NOR2_X1 U11940 ( .A1(n13689), .A2(n10404), .ZN(n10394) );
  INV_X1 U11941 ( .A(n10392), .ZN(n10379) );
  AND3_X1 U11942 ( .A1(n10244), .A2(n10243), .A3(n10261), .ZN(n10246) );
  NAND2_X1 U11943 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10248) );
  AOI21_X1 U11944 ( .B1(n9692), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A(n9919), 
        .ZN(n10251) );
  AND2_X1 U11945 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n9919) );
  NAND3_X1 U11946 ( .A1(n19989), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20039), 
        .ZN(n19518) );
  AND2_X1 U11947 ( .A1(n20208), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10682) );
  INV_X1 U11948 ( .A(n17807), .ZN(n9938) );
  NAND2_X1 U11949 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n17147), .ZN(
        n12178) );
  INV_X1 U11950 ( .A(n12179), .ZN(n9849) );
  INV_X1 U11951 ( .A(n12180), .ZN(n9848) );
  OR2_X1 U11952 ( .A1(n17176), .A2(n14265), .ZN(n9721) );
  NOR2_X1 U11953 ( .A1(n12181), .A2(n17175), .ZN(n12335) );
  NOR2_X1 U11954 ( .A1(n9949), .A2(n9951), .ZN(n9948) );
  INV_X1 U11955 ( .A(n10174), .ZN(n9951) );
  INV_X1 U11956 ( .A(n9950), .ZN(n9949) );
  NOR2_X1 U11957 ( .A1(n21234), .A2(n18121), .ZN(n9950) );
  NAND2_X1 U11958 ( .A1(n10152), .A2(n9892), .ZN(n9893) );
  AND2_X1 U11959 ( .A1(n12086), .A2(n12085), .ZN(n14775) );
  AND2_X1 U11960 ( .A1(n11928), .A2(n15145), .ZN(n11650) );
  NAND2_X1 U11961 ( .A1(n12472), .A2(n12105), .ZN(n13325) );
  INV_X1 U11962 ( .A(n13110), .ZN(n13388) );
  NOR2_X1 U11963 ( .A1(n10033), .A2(n10031), .ZN(n10030) );
  INV_X1 U11964 ( .A(n14317), .ZN(n10033) );
  INV_X1 U11965 ( .A(n12140), .ZN(n10028) );
  INV_X1 U11966 ( .A(n12021), .ZN(n11955) );
  OAI21_X1 U11967 ( .B1(n10196), .B2(n15076), .A(n11850), .ZN(n14692) );
  AND2_X1 U11968 ( .A1(n10015), .A2(n10014), .ZN(n10013) );
  INV_X1 U11969 ( .A(n14717), .ZN(n10014) );
  AND2_X1 U11970 ( .A1(n11720), .A2(n11719), .ZN(n14758) );
  OR2_X1 U11971 ( .A1(n15121), .A2(n10196), .ZN(n11719) );
  NOR2_X1 U11972 ( .A1(n11649), .A2(n16277), .ZN(n11670) );
  OR2_X1 U11973 ( .A1(n11629), .A2(n15167), .ZN(n11649) );
  NAND2_X1 U11974 ( .A1(n11613), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11629) );
  NOR2_X1 U11975 ( .A1(n21218), .A2(n11557), .ZN(n11613) );
  NOR2_X1 U11976 ( .A1(n11538), .A2(n16293), .ZN(n11556) );
  INV_X1 U11977 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16293) );
  AND2_X1 U11978 ( .A1(n14980), .A2(n14981), .ZN(n14982) );
  NOR2_X1 U11979 ( .A1(n11504), .A2(n15200), .ZN(n11505) );
  NAND2_X1 U11980 ( .A1(n11505), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11538) );
  AND3_X1 U11981 ( .A1(n11483), .A2(n11482), .A3(n11481), .ZN(n13944) );
  AND2_X1 U11982 ( .A1(n11462), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11498) );
  AND2_X1 U11983 ( .A1(n11442), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11462) );
  AOI21_X1 U11984 ( .B1(n13996), .B2(n11590), .A(n11434), .ZN(n13837) );
  INV_X1 U11985 ( .A(n11409), .ZN(n11410) );
  INV_X1 U11986 ( .A(n13706), .ZN(n11413) );
  INV_X1 U11987 ( .A(n13444), .ZN(n11414) );
  NAND2_X1 U11988 ( .A1(n11384), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11409) );
  NAND2_X1 U11989 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11356) );
  NOR2_X1 U11990 ( .A1(n11356), .A2(n11355), .ZN(n11384) );
  INV_X1 U11991 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11355) );
  NOR3_X1 U11992 ( .A1(n14720), .A2(n9882), .A3(n14319), .ZN(n14318) );
  OR2_X1 U11993 ( .A1(n9685), .A2(n15251), .ZN(n15021) );
  NOR2_X1 U11994 ( .A1(n14720), .A2(n9881), .ZN(n14690) );
  INV_X1 U11995 ( .A(n9883), .ZN(n9881) );
  OR2_X1 U11996 ( .A1(n14728), .A2(n14718), .ZN(n14720) );
  NOR2_X1 U11997 ( .A1(n14720), .A2(n14704), .ZN(n14703) );
  NOR2_X1 U11998 ( .A1(n14761), .A2(n14744), .ZN(n14745) );
  NAND2_X1 U11999 ( .A1(n14745), .A2(n14729), .ZN(n14728) );
  NAND2_X1 U12000 ( .A1(n15013), .A2(n15011), .ZN(n15107) );
  NAND2_X1 U12001 ( .A1(n14788), .A2(n14775), .ZN(n14774) );
  OR2_X1 U12002 ( .A1(n14774), .A2(n14759), .ZN(n14761) );
  AND2_X1 U12003 ( .A1(n12083), .A2(n12082), .ZN(n14789) );
  NOR2_X1 U12004 ( .A1(n14801), .A2(n14789), .ZN(n14788) );
  OAI21_X1 U12005 ( .B1(n15010), .B2(n9978), .A(n9976), .ZN(n15014) );
  AND2_X1 U12006 ( .A1(n12078), .A2(n12077), .ZN(n15365) );
  AND2_X1 U12007 ( .A1(n14879), .A2(n14878), .ZN(n14881) );
  OR2_X1 U12008 ( .A1(n9685), .A2(n15008), .ZN(n15173) );
  NOR2_X1 U12009 ( .A1(n14851), .A2(n14836), .ZN(n14879) );
  NAND2_X1 U12010 ( .A1(n10175), .A2(n9885), .ZN(n14851) );
  AND2_X1 U12011 ( .A1(n9765), .A2(n9886), .ZN(n9885) );
  INV_X1 U12012 ( .A(n14849), .ZN(n9886) );
  NAND2_X1 U12013 ( .A1(n10175), .A2(n9765), .ZN(n15399) );
  AND2_X1 U12014 ( .A1(n10175), .A2(n14893), .ZN(n15401) );
  AND2_X1 U12015 ( .A1(n14023), .A2(n12060), .ZN(n10175) );
  INV_X1 U12016 ( .A(n14031), .ZN(n12060) );
  AND2_X1 U12017 ( .A1(n12052), .A2(n12051), .ZN(n13822) );
  NOR2_X1 U12018 ( .A1(n9879), .A2(n13825), .ZN(n9878) );
  INV_X1 U12019 ( .A(n9880), .ZN(n9879) );
  NAND2_X1 U12020 ( .A1(n12043), .A2(n9880), .ZN(n16401) );
  NAND2_X1 U12021 ( .A1(n12043), .A2(n12042), .ZN(n16399) );
  NAND2_X1 U12022 ( .A1(n20361), .A2(n13985), .ZN(n16343) );
  NAND2_X1 U12023 ( .A1(n16343), .A2(n16342), .ZN(n16341) );
  NAND2_X1 U12024 ( .A1(n13471), .A2(n13448), .ZN(n13737) );
  NAND4_X1 U12025 ( .A1(n9958), .A2(n9961), .A3(n9956), .A4(n9955), .ZN(n13673) );
  NAND2_X1 U12026 ( .A1(n9962), .A2(n20387), .ZN(n9961) );
  NAND2_X1 U12027 ( .A1(n13673), .A2(n13672), .ZN(n13978) );
  NAND2_X1 U12028 ( .A1(n12032), .A2(n12031), .ZN(n13469) );
  AND2_X1 U12029 ( .A1(n16364), .A2(n14016), .ZN(n20372) );
  NAND2_X1 U12030 ( .A1(n11317), .A2(n11316), .ZN(n11318) );
  NAND2_X1 U12031 ( .A1(n20522), .A2(n11289), .ZN(n20467) );
  NAND2_X1 U12032 ( .A1(n11297), .A2(n11296), .ZN(n11299) );
  AND2_X1 U12033 ( .A1(n13200), .A2(n13199), .ZN(n13583) );
  NAND2_X1 U12034 ( .A1(n13626), .A2(n13627), .ZN(n20526) );
  INV_X1 U12035 ( .A(n20721), .ZN(n20850) );
  OR2_X1 U12036 ( .A1(n13627), .A2(n11352), .ZN(n20641) );
  OR2_X1 U12037 ( .A1(n13626), .A2(n13628), .ZN(n20697) );
  INV_X1 U12038 ( .A(n13302), .ZN(n20784) );
  INV_X1 U12039 ( .A(n20700), .ZN(n20819) );
  OR2_X1 U12040 ( .A1(n13627), .A2(n13629), .ZN(n20851) );
  AOI21_X1 U12041 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20820), .A(n20557), 
        .ZN(n20908) );
  OR2_X1 U12042 ( .A1(n20851), .A2(n20850), .ZN(n20859) );
  NAND3_X1 U12043 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20963), .A3(n20423), 
        .ZN(n20458) );
  INV_X1 U12044 ( .A(n16615), .ZN(n20220) );
  INV_X1 U12045 ( .A(n12963), .ZN(n13082) );
  NOR2_X1 U12046 ( .A1(n10979), .A2(n10978), .ZN(n12519) );
  NAND2_X1 U12047 ( .A1(n10970), .A2(n10975), .ZN(n10979) );
  NAND2_X1 U12048 ( .A1(n10932), .A2(n10817), .ZN(n10956) );
  OR2_X1 U12049 ( .A1(n10931), .A2(n10932), .ZN(n19161) );
  AND2_X1 U12050 ( .A1(n10896), .A2(n10898), .ZN(n19201) );
  NAND2_X1 U12051 ( .A1(n10916), .A2(n10815), .ZN(n10920) );
  AND2_X1 U12052 ( .A1(n10917), .A2(n10919), .ZN(n19227) );
  NAND2_X1 U12053 ( .A1(n9923), .A2(n10868), .ZN(n9922) );
  INV_X1 U12054 ( .A(n9924), .ZN(n9923) );
  NAND2_X1 U12055 ( .A1(n10074), .A2(n10073), .ZN(n10786) );
  NAND2_X1 U12056 ( .A1(n10070), .A2(n10069), .ZN(n10775) );
  INV_X1 U12057 ( .A(n19506), .ZN(n10404) );
  NAND2_X1 U12058 ( .A1(n10081), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10080) );
  NAND2_X1 U12059 ( .A1(n15472), .A2(n9783), .ZN(n15611) );
  XNOR2_X1 U12060 ( .A(n14503), .B(n14504), .ZN(n15552) );
  NAND2_X1 U12061 ( .A1(n15472), .A2(n10104), .ZN(n15627) );
  NAND2_X1 U12062 ( .A1(n9984), .A2(n10178), .ZN(n15555) );
  INV_X1 U12063 ( .A(n15566), .ZN(n9984) );
  NAND2_X1 U12064 ( .A1(n15472), .A2(n12754), .ZN(n15625) );
  OAI211_X1 U12065 ( .C1(n14368), .C2(n14461), .A(n10003), .B(n10001), .ZN(
        n15568) );
  NAND2_X1 U12066 ( .A1(n14482), .A2(n10004), .ZN(n10003) );
  NOR2_X1 U12067 ( .A1(n14482), .A2(n10004), .ZN(n10002) );
  AND2_X1 U12068 ( .A1(n12746), .A2(n12745), .ZN(n15667) );
  CLKBUF_X1 U12069 ( .A(n14127), .Z(n13912) );
  NOR2_X1 U12070 ( .A1(n9995), .A2(n9993), .ZN(n9992) );
  INV_X1 U12071 ( .A(n13928), .ZN(n9993) );
  NOR2_X1 U12072 ( .A1(n16125), .A2(n10108), .ZN(n16099) );
  AND2_X1 U12073 ( .A1(n16564), .A2(n10101), .ZN(n16166) );
  OAI21_X1 U12074 ( .B1(n12808), .B2(n12807), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12872) );
  OR2_X1 U12075 ( .A1(n12529), .A2(n12528), .ZN(n13957) );
  NOR2_X1 U12076 ( .A1(n13681), .A2(n10097), .ZN(n13956) );
  NAND2_X1 U12077 ( .A1(n10096), .A2(n9709), .ZN(n10097) );
  INV_X1 U12078 ( .A(n12872), .ZN(n19519) );
  NOR2_X1 U12079 ( .A1(n12511), .A2(n15714), .ZN(n12513) );
  NAND2_X1 U12080 ( .A1(n9834), .A2(n9833), .ZN(n9832) );
  NOR2_X1 U12081 ( .A1(n9835), .A2(n15736), .ZN(n9833) );
  INV_X1 U12082 ( .A(n10796), .ZN(n9834) );
  NAND2_X1 U12083 ( .A1(n10068), .A2(n10067), .ZN(n10772) );
  NOR2_X1 U12084 ( .A1(n15485), .A2(n10125), .ZN(n15563) );
  INV_X1 U12085 ( .A(n10127), .ZN(n10125) );
  INV_X1 U12086 ( .A(n10123), .ZN(n14104) );
  AND2_X1 U12087 ( .A1(n13931), .A2(n13930), .ZN(n13933) );
  NAND2_X1 U12088 ( .A1(n10064), .A2(n10063), .ZN(n10752) );
  NOR2_X1 U12089 ( .A1(n13620), .A2(n12816), .ZN(n13931) );
  NAND2_X1 U12090 ( .A1(n10060), .A2(n10059), .ZN(n10740) );
  AND2_X1 U12091 ( .A1(n9711), .A2(n13352), .ZN(n10116) );
  NAND2_X1 U12092 ( .A1(n10118), .A2(n10119), .ZN(n13526) );
  NAND2_X1 U12093 ( .A1(n10058), .A2(n10057), .ZN(n10724) );
  INV_X1 U12094 ( .A(n10636), .ZN(n13952) );
  XNOR2_X1 U12095 ( .A(n10514), .B(n10696), .ZN(n14631) );
  INV_X1 U12096 ( .A(n10163), .ZN(n10162) );
  NAND2_X1 U12097 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10161) );
  NAND2_X1 U12098 ( .A1(n10163), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10159) );
  NOR2_X2 U12099 ( .A1(n15720), .A2(n9830), .ZN(n15713) );
  NAND2_X1 U12100 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9830) );
  OR2_X1 U12101 ( .A1(n15699), .A2(n9915), .ZN(n9913) );
  INV_X1 U12102 ( .A(n10092), .ZN(n15734) );
  NAND2_X1 U12103 ( .A1(n9851), .A2(n9854), .ZN(n15758) );
  NOR2_X1 U12104 ( .A1(n15485), .A2(n15469), .ZN(n15561) );
  NAND2_X1 U12105 ( .A1(n10066), .A2(n10065), .ZN(n10764) );
  NAND2_X1 U12106 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10065) );
  OAI21_X1 U12107 ( .B1(n19161), .B2(n10869), .A(n15781), .ZN(n15775) );
  NAND2_X1 U12108 ( .A1(n10123), .A2(n10122), .ZN(n15588) );
  INV_X1 U12109 ( .A(n14103), .ZN(n10122) );
  NAND2_X1 U12110 ( .A1(n10130), .A2(n10129), .ZN(n13620) );
  INV_X1 U12111 ( .A(n13617), .ZN(n10129) );
  NAND2_X1 U12112 ( .A1(n14233), .A2(n16519), .ZN(n15872) );
  NAND2_X1 U12113 ( .A1(n14231), .A2(n10877), .ZN(n9820) );
  NAND2_X1 U12114 ( .A1(n10052), .A2(n10051), .ZN(n10728) );
  NOR2_X1 U12115 ( .A1(n13277), .A2(n13256), .ZN(n13527) );
  NAND2_X1 U12116 ( .A1(n10637), .A2(n10819), .ZN(n9822) );
  NAND2_X1 U12117 ( .A1(n10039), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10860) );
  OAI21_X1 U12118 ( .B1(n10859), .B2(n14277), .A(n19301), .ZN(n10039) );
  NAND2_X1 U12119 ( .A1(n10054), .A2(n10053), .ZN(n10720) );
  AND2_X1 U12120 ( .A1(n13091), .A2(n13080), .ZN(n16046) );
  OR2_X1 U12121 ( .A1(n13681), .A2(n10099), .ZN(n13553) );
  NAND2_X1 U12122 ( .A1(n10096), .A2(n13455), .ZN(n10099) );
  NAND2_X1 U12123 ( .A1(n13240), .A2(n13174), .ZN(n13260) );
  CLKBUF_X1 U12124 ( .A(n10339), .Z(n13696) );
  NAND2_X1 U12125 ( .A1(n13057), .A2(n12979), .ZN(n16597) );
  NOR2_X1 U12126 ( .A1(n13689), .A2(n19506), .ZN(n10395) );
  AND2_X1 U12127 ( .A1(n20177), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19749) );
  AND2_X1 U12128 ( .A1(n20177), .A2(n20203), .ZN(n19719) );
  NAND2_X1 U12129 ( .A1(n19520), .A2(n19657), .ZN(n19831) );
  INV_X1 U12130 ( .A(n12989), .ZN(n19549) );
  AND2_X1 U12131 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19987), .ZN(
        n13161) );
  NAND2_X1 U12132 ( .A1(n19521), .A2(n19784), .ZN(n19962) );
  NOR2_X1 U12133 ( .A1(n20177), .A2(n19784), .ZN(n19986) );
  NAND2_X1 U12134 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20039), .ZN(n19565) );
  NOR2_X2 U12135 ( .A1(n19517), .A2(n19518), .ZN(n19564) );
  AND2_X1 U12136 ( .A1(n9934), .A2(n9932), .ZN(n16895) );
  NOR2_X1 U12137 ( .A1(n9933), .A2(n17144), .ZN(n9932) );
  INV_X1 U12138 ( .A(n9935), .ZN(n9933) );
  NAND2_X1 U12139 ( .A1(n17144), .A2(n9938), .ZN(n9935) );
  OR2_X1 U12140 ( .A1(n16915), .A2(n9936), .ZN(n9934) );
  NAND2_X1 U12141 ( .A1(n9938), .A2(n9937), .ZN(n9936) );
  INV_X1 U12142 ( .A(n17827), .ZN(n9937) );
  NOR2_X1 U12143 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17029), .ZN(n17016) );
  INV_X1 U12144 ( .A(n12372), .ZN(n9799) );
  NOR2_X1 U12145 ( .A1(n9798), .A2(n9796), .ZN(n9795) );
  NOR2_X1 U12146 ( .A1(n17641), .A2(n17640), .ZN(n17672) );
  NAND2_X1 U12147 ( .A1(n12458), .A2(n9948), .ZN(n16810) );
  NAND2_X1 U12148 ( .A1(n12458), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17758) );
  NAND2_X1 U12149 ( .A1(n17903), .A2(n9945), .ZN(n17794) );
  AND2_X1 U12150 ( .A1(n9716), .A2(n9776), .ZN(n9945) );
  NOR2_X1 U12151 ( .A1(n18265), .A2(n17806), .ZN(n17828) );
  NOR2_X1 U12152 ( .A1(n18126), .A2(n18079), .ZN(n17841) );
  NOR2_X1 U12153 ( .A1(n17906), .A2(n16996), .ZN(n17877) );
  INV_X1 U12154 ( .A(n17876), .ZN(n17879) );
  INV_X1 U12155 ( .A(n17880), .ZN(n17976) );
  NOR2_X1 U12156 ( .A1(n18061), .A2(n18062), .ZN(n18029) );
  NOR2_X1 U12157 ( .A1(n17819), .A2(n9889), .ZN(n17815) );
  INV_X1 U12158 ( .A(n12299), .ZN(n9889) );
  OAI21_X1 U12159 ( .B1(n17914), .B2(n17806), .A(n12298), .ZN(n12299) );
  NOR2_X1 U12160 ( .A1(n18322), .A2(n18267), .ZN(n17950) );
  INV_X1 U12161 ( .A(n18323), .ZN(n18301) );
  INV_X1 U12162 ( .A(n17939), .ZN(n18324) );
  NAND2_X1 U12163 ( .A1(n9893), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9894) );
  NAND2_X1 U12164 ( .A1(n12290), .A2(n9890), .ZN(n18037) );
  OAI21_X1 U12165 ( .B1(n9892), .B2(n18360), .A(n18038), .ZN(n9891) );
  INV_X1 U12166 ( .A(n10149), .ZN(n12276) );
  NOR2_X1 U12167 ( .A1(n18108), .A2(n18107), .ZN(n18106) );
  INV_X1 U12168 ( .A(n18303), .ZN(n18906) );
  NAND2_X1 U12169 ( .A1(n12419), .A2(n12422), .ZN(n14250) );
  INV_X1 U12170 ( .A(n12408), .ZN(n12416) );
  OAI21_X1 U12171 ( .B1(n12332), .B2(n12426), .A(n12427), .ZN(n16786) );
  INV_X1 U12172 ( .A(n18924), .ZN(n18933) );
  AND2_X1 U12173 ( .A1(n9845), .A2(n14249), .ZN(n16822) );
  INV_X1 U12174 ( .A(n14250), .ZN(n9845) );
  NOR2_X1 U12175 ( .A1(n12355), .A2(n12354), .ZN(n18491) );
  NOR2_X1 U12176 ( .A1(n12345), .A2(n12344), .ZN(n18497) );
  NOR2_X1 U12177 ( .A1(n12394), .A2(n12393), .ZN(n18503) );
  NOR2_X1 U12178 ( .A1(n12384), .A2(n12383), .ZN(n18510) );
  NAND2_X1 U12179 ( .A1(n21075), .A2(n18473), .ZN(n18597) );
  INV_X1 U12180 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19123) );
  NOR2_X1 U12181 ( .A1(n18970), .A2(n19123), .ZN(n19107) );
  AND2_X1 U12182 ( .A1(n20261), .A2(n12134), .ZN(n20339) );
  NAND2_X1 U12183 ( .A1(n12133), .A2(n12132), .ZN(n20308) );
  INV_X1 U12184 ( .A(n14896), .ZN(n20351) );
  INV_X1 U12185 ( .A(n20356), .ZN(n14885) );
  NAND2_X1 U12186 ( .A1(n20356), .A2(n20457), .ZN(n14896) );
  AND2_X2 U12187 ( .A1(n13106), .A2(n13290), .ZN(n20356) );
  OR2_X1 U12188 ( .A1(n12171), .A2(n20421), .ZN(n14962) );
  INV_X1 U12189 ( .A(n14995), .ZN(n14964) );
  INV_X1 U12190 ( .A(n14962), .ZN(n14969) );
  AND2_X1 U12191 ( .A1(n12158), .A2(n13290), .ZN(n14988) );
  NAND2_X1 U12192 ( .A1(n13188), .A2(n12157), .ZN(n12158) );
  OAI21_X1 U12193 ( .B1(n13269), .B2(n13268), .A(n13758), .ZN(n13512) );
  NOR2_X1 U12194 ( .A1(n13512), .A2(n21051), .ZN(n16264) );
  INV_X1 U12195 ( .A(n13512), .ZN(n13783) );
  INV_X1 U12196 ( .A(n13357), .ZN(n13400) );
  OAI21_X1 U12197 ( .B1(n14316), .B2(n14317), .A(n12141), .ZN(n15047) );
  AND2_X1 U12198 ( .A1(n11876), .A2(n11853), .ZN(n15065) );
  AND2_X1 U12199 ( .A1(n11717), .A2(n11695), .ZN(n15130) );
  INV_X1 U12200 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21227) );
  INV_X1 U12201 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16277) );
  INV_X1 U12202 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15167) );
  INV_X1 U12203 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n21218) );
  INV_X1 U12204 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15200) );
  NAND2_X1 U12205 ( .A1(n10012), .A2(n10010), .ZN(n13427) );
  OR2_X1 U12206 ( .A1(n13332), .A2(n16229), .ZN(n20363) );
  INV_X1 U12207 ( .A(n20363), .ZN(n16345) );
  NAND2_X1 U12208 ( .A1(n9669), .A2(n9805), .ZN(n9804) );
  XNOR2_X1 U12209 ( .A(n9964), .B(n15023), .ZN(n15235) );
  NAND2_X1 U12210 ( .A1(n9967), .A2(n9965), .ZN(n9964) );
  NAND2_X1 U12211 ( .A1(n15022), .A2(n9708), .ZN(n9967) );
  OR3_X1 U12212 ( .A1(n15288), .A2(n15270), .A3(n15210), .ZN(n15260) );
  NOR2_X1 U12213 ( .A1(n15309), .A2(n15314), .ZN(n20411) );
  AND2_X1 U12214 ( .A1(n13324), .A2(n13323), .ZN(n20406) );
  INV_X1 U12215 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20820) );
  INV_X1 U12216 ( .A(n16247), .ZN(n15422) );
  INV_X1 U12217 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16422) );
  INV_X1 U12218 ( .A(n20960), .ZN(n20460) );
  OR2_X1 U12219 ( .A1(n20526), .A2(n20700), .ZN(n20513) );
  INV_X1 U12220 ( .A(n20572), .ZN(n20577) );
  INV_X1 U12221 ( .A(n20600), .ZN(n20603) );
  INV_X1 U12222 ( .A(n20629), .ZN(n20630) );
  OAI211_X1 U12223 ( .C1(n20689), .C2(n20674), .A(n20727), .B(n20673), .ZN(
        n20692) );
  OAI22_X1 U12224 ( .A1(n20731), .A2(n20730), .B1(n20729), .B2(n20847), .ZN(
        n20748) );
  INV_X1 U12225 ( .A(n20818), .ZN(n20779) );
  OAI22_X1 U12226 ( .A1(n20798), .A2(n20797), .B1(n20796), .B2(n20846), .ZN(
        n20814) );
  NOR2_X2 U12227 ( .A1(n20785), .A2(n20784), .ZN(n20842) );
  INV_X1 U12228 ( .A(n20859), .ZN(n20956) );
  NAND2_X1 U12229 ( .A1(n10292), .A2(n13056), .ZN(n10298) );
  NOR2_X1 U12230 ( .A1(n9722), .A2(n10131), .ZN(n14288) );
  NAND2_X1 U12231 ( .A1(n19183), .A2(n10182), .ZN(n19175) );
  INV_X1 U12232 ( .A(n19215), .ZN(n9843) );
  INV_X1 U12233 ( .A(n12505), .ZN(n19198) );
  AND2_X1 U12234 ( .A1(n20221), .A2(n12522), .ZN(n19317) );
  INV_X1 U12235 ( .A(n19318), .ZN(n19260) );
  INV_X1 U12236 ( .A(n19326), .ZN(n19298) );
  NAND2_X1 U12237 ( .A1(n19260), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19326) );
  OR2_X1 U12238 ( .A1(n15439), .A2(n15438), .ZN(n15703) );
  AND2_X1 U12239 ( .A1(n12739), .A2(n12738), .ZN(n13831) );
  NAND2_X1 U12240 ( .A1(n10714), .A2(n10713), .ZN(n13183) );
  INV_X1 U12241 ( .A(n19314), .ZN(n13699) );
  INV_X1 U12242 ( .A(n9989), .ZN(n9988) );
  OAI21_X1 U12243 ( .B1(n15526), .B2(n9990), .A(n9719), .ZN(n9989) );
  NAND2_X1 U12244 ( .A1(n19371), .A2(n10322), .ZN(n19342) );
  NOR2_X1 U12245 ( .A1(n16125), .A2(n16124), .ZN(n16107) );
  NOR2_X1 U12246 ( .A1(n19404), .A2(n19400), .ZN(n19379) );
  INV_X1 U12247 ( .A(n16479), .ZN(n19404) );
  INV_X1 U12248 ( .A(n19342), .ZN(n19400) );
  OR2_X1 U12249 ( .A1(n19338), .A2(n13006), .ZN(n19365) );
  AND2_X1 U12250 ( .A1(n12837), .A2(n12774), .ZN(n19480) );
  AND2_X1 U12251 ( .A1(n19410), .A2(n12849), .ZN(n19481) );
  INV_X1 U12252 ( .A(n19480), .ZN(n19410) );
  OR2_X1 U12253 ( .A1(n15435), .A2(n16526), .ZN(n14661) );
  INV_X1 U12254 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15864) );
  INV_X1 U12255 ( .A(n19486), .ZN(n16526) );
  AND2_X1 U12256 ( .A1(n16541), .A2(n10798), .ZN(n16533) );
  INV_X1 U12257 ( .A(n16541), .ZN(n19484) );
  AND2_X1 U12258 ( .A1(n10702), .A2(n10292), .ZN(n16529) );
  OAI21_X1 U12259 ( .B1(n15684), .B2(n15687), .A(n10179), .ZN(n14280) );
  NAND2_X1 U12260 ( .A1(n14616), .A2(n19505), .ZN(n14617) );
  XNOR2_X1 U12261 ( .A(n9914), .B(n9736), .ZN(n15906) );
  NAND2_X1 U12262 ( .A1(n9855), .A2(n15757), .ZN(n9852) );
  NAND2_X1 U12263 ( .A1(n15757), .A2(n15973), .ZN(n9853) );
  CLKBUF_X1 U12264 ( .A(n15779), .Z(n15780) );
  NAND2_X1 U12265 ( .A1(n14233), .A2(n10090), .ZN(n10085) );
  CLKBUF_X1 U12266 ( .A(n14069), .Z(n14070) );
  INV_X1 U12267 ( .A(n19502), .ZN(n16568) );
  AND2_X1 U12268 ( .A1(n13091), .A2(n13090), .ZN(n19505) );
  INV_X1 U12269 ( .A(n19515), .ZN(n16550) );
  INV_X1 U12270 ( .A(n19505), .ZN(n16547) );
  AND2_X1 U12271 ( .A1(n13091), .A2(n13404), .ZN(n16045) );
  OR2_X1 U12272 ( .A1(n16045), .A2(n16046), .ZN(n19499) );
  INV_X1 U12273 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20208) );
  INV_X1 U12274 ( .A(n19784), .ZN(n20203) );
  INV_X1 U12275 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20199) );
  INV_X1 U12276 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20190) );
  NAND2_X1 U12277 ( .A1(n13262), .A2(n13261), .ZN(n20177) );
  OR2_X1 U12278 ( .A1(n13260), .A2(n13259), .ZN(n13262) );
  NAND2_X1 U12279 ( .A1(n13159), .A2(n13046), .ZN(n20193) );
  AND2_X1 U12280 ( .A1(n13241), .A2(n13240), .ZN(n20184) );
  NAND2_X1 U12281 ( .A1(n13159), .A2(n13158), .ZN(n13239) );
  INV_X1 U12282 ( .A(n20177), .ZN(n19521) );
  INV_X1 U12283 ( .A(n19666), .ZN(n19684) );
  AND2_X1 U12284 ( .A1(n19723), .A2(n19722), .ZN(n19729) );
  INV_X1 U12285 ( .A(n19729), .ZN(n19746) );
  AOI22_X1 U12286 ( .A1(n19793), .A2(n19792), .B1(n19791), .B2(n19953), .ZN(
        n19817) );
  INV_X1 U12287 ( .A(n19910), .ZN(n19920) );
  INV_X1 U12288 ( .A(n20051), .ZN(n19932) );
  INV_X1 U12289 ( .A(n20045), .ZN(n19988) );
  INV_X1 U12290 ( .A(n20057), .ZN(n20004) );
  INV_X1 U12291 ( .A(n20065), .ZN(n20008) );
  OAI22_X1 U12292 ( .A1(n19559), .A2(n19558), .B1(n19557), .B2(n19556), .ZN(
        n20017) );
  OAI21_X1 U12293 ( .B1(n19998), .B2(n19997), .A(n19996), .ZN(n20023) );
  INV_X1 U12294 ( .A(n19935), .ZN(n20048) );
  INV_X1 U12295 ( .A(n20093), .ZN(n20061) );
  OAI22_X1 U12296 ( .A1(n19544), .A2(n19558), .B1(n19543), .B2(n19556), .ZN(
        n20060) );
  INV_X1 U12297 ( .A(n19974), .ZN(n20068) );
  INV_X1 U12298 ( .A(n19978), .ZN(n20074) );
  INV_X1 U12299 ( .A(n20020), .ZN(n20080) );
  AND2_X1 U12300 ( .A1(n13161), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20085) );
  AND2_X1 U12301 ( .A1(n19986), .A2(n20174), .ZN(n20089) );
  INV_X1 U12302 ( .A(n20028), .ZN(n20088) );
  AND2_X1 U12303 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10700), .ZN(n20095) );
  INV_X1 U12304 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20041) );
  NOR3_X1 U12305 ( .A1(n16615), .A2(n19953), .A3(n16614), .ZN(n20101) );
  NOR2_X1 U12306 ( .A1(n12418), .A2(n18485), .ZN(n16792) );
  NOR3_X2 U12307 ( .A1(n18475), .A2(n17495), .A3(n14255), .ZN(n17706) );
  NAND2_X1 U12308 ( .A1(n9931), .A2(n9942), .ZN(n16842) );
  INV_X1 U12309 ( .A(n9931), .ZN(n16854) );
  NOR2_X1 U12310 ( .A1(n16915), .A2(n17827), .ZN(n16914) );
  INV_X1 U12311 ( .A(n9941), .ZN(n16946) );
  AND2_X1 U12312 ( .A1(n17903), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17876) );
  NOR2_X1 U12313 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17003), .ZN(n16990) );
  INV_X1 U12314 ( .A(n17146), .ZN(n17178) );
  NOR2_X1 U12315 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17096), .ZN(n17083) );
  OR3_X1 U12316 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .A3(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17169) );
  INV_X1 U12317 ( .A(n17168), .ZN(n17182) );
  INV_X1 U12318 ( .A(n17191), .ZN(n17181) );
  OAI211_X1 U12319 ( .C1(n18970), .C2(n18964), .A(n16825), .B(n19126), .ZN(
        n17190) );
  AND3_X1 U12320 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17278), .ZN(n17265) );
  NOR3_X1 U12321 ( .A1(n14135), .A2(n17403), .A3(n17333), .ZN(n17331) );
  NAND2_X1 U12322 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17404), .ZN(n17403) );
  OR2_X1 U12323 ( .A1(n12364), .A2(n12365), .ZN(n17597) );
  INV_X1 U12324 ( .A(n17418), .ZN(n17435) );
  INV_X1 U12325 ( .A(n17597), .ZN(n18518) );
  NAND2_X1 U12326 ( .A1(n17512), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n17506) );
  NAND2_X1 U12327 ( .A1(n17521), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17517) );
  NOR2_X1 U12328 ( .A1(n17527), .A2(n17653), .ZN(n17521) );
  INV_X1 U12329 ( .A(n17548), .ZN(n17544) );
  INV_X1 U12330 ( .A(n17562), .ZN(n17558) );
  AND2_X1 U12331 ( .A1(n17577), .A2(n9846), .ZN(n17579) );
  NOR2_X1 U12332 ( .A1(n17488), .A2(n9847), .ZN(n9846) );
  INV_X1 U12333 ( .A(n17635), .ZN(n17614) );
  NOR2_X1 U12334 ( .A1(n12211), .A2(n12210), .ZN(n17623) );
  INV_X1 U12335 ( .A(n17580), .ZN(n17622) );
  INV_X1 U12336 ( .A(n17630), .ZN(n17635) );
  NOR2_X1 U12337 ( .A1(n18936), .A2(n17622), .ZN(n17636) );
  NOR2_X1 U12338 ( .A1(n12264), .A2(n9896), .ZN(n12271) );
  INV_X1 U12339 ( .A(n17636), .ZN(n17633) );
  CLKBUF_X1 U12340 ( .A(n17688), .Z(n17700) );
  CLKBUF_X1 U12341 ( .A(n17747), .Z(n17750) );
  NOR2_X1 U12342 ( .A1(n17750), .A2(n19112), .ZN(n17751) );
  NAND2_X1 U12343 ( .A1(n17903), .A2(n9714), .ZN(n17864) );
  NAND2_X1 U12344 ( .A1(n18020), .A2(n18237), .ZN(n17927) );
  NAND2_X1 U12345 ( .A1(n17977), .A2(n9771), .ZN(n17946) );
  INV_X1 U12346 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17947) );
  NAND2_X1 U12347 ( .A1(n9802), .A2(n9801), .ZN(n9800) );
  INV_X1 U12348 ( .A(n18322), .ZN(n9801) );
  INV_X1 U12349 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18031) );
  INV_X1 U12350 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18048) );
  NAND2_X1 U12351 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n18073), .ZN(
        n18061) );
  INV_X1 U12352 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18062) );
  NOR2_X1 U12353 ( .A1(n18085), .A2(n18093), .ZN(n18073) );
  INV_X1 U12354 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18093) );
  NAND2_X1 U12355 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18085) );
  INV_X1 U12356 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19075) );
  INV_X1 U12357 ( .A(n18118), .ZN(n18129) );
  INV_X1 U12358 ( .A(n18115), .ZN(n18130) );
  NAND2_X1 U12359 ( .A1(n16639), .A2(n16638), .ZN(n16678) );
  INV_X1 U12360 ( .A(n10140), .ZN(n10139) );
  OAI22_X1 U12361 ( .A1(n9784), .A2(n12305), .B1(n16686), .B2(n10145), .ZN(
        n10140) );
  NAND2_X1 U12362 ( .A1(n10148), .A2(n16683), .ZN(n9904) );
  AND2_X1 U12363 ( .A1(n12301), .A2(n12300), .ZN(n17788) );
  NOR2_X1 U12364 ( .A1(n18921), .A2(n18933), .ZN(n18337) );
  NAND2_X1 U12365 ( .A1(n9901), .A2(n9900), .ZN(n18058) );
  INV_X1 U12366 ( .A(n18455), .ZN(n18441) );
  NOR2_X1 U12367 ( .A1(n18385), .A2(n18451), .ZN(n18445) );
  INV_X1 U12368 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18951) );
  INV_X1 U12369 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18478) );
  INV_X1 U12370 ( .A(n19107), .ZN(n18967) );
  INV_X1 U12371 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19068) );
  CLKBUF_X1 U12372 ( .A(n16778), .Z(n21255) );
  NAND2_X1 U12373 ( .A1(n12138), .A2(n12137), .ZN(n12139) );
  NOR2_X1 U12374 ( .A1(n15040), .A2(n20287), .ZN(n9870) );
  AND2_X1 U12375 ( .A1(n12795), .A2(n12794), .ZN(n12796) );
  NAND2_X1 U12376 ( .A1(n12793), .A2(n19313), .ZN(n12794) );
  OAI21_X1 U12377 ( .B1(n15427), .B2(n16444), .A(n16443), .ZN(n16445) );
  CLKBUF_X3 U12378 ( .A(n14166), .Z(n17411) );
  NAND2_X1 U12379 ( .A1(n10037), .A2(n10176), .ZN(n13821) );
  AND2_X1 U12380 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10417) );
  AND2_X1 U12381 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11008) );
  AND3_X1 U12382 ( .A1(n12303), .A2(n17786), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9705) );
  AND2_X1 U12383 ( .A1(n16147), .A2(n16150), .ZN(n9706) );
  NAND2_X1 U12384 ( .A1(n12497), .A2(n9748), .ZN(n12493) );
  NAND2_X1 U12385 ( .A1(n12497), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12494) );
  NAND2_X1 U12386 ( .A1(n14757), .A2(n10015), .ZN(n14716) );
  NAND2_X1 U12387 ( .A1(n14757), .A2(n14758), .ZN(n14742) );
  NAND2_X1 U12388 ( .A1(n14368), .A2(n10007), .ZN(n15573) );
  OR2_X1 U12389 ( .A1(n12489), .A2(n9762), .ZN(n9707) );
  NAND2_X1 U12390 ( .A1(n15850), .A2(n9788), .ZN(n15793) );
  NAND2_X1 U12391 ( .A1(n10229), .A2(n10228), .ZN(n10302) );
  NAND2_X1 U12392 ( .A1(n18118), .A2(n17605), .ZN(n17971) );
  INV_X1 U12393 ( .A(n17971), .ZN(n9802) );
  AND2_X1 U12394 ( .A1(n9773), .A2(n15021), .ZN(n9708) );
  AND2_X1 U12395 ( .A1(n13455), .A2(n13556), .ZN(n9709) );
  INV_X1 U12396 ( .A(n9864), .ZN(n14233) );
  AND4_X1 U12397 ( .A1(n10321), .A2(n10306), .A3(n10307), .A4(n10322), .ZN(
        n10315) );
  NAND2_X1 U12398 ( .A1(n15751), .A2(n9791), .ZN(n9710) );
  AND2_X1 U12399 ( .A1(n10119), .A2(n10117), .ZN(n9711) );
  NAND2_X1 U12400 ( .A1(n18330), .A2(n18337), .ZN(n18359) );
  INV_X1 U12401 ( .A(n18359), .ZN(n9803) );
  INV_X1 U12402 ( .A(n13736), .ZN(n12042) );
  INV_X1 U12403 ( .A(n14811), .ZN(n10024) );
  OR2_X1 U12404 ( .A1(n10093), .A2(n9759), .ZN(n9713) );
  OR2_X1 U12405 ( .A1(n13621), .A2(n13622), .ZN(n13830) );
  AND2_X1 U12406 ( .A1(n12457), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9714) );
  NOR3_X1 U12407 ( .A1(n12487), .A2(n10796), .A3(n15754), .ZN(n12509) );
  AND2_X1 U12408 ( .A1(n13346), .A2(n13350), .ZN(n9715) );
  AND2_X1 U12409 ( .A1(n9714), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9716) );
  AND2_X1 U12410 ( .A1(n10104), .A2(n10103), .ZN(n9717) );
  NOR2_X1 U12411 ( .A1(n12304), .A2(n9792), .ZN(n9718) );
  OR2_X1 U12412 ( .A1(n14582), .A2(n14604), .ZN(n9719) );
  AND2_X1 U12413 ( .A1(n16002), .A2(n10154), .ZN(n9720) );
  INV_X1 U12414 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12320) );
  OR3_X1 U12415 ( .A1(n15485), .A2(n10126), .A3(n15546), .ZN(n9722) );
  OR2_X1 U12416 ( .A1(n15611), .A2(n12830), .ZN(n9723) );
  AND2_X1 U12417 ( .A1(n12472), .A2(n13107), .ZN(n9724) );
  NAND2_X1 U12418 ( .A1(n15850), .A2(n16002), .ZN(n15816) );
  NAND2_X1 U12419 ( .A1(n15197), .A2(n14998), .ZN(n15149) );
  NAND2_X1 U12420 ( .A1(n9860), .A2(n10083), .ZN(n15763) );
  NOR2_X1 U12421 ( .A1(n12498), .A2(n10719), .ZN(n12496) );
  INV_X1 U12422 ( .A(n12811), .ZN(n19289) );
  INV_X1 U12423 ( .A(n10300), .ZN(n10306) );
  AND2_X1 U12424 ( .A1(n14757), .A2(n10017), .ZN(n9725) );
  AND3_X1 U12425 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12500) );
  AND2_X1 U12426 ( .A1(n12497), .A2(n9837), .ZN(n12495) );
  AND2_X1 U12427 ( .A1(n15751), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15742) );
  AND2_X1 U12428 ( .A1(n10141), .A2(n10139), .ZN(n9726) );
  INV_X1 U12429 ( .A(n15701), .ZN(n9915) );
  NOR2_X1 U12430 ( .A1(n12827), .A2(n10869), .ZN(n15701) );
  AND4_X1 U12431 ( .A1(n12215), .A2(n12214), .A3(n12213), .A4(n12212), .ZN(
        n9727) );
  AND2_X1 U12432 ( .A1(n15850), .A2(n9720), .ZN(n15800) );
  NAND2_X1 U12433 ( .A1(n10024), .A2(n10025), .ZN(n14795) );
  NOR2_X1 U12434 ( .A1(n14811), .A2(n14813), .ZN(n14812) );
  AND2_X1 U12435 ( .A1(n12043), .A2(n9878), .ZN(n9728) );
  AND3_X1 U12436 ( .A1(n10256), .A2(n10255), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9729) );
  OR2_X1 U12437 ( .A1(n14720), .A2(n9882), .ZN(n9730) );
  NAND2_X1 U12438 ( .A1(n10950), .A2(n10949), .ZN(n15975) );
  AND2_X1 U12439 ( .A1(n20446), .A2(n13642), .ZN(n9731) );
  NAND2_X1 U12440 ( .A1(n10085), .A2(n10089), .ZN(n15862) );
  NAND2_X1 U12441 ( .A1(n9849), .A2(n9848), .ZN(n17209) );
  OR2_X1 U12442 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n10971), .ZN(n9732) );
  AND2_X1 U12443 ( .A1(n10086), .A2(n14234), .ZN(n9733) );
  NAND2_X1 U12444 ( .A1(n9669), .A2(n15021), .ZN(n15041) );
  NAND2_X1 U12445 ( .A1(n9821), .A2(n9820), .ZN(n16515) );
  AND3_X1 U12446 ( .A1(n18027), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n9734) );
  NOR2_X1 U12447 ( .A1(n10847), .A2(n9924), .ZN(n9735) );
  XOR2_X1 U12448 ( .A(n15702), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .Z(
        n9736) );
  AND3_X1 U12450 ( .A1(n10200), .A2(n10199), .A3(n10261), .ZN(n9737) );
  AND2_X1 U12451 ( .A1(n12496), .A2(n10792), .ZN(n12497) );
  NAND2_X1 U12452 ( .A1(n15699), .A2(n9915), .ZN(n9912) );
  NAND2_X1 U12453 ( .A1(n15713), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15707) );
  AND2_X1 U12454 ( .A1(n14368), .A2(n10005), .ZN(n9738) );
  OR2_X1 U12455 ( .A1(n14231), .A2(n10877), .ZN(n9739) );
  OR2_X1 U12456 ( .A1(n15485), .A2(n10126), .ZN(n9740) );
  NAND2_X1 U12457 ( .A1(n10024), .A2(n10022), .ZN(n9741) );
  AND2_X1 U12458 ( .A1(n13107), .A2(n12025), .ZN(n9742) );
  AND3_X1 U12459 ( .A1(n10204), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10202), .ZN(n9743) );
  AND2_X1 U12460 ( .A1(n15150), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9744) );
  OR2_X1 U12461 ( .A1(n12274), .A2(n12275), .ZN(n9745) );
  NAND2_X1 U12462 ( .A1(n14237), .A2(n14234), .ZN(n9864) );
  AND2_X1 U12463 ( .A1(n11125), .A2(n11124), .ZN(n9746) );
  INV_X1 U12464 ( .A(n15720), .ZN(n9829) );
  NAND2_X1 U12465 ( .A1(n11130), .A2(n13293), .ZN(n9747) );
  AND2_X1 U12466 ( .A1(n9837), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9748) );
  AND3_X1 U12467 ( .A1(n10276), .A2(n10274), .A3(n10261), .ZN(n9749) );
  AND2_X1 U12468 ( .A1(n10269), .A2(n10268), .ZN(n9750) );
  AND2_X1 U12469 ( .A1(n9810), .A2(n14998), .ZN(n9751) );
  INV_X1 U12470 ( .A(n15973), .ZN(n9856) );
  AND2_X1 U12471 ( .A1(n10321), .A2(n10305), .ZN(n9752) );
  INV_X1 U12472 ( .A(n10147), .ZN(n16626) );
  NAND2_X1 U12473 ( .A1(n10148), .A2(n9718), .ZN(n10147) );
  NAND2_X1 U12474 ( .A1(n9829), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15712) );
  NAND2_X1 U12475 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12285), .ZN(
        n9753) );
  XNOR2_X1 U12476 ( .A(n10638), .B(n10869), .ZN(n14231) );
  OR2_X1 U12477 ( .A1(n10847), .A2(n10846), .ZN(n9928) );
  NAND2_X1 U12478 ( .A1(n13307), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13646) );
  INV_X1 U12479 ( .A(n12284), .ZN(n10137) );
  NAND3_X1 U12480 ( .A1(n16146), .A2(n15871), .A3(n16151), .ZN(n9754) );
  INV_X1 U12481 ( .A(n10091), .ZN(n10090) );
  NAND2_X1 U12482 ( .A1(n9706), .A2(n16519), .ZN(n10091) );
  INV_X1 U12483 ( .A(n9855), .ZN(n9854) );
  OAI21_X1 U12484 ( .B1(n10949), .B2(n9856), .A(n15974), .ZN(n9855) );
  NAND2_X1 U12486 ( .A1(n10151), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10152) );
  NAND2_X1 U12487 ( .A1(n9820), .A2(n9819), .ZN(n9755) );
  OR2_X1 U12488 ( .A1(n15701), .A2(n15894), .ZN(n9756) );
  AND3_X1 U12489 ( .A1(n12371), .A2(n12370), .A3(n9797), .ZN(n9757) );
  AND3_X1 U12490 ( .A1(n10465), .A2(n10464), .A3(n10467), .ZN(n9758) );
  NOR2_X1 U12491 ( .A1(n15701), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9759) );
  AND2_X1 U12492 ( .A1(n15773), .A2(n9917), .ZN(n9760) );
  OR2_X1 U12493 ( .A1(n9942), .A2(n17859), .ZN(n9761) );
  NAND2_X1 U12494 ( .A1(n14881), .A2(n14823), .ZN(n14799) );
  AND2_X1 U12495 ( .A1(n9894), .A2(n12290), .ZN(n18036) );
  NOR2_X1 U12496 ( .A1(n12493), .A2(n15864), .ZN(n12491) );
  OR2_X1 U12497 ( .A1(n15840), .A2(n15826), .ZN(n9762) );
  NAND2_X1 U12498 ( .A1(n12569), .A2(n12568), .ZN(n16564) );
  NAND2_X1 U12499 ( .A1(n16564), .A2(n16563), .ZN(n13599) );
  NOR3_X1 U12500 ( .A1(n12489), .A2(n9762), .A3(n15817), .ZN(n12488) );
  NOR2_X1 U12501 ( .A1(n12489), .A2(n15840), .ZN(n12490) );
  AND2_X1 U12502 ( .A1(n12491), .A2(n10793), .ZN(n12492) );
  NAND2_X1 U12503 ( .A1(n15590), .A2(n15581), .ZN(n15482) );
  AND2_X1 U12504 ( .A1(n13219), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11780) );
  AND2_X1 U12505 ( .A1(n15658), .A2(n15659), .ZN(n15657) );
  AND2_X1 U12506 ( .A1(n10037), .A2(n10035), .ZN(n9763) );
  AND2_X1 U12507 ( .A1(n14368), .A2(n15585), .ZN(n15579) );
  NAND2_X1 U12508 ( .A1(n11414), .A2(n11413), .ZN(n13704) );
  NAND2_X1 U12509 ( .A1(n13261), .A2(n13177), .ZN(n13347) );
  AND2_X1 U12510 ( .A1(n15472), .A2(n9717), .ZN(n9764) );
  AND2_X1 U12511 ( .A1(n14893), .A2(n15400), .ZN(n9765) );
  NAND2_X1 U12512 ( .A1(n14217), .A2(n14216), .ZN(n14997) );
  NAND2_X1 U12513 ( .A1(n9814), .A2(n14004), .ZN(n14088) );
  NAND2_X1 U12514 ( .A1(n16341), .A2(n13995), .ZN(n16336) );
  NAND2_X1 U12515 ( .A1(n14071), .A2(n9822), .ZN(n14230) );
  AND2_X1 U12516 ( .A1(n16001), .A2(n15645), .ZN(n15472) );
  INV_X1 U12517 ( .A(n19112), .ZN(n16828) );
  NOR2_X2 U12518 ( .A1(n12317), .A2(n12316), .ZN(n19112) );
  AND2_X1 U12519 ( .A1(n16122), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9766) );
  AND2_X1 U12520 ( .A1(n14127), .A2(n10188), .ZN(n14368) );
  NOR2_X1 U12521 ( .A1(n16125), .A2(n10110), .ZN(n16097) );
  NAND2_X1 U12522 ( .A1(n14069), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14071) );
  AND2_X1 U12523 ( .A1(n10537), .A2(n13788), .ZN(n13949) );
  AND2_X1 U12524 ( .A1(n13505), .A2(n13436), .ZN(n9767) );
  NOR2_X1 U12525 ( .A1(n16914), .A2(n17144), .ZN(n9768) );
  AND2_X1 U12526 ( .A1(n10101), .A2(n16167), .ZN(n9769) );
  NAND2_X1 U12527 ( .A1(n11351), .A2(n11350), .ZN(n11352) );
  INV_X1 U12528 ( .A(n13801), .ZN(n10037) );
  AND2_X1 U12529 ( .A1(n13642), .A2(n13637), .ZN(n14005) );
  INV_X1 U12530 ( .A(n14005), .ZN(n9971) );
  AND3_X1 U12531 ( .A1(n10816), .A2(n10910), .A3(n9929), .ZN(n9770) );
  AND2_X1 U12532 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n9771) );
  AND2_X1 U12533 ( .A1(n15555), .A2(n14479), .ZN(n9772) );
  NOR2_X1 U12534 ( .A1(n15011), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9773) );
  OR2_X1 U12535 ( .A1(n10532), .A2(n10531), .ZN(n12532) );
  NAND2_X1 U12536 ( .A1(n9656), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n9774) );
  AND2_X1 U12537 ( .A1(n9715), .A2(n9767), .ZN(n9775) );
  AND3_X1 U12538 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U12539 ( .A1(n13347), .A2(n9715), .ZN(n13437) );
  INV_X1 U12540 ( .A(n13277), .ZN(n10118) );
  AND2_X1 U12541 ( .A1(n12458), .A2(n9950), .ZN(n9777) );
  AND2_X2 U12542 ( .A1(n11068), .A2(n11067), .ZN(n20438) );
  XNOR2_X1 U12543 ( .A(n16640), .B(n16830), .ZN(n16820) );
  NAND2_X1 U12544 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  AND2_X1 U12545 ( .A1(n13347), .A2(n9775), .ZN(n13476) );
  OR2_X1 U12546 ( .A1(n12487), .A2(n10796), .ZN(n9778) );
  NAND2_X1 U12547 ( .A1(n9994), .A2(n9992), .ZN(n13911) );
  NAND2_X1 U12548 ( .A1(n12531), .A2(n12530), .ZN(n12740) );
  INV_X1 U12549 ( .A(n12740), .ZN(n9916) );
  AND2_X1 U12550 ( .A1(n14823), .A2(n9887), .ZN(n9779) );
  NOR3_X1 U12551 ( .A1(n14482), .A2(n14481), .A3(n15559), .ZN(n9780) );
  AND2_X1 U12552 ( .A1(n10816), .A2(n10910), .ZN(n9781) );
  AND2_X1 U12553 ( .A1(n9941), .A2(n9942), .ZN(n9782) );
  CLKBUF_X3 U12554 ( .A(n16820), .Z(n17144) );
  INV_X1 U12555 ( .A(n15436), .ZN(n10136) );
  AND2_X1 U12556 ( .A1(n9717), .A2(n15612), .ZN(n9783) );
  NAND2_X1 U12557 ( .A1(n10118), .A2(n9711), .ZN(n10121) );
  AND2_X1 U12558 ( .A1(n10145), .A2(n10144), .ZN(n9784) );
  OR3_X1 U12559 ( .A1(n12487), .A2(n10796), .A3(n9835), .ZN(n9785) );
  INV_X1 U12560 ( .A(n10345), .ZN(n12775) );
  AND2_X1 U12561 ( .A1(n10138), .A2(n10137), .ZN(n9786) );
  INV_X2 U12562 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17147) );
  AND2_X1 U12563 ( .A1(n17903), .A2(n9716), .ZN(n9787) );
  INV_X1 U12564 ( .A(n13455), .ZN(n10100) );
  AND2_X1 U12565 ( .A1(n9720), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9788) );
  OR2_X1 U12566 ( .A1(n12511), .A2(n9839), .ZN(n9789) );
  INV_X1 U12567 ( .A(n16332), .ZN(n20422) );
  NOR3_X1 U12568 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12318), .A3(
        n14265), .ZN(n12191) );
  AND2_X1 U12569 ( .A1(n18385), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n9790) );
  AND2_X1 U12570 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9791) );
  INV_X1 U12571 ( .A(n16008), .ZN(n10154) );
  AND2_X1 U12572 ( .A1(n12632), .A2(n12631), .ZN(n13349) );
  OR2_X1 U12573 ( .A1(n17755), .A2(n12306), .ZN(n9792) );
  AND2_X1 U12574 ( .A1(n9791), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9793) );
  AND2_X1 U12575 ( .A1(n20333), .A2(n20262), .ZN(n20320) );
  NOR2_X1 U12576 ( .A1(n19109), .A2(n17672), .ZN(n17688) );
  AOI22_X2 U12577 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19563), .ZN(n20077) );
  NOR2_X2 U12578 ( .A1(n19519), .A2(n19518), .ZN(n19563) );
  AOI22_X2 U12579 ( .A1(DATAI_17_), .A2(n20420), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20459), .ZN(n20920) );
  NAND3_X1 U12580 ( .A1(n12407), .A2(n18491), .A3(n18497), .ZN(n9794) );
  NAND3_X1 U12581 ( .A1(n9799), .A2(n9795), .A3(n12369), .ZN(n17642) );
  NAND3_X1 U12582 ( .A1(n12368), .A2(n12374), .A3(n9757), .ZN(n9796) );
  NOR2_X2 U12583 ( .A1(n16794), .A2(n19112), .ZN(n18118) );
  NAND2_X1 U12584 ( .A1(n15024), .A2(n9804), .ZN(n15025) );
  NOR2_X1 U12585 ( .A1(n10996), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9806) );
  INV_X1 U12586 ( .A(n11299), .ZN(n9809) );
  INV_X1 U12587 ( .A(n11298), .ZN(n9808) );
  INV_X1 U12588 ( .A(n11391), .ZN(n11393) );
  NAND2_X2 U12589 ( .A1(n9807), .A2(n11352), .ZN(n11391) );
  INV_X1 U12590 ( .A(n11353), .ZN(n9807) );
  NAND2_X2 U12591 ( .A1(n9809), .A2(n9808), .ZN(n11353) );
  INV_X1 U12592 ( .A(n15010), .ZN(n9972) );
  OAI21_X2 U12593 ( .B1(n15050), .B2(n15051), .A(n15135), .ZN(n15072) );
  NAND2_X2 U12594 ( .A1(n15017), .A2(n15108), .ZN(n15050) );
  OAI21_X2 U12595 ( .B1(n15118), .B2(n15016), .A(n15135), .ZN(n15108) );
  NAND2_X2 U12596 ( .A1(n15107), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15017) );
  NAND4_X1 U12597 ( .A1(n13209), .A2(n20450), .A3(n11172), .A4(n11301), .ZN(
        n13322) );
  NAND3_X1 U12598 ( .A1(n13209), .A2(n20450), .A3(n11172), .ZN(n13213) );
  NAND2_X1 U12599 ( .A1(n9813), .A2(n13104), .ZN(n12156) );
  NAND3_X1 U12600 ( .A1(n14071), .A2(n9822), .A3(n9816), .ZN(n9817) );
  NAND3_X1 U12601 ( .A1(n14071), .A2(n9822), .A3(n9739), .ZN(n9821) );
  NAND2_X1 U12602 ( .A1(n9827), .A2(n9826), .ZN(n10372) );
  AND2_X1 U12603 ( .A1(n9828), .A2(n10364), .ZN(n10371) );
  NAND3_X1 U12604 ( .A1(n9827), .A2(n9826), .A3(n9828), .ZN(n9825) );
  AND2_X2 U12605 ( .A1(n9825), .A2(n9823), .ZN(n10709) );
  NAND2_X1 U12606 ( .A1(n15850), .A2(n9831), .ZN(n15779) );
  INV_X1 U12607 ( .A(n15779), .ZN(n10667) );
  NAND3_X1 U12608 ( .A1(n10508), .A2(n10507), .A3(n12532), .ZN(n10844) );
  INV_X1 U12609 ( .A(n10538), .ZN(n10539) );
  NOR2_X2 U12610 ( .A1(n12487), .A2(n9832), .ZN(n12510) );
  NOR3_X2 U12611 ( .A1(n12489), .A2(n9762), .A3(n9836), .ZN(n12504) );
  NAND2_X1 U12612 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12499) );
  INV_X1 U12613 ( .A(n12499), .ZN(n9841) );
  NAND2_X1 U12614 ( .A1(n9841), .A2(n9840), .ZN(n12498) );
  AND2_X1 U12615 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n9840) );
  NAND2_X1 U12616 ( .A1(n9842), .A2(n16496), .ZN(n12505) );
  NAND3_X1 U12617 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .ZN(n9847) );
  OR2_X1 U12618 ( .A1(n10950), .A2(n9853), .ZN(n9850) );
  OR2_X1 U12619 ( .A1(n10950), .A2(n9856), .ZN(n9851) );
  NAND2_X1 U12620 ( .A1(n9850), .A2(n9852), .ZN(n15967) );
  NAND2_X1 U12621 ( .A1(n10587), .A2(n10586), .ZN(n10851) );
  NAND2_X1 U12622 ( .A1(n10539), .A2(n9857), .ZN(n10626) );
  NAND2_X1 U12623 ( .A1(n14237), .A2(n9733), .ZN(n9860) );
  OAI21_X1 U12624 ( .B1(n14237), .B2(n9863), .A(n9861), .ZN(n10934) );
  NAND3_X1 U12625 ( .A1(n9876), .A2(n9874), .A3(n9873), .ZN(n12026) );
  INV_X1 U12626 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9877) );
  NAND2_X1 U12627 ( .A1(n12303), .A2(n17786), .ZN(n9888) );
  INV_X1 U12628 ( .A(n9893), .ZN(n12455) );
  INV_X1 U12629 ( .A(n9894), .ZN(n17913) );
  OAI211_X1 U12630 ( .C1(n9908), .C2(n15700), .A(n9907), .B(n9905), .ZN(n9914)
         );
  NAND2_X1 U12631 ( .A1(n15699), .A2(n15701), .ZN(n9907) );
  NAND3_X1 U12632 ( .A1(n9910), .A2(n9909), .A3(n9912), .ZN(n15711) );
  NAND2_X1 U12633 ( .A1(n15700), .A2(n9915), .ZN(n9909) );
  OR2_X1 U12634 ( .A1(n15700), .A2(n9913), .ZN(n9910) );
  NOR2_X2 U12635 ( .A1(n10847), .A2(n9922), .ZN(n10871) );
  INV_X1 U12636 ( .A(n9928), .ZN(n10845) );
  NAND2_X1 U12637 ( .A1(n9934), .A2(n9935), .ZN(n16909) );
  NAND2_X1 U12638 ( .A1(n9939), .A2(n9761), .ZN(n16936) );
  NAND3_X1 U12639 ( .A1(n16959), .A2(n9940), .A3(n16818), .ZN(n9939) );
  NAND2_X1 U12640 ( .A1(n16959), .A2(n9944), .ZN(n16947) );
  INV_X1 U12641 ( .A(n17867), .ZN(n9943) );
  AND2_X1 U12642 ( .A1(n9952), .A2(n11231), .ZN(n11288) );
  NAND2_X1 U12643 ( .A1(n11093), .A2(n9953), .ZN(n11132) );
  NAND3_X1 U12644 ( .A1(n9954), .A2(n20446), .A3(n13642), .ZN(n9953) );
  NAND2_X1 U12645 ( .A1(n13662), .A2(n13661), .ZN(n13668) );
  NAND2_X1 U12646 ( .A1(n9712), .A2(n13662), .ZN(n9955) );
  NAND2_X1 U12647 ( .A1(n9959), .A2(n9957), .ZN(n9956) );
  INV_X1 U12648 ( .A(n13661), .ZN(n9957) );
  NAND2_X1 U12649 ( .A1(n9960), .A2(n9959), .ZN(n9958) );
  AND2_X1 U12650 ( .A1(n13667), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9959) );
  NAND2_X1 U12651 ( .A1(n15062), .A2(n9966), .ZN(n9965) );
  NAND2_X1 U12652 ( .A1(n11314), .A2(n11315), .ZN(n9970) );
  NAND2_X1 U12653 ( .A1(n9970), .A2(n9968), .ZN(n13306) );
  OAI21_X1 U12654 ( .B1(n9972), .B2(n9975), .A(n9973), .ZN(n15117) );
  INV_X1 U12655 ( .A(n15117), .ZN(n15012) );
  INV_X1 U12656 ( .A(n10172), .ZN(n9979) );
  INV_X1 U12657 ( .A(n10330), .ZN(n10115) );
  NAND2_X1 U12658 ( .A1(n15566), .A2(n14479), .ZN(n9983) );
  NAND2_X1 U12659 ( .A1(n15527), .A2(n9986), .ZN(n9985) );
  OAI211_X1 U12660 ( .C1(n15527), .C2(n9990), .A(n9988), .B(n9985), .ZN(n14629) );
  NAND2_X1 U12661 ( .A1(n15527), .A2(n15526), .ZN(n15528) );
  OAI21_X1 U12662 ( .B1(n14629), .B2(n15594), .A(n14606), .ZN(P2_U2857) );
  NOR2_X1 U12663 ( .A1(n13621), .A2(n9995), .ZN(n13910) );
  INV_X1 U12664 ( .A(n13621), .ZN(n9994) );
  OAI21_X1 U12665 ( .B1(n15544), .B2(n9998), .A(n9997), .ZN(n14547) );
  NAND2_X1 U12666 ( .A1(n14368), .A2(n10002), .ZN(n10001) );
  NOR2_X4 U12667 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13569) );
  NAND2_X1 U12668 ( .A1(n10008), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11176) );
  NOR2_X1 U12669 ( .A1(n10008), .A2(n13283), .ZN(n13308) );
  NAND3_X1 U12670 ( .A1(n11174), .A2(n11175), .A3(n11173), .ZN(n10008) );
  NAND3_X1 U12671 ( .A1(n11326), .A2(n10012), .A3(n10010), .ZN(n13424) );
  NOR2_X2 U12672 ( .A1(n14811), .A2(n10020), .ZN(n14770) );
  AND2_X1 U12673 ( .A1(n14679), .A2(n10029), .ZN(n14316) );
  NAND2_X1 U12674 ( .A1(n14679), .A2(n14680), .ZN(n14668) );
  NAND2_X2 U12675 ( .A1(n10040), .A2(n10395), .ZN(n10551) );
  NAND2_X1 U12676 ( .A1(n10394), .A2(n10040), .ZN(n10552) );
  INV_X1 U12677 ( .A(n10402), .ZN(n10040) );
  NAND2_X1 U12678 ( .A1(n10374), .A2(n10375), .ZN(n10373) );
  NAND3_X1 U12679 ( .A1(n10374), .A2(n10351), .A3(n10375), .ZN(n10041) );
  NAND2_X1 U12680 ( .A1(n10310), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10046) );
  NAND2_X1 U12681 ( .A1(n9663), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10050) );
  OAI21_X1 U12682 ( .B1(n15758), .B2(n10959), .A(n10075), .ZN(n10964) );
  OAI21_X1 U12683 ( .B1(n15757), .B2(n10959), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10076) );
  INV_X2 U12684 ( .A(n10305), .ZN(n10322) );
  NAND2_X1 U12685 ( .A1(n10077), .A2(n10261), .ZN(n10082) );
  NAND4_X1 U12686 ( .A1(n10208), .A2(n10209), .A3(n10207), .A4(n10210), .ZN(
        n10077) );
  NAND2_X2 U12687 ( .A1(n10079), .A2(n10078), .ZN(n10300) );
  NAND3_X1 U12688 ( .A1(n10251), .A2(n10252), .A3(n10190), .ZN(n10078) );
  NAND3_X1 U12689 ( .A1(n10246), .A2(n10245), .A3(n10247), .ZN(n10079) );
  NAND2_X2 U12690 ( .A1(n10082), .A2(n10080), .ZN(n10305) );
  NAND4_X1 U12691 ( .A1(n10215), .A2(n10213), .A3(n10212), .A4(n10214), .ZN(
        n10081) );
  NAND2_X1 U12692 ( .A1(n15734), .A2(n15732), .ZN(n15726) );
  NAND3_X1 U12693 ( .A1(n10096), .A2(n9709), .A3(n13957), .ZN(n10095) );
  INV_X1 U12694 ( .A(n12558), .ZN(n10096) );
  OR2_X1 U12695 ( .A1(n13681), .A2(n12558), .ZN(n10098) );
  NAND3_X1 U12696 ( .A1(n10463), .A2(n10466), .A3(n9758), .ZN(n10112) );
  NAND4_X1 U12697 ( .A1(n10114), .A2(n12898), .A3(n20220), .A4(n10113), .ZN(
        n10311) );
  NAND2_X1 U12698 ( .A1(n10310), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10113) );
  NAND2_X1 U12699 ( .A1(n10703), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10114) );
  NOR2_X2 U12700 ( .A1(n10345), .A2(n14477), .ZN(n10703) );
  NAND2_X1 U12701 ( .A1(n10118), .A2(n10116), .ZN(n13507) );
  INV_X1 U12702 ( .A(n10121), .ZN(n13419) );
  NOR2_X2 U12703 ( .A1(n15588), .A2(n15587), .ZN(n15590) );
  NOR2_X2 U12704 ( .A1(n13869), .A2(n14062), .ZN(n10123) );
  NAND2_X1 U12705 ( .A1(n10714), .A2(n10124), .ZN(n13181) );
  INV_X1 U12706 ( .A(n15560), .ZN(n10128) );
  NOR2_X2 U12707 ( .A1(n13433), .A2(n13474), .ZN(n10130) );
  OR3_X1 U12708 ( .A1(n9722), .A2(n12828), .A3(n10135), .ZN(n14282) );
  NOR3_X1 U12709 ( .A1(n9722), .A2(n10136), .A3(n12828), .ZN(n15439) );
  NOR2_X1 U12710 ( .A1(n9722), .A2(n12828), .ZN(n15437) );
  NAND3_X1 U12711 ( .A1(n10134), .A2(n10133), .A3(n10132), .ZN(n10131) );
  INV_X1 U12712 ( .A(n10138), .ZN(n18070) );
  XNOR2_X1 U12713 ( .A(n12282), .B(n12283), .ZN(n18071) );
  NOR2_X1 U12714 ( .A1(n18087), .A2(n12280), .ZN(n12282) );
  NAND2_X1 U12715 ( .A1(n16686), .A2(n12305), .ZN(n10148) );
  NAND3_X1 U12716 ( .A1(n10142), .A2(n10147), .A3(n16628), .ZN(n10141) );
  INV_X1 U12717 ( .A(n18051), .ZN(n10151) );
  NAND2_X1 U12718 ( .A1(n10152), .A2(n10150), .ZN(n12290) );
  INV_X1 U12719 ( .A(n10152), .ZN(n18050) );
  NAND3_X1 U12720 ( .A1(n12300), .A2(n12301), .A3(n17787), .ZN(n17786) );
  AND2_X4 U12721 ( .A1(n10431), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10284) );
  AND3_X2 U12722 ( .A1(n10339), .A2(n10153), .A3(n13840), .ZN(n10211) );
  NAND2_X2 U12723 ( .A1(n10156), .A2(n10155), .ZN(n13056) );
  NAND3_X1 U12724 ( .A1(n9749), .A2(n10277), .A3(n10275), .ZN(n10155) );
  NAND3_X1 U12725 ( .A1(n21259), .A2(n9750), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10156) );
  NAND2_X1 U12727 ( .A1(n15751), .A2(n9793), .ZN(n15720) );
  INV_X1 U12728 ( .A(n15712), .ZN(n10158) );
  NOR2_X1 U12729 ( .A1(n15712), .A2(n10159), .ZN(n15691) );
  NAND2_X1 U12730 ( .A1(n10158), .A2(n10160), .ZN(n14313) );
  NOR2_X1 U12731 ( .A1(n10162), .A2(n10161), .ZN(n10160) );
  NAND2_X1 U12732 ( .A1(n10991), .A2(n10990), .ZN(n10992) );
  INV_X1 U12733 ( .A(n14623), .ZN(n10991) );
  NAND2_X1 U12734 ( .A1(n11197), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11183) );
  AND2_X1 U12735 ( .A1(n13176), .A2(n13175), .ZN(n13177) );
  CLKBUF_X1 U12736 ( .A(n14842), .Z(n14844) );
  NAND2_X1 U12737 ( .A1(n14842), .A2(n11521), .ZN(n11555) );
  NAND2_X1 U12738 ( .A1(n13424), .A2(n11327), .ZN(n13466) );
  NAND4_X4 U12739 ( .A1(n11091), .A2(n11090), .A3(n11089), .A4(n11088), .ZN(
        n12155) );
  XNOR2_X1 U12740 ( .A(n13155), .B(n13156), .ZN(n13044) );
  NOR2_X1 U12741 ( .A1(n13155), .A2(n12952), .ZN(n19784) );
  AND2_X1 U12742 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10260) );
  AOI22_X1 U12743 ( .A1(n9692), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U12744 ( .A1(n9691), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10201) );
  INV_X1 U12745 ( .A(n13154), .ZN(n13259) );
  AND2_X1 U12746 ( .A1(n13012), .A2(n13011), .ZN(n13693) );
  NAND2_X1 U12747 ( .A1(n13949), .A2(n13950), .ZN(n10635) );
  INV_X1 U12748 ( .A(n10819), .ZN(n10628) );
  CLKBUF_X1 U12749 ( .A(n13146), .Z(n13454) );
  MUX2_X1 U12751 ( .A(n10322), .B(n10300), .S(n10321), .Z(n10323) );
  CLKBUF_X1 U12752 ( .A(n12980), .Z(n12988) );
  AOI21_X1 U12753 ( .B1(n10423), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n10261), .ZN(n10249) );
  AOI22_X1 U12754 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10202) );
  AND4_X1 U12755 ( .A1(n10412), .A2(n10411), .A3(n10410), .A4(n10409), .ZN(
        n10413) );
  AND2_X1 U12756 ( .A1(n12718), .A2(n12717), .ZN(n13622) );
  AND2_X1 U12757 ( .A1(n20363), .A2(n13334), .ZN(n20357) );
  INV_X1 U12758 ( .A(n13164), .ZN(n13167) );
  NAND2_X1 U12759 ( .A1(n14440), .A2(n10431), .ZN(n10164) );
  AND2_X1 U12760 ( .A1(n14522), .A2(n10185), .ZN(n10165) );
  AND4_X1 U12761 ( .A1(n12578), .A2(n12577), .A3(n12576), .A4(n12575), .ZN(
        n10166) );
  AND3_X1 U12762 ( .A1(n12467), .A2(n10177), .A3(n12466), .ZN(n10167) );
  AND3_X1 U12763 ( .A1(n12218), .A2(n12217), .A3(n12216), .ZN(n10168) );
  AND4_X1 U12764 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(
        n10169) );
  NAND2_X1 U12765 ( .A1(n11135), .A2(n13310), .ZN(n12942) );
  INV_X1 U12766 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20966) );
  NOR2_X1 U12767 ( .A1(n20753), .A2(n20786), .ZN(n10170) );
  AND4_X1 U12768 ( .A1(n12229), .A2(n12228), .A3(n12227), .A4(n12226), .ZN(
        n10171) );
  OR2_X1 U12769 ( .A1(n15011), .A2(n15007), .ZN(n10172) );
  INV_X1 U12770 ( .A(n15252), .ZN(n15019) );
  OR2_X1 U12771 ( .A1(n20220), .A2(n20199), .ZN(n10173) );
  AND2_X1 U12772 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10174) );
  NAND2_X1 U12773 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17881) );
  INV_X1 U12774 ( .A(n17881), .ZN(n12457) );
  NAND2_X1 U12775 ( .A1(n11467), .A2(n11466), .ZN(n10176) );
  INV_X1 U12776 ( .A(n10430), .ZN(n10646) );
  NOR2_X1 U12777 ( .A1(n12464), .A2(n12463), .ZN(n10177) );
  INV_X1 U12778 ( .A(n19055), .ZN(n19120) );
  NAND2_X1 U12779 ( .A1(n9738), .A2(n14461), .ZN(n10178) );
  AND2_X1 U12780 ( .A1(n15685), .A2(n15683), .ZN(n10179) );
  OR2_X1 U12781 ( .A1(n13325), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10180) );
  OR2_X1 U12782 ( .A1(n15011), .A2(n16384), .ZN(n10181) );
  NAND2_X1 U12783 ( .A1(n12811), .A2(n19186), .ZN(n10182) );
  AND2_X1 U12784 ( .A1(n10262), .A2(n10261), .ZN(n10183) );
  AND2_X1 U12785 ( .A1(n15316), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10184) );
  INV_X1 U12786 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15023) );
  INV_X1 U12787 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12306) );
  INV_X1 U12788 ( .A(n15789), .ZN(n10945) );
  AND2_X1 U12789 ( .A1(n14521), .A2(n14541), .ZN(n10185) );
  NOR2_X1 U12790 ( .A1(n20753), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10186) );
  OR2_X1 U12791 ( .A1(n13325), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10187) );
  OR2_X1 U12792 ( .A1(n12847), .A2(n10292), .ZN(n16537) );
  INV_X1 U12793 ( .A(n16537), .ZN(n10990) );
  NOR2_X1 U12794 ( .A1(n14129), .A2(n14126), .ZN(n10188) );
  AND4_X1 U12795 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(
        n10189) );
  AND3_X1 U12796 ( .A1(n10250), .A2(n10249), .A3(n10248), .ZN(n10190) );
  INV_X1 U12797 ( .A(n11352), .ZN(n13629) );
  OR2_X1 U12798 ( .A1(n17933), .A2(n18135), .ZN(n10191) );
  AND2_X1 U12799 ( .A1(n16693), .A2(n16692), .ZN(n10192) );
  CLKBUF_X3 U12800 ( .A(n12239), .Z(n17348) );
  CLKBUF_X3 U12801 ( .A(n12335), .Z(n16181) );
  NOR2_X1 U12802 ( .A1(n12178), .A2(n12181), .ZN(n12307) );
  NOR2_X1 U12803 ( .A1(n19506), .A2(n19314), .ZN(n10193) );
  AND3_X1 U12804 ( .A1(n10460), .A2(n10459), .A3(n10458), .ZN(n10194) );
  OR2_X1 U12805 ( .A1(n12552), .A2(n12551), .ZN(n10195) );
  NAND2_X1 U12806 ( .A1(n13049), .A2(n20095), .ZN(n15578) );
  OR2_X1 U12807 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n10196) );
  INV_X1 U12808 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10442) );
  INV_X1 U12809 ( .A(n11990), .ZN(n11987) );
  NOR2_X1 U12810 ( .A1(n12942), .A2(n11158), .ZN(n11160) );
  AOI22_X1 U12811 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10559), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10409) );
  INV_X1 U12812 ( .A(n11213), .ZN(n11830) );
  NAND2_X1 U12813 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10254) );
  AND2_X1 U12814 ( .A1(n12999), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10319) );
  NAND2_X1 U12815 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10464) );
  INV_X1 U12816 ( .A(n10323), .ZN(n10326) );
  AOI22_X1 U12817 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10199) );
  OR2_X1 U12818 ( .A1(n11378), .A2(n11377), .ZN(n13987) );
  AND2_X1 U12819 ( .A1(n11283), .A2(n10189), .ZN(n13639) );
  INV_X1 U12820 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11003) );
  NOR2_X1 U12821 ( .A1(n10332), .A2(n10312), .ZN(n12980) );
  AND2_X1 U12822 ( .A1(n10673), .A2(n10672), .ZN(n10675) );
  NAND2_X1 U12823 ( .A1(n11148), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11045) );
  NOR2_X1 U12824 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10995) );
  INV_X1 U12825 ( .A(n14877), .ZN(n11595) );
  OAI21_X1 U12826 ( .B1(n11902), .B2(n13805), .A(n11447), .ZN(n11448) );
  NAND2_X1 U12827 ( .A1(n9685), .A2(n15019), .ZN(n15020) );
  INV_X1 U12828 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12025) );
  OAI211_X1 U12829 ( .C1(n9694), .C2(n11003), .A(n11002), .B(n11001), .ZN(
        n11004) );
  INV_X1 U12830 ( .A(n14503), .ZN(n14505) );
  INV_X1 U12831 ( .A(n10344), .ZN(n10370) );
  INV_X1 U12832 ( .A(n19535), .ZN(n10292) );
  AOI21_X1 U12833 ( .B1(n20786), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11962), .ZN(n11961) );
  OAI211_X1 U12834 ( .C1(n9694), .C2(n11047), .A(n11046), .B(n11045), .ZN(
        n11048) );
  INV_X1 U12835 ( .A(n13445), .ZN(n11389) );
  NOR2_X1 U12836 ( .A1(n11852), .A2(n11854), .ZN(n11924) );
  OR2_X1 U12837 ( .A1(n11741), .A2(n11740), .ZN(n11742) );
  NAND2_X1 U12838 ( .A1(n14027), .A2(n14843), .ZN(n14842) );
  NOR2_X1 U12839 ( .A1(n11227), .A2(n11226), .ZN(n13669) );
  INV_X1 U12840 ( .A(n13429), .ZN(n12031) );
  NOR2_X1 U12841 ( .A1(n12972), .A2(n12967), .ZN(n12971) );
  AND2_X1 U12842 ( .A1(n12525), .A2(n10810), .ZN(n10846) );
  INV_X1 U12843 ( .A(n13622), .ZN(n13623) );
  INV_X1 U12844 ( .A(n13182), .ZN(n10718) );
  AOI22_X1 U12845 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10423), .B1(
        n10424), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10210) );
  OR2_X1 U12846 ( .A1(n14505), .A2(n14504), .ZN(n14506) );
  AOI22_X1 U12847 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10285) );
  NAND2_X1 U12848 ( .A1(n10365), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10354) );
  INV_X1 U12849 ( .A(n10638), .ZN(n10662) );
  NAND2_X1 U12850 ( .A1(n12307), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12216) );
  AOI21_X1 U12851 ( .B1(n16691), .B2(n18906), .A(n16690), .ZN(n16692) );
  NOR2_X1 U12852 ( .A1(n17623), .A2(n12277), .ZN(n12261) );
  NOR2_X1 U12853 ( .A1(n11049), .A2(n11048), .ZN(n11050) );
  AND2_X1 U12854 ( .A1(n20261), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20340) );
  AND2_X1 U12855 ( .A1(n13224), .A2(n12151), .ZN(n12152) );
  AND2_X1 U12856 ( .A1(n11925), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12021) );
  OR2_X1 U12857 ( .A1(n11742), .A2(n14731), .ZN(n11776) );
  NAND2_X1 U12858 ( .A1(n11671), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11694) );
  NAND2_X1 U12859 ( .A1(n11556), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11557) );
  INV_X1 U12860 ( .A(n11359), .ZN(n11902) );
  INV_X1 U12861 ( .A(n11503), .ZN(n11590) );
  NAND2_X1 U12862 ( .A1(n15017), .A2(n15011), .ZN(n15081) );
  AND2_X1 U12863 ( .A1(n12065), .A2(n12064), .ZN(n15400) );
  AND2_X1 U12864 ( .A1(n20966), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12142) );
  NOR2_X1 U12865 ( .A1(n20667), .A2(n20666), .ZN(n20754) );
  OR2_X1 U12866 ( .A1(n10685), .A2(n12956), .ZN(n10681) );
  AND2_X1 U12867 ( .A1(n10874), .A2(n10873), .ZN(n19261) );
  NAND2_X1 U12868 ( .A1(n10840), .A2(n10839), .ZN(n10847) );
  NAND2_X1 U12869 ( .A1(n10830), .A2(n10833), .ZN(n10829) );
  INV_X1 U12870 ( .A(n14482), .ZN(n14461) );
  INV_X1 U12871 ( .A(n12773), .ZN(n12774) );
  NAND2_X1 U12872 ( .A1(n12510), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12511) );
  NOR2_X1 U12873 ( .A1(n14613), .A2(n15882), .ZN(n14614) );
  INV_X1 U12874 ( .A(n10869), .ZN(n14277) );
  OAI21_X1 U12875 ( .B1(n13537), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13535), .ZN(n10838) );
  AND2_X1 U12876 ( .A1(n12260), .A2(n17609), .ZN(n12286) );
  INV_X1 U12877 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12274) );
  AND2_X1 U12878 ( .A1(n20962), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16243) );
  INV_X1 U12879 ( .A(n12136), .ZN(n12137) );
  INV_X1 U12880 ( .A(n20333), .ZN(n14817) );
  INV_X1 U12881 ( .A(n20340), .ZN(n20279) );
  NAND2_X1 U12882 ( .A1(n21047), .A2(n12020), .ZN(n20261) );
  AND2_X1 U12883 ( .A1(n11955), .A2(n11927), .ZN(n14320) );
  OR2_X1 U12884 ( .A1(n14991), .A2(n13293), .ZN(n12171) );
  AND2_X1 U12885 ( .A1(n13195), .A2(n12156), .ZN(n12157) );
  OAI21_X1 U12886 ( .B1(n10196), .B2(n15058), .A(n11903), .ZN(n14669) );
  AND3_X1 U12887 ( .A1(n11594), .A2(n11593), .A3(n11592), .ZN(n14877) );
  INV_X1 U12888 ( .A(n20357), .ZN(n15201) );
  AND2_X1 U12889 ( .A1(n12068), .A2(n12067), .ZN(n14849) );
  AND2_X1 U12890 ( .A1(n13318), .A2(n13317), .ZN(n20371) );
  OAI21_X1 U12891 ( .B1(n21054), .B2(n16427), .A(n15422), .ZN(n20423) );
  NOR2_X1 U12892 ( .A1(n20424), .A2(n20557), .ZN(n20727) );
  NOR2_X1 U12893 ( .A1(n20558), .A2(n20557), .ZN(n20857) );
  INV_X1 U12894 ( .A(n10366), .ZN(n14286) );
  NOR2_X1 U12895 ( .A1(n15466), .A2(n15756), .ZN(n15467) );
  INV_X1 U12896 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19262) );
  INV_X1 U12897 ( .A(n15472), .ZN(n15646) );
  INV_X1 U12898 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15690) );
  OR2_X1 U12899 ( .A1(n10692), .A2(n12981), .ZN(n13081) );
  AND3_X1 U12900 ( .A1(n13021), .A2(n13020), .A3(n13019), .ZN(n16589) );
  NAND2_X1 U12901 ( .A1(n20177), .A2(n19784), .ZN(n19760) );
  NOR2_X1 U12902 ( .A1(n20184), .A2(n19657), .ZN(n19898) );
  INV_X1 U12903 ( .A(n19986), .ZN(n19856) );
  INV_X1 U12904 ( .A(n19956), .ZN(n20039) );
  INV_X1 U12905 ( .A(n17916), .ZN(n17919) );
  NOR2_X1 U12906 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17055), .ZN(n17037) );
  NOR2_X1 U12907 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17118), .ZN(n17109) );
  NOR2_X1 U12908 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17133), .ZN(n17132) );
  NOR2_X1 U12909 ( .A1(n12415), .A2(n18918), .ZN(n14134) );
  NOR2_X1 U12910 ( .A1(n17657), .A2(n17533), .ZN(n17532) );
  INV_X1 U12911 ( .A(n12231), .ZN(n12236) );
  OAI21_X1 U12912 ( .B1(n16271), .B2(n16270), .A(n19107), .ZN(n17487) );
  OR2_X1 U12913 ( .A1(n12465), .A2(n16628), .ZN(n12466) );
  NOR2_X1 U12914 ( .A1(n16203), .A2(n17792), .ZN(n18131) );
  NOR2_X1 U12915 ( .A1(n17844), .A2(n16817), .ZN(n17823) );
  INV_X1 U12916 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17917) );
  NAND2_X1 U12917 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17934), .ZN(
        n18322) );
  NOR2_X1 U12918 ( .A1(n18048), .A2(n18031), .ZN(n18027) );
  INV_X1 U12919 ( .A(n16635), .ZN(n16636) );
  NOR2_X1 U12920 ( .A1(n17799), .A2(n16203), .ZN(n18139) );
  NAND2_X1 U12921 ( .A1(n16681), .A2(n12286), .ZN(n17933) );
  NAND2_X1 U12922 ( .A1(n12454), .A2(n18025), .ZN(n17939) );
  NAND2_X1 U12923 ( .A1(n19125), .A2(n14259), .ZN(n18924) );
  NOR2_X1 U12924 ( .A1(n12404), .A2(n12403), .ZN(n18485) );
  INV_X1 U12925 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18916) );
  OR2_X1 U12926 ( .A1(n13332), .A2(n13028), .ZN(n13268) );
  OAI21_X1 U12927 ( .B1(n15231), .B2(n20325), .A(n12481), .ZN(n12482) );
  OR2_X1 U12928 ( .A1(n20333), .A2(n20332), .ZN(n20292) );
  AND2_X1 U12929 ( .A1(n20261), .A2(n12023), .ZN(n20317) );
  NOR2_X1 U12930 ( .A1(n12128), .A2(n12131), .ZN(n20333) );
  NOR2_X1 U12931 ( .A1(n14962), .A2(n16701), .ZN(n12172) );
  NOR2_X2 U12932 ( .A1(n12171), .A2(n20419), .ZN(n14970) );
  NOR2_X1 U12933 ( .A1(n14991), .A2(n13249), .ZN(n14993) );
  INV_X1 U12934 ( .A(n20368), .ZN(n16321) );
  NAND2_X1 U12935 ( .A1(n11410), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11431) );
  AND2_X1 U12936 ( .A1(n13330), .A2(n20909), .ZN(n16332) );
  OR2_X1 U12937 ( .A1(n15302), .A2(n15220), .ZN(n15293) );
  NOR2_X1 U12939 ( .A1(n16396), .A2(n15214), .ZN(n16355) );
  INV_X1 U12940 ( .A(n20408), .ZN(n20399) );
  INV_X1 U12941 ( .A(n20370), .ZN(n20390) );
  NOR2_X1 U12942 ( .A1(n20674), .A2(n13285), .ZN(n16247) );
  NOR2_X1 U12943 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16419) );
  INV_X1 U12944 ( .A(n20513), .ZN(n20517) );
  INV_X1 U12945 ( .A(n20546), .ZN(n20547) );
  OR2_X1 U12946 ( .A1(n9702), .A2(n20784), .ZN(n20664) );
  OR2_X1 U12947 ( .A1(n9702), .A2(n13302), .ZN(n20700) );
  INV_X1 U12948 ( .A(n20663), .ZN(n20654) );
  INV_X1 U12949 ( .A(n20657), .ZN(n20691) );
  INV_X1 U12950 ( .A(n20752), .ZN(n20744) );
  AND2_X1 U12951 ( .A1(n9702), .A2(n13302), .ZN(n20721) );
  INV_X1 U12952 ( .A(n20697), .ZN(n20762) );
  OAI211_X1 U12953 ( .C1(n20888), .C2(n20858), .A(n20857), .B(n20856), .ZN(
        n20891) );
  INV_X1 U12954 ( .A(n21011), .ZN(n21026) );
  INV_X1 U12955 ( .A(n19292), .ZN(n19313) );
  INV_X1 U12956 ( .A(n15827), .ZN(n16062) );
  INV_X1 U12957 ( .A(n15594), .ZN(n15575) );
  INV_X1 U12958 ( .A(n19371), .ZN(n19399) );
  INV_X1 U12959 ( .A(n12946), .ZN(n12884) );
  INV_X1 U12960 ( .A(n12504), .ZN(n12507) );
  AND2_X1 U12961 ( .A1(n16541), .A2(n20192), .ZN(n19486) );
  INV_X1 U12962 ( .A(n13168), .ZN(n13147) );
  OAI21_X1 U12963 ( .B1(n19531), .B2(n19530), .A(n19529), .ZN(n19568) );
  NOR2_X1 U12964 ( .A1(n19658), .A2(n19886), .ZN(n19647) );
  NOR2_X1 U12965 ( .A1(n19658), .A2(n19961), .ZN(n19705) );
  INV_X1 U12966 ( .A(n19783), .ZN(n19765) );
  NOR2_X2 U12967 ( .A1(n19761), .A2(n19760), .ZN(n19816) );
  NOR2_X2 U12968 ( .A1(n19856), .A2(n19831), .ZN(n19851) );
  NOR2_X1 U12969 ( .A1(n19856), .A2(n19886), .ZN(n19910) );
  AND2_X1 U12970 ( .A1(n20184), .A2(n19657), .ZN(n19959) );
  INV_X1 U12971 ( .A(n20027), .ZN(n20014) );
  INV_X1 U12972 ( .A(n20174), .ZN(n19761) );
  INV_X1 U12973 ( .A(n17705), .ZN(n17641) );
  NOR2_X1 U12974 ( .A1(n16822), .A2(n16821), .ZN(n18909) );
  NOR2_X1 U12975 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16940), .ZN(n16927) );
  NOR2_X1 U12976 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16962), .ZN(n16948) );
  NOR2_X1 U12977 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16985), .ZN(n16969) );
  INV_X1 U12978 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17918) );
  NOR2_X1 U12979 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17077), .ZN(n17059) );
  NOR2_X2 U12980 ( .A1(n18959), .A2(n16826), .ZN(n17168) );
  NAND2_X1 U12981 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17291), .ZN(n17262) );
  NAND2_X1 U12982 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17318), .ZN(n17303) );
  NOR2_X1 U12983 ( .A1(n17419), .A2(n17435), .ZN(n17404) );
  INV_X1 U12984 ( .A(n17506), .ZN(n17501) );
  OR2_X1 U12985 ( .A1(n17655), .A2(n17526), .ZN(n17527) );
  NOR2_X1 U12986 ( .A1(n17665), .A2(n17557), .ZN(n17552) );
  NAND2_X1 U12987 ( .A1(n17597), .A2(n16272), .ZN(n17627) );
  OAI21_X1 U12988 ( .B1(n9705), .B2(n17933), .A(n16682), .ZN(n17767) );
  INV_X1 U12989 ( .A(n17965), .ZN(n17979) );
  NAND2_X1 U12990 ( .A1(n18237), .A2(n17939), .ZN(n18272) );
  NAND2_X1 U12991 ( .A1(n17950), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18265) );
  OAI21_X1 U12992 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19106), .A(n16794), 
        .ZN(n18125) );
  NOR2_X1 U12993 ( .A1(n16681), .A2(n18912), .ZN(n18323) );
  NOR2_X1 U12994 ( .A1(n18313), .A2(n18433), .ZN(n18344) );
  INV_X1 U12995 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18942) );
  INV_X1 U12996 ( .A(n18847), .ZN(n18827) );
  INV_X1 U12997 ( .A(n18574), .ZN(n18637) );
  INV_X1 U12998 ( .A(n18664), .ZN(n18729) );
  INV_X1 U12999 ( .A(n18756), .ZN(n18817) );
  OAI22_X1 U13000 ( .A1(n12430), .A2(n18912), .B1(n16198), .B2(n18303), .ZN(
        n18957) );
  INV_X1 U13001 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18982) );
  INV_X1 U13002 ( .A(n19519), .ZN(n19517) );
  OR2_X1 U13003 ( .A1(n13332), .A2(n12942), .ZN(n13098) );
  INV_X1 U13004 ( .A(n12482), .ZN(n12483) );
  INV_X1 U13005 ( .A(n20334), .ZN(n20325) );
  INV_X1 U13006 ( .A(n20317), .ZN(n20287) );
  AND2_X1 U13007 ( .A1(n20287), .A2(n13855), .ZN(n13975) );
  NAND2_X1 U13008 ( .A1(n14988), .A2(n13249), .ZN(n14995) );
  INV_X1 U13009 ( .A(n14993), .ZN(n14987) );
  NAND3_X1 U13010 ( .A1(n13267), .A2(n16235), .A3(n13282), .ZN(n13758) );
  NOR2_X1 U13011 ( .A1(n13098), .A2(n13097), .ZN(n13114) );
  NAND2_X1 U13012 ( .A1(n13114), .A2(n11968), .ZN(n13357) );
  OR2_X1 U13013 ( .A1(n20357), .A2(n13648), .ZN(n20368) );
  INV_X1 U13014 ( .A(n20406), .ZN(n16412) );
  NAND2_X1 U13015 ( .A1(n13324), .A2(n13301), .ZN(n20408) );
  INV_X1 U13016 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16215) );
  OR2_X1 U13017 ( .A1(n20526), .A2(n20664), .ZN(n20492) );
  OR2_X1 U13018 ( .A1(n20526), .A2(n20850), .ZN(n20546) );
  OR2_X1 U13019 ( .A1(n20526), .A2(n20760), .ZN(n20572) );
  OR2_X1 U13020 ( .A1(n20641), .A2(n20664), .ZN(n20600) );
  OR2_X1 U13021 ( .A1(n20641), .A2(n20700), .ZN(n20629) );
  OR2_X1 U13022 ( .A1(n20641), .A2(n20850), .ZN(n20663) );
  NAND2_X1 U13023 ( .A1(n20762), .A2(n20665), .ZN(n20720) );
  NAND2_X1 U13024 ( .A1(n20762), .A2(n20721), .ZN(n20783) );
  NAND2_X1 U13025 ( .A1(n20762), .A2(n20761), .ZN(n20818) );
  NAND2_X1 U13026 ( .A1(n20904), .A2(n20819), .ZN(n20894) );
  OR2_X1 U13027 ( .A1(n20851), .A2(n20760), .ZN(n20960) );
  INV_X1 U13028 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20962) );
  INV_X1 U13029 ( .A(n21036), .ZN(n20968) );
  INV_X1 U13030 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n16263) );
  NAND2_X1 U13031 ( .A1(n20041), .A2(n19953), .ZN(n20183) );
  NAND2_X1 U13032 ( .A1(n13051), .A2(n10701), .ZN(n12847) );
  INV_X1 U13033 ( .A(n19317), .ZN(n19300) );
  INV_X1 U13034 ( .A(n19319), .ZN(n19312) );
  INV_X1 U13035 ( .A(n15578), .ZN(n15572) );
  NAND2_X1 U13036 ( .A1(n19371), .A2(n10293), .ZN(n16479) );
  AND2_X1 U13037 ( .A1(n13000), .A2(n20095), .ZN(n19371) );
  INV_X1 U13038 ( .A(n19365), .ZN(n19408) );
  OR2_X1 U13039 ( .A1(n19456), .A2(n20223), .ZN(n19459) );
  INV_X1 U13040 ( .A(n19456), .ZN(n19478) );
  INV_X1 U13041 ( .A(n19481), .ZN(n12947) );
  INV_X1 U13042 ( .A(n16529), .ZN(n19490) );
  INV_X1 U13043 ( .A(n16533), .ZN(n19496) );
  NAND2_X1 U13044 ( .A1(n13091), .A2(n20210), .ZN(n19502) );
  NAND2_X1 U13045 ( .A1(n13091), .A2(n20212), .ZN(n19515) );
  INV_X1 U13046 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13026) );
  OR2_X1 U13047 ( .A1(n19831), .A2(n19658), .ZN(n19597) );
  INV_X1 U13048 ( .A(n19647), .ZN(n19656) );
  INV_X1 U13049 ( .A(n19705), .ZN(n19714) );
  INV_X1 U13050 ( .A(n19745), .ZN(n19738) );
  AND2_X1 U13051 ( .A1(n19755), .A2(n19754), .ZN(n19768) );
  NAND2_X1 U13052 ( .A1(n19719), .A2(n20174), .ZN(n19783) );
  AOI211_X2 U13053 ( .C1(n19790), .C2(n19791), .A(n19956), .B(n19789), .ZN(
        n19821) );
  AOI21_X1 U13054 ( .B1(n19827), .B2(n19829), .A(n19826), .ZN(n19855) );
  INV_X1 U13055 ( .A(n19948), .ZN(n19925) );
  NAND2_X1 U13056 ( .A1(n19986), .A2(n19959), .ZN(n19985) );
  OR2_X1 U13057 ( .A1(n19962), .A2(n19961), .ZN(n20027) );
  INV_X1 U13058 ( .A(n20089), .ZN(n20064) );
  OR2_X1 U13059 ( .A1(n19962), .A2(n19761), .ZN(n20093) );
  NAND2_X1 U13060 ( .A1(n19107), .A2(n18957), .ZN(n16794) );
  INV_X1 U13061 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17995) );
  INV_X1 U13062 ( .A(n17192), .ZN(n17157) );
  NOR2_X1 U13063 ( .A1(n16902), .A2(n17238), .ZN(n17243) );
  NOR2_X1 U13064 ( .A1(n17305), .A2(n17330), .ZN(n17318) );
  NOR2_X2 U13065 ( .A1(n17481), .A2(n18518), .ZN(n17482) );
  INV_X1 U13066 ( .A(n17627), .ZN(n17580) );
  INV_X1 U13067 ( .A(n16681), .ZN(n17605) );
  NOR2_X1 U13068 ( .A1(n12201), .A2(n12200), .ZN(n17613) );
  NAND2_X1 U13069 ( .A1(n18936), .A2(n16272), .ZN(n17630) );
  INV_X1 U13070 ( .A(n17672), .ZN(n17703) );
  NAND2_X1 U13071 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18122), .ZN(n17965) );
  INV_X1 U13072 ( .A(n18039), .ZN(n18024) );
  NOR2_X1 U13073 ( .A1(n18079), .A2(n18080), .ZN(n18122) );
  XNOR2_X1 U13074 ( .A(n17774), .B(n17933), .ZN(n18144) );
  INV_X1 U13075 ( .A(n18451), .ZN(n18433) );
  INV_X1 U13076 ( .A(n18367), .ZN(n18352) );
  INV_X1 U13077 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18940) );
  INV_X1 U13078 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18947) );
  INV_X1 U13079 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18500) );
  INV_X1 U13080 ( .A(n18523), .ZN(n18858) );
  INV_X1 U13081 ( .A(n18539), .ZN(n18888) );
  INV_X1 U13082 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19000) );
  NOR2_X1 U13083 ( .A1(n18982), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n19055) );
  INV_X1 U13084 ( .A(n16744), .ZN(n16750) );
  NAND2_X1 U13085 ( .A1(n12468), .A2(n10167), .ZN(P3_U2800) );
  INV_X1 U13086 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15882) );
  AND2_X4 U13087 ( .A1(n10418), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10416) );
  AOI22_X1 U13088 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10200) );
  AND2_X4 U13089 ( .A1(n10431), .A2(n16575), .ZN(n10424) );
  AND2_X4 U13090 ( .A1(n10417), .A2(n10339), .ZN(n10423) );
  AND3_X4 U13091 ( .A1(n13840), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13092 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U13093 ( .A1(n9691), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U13094 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10204) );
  AOI22_X1 U13095 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U13096 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U13097 ( .A1(n9692), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U13098 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U13099 ( .A1(n9691), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U13100 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10214) );
  CLKBUF_X1 U13101 ( .A(n10211), .Z(n10278) );
  AOI22_X1 U13102 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U13103 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U13104 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9680), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10220) );
  AOI21_X1 U13105 ( .B1(n9692), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A(n10216), .ZN(n10219) );
  AOI22_X1 U13106 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10218) );
  AOI22_X1 U13107 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10217) );
  NAND4_X1 U13108 ( .A1(n10220), .A2(n10219), .A3(n10218), .A4(n10217), .ZN(
        n10221) );
  NAND2_X1 U13109 ( .A1(n10221), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10229) );
  AOI22_X1 U13110 ( .A1(n9692), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10224) );
  AOI22_X1 U13111 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U13112 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10222) );
  NAND3_X1 U13113 ( .A1(n10224), .A2(n10223), .A3(n10222), .ZN(n10227) );
  AOI22_X1 U13114 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10225) );
  INV_X1 U13115 ( .A(n10225), .ZN(n10226) );
  OAI21_X1 U13116 ( .B1(n10227), .B2(n10226), .A(n10261), .ZN(n10228) );
  AOI22_X1 U13117 ( .A1(n14590), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10235) );
  AOI22_X1 U13118 ( .A1(n9692), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10234) );
  AOI22_X1 U13119 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10232) );
  NAND2_X1 U13120 ( .A1(n10423), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10230) );
  NAND3_X1 U13121 ( .A1(n10235), .A2(n10234), .A3(n10233), .ZN(n10242) );
  AOI22_X1 U13122 ( .A1(n9691), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U13123 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U13124 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10238) );
  NAND3_X1 U13125 ( .A1(n10240), .A2(n10239), .A3(n10238), .ZN(n10241) );
  AOI22_X1 U13126 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10247) );
  AOI22_X1 U13127 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U13128 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U13129 ( .A1(n9695), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U13130 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U13131 ( .A1(n10423), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10253) );
  AOI22_X1 U13132 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U13133 ( .A1(n14590), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U13134 ( .A1(n9691), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U13135 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U13136 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U13137 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10263) );
  NAND4_X1 U13138 ( .A1(n10265), .A2(n10264), .A3(n10183), .A4(n10263), .ZN(
        n10266) );
  AOI22_X1 U13139 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10269) );
  AOI22_X1 U13140 ( .A1(n9691), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10268) );
  AOI22_X1 U13141 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10272) );
  NAND2_X1 U13142 ( .A1(n9695), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10270) );
  AOI22_X1 U13144 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13145 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13146 ( .A1(n9691), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U13147 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10274) );
  AOI22_X1 U13148 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9680), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U13149 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U13150 ( .A1(n9692), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U13151 ( .A1(n10424), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10423), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10279) );
  NAND4_X1 U13152 ( .A1(n10282), .A2(n10281), .A3(n10280), .A4(n10279), .ZN(
        n10283) );
  AOI22_X1 U13153 ( .A1(n9691), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13154 ( .A1(n14442), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U13155 ( .A1(n10211), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9679), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10286) );
  NAND4_X1 U13156 ( .A1(n10288), .A2(n10287), .A3(n10286), .A4(n10285), .ZN(
        n10289) );
  NAND2_X1 U13157 ( .A1(n10289), .A2(n10261), .ZN(n10290) );
  NAND2_X1 U13158 ( .A1(n12775), .A2(n10292), .ZN(n12773) );
  NAND2_X1 U13159 ( .A1(n10312), .A2(n10452), .ZN(n10295) );
  INV_X1 U13160 ( .A(n12984), .ZN(n10293) );
  NAND3_X1 U13161 ( .A1(n13012), .A2(n13073), .A3(n13011), .ZN(n13088) );
  NAND3_X1 U13162 ( .A1(n10452), .A2(n13056), .A3(n10306), .ZN(n10301) );
  NAND2_X1 U13163 ( .A1(n12998), .A2(n13004), .ZN(n10347) );
  AND2_X2 U13164 ( .A1(n9661), .A2(n10306), .ZN(n10332) );
  INV_X1 U13165 ( .A(n10296), .ZN(n13069) );
  INV_X1 U13166 ( .A(n10302), .ZN(n19545) );
  AND2_X1 U13167 ( .A1(n13069), .A2(n19545), .ZN(n10303) );
  NAND4_X1 U13168 ( .A1(n12773), .A2(n13088), .A3(n10347), .A4(n12987), .ZN(
        n10304) );
  AND2_X2 U13169 ( .A1(n10304), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10365) );
  NOR2_X1 U13170 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16615) );
  NAND2_X1 U13171 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12898) );
  AOI21_X1 U13172 ( .B1(n10365), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n10311), .ZN(n10338) );
  NAND2_X1 U13173 ( .A1(n12980), .A2(n19549), .ZN(n10314) );
  OAI21_X1 U13174 ( .B1(n13066), .B2(n19545), .A(n10316), .ZN(n10320) );
  INV_X1 U13175 ( .A(n10315), .ZN(n10318) );
  NAND2_X1 U13176 ( .A1(n12984), .A2(n10452), .ZN(n13072) );
  NAND2_X1 U13177 ( .A1(n10320), .A2(n10319), .ZN(n10337) );
  NAND2_X1 U13178 ( .A1(n12984), .A2(n13078), .ZN(n10325) );
  INV_X1 U13179 ( .A(n10332), .ZN(n10324) );
  NAND4_X1 U13180 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n19539), .ZN(
        n10329) );
  INV_X1 U13181 ( .A(n10327), .ZN(n10328) );
  NAND3_X1 U13182 ( .A1(n10329), .A2(n10328), .A3(n13056), .ZN(n13068) );
  NAND2_X1 U13183 ( .A1(n10331), .A2(n10332), .ZN(n10692) );
  AND2_X1 U13184 ( .A1(n19539), .A2(n9676), .ZN(n10333) );
  NAND2_X1 U13185 ( .A1(n10692), .A2(n10333), .ZN(n13013) );
  NAND3_X1 U13186 ( .A1(n10330), .A2(n13013), .A3(n10297), .ZN(n10334) );
  NAND2_X1 U13187 ( .A1(n13068), .A2(n10334), .ZN(n10335) );
  NAND2_X1 U13188 ( .A1(n10335), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10336) );
  NAND2_X1 U13189 ( .A1(n10338), .A2(n10370), .ZN(n10374) );
  NAND2_X1 U13190 ( .A1(n10344), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10343) );
  INV_X1 U13191 ( .A(n13088), .ZN(n10341) );
  NAND2_X2 U13192 ( .A1(n10346), .A2(n12987), .ZN(n16591) );
  INV_X1 U13193 ( .A(n10347), .ZN(n10348) );
  OR2_X2 U13194 ( .A1(n16591), .A2(n10348), .ZN(n13087) );
  NAND2_X1 U13195 ( .A1(n13087), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10349) );
  NAND3_X1 U13196 ( .A1(n10350), .A2(n10173), .A3(n10349), .ZN(n10351) );
  NAND2_X1 U13197 ( .A1(n10703), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U13198 ( .A1(n10310), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10352) );
  INV_X1 U13199 ( .A(n10377), .ZN(n10356) );
  AOI21_X1 U13200 ( .B1(n16267), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10357) );
  NAND2_X1 U13201 ( .A1(n10365), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10361) );
  INV_X1 U13202 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10358) );
  AOI21_X1 U13203 ( .B1(n10703), .B2(P2_REIP_REG_2__SCAN_IN), .A(n10359), .ZN(
        n10360) );
  NAND2_X1 U13204 ( .A1(n10361), .A2(n10360), .ZN(n10362) );
  NAND2_X1 U13205 ( .A1(n10363), .A2(n10362), .ZN(n10364) );
  INV_X1 U13206 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13457) );
  INV_X1 U13207 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12501) );
  AOI21_X1 U13208 ( .B1(n10703), .B2(P2_REIP_REG_3__SCAN_IN), .A(n10367), .ZN(
        n10368) );
  INV_X1 U13209 ( .A(n10368), .ZN(n10369) );
  XNOR2_X2 U13210 ( .A(n10709), .B(n10708), .ZN(n10391) );
  BUF_X2 U13211 ( .A(n10391), .Z(n13146) );
  XNOR2_X1 U13212 ( .A(n10372), .B(n10371), .ZN(n10380) );
  AND2_X2 U13213 ( .A1(n13146), .A2(n13689), .ZN(n10407) );
  OR2_X1 U13214 ( .A1(n10375), .A2(n10374), .ZN(n10376) );
  AND2_X2 U13215 ( .A1(n10407), .A2(n10389), .ZN(n10541) );
  AOI22_X1 U13216 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10540), .B1(
        n10541), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10401) );
  INV_X1 U13217 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10384) );
  INV_X1 U13218 ( .A(n10380), .ZN(n14655) );
  AND2_X1 U13219 ( .A1(n14655), .A2(n10389), .ZN(n10381) );
  INV_X1 U13220 ( .A(n10391), .ZN(n13263) );
  NAND2_X2 U13221 ( .A1(n10381), .A2(n13263), .ZN(n19630) );
  NAND2_X2 U13222 ( .A1(n13263), .A2(n10382), .ZN(n19572) );
  INV_X1 U13223 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10383) );
  OAI22_X1 U13224 ( .A1(n10384), .A2(n19630), .B1(n19572), .B2(n10383), .ZN(
        n10388) );
  INV_X1 U13225 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14114) );
  AND2_X1 U13226 ( .A1(n13689), .A2(n10390), .ZN(n10385) );
  NAND2_X2 U13227 ( .A1(n13263), .A2(n10385), .ZN(n10546) );
  AND2_X1 U13228 ( .A1(n13689), .A2(n10389), .ZN(n10386) );
  INV_X1 U13229 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14107) );
  NOR2_X1 U13230 ( .A1(n10388), .A2(n10387), .ZN(n10400) );
  AND2_X2 U13231 ( .A1(n13146), .A2(n14655), .ZN(n10408) );
  AND2_X2 U13232 ( .A1(n10408), .A2(n10390), .ZN(n10543) );
  OR2_X2 U13233 ( .A1(n10391), .A2(n19314), .ZN(n10402) );
  XNOR2_X2 U13234 ( .A(n10393), .B(n10392), .ZN(n19506) );
  INV_X1 U13235 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10396) );
  INV_X1 U13236 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13145) );
  INV_X1 U13237 ( .A(n10397), .ZN(n10398) );
  INV_X1 U13238 ( .A(n10402), .ZN(n10403) );
  NAND2_X2 U13239 ( .A1(n10403), .A2(n13689), .ZN(n10405) );
  NOR2_X4 U13240 ( .A1(n10405), .A2(n19506), .ZN(n10564) );
  NAND2_X1 U13241 ( .A1(n10564), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10412) );
  AND2_X1 U13242 ( .A1(n19506), .A2(n13699), .ZN(n10406) );
  AND2_X2 U13244 ( .A1(n10407), .A2(n10193), .ZN(n10561) );
  NOR2_X4 U13245 ( .A1(n10405), .A2(n13845), .ZN(n10563) );
  NAND2_X1 U13246 ( .A1(n10563), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10410) );
  AND2_X2 U13247 ( .A1(n10408), .A2(n10193), .ZN(n10560) );
  NAND2_X1 U13248 ( .A1(n10414), .A2(n10413), .ZN(n10415) );
  NAND2_X1 U13249 ( .A1(n10415), .A2(n9676), .ZN(n10441) );
  AOI22_X1 U13250 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10604), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13251 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10605), .B1(
        n10606), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10427) );
  AND2_X1 U13252 ( .A1(n10417), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10687) );
  AND2_X2 U13253 ( .A1(n10687), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14420) );
  INV_X1 U13254 ( .A(n14420), .ZN(n13411) );
  NAND2_X1 U13255 ( .A1(n14421), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10421) );
  AND2_X1 U13256 ( .A1(n13696), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10419) );
  NAND2_X1 U13257 ( .A1(n14431), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10420) );
  OAI211_X1 U13258 ( .C1(n13411), .C2(n13145), .A(n10421), .B(n10420), .ZN(
        n10422) );
  INV_X1 U13259 ( .A(n10422), .ZN(n10426) );
  CLKBUF_X3 U13260 ( .A(n10423), .Z(n14593) );
  INV_X1 U13261 ( .A(n10424), .ZN(n14588) );
  AND2_X2 U13262 ( .A1(n10424), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10494) );
  AOI22_X1 U13263 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10468), .B1(
        n10494), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10425) );
  NAND4_X1 U13264 ( .A1(n10428), .A2(n10427), .A3(n10426), .A4(n10425), .ZN(
        n10438) );
  AND2_X2 U13265 ( .A1(n14593), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10578) );
  AOI22_X1 U13266 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14430), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10436) );
  AND2_X2 U13267 ( .A1(n14442), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10645) );
  INV_X1 U13268 ( .A(n10429), .ZN(n14445) );
  AND2_X2 U13269 ( .A1(n10429), .A2(n10261), .ZN(n10430) );
  AOI22_X1 U13270 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10645), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10435) );
  AND2_X1 U13271 ( .A1(n13840), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10432) );
  AND2_X2 U13272 ( .A1(n14440), .A2(n10432), .ZN(n14432) );
  AOI22_X1 U13273 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14404), .B1(
        n14432), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10434) );
  AND2_X2 U13274 ( .A1(n10429), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14433) );
  NAND2_X1 U13275 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10433) );
  NAND4_X1 U13276 ( .A1(n10436), .A2(n10435), .A3(n10434), .A4(n10433), .ZN(
        n10437) );
  NOR2_X1 U13277 ( .A1(n10438), .A2(n10437), .ZN(n12561) );
  INV_X1 U13278 ( .A(n12561), .ZN(n10439) );
  NAND2_X1 U13279 ( .A1(n10439), .A2(n10452), .ZN(n10440) );
  NAND2_X1 U13280 ( .A1(n10441), .A2(n10440), .ZN(n10507) );
  INV_X1 U13281 ( .A(n10507), .ZN(n10505) );
  NOR2_X1 U13282 ( .A1(n10551), .A2(n10442), .ZN(n10443) );
  INV_X1 U13283 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10444) );
  NOR2_X1 U13284 ( .A1(n10552), .A2(n10444), .ZN(n10447) );
  INV_X1 U13285 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10445) );
  INV_X1 U13286 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n21236) );
  OAI22_X1 U13287 ( .A1(n19630), .A2(n10445), .B1(n10547), .B2(n21236), .ZN(
        n10446) );
  NOR2_X1 U13288 ( .A1(n10447), .A2(n10446), .ZN(n10450) );
  AOI22_X1 U13289 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10561), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10449) );
  AOI22_X1 U13290 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10542), .B1(
        n10541), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10448) );
  AND4_X1 U13291 ( .A1(n10451), .A2(n10450), .A3(n10449), .A4(n10448), .ZN(
        n10462) );
  INV_X1 U13292 ( .A(n10559), .ZN(n19993) );
  INV_X1 U13293 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12597) );
  INV_X1 U13294 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10453) );
  OAI21_X1 U13295 ( .B1(n19572), .B2(n10453), .A(n9676), .ZN(n10454) );
  INV_X1 U13296 ( .A(n10454), .ZN(n10456) );
  INV_X1 U13297 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13879) );
  OR2_X1 U13298 ( .A1(n10546), .A2(n13879), .ZN(n10455) );
  INV_X1 U13299 ( .A(n10457), .ZN(n10461) );
  NAND2_X1 U13300 ( .A1(n10563), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10460) );
  AOI22_X1 U13301 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10560), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10459) );
  NAND2_X1 U13302 ( .A1(n10564), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10458) );
  NAND3_X1 U13303 ( .A1(n10462), .A2(n10461), .A3(n10194), .ZN(n10504) );
  AOI22_X1 U13304 ( .A1(n14430), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14420), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13305 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14433), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13306 ( .A1(n10607), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13307 ( .A1(n14431), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13308 ( .A1(n14432), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14404), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13309 ( .A1(n10578), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U13310 ( .A1(n10606), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10605), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10469) );
  NAND4_X1 U13311 ( .A1(n10472), .A2(n10471), .A3(n10470), .A4(n10469), .ZN(
        n10473) );
  OR2_X1 U13312 ( .A1(n12540), .A2(n9676), .ZN(n12897) );
  AOI22_X1 U13313 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14430), .B1(
        n14433), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10477) );
  AOI22_X1 U13314 ( .A1(n10604), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n14420), .ZN(n10476) );
  AOI22_X1 U13315 ( .A1(n10606), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10494), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U13316 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10605), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10474) );
  NAND4_X1 U13317 ( .A1(n10477), .A2(n10476), .A3(n10475), .A4(n10474), .ZN(
        n10483) );
  AOI22_X1 U13318 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14432), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U13319 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14404), .B1(
        n14431), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10480) );
  AOI22_X1 U13320 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10468), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13321 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10578), .B1(
        n10645), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10478) );
  NAND4_X1 U13322 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10482) );
  NOR2_X1 U13323 ( .A1(n10483), .A2(n10482), .ZN(n12546) );
  NOR2_X1 U13324 ( .A1(n12897), .A2(n12546), .ZN(n10514) );
  AOI22_X1 U13325 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n14430), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13326 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10645), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13327 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n14432), .B1(
        n14431), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10485) );
  NAND2_X1 U13328 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10484) );
  AND4_X1 U13329 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10502) );
  AOI22_X1 U13330 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14404), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10492) );
  NAND2_X1 U13331 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10491) );
  INV_X1 U13332 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14049) );
  OR2_X1 U13333 ( .A1(n14417), .A2(n14049), .ZN(n10490) );
  INV_X1 U13334 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10488) );
  OR2_X1 U13335 ( .A1(n14412), .A2(n10488), .ZN(n10489) );
  NAND4_X1 U13336 ( .A1(n10492), .A2(n10491), .A3(n10490), .A4(n10489), .ZN(
        n10500) );
  INV_X1 U13337 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12618) );
  OR2_X1 U13338 ( .A1(n14416), .A2(n12618), .ZN(n10498) );
  INV_X1 U13339 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10493) );
  OR2_X1 U13340 ( .A1(n14411), .A2(n10493), .ZN(n10497) );
  NAND2_X1 U13341 ( .A1(n10468), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10496) );
  NAND2_X1 U13342 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10495) );
  NAND4_X1 U13343 ( .A1(n10498), .A2(n10497), .A3(n10496), .A4(n10495), .ZN(
        n10499) );
  NOR2_X1 U13344 ( .A1(n10500), .A2(n10499), .ZN(n10501) );
  OR2_X1 U13345 ( .A1(n10514), .A2(n10696), .ZN(n10503) );
  NAND2_X1 U13346 ( .A1(n10504), .A2(n10503), .ZN(n10506) );
  NAND2_X1 U13347 ( .A1(n10505), .A2(n10506), .ZN(n10509) );
  INV_X1 U13348 ( .A(n10506), .ZN(n10508) );
  AND2_X2 U13349 ( .A1(n10509), .A2(n10538), .ZN(n13538) );
  INV_X1 U13350 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14633) );
  NAND2_X1 U13351 ( .A1(n12897), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12896) );
  INV_X1 U13352 ( .A(n12896), .ZN(n10511) );
  INV_X1 U13353 ( .A(n12546), .ZN(n10510) );
  XNOR2_X1 U13354 ( .A(n12540), .B(n10510), .ZN(n10512) );
  NAND2_X1 U13355 ( .A1(n10511), .A2(n10512), .ZN(n10513) );
  XOR2_X1 U13356 ( .A(n10512), .B(n10511), .Z(n14340) );
  NAND2_X1 U13357 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14340), .ZN(
        n14339) );
  NAND2_X1 U13358 ( .A1(n10513), .A2(n14339), .ZN(n10515) );
  XNOR2_X1 U13359 ( .A(n14633), .B(n10515), .ZN(n14632) );
  NAND2_X1 U13360 ( .A1(n14632), .A2(n14631), .ZN(n14630) );
  NAND2_X1 U13361 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10515), .ZN(
        n10516) );
  NAND2_X1 U13362 ( .A1(n14630), .A2(n10516), .ZN(n10517) );
  INV_X1 U13363 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14291) );
  XNOR2_X1 U13364 ( .A(n10517), .B(n14291), .ZN(n13539) );
  NAND2_X1 U13365 ( .A1(n13538), .A2(n13539), .ZN(n10519) );
  NAND2_X1 U13366 ( .A1(n10517), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10518) );
  AOI22_X1 U13367 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10604), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13368 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10605), .B1(
        n10606), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10525) );
  INV_X1 U13369 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13178) );
  NAND2_X1 U13370 ( .A1(n14404), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10521) );
  NAND2_X1 U13371 ( .A1(n14421), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10520) );
  OAI211_X1 U13372 ( .C1(n13411), .C2(n13178), .A(n10521), .B(n10520), .ZN(
        n10522) );
  INV_X1 U13373 ( .A(n10522), .ZN(n10524) );
  AOI22_X1 U13374 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10494), .B1(
        n14430), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10523) );
  NAND4_X1 U13375 ( .A1(n10526), .A2(n10525), .A3(n10524), .A4(n10523), .ZN(
        n10532) );
  AOI22_X1 U13376 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10468), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13377 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10645), .B1(
        n14433), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13378 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14432), .B1(
        n14431), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10528) );
  NAND2_X1 U13379 ( .A1(n10430), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10527) );
  NAND4_X1 U13380 ( .A1(n10530), .A2(n10529), .A3(n10528), .A4(n10527), .ZN(
        n10531) );
  XNOR2_X1 U13381 ( .A(n10538), .B(n12532), .ZN(n10534) );
  NAND2_X1 U13382 ( .A1(n10533), .A2(n10534), .ZN(n13787) );
  INV_X1 U13383 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13954) );
  NAND2_X1 U13384 ( .A1(n13787), .A2(n13954), .ZN(n10537) );
  INV_X1 U13385 ( .A(n10533), .ZN(n10536) );
  INV_X1 U13386 ( .A(n10534), .ZN(n10535) );
  NAND2_X1 U13387 ( .A1(n10536), .A2(n10535), .ZN(n13788) );
  AOI22_X1 U13388 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n10540), .B1(
        n10541), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13389 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n10542), .B1(
        n10543), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10557) );
  INV_X1 U13390 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10545) );
  INV_X1 U13391 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10544) );
  OAI22_X1 U13392 ( .A1(n10545), .A2(n19630), .B1(n19572), .B2(n10544), .ZN(
        n10550) );
  INV_X1 U13393 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10548) );
  INV_X1 U13394 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14373) );
  OAI22_X1 U13395 ( .A1(n10548), .A2(n10546), .B1(n19752), .B2(n14373), .ZN(
        n10549) );
  NOR2_X1 U13396 ( .A1(n10550), .A2(n10549), .ZN(n10556) );
  INV_X1 U13397 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13271) );
  INV_X1 U13398 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10553) );
  OAI22_X1 U13399 ( .A1(n13271), .A2(n10551), .B1(n19600), .B2(n10553), .ZN(
        n10554) );
  INV_X1 U13400 ( .A(n10554), .ZN(n10555) );
  NAND4_X1 U13401 ( .A1(n10558), .A2(n10557), .A3(n10556), .A4(n10555), .ZN(
        n10570) );
  AOI22_X1 U13402 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n10559), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13403 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n10561), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10567) );
  NAND2_X1 U13404 ( .A1(n10563), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10566) );
  NAND2_X1 U13405 ( .A1(n10564), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10565) );
  NAND4_X1 U13406 ( .A1(n10568), .A2(n10567), .A3(n10566), .A4(n10565), .ZN(
        n10569) );
  AOI22_X1 U13407 ( .A1(n10604), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10606), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10577) );
  AOI22_X1 U13408 ( .A1(n10607), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10605), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10576) );
  NAND2_X1 U13409 ( .A1(n14404), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10572) );
  NAND2_X1 U13410 ( .A1(n14421), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10571) );
  OAI211_X1 U13411 ( .C1(n13411), .C2(n13271), .A(n10572), .B(n10571), .ZN(
        n10573) );
  INV_X1 U13412 ( .A(n10573), .ZN(n10575) );
  AOI22_X1 U13413 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10574) );
  NAND4_X1 U13414 ( .A1(n10577), .A2(n10576), .A3(n10575), .A4(n10574), .ZN(
        n10584) );
  AOI22_X1 U13415 ( .A1(n14430), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10582) );
  AOI22_X1 U13416 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14433), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10581) );
  AOI22_X1 U13417 ( .A1(n14432), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14431), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10580) );
  NAND2_X1 U13418 ( .A1(n10430), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10579) );
  NAND4_X1 U13419 ( .A1(n10582), .A2(n10581), .A3(n10580), .A4(n10579), .ZN(
        n10583) );
  INV_X1 U13420 ( .A(n10809), .ZN(n10585) );
  NAND2_X1 U13421 ( .A1(n10585), .A2(n10452), .ZN(n10586) );
  INV_X1 U13422 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13955) );
  NAND2_X1 U13423 ( .A1(n10859), .A2(n13955), .ZN(n13950) );
  INV_X1 U13424 ( .A(n10635), .ZN(n10629) );
  AOI22_X1 U13425 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10541), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U13426 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10543), .B1(
        n10560), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10596) );
  INV_X1 U13427 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10589) );
  INV_X1 U13428 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10588) );
  OAI22_X1 U13429 ( .A1(n10589), .A2(n19630), .B1(n19572), .B2(n10588), .ZN(
        n10591) );
  INV_X1 U13430 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14397) );
  INV_X1 U13431 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14390) );
  OAI22_X1 U13432 ( .A1(n14397), .A2(n10546), .B1(n19752), .B2(n14390), .ZN(
        n10590) );
  NOR2_X1 U13433 ( .A1(n10591), .A2(n10590), .ZN(n10595) );
  INV_X1 U13434 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10610) );
  INV_X1 U13435 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10592) );
  OAI22_X1 U13436 ( .A1(n10610), .A2(n10551), .B1(n19600), .B2(n10592), .ZN(
        n10593) );
  INV_X1 U13437 ( .A(n10593), .ZN(n10594) );
  NAND4_X1 U13438 ( .A1(n10597), .A2(n10596), .A3(n10595), .A4(n10594), .ZN(
        n10603) );
  AOI22_X1 U13439 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10542), .B1(
        n10559), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U13440 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10561), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10600) );
  NAND2_X1 U13441 ( .A1(n10563), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10599) );
  NAND2_X1 U13442 ( .A1(n10564), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10598) );
  NAND4_X1 U13443 ( .A1(n10601), .A2(n10600), .A3(n10599), .A4(n10598), .ZN(
        n10602) );
  AOI22_X1 U13444 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10605), .B1(
        n10604), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13445 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10607), .B1(
        n10606), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10614) );
  NAND2_X1 U13446 ( .A1(n14421), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10609) );
  NAND2_X1 U13447 ( .A1(n14431), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10608) );
  OAI211_X1 U13448 ( .C1(n13411), .C2(n10610), .A(n10609), .B(n10608), .ZN(
        n10611) );
  INV_X1 U13449 ( .A(n10611), .ZN(n10613) );
  AOI22_X1 U13450 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10494), .B1(
        n14430), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10612) );
  NAND4_X1 U13451 ( .A1(n10615), .A2(n10614), .A3(n10613), .A4(n10612), .ZN(
        n10621) );
  AOI22_X1 U13452 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10468), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13453 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10645), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13454 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14404), .B1(
        n14432), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U13455 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10616) );
  NAND4_X1 U13456 ( .A1(n10619), .A2(n10618), .A3(n10617), .A4(n10616), .ZN(
        n10620) );
  INV_X1 U13457 ( .A(n10811), .ZN(n12564) );
  NAND2_X1 U13458 ( .A1(n12564), .A2(n10452), .ZN(n10622) );
  NAND2_X1 U13459 ( .A1(n10626), .A2(n10631), .ZN(n10627) );
  AND2_X2 U13460 ( .A1(n10638), .A2(n10627), .ZN(n10819) );
  NAND2_X1 U13461 ( .A1(n10629), .A2(n10628), .ZN(n10634) );
  INV_X1 U13462 ( .A(n10859), .ZN(n10630) );
  NAND3_X1 U13463 ( .A1(n10635), .A2(n10819), .A3(n10636), .ZN(n10633) );
  NAND2_X1 U13464 ( .A1(n13952), .A2(n10631), .ZN(n10632) );
  NAND3_X1 U13465 ( .A1(n10634), .A2(n10633), .A3(n10632), .ZN(n14069) );
  NAND2_X1 U13466 ( .A1(n13953), .A2(n10636), .ZN(n10637) );
  AOI22_X1 U13467 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14431), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10644) );
  NAND2_X1 U13468 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10643) );
  INV_X1 U13469 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10639) );
  OR2_X1 U13470 ( .A1(n14417), .A2(n10639), .ZN(n10642) );
  INV_X1 U13471 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10640) );
  OR2_X1 U13472 ( .A1(n14411), .A2(n10640), .ZN(n10641) );
  INV_X1 U13473 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14413) );
  INV_X1 U13474 ( .A(n10645), .ZN(n10647) );
  INV_X1 U13475 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14424) );
  OAI22_X1 U13476 ( .A1(n14413), .A2(n10647), .B1(n10646), .B2(n14424), .ZN(
        n10651) );
  INV_X1 U13477 ( .A(n14433), .ZN(n10690) );
  INV_X1 U13478 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12726) );
  NAND2_X1 U13479 ( .A1(n14404), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10649) );
  NAND2_X1 U13480 ( .A1(n14432), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10648) );
  OAI211_X1 U13481 ( .C1(n10690), .C2(n12726), .A(n10649), .B(n10648), .ZN(
        n10650) );
  NOR2_X1 U13482 ( .A1(n10651), .A2(n10650), .ZN(n10659) );
  INV_X1 U13483 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10652) );
  OR2_X1 U13484 ( .A1(n14412), .A2(n10652), .ZN(n10656) );
  INV_X1 U13485 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12731) );
  OR2_X1 U13486 ( .A1(n14416), .A2(n12731), .ZN(n10655) );
  NAND2_X1 U13487 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10654) );
  NAND2_X1 U13488 ( .A1(n14430), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10653) );
  AOI22_X1 U13489 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10468), .B1(
        n10578), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10657) );
  NAND4_X1 U13490 ( .A1(n10660), .A2(n10659), .A3(n10658), .A4(n10657), .ZN(
        n10814) );
  INV_X1 U13491 ( .A(n10814), .ZN(n10869) );
  INV_X1 U13492 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10877) );
  AND2_X1 U13493 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10661) );
  INV_X1 U13494 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16557) );
  OAI21_X1 U13495 ( .B1(n10638), .B2(n10869), .A(n16557), .ZN(n10663) );
  NAND2_X1 U13496 ( .A1(n10664), .A2(n10663), .ZN(n16516) );
  INV_X1 U13497 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16156) );
  INV_X1 U13498 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16137) );
  NOR2_X1 U13499 ( .A1(n16156), .A2(n16137), .ZN(n16138) );
  AND4_X1 U13500 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(n16138), .ZN(n16002) );
  NAND2_X1 U13501 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16055) );
  INV_X1 U13502 ( .A(n16055), .ZN(n10666) );
  AND2_X1 U13503 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10665) );
  NAND2_X1 U13504 ( .A1(n10666), .A2(n10665), .ZN(n16008) );
  INV_X1 U13505 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16010) );
  INV_X1 U13506 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15781) );
  NAND2_X1 U13507 ( .A1(n10667), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15778) );
  INV_X1 U13508 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15977) );
  NOR2_X2 U13509 ( .A1(n15778), .A2(n15977), .ZN(n15751) );
  INV_X1 U13510 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15922) );
  INV_X1 U13511 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15894) );
  AOI21_X1 U13512 ( .B1(n15882), .B2(n15707), .A(n15691), .ZN(n14621) );
  XNOR2_X1 U13513 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10693) );
  NAND2_X1 U13514 ( .A1(n10693), .A2(n10682), .ZN(n10669) );
  NAND2_X1 U13515 ( .A1(n20199), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10668) );
  NAND2_X1 U13516 ( .A1(n10669), .A2(n10668), .ZN(n10678) );
  XNOR2_X1 U13517 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10676) );
  NAND2_X1 U13518 ( .A1(n10678), .A2(n10676), .ZN(n10671) );
  NAND2_X1 U13519 ( .A1(n20190), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10670) );
  NAND2_X1 U13520 ( .A1(n10671), .A2(n10670), .ZN(n10673) );
  XNOR2_X1 U13521 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10672) );
  NOR2_X1 U13522 ( .A1(n10673), .A2(n10672), .ZN(n10674) );
  INV_X1 U13523 ( .A(n10676), .ZN(n10677) );
  XNOR2_X1 U13524 ( .A(n10678), .B(n10677), .ZN(n12954) );
  NAND2_X1 U13525 ( .A1(n12971), .A2(n12954), .ZN(n10685) );
  XNOR2_X1 U13526 ( .A(n10693), .B(n10682), .ZN(n12956) );
  INV_X1 U13527 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16268) );
  NOR2_X1 U13528 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16268), .ZN(
        n10680) );
  OAI22_X1 U13529 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13026), .B1(
        n10680), .B2(n10679), .ZN(n12978) );
  INV_X1 U13530 ( .A(n12978), .ZN(n12974) );
  INV_X1 U13531 ( .A(n10682), .ZN(n10684) );
  NAND2_X1 U13532 ( .A1(n13696), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10683) );
  NAND2_X1 U13533 ( .A1(n10684), .A2(n10683), .ZN(n12955) );
  OR2_X1 U13534 ( .A1(n10685), .A2(n12955), .ZN(n10686) );
  NAND2_X1 U13535 ( .A1(n16590), .A2(n10686), .ZN(n10691) );
  NOR2_X1 U13536 ( .A1(n10687), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13023) );
  INV_X1 U13537 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n10688) );
  NAND2_X1 U13538 ( .A1(n10688), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10689) );
  AOI21_X1 U13539 ( .B1(n10690), .B2(n13023), .A(n10689), .ZN(n20201) );
  AOI21_X1 U13540 ( .B1(n10691), .B2(n10785), .A(n20201), .ZN(n20217) );
  INV_X1 U13541 ( .A(n10692), .ZN(n16598) );
  NAND3_X1 U13542 ( .A1(n20217), .A2(n16598), .A3(n9676), .ZN(n10699) );
  INV_X1 U13543 ( .A(n10693), .ZN(n10694) );
  NOR2_X1 U13544 ( .A1(n12955), .A2(n10694), .ZN(n12964) );
  MUX2_X1 U13545 ( .A(n10696), .B(n12954), .S(n12963), .Z(n10805) );
  OAI21_X1 U13546 ( .B1(n12964), .B2(n10805), .A(n12971), .ZN(n10697) );
  NAND2_X1 U13547 ( .A1(n10697), .A2(n12974), .ZN(n20213) );
  NAND2_X1 U13548 ( .A1(n10297), .A2(n10452), .ZN(n12981) );
  NAND2_X1 U13549 ( .A1(n10699), .A2(n10698), .ZN(n13051) );
  NAND2_X1 U13550 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n10785), .ZN(n19133) );
  INV_X1 U13551 ( .A(n19133), .ZN(n10700) );
  INV_X1 U13552 ( .A(n20095), .ZN(n16622) );
  NOR2_X1 U13553 ( .A1(n13056), .A2(n16622), .ZN(n10701) );
  INV_X1 U13554 ( .A(n12847), .ZN(n10702) );
  NAND2_X1 U13555 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10707) );
  INV_X1 U13556 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10704) );
  INV_X1 U13557 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15515) );
  AOI21_X1 U13558 ( .B1(n10736), .B2(P2_REIP_REG_10__SCAN_IN), .A(n10705), 
        .ZN(n10706) );
  NAND2_X1 U13559 ( .A1(n10707), .A2(n10706), .ZN(n13352) );
  NAND2_X1 U13560 ( .A1(n10709), .A2(n10708), .ZN(n10714) );
  INV_X1 U13561 ( .A(n10710), .ZN(n10711) );
  OR2_X1 U13562 ( .A1(n10712), .A2(n10711), .ZN(n10713) );
  CLKBUF_X3 U13563 ( .A(n10366), .Z(n12790) );
  NAND2_X1 U13564 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10717) );
  INV_X1 U13565 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13185) );
  AOI21_X1 U13566 ( .B1(n10736), .B2(P2_REIP_REG_4__SCAN_IN), .A(n10715), .ZN(
        n10716) );
  NAND2_X1 U13567 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10722) );
  INV_X1 U13568 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13245) );
  INV_X1 U13569 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10719) );
  AOI21_X1 U13570 ( .B1(n10736), .B2(P2_REIP_REG_5__SCAN_IN), .A(n10720), .ZN(
        n10721) );
  NAND2_X1 U13571 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10726) );
  INV_X1 U13572 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19284) );
  INV_X1 U13573 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10723) );
  AOI21_X1 U13574 ( .B1(n10736), .B2(P2_REIP_REG_6__SCAN_IN), .A(n10724), .ZN(
        n10725) );
  NAND2_X1 U13575 ( .A1(n10726), .A2(n10725), .ZN(n13275) );
  NAND2_X1 U13576 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10730) );
  INV_X1 U13577 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10813) );
  INV_X1 U13578 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10727) );
  AOI21_X1 U13579 ( .B1(n10736), .B2(P2_REIP_REG_7__SCAN_IN), .A(n10728), .ZN(
        n10729) );
  AOI22_X1 U13580 ( .A1(n9663), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10732) );
  NAND2_X1 U13581 ( .A1(n10736), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10731) );
  OAI211_X1 U13582 ( .C1(n14286), .C2(n16557), .A(n10732), .B(n10731), .ZN(
        n13528) );
  NAND2_X1 U13583 ( .A1(n10736), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13584 ( .A1(n9663), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10733) );
  NAND2_X1 U13585 ( .A1(n10734), .A2(n10733), .ZN(n10735) );
  AOI21_X1 U13586 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10735), .ZN(n13418) );
  INV_X1 U13587 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U13588 ( .A1(n9663), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n10737) );
  OAI21_X1 U13589 ( .B1(n12788), .B2(n10738), .A(n10737), .ZN(n10739) );
  AOI21_X1 U13590 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10739), .ZN(n13506) );
  NOR2_X2 U13591 ( .A1(n13507), .A2(n13506), .ZN(n13509) );
  NAND2_X1 U13592 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10742) );
  AOI21_X1 U13593 ( .B1(n10736), .B2(P2_REIP_REG_12__SCAN_IN), .A(n10740), 
        .ZN(n10741) );
  NAND2_X1 U13594 ( .A1(n10742), .A2(n10741), .ZN(n13434) );
  NAND2_X1 U13595 ( .A1(n13509), .A2(n13434), .ZN(n13433) );
  INV_X1 U13596 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n16109) );
  AOI22_X1 U13597 ( .A1(n9663), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10743) );
  OAI21_X1 U13598 ( .B1(n12788), .B2(n16109), .A(n10743), .ZN(n10744) );
  AOI21_X1 U13599 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10744), .ZN(n13474) );
  INV_X1 U13600 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U13601 ( .A1(n9663), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10745) );
  OAI21_X1 U13602 ( .B1(n12788), .B2(n12721), .A(n10745), .ZN(n10746) );
  AOI21_X1 U13603 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n10746), .ZN(n13617) );
  INV_X1 U13604 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n15841) );
  AOI22_X1 U13605 ( .A1(n9663), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10747) );
  OAI21_X1 U13606 ( .B1(n12788), .B2(n15841), .A(n10747), .ZN(n10748) );
  AOI21_X1 U13607 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10748), .ZN(n12816) );
  NAND2_X1 U13608 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10751) );
  INV_X1 U13609 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n13936) );
  INV_X1 U13610 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15826) );
  AOI21_X1 U13611 ( .B1(n10736), .B2(P2_REIP_REG_16__SCAN_IN), .A(n10749), 
        .ZN(n10750) );
  NAND2_X1 U13612 ( .A1(n10751), .A2(n10750), .ZN(n13930) );
  NAND2_X1 U13613 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10754) );
  INV_X1 U13614 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15817) );
  AOI21_X1 U13615 ( .B1(n10736), .B2(P2_REIP_REG_17__SCAN_IN), .A(n10752), 
        .ZN(n10753) );
  NAND2_X1 U13616 ( .A1(n10754), .A2(n10753), .ZN(n13870) );
  NAND2_X1 U13617 ( .A1(n13933), .A2(n13870), .ZN(n13869) );
  INV_X1 U13618 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13619 ( .A1(n9663), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10755) );
  OAI21_X1 U13620 ( .B1(n12788), .B2(n10756), .A(n10755), .ZN(n10757) );
  AOI21_X1 U13621 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n10757), .ZN(n14062) );
  INV_X1 U13622 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13623 ( .A1(n9663), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10758) );
  OAI21_X1 U13624 ( .B1(n12788), .B2(n10759), .A(n10758), .ZN(n10760) );
  AOI21_X1 U13625 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10760), .ZN(n14103) );
  INV_X1 U13626 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U13627 ( .A1(n9663), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10761) );
  OAI21_X1 U13628 ( .B1(n12788), .B2(n12749), .A(n10761), .ZN(n10762) );
  AOI21_X1 U13629 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10762), .ZN(n15587) );
  INV_X1 U13630 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15583) );
  INV_X1 U13631 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10763) );
  AOI21_X1 U13632 ( .B1(n10736), .B2(P2_REIP_REG_21__SCAN_IN), .A(n10764), 
        .ZN(n10765) );
  OAI21_X1 U13633 ( .B1(n14286), .B2(n15781), .A(n10765), .ZN(n15581) );
  INV_X1 U13634 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U13635 ( .A1(n9663), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10766) );
  OAI21_X1 U13636 ( .B1(n12788), .B2(n10767), .A(n10766), .ZN(n10768) );
  AOI21_X1 U13637 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10768), .ZN(n15483) );
  OR2_X2 U13638 ( .A1(n15482), .A2(n15483), .ZN(n15485) );
  INV_X1 U13639 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13640 ( .A1(n9663), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10769) );
  OAI21_X1 U13641 ( .B1(n12788), .B2(n10770), .A(n10769), .ZN(n10771) );
  AOI21_X1 U13642 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10771), .ZN(n15469) );
  NAND2_X1 U13643 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10774) );
  INV_X1 U13644 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16464) );
  AOI21_X1 U13645 ( .B1(n10736), .B2(P2_REIP_REG_24__SCAN_IN), .A(n10772), 
        .ZN(n10773) );
  NAND2_X1 U13646 ( .A1(n10774), .A2(n10773), .ZN(n15560) );
  NAND2_X1 U13647 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10777) );
  INV_X1 U13648 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15553) );
  INV_X1 U13649 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15736) );
  AOI21_X1 U13650 ( .B1(n10736), .B2(P2_REIP_REG_25__SCAN_IN), .A(n10775), 
        .ZN(n10776) );
  NAND2_X1 U13651 ( .A1(n10777), .A2(n10776), .ZN(n15453) );
  INV_X1 U13652 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n16455) );
  AOI22_X1 U13653 ( .A1(n9663), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10778) );
  OAI21_X1 U13654 ( .B1(n12788), .B2(n16455), .A(n10778), .ZN(n10779) );
  AOI21_X1 U13655 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10779), .ZN(n15546) );
  INV_X1 U13656 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20157) );
  AOI22_X1 U13657 ( .A1(n9663), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n10780) );
  OAI21_X1 U13658 ( .B1(n12788), .B2(n20157), .A(n10780), .ZN(n10781) );
  AOI21_X1 U13659 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10781), .ZN(n12828) );
  NAND2_X1 U13660 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10784) );
  INV_X1 U13661 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n10785) );
  INV_X1 U13662 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15706) );
  AOI21_X1 U13663 ( .B1(n10736), .B2(P2_REIP_REG_28__SCAN_IN), .A(n10782), 
        .ZN(n10783) );
  NAND2_X1 U13664 ( .A1(n10784), .A2(n10783), .ZN(n15436) );
  NAND2_X1 U13665 ( .A1(n12790), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10788) );
  INV_X1 U13666 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10799) );
  AOI21_X1 U13667 ( .B1(n10736), .B2(P2_REIP_REG_29__SCAN_IN), .A(n10786), 
        .ZN(n10787) );
  NAND2_X1 U13668 ( .A1(n10788), .A2(n10787), .ZN(n10789) );
  OR2_X1 U13669 ( .A1(n15439), .A2(n10789), .ZN(n10790) );
  NAND2_X1 U13670 ( .A1(n14282), .A2(n10790), .ZN(n16441) );
  NAND2_X1 U13671 ( .A1(n10785), .A2(n20041), .ZN(n13403) );
  NAND2_X1 U13672 ( .A1(n20183), .A2(n13403), .ZN(n20191) );
  NAND2_X1 U13673 ( .A1(n20191), .A2(n16267), .ZN(n10791) );
  AND2_X1 U13674 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20192) );
  AND2_X1 U13675 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10792) );
  AND2_X1 U13676 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10793) );
  NAND2_X1 U13677 ( .A1(n12492), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12489) );
  INV_X1 U13678 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15840) );
  AND2_X1 U13679 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10794) );
  NAND2_X1 U13680 ( .A1(n12504), .A2(n10794), .ZN(n12487) );
  INV_X1 U13681 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10795) );
  OR2_X1 U13682 ( .A1(n10795), .A2(n10763), .ZN(n10796) );
  INV_X1 U13683 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15754) );
  INV_X1 U13684 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15723) );
  INV_X1 U13685 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15714) );
  INV_X1 U13686 ( .A(n12485), .ZN(n12515) );
  NAND2_X1 U13687 ( .A1(n9789), .A2(n10799), .ZN(n10797) );
  AND2_X1 U13688 ( .A1(n12515), .A2(n10797), .ZN(n16434) );
  NAND2_X1 U13689 ( .A1(n16267), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13168) );
  OAI21_X1 U13690 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n10785), .A(n13168), 
        .ZN(n10798) );
  NOR2_X1 U13691 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16617) );
  NAND2_X1 U13692 ( .A1(n16617), .A2(n20041), .ZN(n12841) );
  INV_X2 U13693 ( .A(n19277), .ZN(n19303) );
  NAND2_X1 U13694 ( .A1(n19303), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n14610) );
  OAI21_X1 U13695 ( .B1(n16541), .B2(n10799), .A(n14610), .ZN(n10800) );
  AOI21_X1 U13696 ( .B1(n16434), .B2(n16533), .A(n10800), .ZN(n10801) );
  OAI21_X1 U13697 ( .B1(n16441), .B2(n16526), .A(n10801), .ZN(n10802) );
  AOI21_X1 U13698 ( .B1(n14621), .B2(n16529), .A(n10802), .ZN(n10993) );
  INV_X1 U13699 ( .A(n12972), .ZN(n10803) );
  MUX2_X1 U13700 ( .A(n12532), .B(n10803), .S(n12963), .Z(n10804) );
  INV_X4 U13701 ( .A(n12530), .ZN(n10812) );
  MUX2_X1 U13702 ( .A(n10804), .B(n13185), .S(n10812), .Z(n10840) );
  MUX2_X1 U13703 ( .A(n10805), .B(n10358), .S(n10812), .Z(n10830) );
  OR2_X1 U13704 ( .A1(n12546), .A2(n10812), .ZN(n10807) );
  INV_X1 U13705 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13235) );
  INV_X1 U13706 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13708) );
  NAND2_X1 U13707 ( .A1(n10831), .A2(n13708), .ZN(n10806) );
  NAND2_X1 U13708 ( .A1(n10807), .A2(n10806), .ZN(n10833) );
  MUX2_X1 U13709 ( .A(n12561), .B(n12967), .S(n12963), .Z(n10808) );
  MUX2_X1 U13710 ( .A(n10808), .B(P2_EBX_REG_3__SCAN_IN), .S(n10812), .Z(
        n10825) );
  NOR2_X2 U13711 ( .A1(n10829), .A2(n10825), .ZN(n10839) );
  NAND2_X1 U13712 ( .A1(n12530), .A2(n10809), .ZN(n12525) );
  NAND2_X1 U13713 ( .A1(n10812), .A2(n13245), .ZN(n10810) );
  MUX2_X1 U13714 ( .A(n10811), .B(n19284), .S(n10812), .Z(n10820) );
  MUX2_X1 U13715 ( .A(n10814), .B(n10813), .S(n10812), .Z(n10864) );
  INV_X1 U13716 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n21083) );
  NAND2_X1 U13717 ( .A1(n10812), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10868) );
  INV_X1 U13718 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13423) );
  NAND2_X1 U13719 ( .A1(n10812), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10893) );
  NAND2_X1 U13720 ( .A1(n10812), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10923) );
  OAI21_X1 U13721 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n10812), .ZN(n10815) );
  NAND2_X1 U13722 ( .A1(n10812), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10910) );
  OAI21_X1 U13723 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(P2_EBX_REG_18__SCAN_IN), 
        .A(n10812), .ZN(n10816) );
  NAND2_X1 U13724 ( .A1(n10812), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10817) );
  AND2_X1 U13725 ( .A1(n10812), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10954) );
  NAND2_X1 U13726 ( .A1(n10812), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10975) );
  AND2_X1 U13727 ( .A1(n10812), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10978) );
  NAND2_X1 U13728 ( .A1(n10812), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12518) );
  XNOR2_X1 U13729 ( .A(n12519), .B(n12518), .ZN(n10818) );
  INV_X1 U13730 ( .A(n10818), .ZN(n16439) );
  NAND3_X1 U13731 ( .A1(n16439), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14277), .ZN(n15683) );
  OAI21_X1 U13732 ( .B1(n10818), .B2(n10869), .A(n15882), .ZN(n14270) );
  NAND2_X1 U13733 ( .A1(n15683), .A2(n14270), .ZN(n10989) );
  NAND2_X1 U13734 ( .A1(n10819), .A2(n10869), .ZN(n10823) );
  INV_X1 U13735 ( .A(n10866), .ZN(n10822) );
  OR2_X1 U13736 ( .A1(n10845), .A2(n10820), .ZN(n10821) );
  NAND2_X1 U13737 ( .A1(n10822), .A2(n10821), .ZN(n19286) );
  INV_X1 U13738 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10824) );
  NAND2_X1 U13739 ( .A1(n13538), .A2(n10869), .ZN(n10828) );
  INV_X1 U13740 ( .A(n10839), .ZN(n10827) );
  NAND2_X1 U13741 ( .A1(n10829), .A2(n10825), .ZN(n10826) );
  NAND2_X1 U13742 ( .A1(n10827), .A2(n10826), .ZN(n13461) );
  NAND2_X1 U13743 ( .A1(n10828), .A2(n13461), .ZN(n13537) );
  OAI21_X1 U13744 ( .B1(n10833), .B2(n10830), .A(n10829), .ZN(n13687) );
  MUX2_X1 U13745 ( .A(n12955), .B(n12540), .S(n13082), .Z(n10832) );
  AOI21_X1 U13746 ( .B1(n10832), .B2(n12530), .A(n10831), .ZN(n19316) );
  NAND2_X1 U13747 ( .A1(n19316), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14336) );
  INV_X1 U13748 ( .A(n10833), .ZN(n10835) );
  NAND3_X1 U13749 ( .A1(n10812), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n10834) );
  NAND2_X1 U13750 ( .A1(n10835), .A2(n10834), .ZN(n14335) );
  NOR2_X1 U13751 ( .A1(n14336), .A2(n14335), .ZN(n10836) );
  NAND2_X1 U13752 ( .A1(n14336), .A2(n14335), .ZN(n14334) );
  OAI21_X1 U13753 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10836), .A(
        n14334), .ZN(n14635) );
  XNOR2_X1 U13754 ( .A(n13687), .B(n14633), .ZN(n14634) );
  OR2_X1 U13755 ( .A1(n14635), .A2(n14634), .ZN(n14652) );
  OAI21_X1 U13756 ( .B1(n13687), .B2(n14633), .A(n14652), .ZN(n13535) );
  NAND2_X1 U13757 ( .A1(n13537), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10837) );
  NAND2_X1 U13758 ( .A1(n10838), .A2(n10837), .ZN(n13792) );
  OAI21_X1 U13759 ( .B1(n10840), .B2(n10839), .A(n10847), .ZN(n13560) );
  XNOR2_X1 U13760 ( .A(n13560), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13790) );
  NAND2_X1 U13761 ( .A1(n13792), .A2(n13790), .ZN(n10843) );
  INV_X1 U13762 ( .A(n13560), .ZN(n10841) );
  NAND2_X1 U13763 ( .A1(n10841), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10842) );
  NAND2_X1 U13764 ( .A1(n10843), .A2(n10842), .ZN(n13947) );
  NAND2_X1 U13765 ( .A1(n10847), .A2(n10846), .ZN(n10848) );
  NAND2_X1 U13766 ( .A1(n9928), .A2(n10848), .ZN(n19301) );
  AND2_X1 U13767 ( .A1(n19301), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10852) );
  INV_X1 U13768 ( .A(n10852), .ZN(n10850) );
  NOR2_X1 U13769 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10853) );
  INV_X1 U13770 ( .A(n10853), .ZN(n10849) );
  MUX2_X1 U13771 ( .A(n10850), .B(n10849), .S(n10851), .Z(n10858) );
  MUX2_X1 U13772 ( .A(n10853), .B(n10852), .S(n10851), .Z(n10854) );
  NAND2_X1 U13773 ( .A1(n10844), .A2(n10854), .ZN(n10857) );
  OAI21_X1 U13774 ( .B1(n10869), .B2(n13955), .A(n19301), .ZN(n10855) );
  OAI21_X1 U13775 ( .B1(n19301), .B2(n13955), .A(n10855), .ZN(n10856) );
  OAI211_X1 U13776 ( .C1(n10844), .C2(n10858), .A(n10857), .B(n10856), .ZN(
        n13948) );
  NAND2_X1 U13777 ( .A1(n13947), .A2(n13948), .ZN(n10861) );
  INV_X1 U13778 ( .A(n10864), .ZN(n10865) );
  XNOR2_X1 U13779 ( .A(n10866), .B(n10865), .ZN(n19276) );
  NAND2_X1 U13780 ( .A1(n19276), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14234) );
  INV_X1 U13781 ( .A(n10871), .ZN(n10867) );
  OAI21_X1 U13782 ( .B1(n9735), .B2(n10868), .A(n10867), .ZN(n13608) );
  OR2_X1 U13783 ( .A1(n13608), .A2(n10869), .ZN(n10876) );
  INV_X1 U13784 ( .A(n10876), .ZN(n10870) );
  NAND2_X1 U13785 ( .A1(n10870), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16519) );
  NAND2_X1 U13786 ( .A1(n10812), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10872) );
  MUX2_X1 U13787 ( .A(n10872), .B(n10812), .S(n10871), .Z(n10874) );
  INV_X1 U13788 ( .A(n10879), .ZN(n10873) );
  NAND2_X1 U13789 ( .A1(n19261), .A2(n14277), .ZN(n10875) );
  INV_X1 U13790 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16171) );
  NAND2_X1 U13791 ( .A1(n10875), .A2(n16171), .ZN(n16146) );
  NAND2_X1 U13792 ( .A1(n10876), .A2(n16557), .ZN(n16518) );
  INV_X1 U13793 ( .A(n19276), .ZN(n10878) );
  NAND2_X1 U13794 ( .A1(n10878), .A2(n10877), .ZN(n14235) );
  AND2_X1 U13795 ( .A1(n16518), .A2(n14235), .ZN(n15871) );
  NAND2_X1 U13796 ( .A1(n10879), .A2(n10704), .ZN(n10883) );
  NOR2_X1 U13797 ( .A1(n10879), .A2(n10704), .ZN(n10880) );
  NAND2_X1 U13798 ( .A1(n10812), .A2(n10880), .ZN(n10881) );
  AND2_X1 U13799 ( .A1(n10967), .A2(n10881), .ZN(n10882) );
  NAND2_X1 U13800 ( .A1(n10883), .A2(n10882), .ZN(n15516) );
  OR2_X1 U13801 ( .A1(n15516), .A2(n10869), .ZN(n10884) );
  NAND2_X1 U13802 ( .A1(n10884), .A2(n16156), .ZN(n16151) );
  AND2_X1 U13803 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10885) );
  NAND2_X1 U13804 ( .A1(n19261), .A2(n10885), .ZN(n16147) );
  NAND2_X1 U13805 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10886) );
  OR2_X1 U13806 ( .A1(n15516), .A2(n10886), .ZN(n16150) );
  AND3_X1 U13807 ( .A1(n10812), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10883), .ZN(
        n10887) );
  OR2_X1 U13808 ( .A1(n10888), .A2(n10887), .ZN(n13728) );
  NOR2_X1 U13809 ( .A1(n13728), .A2(n10869), .ZN(n10889) );
  NAND2_X1 U13810 ( .A1(n10889), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15861) );
  INV_X1 U13811 ( .A(n10889), .ZN(n10890) );
  NAND2_X1 U13812 ( .A1(n10890), .A2(n16137), .ZN(n15860) );
  INV_X1 U13813 ( .A(n10891), .ZN(n10892) );
  NOR2_X1 U13814 ( .A1(n10893), .A2(n10892), .ZN(n10894) );
  OR2_X1 U13815 ( .A1(n10925), .A2(n10894), .ZN(n19252) );
  NOR2_X1 U13816 ( .A1(n19252), .A2(n10869), .ZN(n16122) );
  NAND2_X1 U13817 ( .A1(n10812), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10895) );
  MUX2_X1 U13818 ( .A(n10895), .B(n10812), .S(n10913), .Z(n10896) );
  INV_X1 U13819 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n14066) );
  NAND2_X1 U13820 ( .A1(n10913), .A2(n14066), .ZN(n10898) );
  NAND2_X1 U13821 ( .A1(n19201), .A2(n14277), .ZN(n10897) );
  INV_X1 U13822 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16040) );
  NAND2_X1 U13823 ( .A1(n10897), .A2(n16040), .ZN(n16028) );
  NAND3_X1 U13824 ( .A1(n10898), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n10812), 
        .ZN(n10899) );
  NAND2_X1 U13825 ( .A1(n10899), .A2(n10901), .ZN(n19188) );
  INV_X1 U13826 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10900) );
  NAND2_X1 U13827 ( .A1(n10941), .A2(n10900), .ZN(n15802) );
  AND2_X1 U13828 ( .A1(n16028), .A2(n15802), .ZN(n15787) );
  INV_X1 U13829 ( .A(n10930), .ZN(n10904) );
  NAND2_X1 U13830 ( .A1(n10812), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10902) );
  MUX2_X1 U13831 ( .A(n10812), .B(n10902), .S(n10901), .Z(n10903) );
  NAND2_X1 U13832 ( .A1(n10904), .A2(n10903), .ZN(n19178) );
  OAI21_X1 U13833 ( .B1(n19178), .B2(n10869), .A(n16010), .ZN(n15790) );
  AND2_X1 U13834 ( .A1(n15787), .A2(n15790), .ZN(n15773) );
  AND2_X1 U13835 ( .A1(n10812), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10906) );
  INV_X1 U13836 ( .A(n10967), .ZN(n10905) );
  AOI21_X1 U13837 ( .B1(n10920), .B2(n10906), .A(n10905), .ZN(n10908) );
  AND2_X1 U13838 ( .A1(n10908), .A2(n10907), .ZN(n15497) );
  NAND2_X1 U13839 ( .A1(n15497), .A2(n14277), .ZN(n10909) );
  XNOR2_X1 U13840 ( .A(n10909), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15824) );
  NOR2_X1 U13841 ( .A1(n10911), .A2(n10910), .ZN(n10912) );
  OR2_X1 U13842 ( .A1(n10913), .A2(n10912), .ZN(n19219) );
  INV_X1 U13843 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16033) );
  OAI21_X1 U13844 ( .B1(n19219), .B2(n10869), .A(n16033), .ZN(n15812) );
  NAND2_X1 U13845 ( .A1(n10812), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10914) );
  MUX2_X1 U13846 ( .A(n10914), .B(n10812), .S(n10916), .Z(n10917) );
  INV_X1 U13847 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10915) );
  NAND2_X1 U13848 ( .A1(n10916), .A2(n10915), .ZN(n10919) );
  AOI21_X1 U13849 ( .B1(n19227), .B2(n14277), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16084) );
  AND2_X1 U13850 ( .A1(n10812), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10918) );
  NAND2_X1 U13851 ( .A1(n10919), .A2(n10918), .ZN(n10921) );
  NAND2_X1 U13852 ( .A1(n10921), .A2(n10920), .ZN(n12815) );
  OR2_X1 U13853 ( .A1(n12815), .A2(n10869), .ZN(n10922) );
  INV_X1 U13854 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16076) );
  NAND2_X1 U13855 ( .A1(n10922), .A2(n16076), .ZN(n15835) );
  INV_X1 U13856 ( .A(n10923), .ZN(n10924) );
  XNOR2_X1 U13857 ( .A(n10925), .B(n10924), .ZN(n19239) );
  NAND2_X1 U13858 ( .A1(n19239), .A2(n14277), .ZN(n10926) );
  INV_X1 U13859 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15853) );
  NAND2_X1 U13860 ( .A1(n10926), .A2(n15853), .ZN(n15847) );
  OAI211_X1 U13861 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16122), .A(
        n15835), .B(n15847), .ZN(n10927) );
  NOR2_X1 U13862 ( .A1(n16084), .A2(n10927), .ZN(n10928) );
  AND2_X1 U13863 ( .A1(n15812), .A2(n10928), .ZN(n10933) );
  NAND2_X1 U13864 ( .A1(n10812), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10929) );
  NOR2_X1 U13865 ( .A1(n10930), .A2(n10929), .ZN(n10931) );
  NAND2_X1 U13866 ( .A1(n10934), .A2(n9760), .ZN(n10950) );
  NAND2_X1 U13867 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10935) );
  OR2_X1 U13868 ( .A1(n19161), .A2(n10935), .ZN(n15774) );
  INV_X1 U13869 ( .A(n19219), .ZN(n10937) );
  AND2_X1 U13870 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10936) );
  NAND2_X1 U13871 ( .A1(n10937), .A2(n10936), .ZN(n15811) );
  AND2_X1 U13872 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10938) );
  NAND2_X1 U13873 ( .A1(n15497), .A2(n10938), .ZN(n15813) );
  AND2_X1 U13874 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10939) );
  NAND2_X1 U13875 ( .A1(n19227), .A2(n10939), .ZN(n16082) );
  OR3_X1 U13876 ( .A1(n12815), .A2(n10869), .A3(n16076), .ZN(n15834) );
  AND2_X1 U13877 ( .A1(n16082), .A2(n15834), .ZN(n15769) );
  AND2_X1 U13878 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10940) );
  NAND2_X1 U13879 ( .A1(n19239), .A2(n10940), .ZN(n15846) );
  NAND4_X1 U13880 ( .A1(n15774), .A2(n15771), .A3(n15769), .A4(n15846), .ZN(
        n10948) );
  INV_X1 U13881 ( .A(n10941), .ZN(n10942) );
  NAND2_X1 U13882 ( .A1(n10942), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15803) );
  AND2_X1 U13883 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10943) );
  NAND2_X1 U13884 ( .A1(n19201), .A2(n10943), .ZN(n16027) );
  NAND2_X1 U13885 ( .A1(n15803), .A2(n16027), .ZN(n15772) );
  INV_X1 U13886 ( .A(n15772), .ZN(n10946) );
  NAND2_X1 U13887 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10944) );
  NOR2_X1 U13888 ( .A1(n19178), .A2(n10944), .ZN(n15789) );
  NAND2_X1 U13889 ( .A1(n10946), .A2(n10945), .ZN(n10947) );
  NAND3_X1 U13890 ( .A1(n10951), .A2(n10812), .A3(P2_EBX_REG_22__SCAN_IN), 
        .ZN(n10952) );
  NAND2_X1 U13891 ( .A1(n10956), .A2(n10952), .ZN(n15487) );
  NAND2_X1 U13892 ( .A1(n10953), .A2(n15977), .ZN(n15973) );
  INV_X1 U13893 ( .A(n10954), .ZN(n10955) );
  XNOR2_X1 U13894 ( .A(n10956), .B(n10955), .ZN(n15465) );
  NAND2_X1 U13895 ( .A1(n15465), .A2(n14277), .ZN(n10957) );
  XNOR2_X1 U13896 ( .A(n10957), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15757) );
  INV_X1 U13897 ( .A(n10957), .ZN(n10958) );
  NAND2_X1 U13898 ( .A1(n10812), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10961) );
  MUX2_X1 U13899 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n10961), .S(n10960), .Z(
        n10962) );
  NAND2_X1 U13900 ( .A1(n10962), .A2(n10967), .ZN(n16465) );
  NOR2_X1 U13901 ( .A1(n16465), .A2(n10869), .ZN(n15743) );
  INV_X1 U13902 ( .A(n15743), .ZN(n10963) );
  INV_X1 U13903 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15947) );
  NOR2_X1 U13904 ( .A1(n10969), .A2(n15553), .ZN(n10965) );
  NAND2_X1 U13905 ( .A1(n10812), .A2(n10965), .ZN(n10966) );
  NAND2_X1 U13906 ( .A1(n10967), .A2(n10966), .ZN(n10968) );
  AOI21_X1 U13907 ( .B1(n10969), .B2(n15553), .A(n10968), .ZN(n15463) );
  AND2_X1 U13908 ( .A1(n15463), .A2(n14277), .ZN(n10983) );
  OR2_X1 U13909 ( .A1(n10983), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15732) );
  INV_X1 U13910 ( .A(n10970), .ZN(n14276) );
  NAND3_X1 U13911 ( .A1(n10812), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n10971), 
        .ZN(n10972) );
  NAND2_X1 U13912 ( .A1(n14276), .A2(n10972), .ZN(n16453) );
  OAI21_X1 U13913 ( .B1(n16453), .B2(n10869), .A(n15922), .ZN(n10974) );
  NAND2_X1 U13914 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10973) );
  NAND2_X1 U13915 ( .A1(n10974), .A2(n10985), .ZN(n15727) );
  INV_X1 U13916 ( .A(n10975), .ZN(n10976) );
  NAND2_X1 U13917 ( .A1(n10976), .A2(n9732), .ZN(n10977) );
  NAND2_X1 U13918 ( .A1(n10979), .A2(n10977), .ZN(n12827) );
  AND2_X1 U13919 ( .A1(n10979), .A2(n10978), .ZN(n10980) );
  NOR2_X1 U13920 ( .A1(n12519), .A2(n10980), .ZN(n15450) );
  OAI21_X1 U13921 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n15702), .ZN(n10981) );
  INV_X1 U13922 ( .A(n15702), .ZN(n10982) );
  INV_X1 U13923 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14612) );
  NAND2_X1 U13924 ( .A1(n10982), .A2(n14612), .ZN(n10986) );
  INV_X1 U13925 ( .A(n10983), .ZN(n10984) );
  INV_X1 U13926 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15937) );
  NAND2_X1 U13927 ( .A1(n15731), .A2(n10985), .ZN(n15699) );
  AOI21_X1 U13928 ( .B1(n10987), .B2(n10986), .A(n15699), .ZN(n10988) );
  INV_X1 U13929 ( .A(n10988), .ZN(n14271) );
  XOR2_X1 U13930 ( .A(n10989), .B(n14271), .Z(n14623) );
  NAND2_X1 U13931 ( .A1(n10993), .A2(n10992), .ZN(P2_U2985) );
  NAND2_X1 U13932 ( .A1(n11780), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11000) );
  AND2_X2 U13933 ( .A1(n13574), .A2(n10995), .ZN(n11214) );
  AOI22_X1 U13934 ( .A1(n9678), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11214), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10999) );
  NAND2_X1 U13935 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10998) );
  NAND2_X1 U13936 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10997) );
  NAND4_X1 U13937 ( .A1(n11000), .A2(n10999), .A3(n10998), .A4(n10997), .ZN(
        n11005) );
  NOR2_X4 U13938 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11010) );
  AND2_X2 U13939 ( .A1(n11007), .A2(n11010), .ZN(n11221) );
  NAND2_X1 U13940 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11002) );
  AND2_X2 U13941 ( .A1(n10996), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11009) );
  AND2_X2 U13942 ( .A1(n11007), .A2(n11009), .ZN(n11069) );
  NAND2_X1 U13943 ( .A1(n11069), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11001) );
  AOI22_X1 U13944 ( .A1(n9662), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9672), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11014) );
  AND2_X2 U13945 ( .A1(n13569), .A2(n11008), .ZN(n11062) );
  AOI22_X1 U13946 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11062), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11013) );
  AND2_X2 U13947 ( .A1(n11009), .A2(n13569), .ZN(n11148) );
  NAND2_X1 U13948 ( .A1(n13569), .A2(n11010), .ZN(n11123) );
  AOI22_X1 U13949 ( .A1(n9699), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9666), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11012) );
  AND2_X2 U13950 ( .A1(n11010), .A2(n13570), .ZN(n11118) );
  AOI22_X1 U13951 ( .A1(n9693), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11118), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U13952 ( .A1(n9678), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11214), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11020) );
  NAND2_X1 U13953 ( .A1(n11780), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11019) );
  NAND2_X1 U13954 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11018) );
  NAND2_X1 U13955 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11017) );
  NAND2_X1 U13956 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11024) );
  NAND2_X1 U13957 ( .A1(n11069), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11023) );
  NAND2_X1 U13958 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11022) );
  NAND2_X1 U13959 ( .A1(n9662), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11021) );
  NAND2_X1 U13960 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11028) );
  NAND2_X1 U13961 ( .A1(n11061), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11027) );
  NAND2_X1 U13962 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11026) );
  NAND2_X1 U13963 ( .A1(n9700), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11025) );
  INV_X1 U13964 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11031) );
  NAND2_X1 U13965 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11030) );
  NAND2_X1 U13966 ( .A1(n9699), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11029) );
  OAI211_X1 U13967 ( .C1(n9694), .C2(n11031), .A(n11030), .B(n11029), .ZN(
        n11032) );
  INV_X1 U13968 ( .A(n9731), .ZN(n13030) );
  AOI22_X1 U13969 ( .A1(n11069), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U13970 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U13971 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9654), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U13972 ( .A1(n11061), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9700), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U13973 ( .A1(n9678), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11214), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11044) );
  NAND2_X1 U13974 ( .A1(n11780), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11043) );
  NAND2_X1 U13975 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11042) );
  NAND2_X1 U13976 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11041) );
  NAND4_X1 U13977 ( .A1(n11044), .A2(n11043), .A3(n11042), .A4(n11041), .ZN(
        n11049) );
  INV_X1 U13978 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U13979 ( .A1(n9678), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11214), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11055) );
  NAND2_X1 U13980 ( .A1(n11780), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11054) );
  NAND2_X1 U13981 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11053) );
  NAND2_X1 U13982 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11052) );
  NAND4_X1 U13983 ( .A1(n11055), .A2(n11054), .A3(n11053), .A4(n11052), .ZN(
        n11060) );
  INV_X1 U13984 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11058) );
  NAND2_X1 U13985 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11057) );
  NAND2_X1 U13986 ( .A1(n11148), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11056) );
  OAI211_X1 U13987 ( .C1(n9694), .C2(n11058), .A(n11057), .B(n11056), .ZN(
        n11059) );
  NOR2_X1 U13988 ( .A1(n11060), .A2(n11059), .ZN(n11068) );
  AOI22_X1 U13989 ( .A1(n11069), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11220), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U13990 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U13991 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9654), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U13992 ( .A1(n11061), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9700), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11063) );
  NAND2_X1 U13993 ( .A1(n11069), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11073) );
  NAND2_X1 U13994 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11072) );
  NAND2_X1 U13995 ( .A1(n11061), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11071) );
  NAND2_X1 U13996 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11070) );
  NAND2_X1 U13997 ( .A1(n9662), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11077) );
  NAND2_X1 U13998 ( .A1(n9699), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11076) );
  NAND2_X1 U13999 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11075) );
  NAND2_X1 U14000 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11074) );
  AOI22_X1 U14001 ( .A1(n9677), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11214), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11082) );
  NAND2_X1 U14002 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11081) );
  NAND2_X1 U14003 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11080) );
  NAND2_X1 U14004 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11079) );
  AND4_X2 U14005 ( .A1(n11082), .A2(n11081), .A3(n11080), .A4(n11079), .ZN(
        n11089) );
  INV_X1 U14006 ( .A(n11780), .ZN(n11086) );
  INV_X1 U14007 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11085) );
  NAND2_X1 U14008 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11084) );
  NAND2_X1 U14009 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11083) );
  OAI211_X1 U14010 ( .C1(n11086), .C2(n11085), .A(n11084), .B(n11083), .ZN(
        n11087) );
  INV_X1 U14011 ( .A(n11087), .ZN(n11088) );
  NAND2_X1 U14012 ( .A1(n13642), .A2(n12155), .ZN(n11092) );
  INV_X1 U14013 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11747) );
  NAND2_X1 U14014 ( .A1(n11148), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11095) );
  NAND2_X1 U14015 ( .A1(n9693), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11094) );
  OAI211_X1 U14016 ( .C1(n9694), .C2(n11747), .A(n11095), .B(n11094), .ZN(
        n11096) );
  INV_X1 U14017 ( .A(n11096), .ZN(n11112) );
  NAND2_X1 U14018 ( .A1(n11069), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11100) );
  NAND2_X1 U14019 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11099) );
  NAND2_X1 U14020 ( .A1(n9662), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11098) );
  NAND2_X1 U14021 ( .A1(n11062), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11097) );
  NAND2_X1 U14022 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11104) );
  NAND2_X1 U14023 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11103) );
  NAND2_X1 U14024 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11102) );
  NAND2_X1 U14025 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11101) );
  NAND2_X1 U14026 ( .A1(n11780), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11108) );
  AOI22_X1 U14027 ( .A1(n9678), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11214), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11107) );
  NAND2_X1 U14028 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11106) );
  NAND2_X1 U14029 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11105) );
  NAND2_X1 U14030 ( .A1(n9662), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11117) );
  NAND2_X1 U14031 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11116) );
  NAND2_X1 U14032 ( .A1(n9677), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11115) );
  NAND2_X1 U14033 ( .A1(n11214), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11114) );
  AND4_X1 U14034 ( .A1(n11117), .A2(n11116), .A3(n11115), .A4(n11114), .ZN(
        n11122) );
  AOI22_X1 U14035 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11118), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11121) );
  NAND2_X1 U14036 ( .A1(n11780), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11120) );
  NAND2_X1 U14037 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11119) );
  AOI22_X1 U14038 ( .A1(n11148), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11127) );
  AOI22_X1 U14039 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9700), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11126) );
  AOI22_X1 U14040 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9693), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11125) );
  AOI22_X1 U14041 ( .A1(n11069), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11124) );
  NAND2_X1 U14042 ( .A1(n11169), .A2(n13303), .ZN(n11131) );
  NAND2_X1 U14043 ( .A1(n12155), .A2(n11165), .ZN(n13293) );
  AND3_X2 U14044 ( .A1(n11132), .A2(n11131), .A3(n9747), .ZN(n11163) );
  NAND2_X1 U14045 ( .A1(n20438), .A2(n13303), .ZN(n12146) );
  INV_X2 U14046 ( .A(n13642), .ZN(n20450) );
  INV_X1 U14047 ( .A(n12149), .ZN(n11135) );
  AOI22_X1 U14048 ( .A1(n9678), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11214), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11139) );
  NAND2_X1 U14049 ( .A1(n11780), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11138) );
  NAND2_X1 U14050 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11137) );
  NAND2_X1 U14051 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11136) );
  NAND2_X1 U14052 ( .A1(n11069), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11143) );
  NAND2_X1 U14053 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11142) );
  NAND2_X1 U14054 ( .A1(n9654), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11141) );
  NAND2_X1 U14055 ( .A1(n11941), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11140) );
  NAND2_X1 U14056 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11147) );
  NAND2_X1 U14057 ( .A1(n11220), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11146) );
  NAND2_X1 U14058 ( .A1(n9662), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11145) );
  NAND2_X1 U14059 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11144) );
  INV_X1 U14060 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11151) );
  NAND2_X1 U14061 ( .A1(n11148), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11150) );
  NAND2_X1 U14062 ( .A1(n11061), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11149) );
  OAI211_X1 U14063 ( .C1(n9694), .C2(n11151), .A(n11150), .B(n11149), .ZN(
        n11152) );
  INV_X1 U14064 ( .A(n11152), .ZN(n11153) );
  NAND4_X4 U14065 ( .A1(n11156), .A2(n11155), .A3(n11154), .A4(n11153), .ZN(
        n13637) );
  NAND2_X1 U14066 ( .A1(n11170), .A2(n13637), .ZN(n13852) );
  NAND2_X1 U14067 ( .A1(n14094), .A2(n13852), .ZN(n13029) );
  INV_X1 U14068 ( .A(n13029), .ZN(n11157) );
  XNOR2_X1 U14069 ( .A(n16263), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n12120) );
  INV_X1 U14070 ( .A(n12120), .ZN(n11158) );
  AND2_X2 U14071 ( .A1(n11968), .A2(n11170), .ZN(n13209) );
  INV_X1 U14072 ( .A(n13293), .ZN(n11301) );
  INV_X1 U14073 ( .A(n13322), .ZN(n11159) );
  NOR2_X1 U14074 ( .A1(n11160), .A2(n11159), .ZN(n11161) );
  NAND2_X1 U14075 ( .A1(n13299), .A2(n11161), .ZN(n11162) );
  INV_X1 U14076 ( .A(n11163), .ZN(n13210) );
  NAND2_X1 U14077 ( .A1(n13210), .A2(n11170), .ZN(n11175) );
  NAND2_X1 U14078 ( .A1(n13248), .A2(n20446), .ZN(n11167) );
  NAND2_X1 U14079 ( .A1(n20450), .A2(n12155), .ZN(n11166) );
  AND2_X1 U14080 ( .A1(n11166), .A2(n11165), .ZN(n11186) );
  NAND2_X1 U14081 ( .A1(n13193), .A2(n15412), .ZN(n11174) );
  NAND2_X1 U14082 ( .A1(n9731), .A2(n13202), .ZN(n13311) );
  OR2_X1 U14083 ( .A1(n11170), .A2(n20438), .ZN(n13203) );
  AND2_X1 U14084 ( .A1(n13203), .A2(n13852), .ZN(n11171) );
  OAI211_X1 U14085 ( .C1(n14094), .C2(n20446), .A(n13311), .B(n11171), .ZN(
        n11191) );
  NOR2_X1 U14086 ( .A1(n11191), .A2(n11172), .ZN(n11173) );
  NAND2_X1 U14087 ( .A1(n11197), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11179) );
  NAND2_X1 U14088 ( .A1(n16419), .A2(n20963), .ZN(n13333) );
  NAND2_X1 U14089 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11200) );
  OAI21_X1 U14090 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11200), .ZN(n20725) );
  OR2_X1 U14091 ( .A1(n16243), .A2(n20722), .ZN(n11195) );
  OAI21_X1 U14092 ( .B1(n13333), .B2(n20725), .A(n11195), .ZN(n11177) );
  INV_X1 U14093 ( .A(n11177), .ZN(n11178) );
  NAND2_X1 U14094 ( .A1(n11179), .A2(n11178), .ZN(n11181) );
  XNOR2_X1 U14095 ( .A(n11181), .B(n11180), .ZN(n11287) );
  MUX2_X1 U14096 ( .A(n13333), .B(n16243), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11182) );
  INV_X1 U14097 ( .A(n13209), .ZN(n13853) );
  INV_X1 U14098 ( .A(n13248), .ZN(n11184) );
  NAND3_X1 U14099 ( .A1(n13853), .A2(n11184), .A3(n13303), .ZN(n11185) );
  NAND2_X1 U14100 ( .A1(n13210), .A2(n11185), .ZN(n11194) );
  INV_X1 U14101 ( .A(n11186), .ZN(n11187) );
  NAND2_X1 U14102 ( .A1(n16235), .A2(n11187), .ZN(n11189) );
  NAND2_X1 U14103 ( .A1(n11172), .A2(n10038), .ZN(n11188) );
  NAND4_X1 U14104 ( .A1(n11189), .A2(n16419), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .A4(n11188), .ZN(n11190) );
  NOR2_X1 U14105 ( .A1(n11191), .A2(n11190), .ZN(n11193) );
  NAND3_X1 U14106 ( .A1(n13193), .A2(n15412), .A3(n13637), .ZN(n11192) );
  NAND3_X1 U14107 ( .A1(n11194), .A2(n11193), .A3(n11192), .ZN(n11231) );
  AND2_X1 U14108 ( .A1(n11195), .A2(n10996), .ZN(n11196) );
  NAND2_X1 U14109 ( .A1(n11290), .A2(n11206), .ZN(n11204) );
  NOR2_X1 U14110 ( .A1(n16243), .A2(n20787), .ZN(n11198) );
  INV_X1 U14111 ( .A(n13333), .ZN(n11202) );
  INV_X1 U14112 ( .A(n11200), .ZN(n11199) );
  NAND2_X1 U14113 ( .A1(n11199), .A2(n20787), .ZN(n20753) );
  NAND2_X1 U14114 ( .A1(n11200), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11201) );
  NAND2_X1 U14115 ( .A1(n20753), .A2(n11201), .ZN(n20430) );
  NAND2_X1 U14116 ( .A1(n11202), .A2(n20430), .ZN(n11205) );
  NAND2_X1 U14117 ( .A1(n11207), .A2(n11205), .ZN(n11203) );
  NAND4_X1 U14118 ( .A1(n11290), .A2(n11207), .A3(n11206), .A4(n11205), .ZN(
        n11208) );
  INV_X1 U14119 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11211) );
  NAND2_X1 U14120 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11210) );
  NAND2_X1 U14121 ( .A1(n11148), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11209) );
  OAI211_X1 U14122 ( .C1(n11934), .C2(n11211), .A(n11210), .B(n11209), .ZN(
        n11212) );
  INV_X1 U14123 ( .A(n11212), .ZN(n11219) );
  INV_X1 U14124 ( .A(n11214), .ZN(n11880) );
  INV_X1 U14125 ( .A(n11880), .ZN(n11339) );
  AOI22_X1 U14126 ( .A1(n9678), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11218) );
  AOI22_X1 U14127 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11217) );
  NAND2_X1 U14128 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11216) );
  NAND4_X1 U14129 ( .A1(n11219), .A2(n11218), .A3(n11217), .A4(n11216), .ZN(
        n11227) );
  AOI22_X1 U14130 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11225) );
  INV_X1 U14131 ( .A(n11221), .ZN(n11882) );
  AOI22_X1 U14132 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11224) );
  AOI22_X1 U14133 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14134 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11222) );
  NAND4_X1 U14135 ( .A1(n11225), .A2(n11224), .A3(n11223), .A4(n11222), .ZN(
        n11226) );
  INV_X1 U14136 ( .A(n11999), .ZN(n11995) );
  INV_X1 U14137 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11228) );
  OAI22_X1 U14138 ( .A1(n11995), .A2(n11228), .B1(n13669), .B2(n11335), .ZN(
        n11229) );
  XNOR2_X1 U14139 ( .A(n11230), .B(n11229), .ZN(n11298) );
  INV_X1 U14140 ( .A(n11231), .ZN(n11232) );
  INV_X1 U14141 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n21070) );
  NAND2_X1 U14142 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11234) );
  NAND2_X1 U14143 ( .A1(n11148), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11233) );
  OAI211_X1 U14144 ( .C1(n11934), .C2(n21070), .A(n11234), .B(n11233), .ZN(
        n11235) );
  INV_X1 U14145 ( .A(n11235), .ZN(n11240) );
  AOI22_X1 U14146 ( .A1(n9678), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11239) );
  AOI22_X1 U14147 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11238) );
  NAND2_X1 U14148 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11237) );
  NAND4_X1 U14149 ( .A1(n11240), .A2(n11239), .A3(n11238), .A4(n11237), .ZN(
        n11246) );
  AOI22_X1 U14150 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14151 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14152 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9654), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U14153 ( .A1(n9693), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11241) );
  NAND4_X1 U14154 ( .A1(n11244), .A2(n11243), .A3(n11242), .A4(n11241), .ZN(
        n11245) );
  NAND2_X1 U14155 ( .A1(n20446), .A2(n14010), .ZN(n11267) );
  INV_X1 U14156 ( .A(n14010), .ZN(n14095) );
  NAND2_X1 U14157 ( .A1(n14095), .A2(n20446), .ZN(n11260) );
  INV_X1 U14158 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11760) );
  NAND2_X1 U14159 ( .A1(n11148), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11248) );
  NAND2_X1 U14160 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11247) );
  OAI211_X1 U14161 ( .C1(n11934), .C2(n11760), .A(n11248), .B(n11247), .ZN(
        n11249) );
  INV_X1 U14162 ( .A(n11249), .ZN(n11253) );
  AOI22_X1 U14163 ( .A1(n9677), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11214), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11252) );
  AOI22_X1 U14164 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11251) );
  NAND2_X1 U14165 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11250) );
  NAND4_X1 U14166 ( .A1(n11253), .A2(n11252), .A3(n11251), .A4(n11250), .ZN(
        n11259) );
  AOI22_X1 U14167 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14168 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14169 ( .A1(n11061), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U14170 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11254) );
  NAND4_X1 U14171 ( .A1(n11257), .A2(n11256), .A3(n11255), .A4(n11254), .ZN(
        n11258) );
  MUX2_X1 U14172 ( .A(n11267), .B(n11260), .S(n13641), .Z(n11261) );
  INV_X1 U14173 ( .A(n11261), .ZN(n11262) );
  NAND2_X1 U14174 ( .A1(n11262), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11315) );
  NAND2_X1 U14175 ( .A1(n11313), .A2(n11315), .ZN(n11266) );
  NAND2_X1 U14176 ( .A1(n11999), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11265) );
  OAI21_X1 U14177 ( .B1(n20963), .B2(n13641), .A(n11970), .ZN(n11263) );
  AND2_X1 U14178 ( .A1(n11263), .A2(n11267), .ZN(n11264) );
  NAND2_X1 U14179 ( .A1(n11265), .A2(n11264), .ZN(n11317) );
  NAND2_X1 U14180 ( .A1(n11266), .A2(n11317), .ZN(n11269) );
  INV_X1 U14181 ( .A(n11267), .ZN(n11268) );
  NAND2_X1 U14182 ( .A1(n11268), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14091) );
  NAND2_X1 U14183 ( .A1(n11999), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11286) );
  AOI22_X1 U14184 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14185 ( .A1(n11221), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14186 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14187 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11271) );
  AND4_X1 U14188 ( .A1(n11274), .A2(n11273), .A3(n11272), .A4(n11271), .ZN(
        n11283) );
  AOI22_X1 U14189 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11148), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11282) );
  NAND2_X1 U14190 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11278) );
  NAND2_X1 U14191 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11277) );
  NAND2_X1 U14192 ( .A1(n9678), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U14193 ( .A1(n11214), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11275) );
  AND4_X1 U14194 ( .A1(n11278), .A2(n11277), .A3(n11276), .A4(n11275), .ZN(
        n11281) );
  NAND2_X1 U14195 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11280) );
  NAND2_X1 U14196 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11279) );
  OAI22_X1 U14197 ( .A1(n13639), .A2(n11335), .B1(n11334), .B2(n14010), .ZN(
        n11284) );
  INV_X1 U14198 ( .A(n11284), .ZN(n11285) );
  INV_X1 U14199 ( .A(n11287), .ZN(n20522) );
  INV_X1 U14200 ( .A(n11288), .ZN(n11289) );
  NAND2_X1 U14201 ( .A1(n20467), .A2(n11290), .ZN(n13937) );
  OR2_X1 U14202 ( .A1(n11334), .A2(n13639), .ZN(n11291) );
  INV_X1 U14203 ( .A(n11292), .ZN(n13638) );
  NAND2_X1 U14204 ( .A1(n11307), .A2(n13638), .ZN(n11297) );
  INV_X1 U14205 ( .A(n11293), .ZN(n11294) );
  NAND2_X1 U14206 ( .A1(n11298), .A2(n11299), .ZN(n11300) );
  NAND2_X1 U14207 ( .A1(n10038), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11503) );
  NAND2_X1 U14208 ( .A1(n11301), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11362) );
  XNOR2_X1 U14209 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20337) );
  AOI21_X1 U14210 ( .B1(n11928), .B2(n20337), .A(n12142), .ZN(n11304) );
  NAND2_X1 U14211 ( .A1(n11359), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11303) );
  OAI211_X1 U14212 ( .C1(n11362), .C2(n11302), .A(n11304), .B(n11303), .ZN(
        n11305) );
  INV_X1 U14213 ( .A(n11305), .ZN(n11306) );
  NAND2_X1 U14214 ( .A1(n12142), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11327) );
  INV_X1 U14215 ( .A(n11307), .ZN(n11308) );
  NAND2_X1 U14216 ( .A1(n13630), .A2(n11590), .ZN(n11312) );
  AOI22_X1 U14217 ( .A1(n11359), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20966), .ZN(n11310) );
  INV_X1 U14218 ( .A(n11362), .ZN(n11381) );
  NAND2_X1 U14219 ( .A1(n11381), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11309) );
  AND2_X1 U14220 ( .A1(n11310), .A2(n11309), .ZN(n11311) );
  NAND2_X1 U14221 ( .A1(n11313), .A2(n11317), .ZN(n11314) );
  INV_X1 U14222 ( .A(n11315), .ZN(n11316) );
  NAND2_X1 U14223 ( .A1(n13302), .A2(n10038), .ZN(n11319) );
  NAND2_X1 U14224 ( .A1(n11319), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13252) );
  NAND2_X1 U14225 ( .A1(n11359), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11322) );
  NAND2_X1 U14226 ( .A1(n20966), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11321) );
  OAI211_X1 U14227 ( .C1(n11362), .C2(n16215), .A(n11322), .B(n11321), .ZN(
        n11323) );
  AOI21_X1 U14228 ( .B1(n11320), .B2(n11590), .A(n11323), .ZN(n11324) );
  OR2_X1 U14229 ( .A1(n13252), .A2(n11324), .ZN(n13253) );
  INV_X1 U14230 ( .A(n11324), .ZN(n13254) );
  OR2_X1 U14231 ( .A1(n13254), .A2(n10196), .ZN(n11325) );
  NAND2_X1 U14232 ( .A1(n13253), .A2(n11325), .ZN(n13102) );
  NAND2_X1 U14233 ( .A1(n11197), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11333) );
  NAND3_X1 U14234 ( .A1(n20786), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20638) );
  INV_X1 U14235 ( .A(n20638), .ZN(n11329) );
  NAND2_X1 U14236 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11329), .ZN(
        n20636) );
  NAND2_X1 U14237 ( .A1(n20786), .A2(n20636), .ZN(n11330) );
  NOR3_X1 U14238 ( .A1(n20786), .A2(n20787), .A3(n20722), .ZN(n20910) );
  NAND2_X1 U14239 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20910), .ZN(
        n20896) );
  NAND2_X1 U14240 ( .A1(n11330), .A2(n20896), .ZN(n20668) );
  OAI22_X1 U14241 ( .A1(n13333), .A2(n20668), .B1(n16243), .B2(n20786), .ZN(
        n11331) );
  INV_X1 U14242 ( .A(n11331), .ZN(n11332) );
  NAND2_X1 U14243 ( .A1(n20426), .A2(n20963), .ZN(n11351) );
  INV_X1 U14244 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11832) );
  NAND2_X1 U14245 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11337) );
  NAND2_X1 U14246 ( .A1(n11148), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11336) );
  OAI211_X1 U14247 ( .C1(n11934), .C2(n11832), .A(n11337), .B(n11336), .ZN(
        n11338) );
  INV_X1 U14248 ( .A(n11338), .ZN(n11343) );
  AOI22_X1 U14249 ( .A1(n9678), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14250 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11341) );
  NAND2_X1 U14251 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11340) );
  NAND4_X1 U14252 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(
        n11349) );
  AOI22_X1 U14253 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14254 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14255 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14256 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11344) );
  NAND4_X1 U14257 ( .A1(n11347), .A2(n11346), .A3(n11345), .A4(n11344), .ZN(
        n11348) );
  AOI22_X1 U14258 ( .A1(n11999), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11990), .B2(n13988), .ZN(n11350) );
  NAND2_X1 U14259 ( .A1(n11353), .A2(n13629), .ZN(n11354) );
  INV_X1 U14260 ( .A(n11356), .ZN(n11358) );
  INV_X1 U14261 ( .A(n11384), .ZN(n11357) );
  OAI21_X1 U14262 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11358), .A(
        n11357), .ZN(n13858) );
  AOI22_X1 U14263 ( .A1(n11928), .A2(n13858), .B1(n12142), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11361) );
  NAND2_X1 U14264 ( .A1(n12143), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11360) );
  OAI211_X1 U14265 ( .C1(n11362), .C2(n13581), .A(n11361), .B(n11360), .ZN(
        n11363) );
  INV_X1 U14266 ( .A(n11363), .ZN(n11364) );
  NAND2_X1 U14267 ( .A1(n13466), .A2(n13467), .ZN(n13446) );
  INV_X1 U14268 ( .A(n13446), .ZN(n11390) );
  NAND2_X1 U14269 ( .A1(n11999), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11380) );
  INV_X1 U14270 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11367) );
  NAND2_X1 U14271 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11366) );
  NAND2_X1 U14272 ( .A1(n11148), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11365) );
  OAI211_X1 U14273 ( .C1(n11934), .C2(n11367), .A(n11366), .B(n11365), .ZN(
        n11368) );
  INV_X1 U14274 ( .A(n11368), .ZN(n11372) );
  AOI22_X1 U14275 ( .A1(n9678), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14276 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11370) );
  NAND2_X1 U14277 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11369) );
  NAND4_X1 U14278 ( .A1(n11372), .A2(n11371), .A3(n11370), .A4(n11369), .ZN(
        n11378) );
  AOI22_X1 U14279 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n9690), .B1(
        n11270), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14280 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14281 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14282 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11373) );
  NAND4_X1 U14283 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n11373), .ZN(
        n11377) );
  NAND2_X1 U14284 ( .A1(n11990), .A2(n13987), .ZN(n11379) );
  NAND2_X1 U14285 ( .A1(n11380), .A2(n11379), .ZN(n11392) );
  XNOR2_X1 U14286 ( .A(n11391), .B(n11392), .ZN(n13979) );
  NAND2_X1 U14287 ( .A1(n11381), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11387) );
  INV_X1 U14288 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11382) );
  AOI21_X1 U14289 ( .B1(n11382), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11383) );
  AOI21_X1 U14290 ( .B1(n12143), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11383), .ZN(
        n11386) );
  OAI21_X1 U14291 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11384), .A(
        n11409), .ZN(n20367) );
  NOR2_X1 U14292 ( .A1(n20367), .A2(n10196), .ZN(n11385) );
  AOI21_X1 U14293 ( .B1(n11387), .B2(n11386), .A(n11385), .ZN(n11388) );
  AOI21_X1 U14294 ( .B1(n13979), .B2(n11590), .A(n11388), .ZN(n13445) );
  NAND2_X1 U14295 ( .A1(n11390), .A2(n11389), .ZN(n13444) );
  NAND2_X1 U14296 ( .A1(n11393), .A2(n11392), .ZN(n11415) );
  NAND2_X1 U14297 ( .A1(n11999), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11408) );
  INV_X1 U14298 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11883) );
  NAND2_X1 U14299 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11395) );
  NAND2_X1 U14300 ( .A1(n11148), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11394) );
  OAI211_X1 U14301 ( .C1(n11934), .C2(n11883), .A(n11395), .B(n11394), .ZN(
        n11396) );
  INV_X1 U14302 ( .A(n11396), .ZN(n11400) );
  AOI22_X1 U14303 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14304 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11398) );
  NAND2_X1 U14305 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11397) );
  NAND4_X1 U14306 ( .A1(n11400), .A2(n11399), .A3(n11398), .A4(n11397), .ZN(
        n11406) );
  AOI22_X1 U14307 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14308 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U14309 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14310 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11401) );
  NAND4_X1 U14311 ( .A1(n11404), .A2(n11403), .A3(n11402), .A4(n11401), .ZN(
        n11405) );
  NAND2_X1 U14312 ( .A1(n11990), .A2(n13997), .ZN(n11407) );
  NAND2_X1 U14313 ( .A1(n11408), .A2(n11407), .ZN(n11416) );
  XNOR2_X1 U14314 ( .A(n11415), .B(n11416), .ZN(n13986) );
  INV_X1 U14315 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13707) );
  OAI21_X1 U14316 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11410), .A(
        n11431), .ZN(n20331) );
  AOI22_X1 U14317 ( .A1(n11928), .A2(n20331), .B1(n12142), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11411) );
  OAI21_X1 U14318 ( .B1(n11902), .B2(n13707), .A(n11411), .ZN(n11412) );
  INV_X1 U14319 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11419) );
  NAND2_X1 U14320 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11418) );
  NAND2_X1 U14321 ( .A1(n11148), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11417) );
  OAI211_X1 U14322 ( .C1(n11934), .C2(n11419), .A(n11418), .B(n11417), .ZN(
        n11420) );
  INV_X1 U14323 ( .A(n11420), .ZN(n11424) );
  AOI22_X1 U14324 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14325 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11422) );
  NAND2_X1 U14326 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11421) );
  NAND4_X1 U14327 ( .A1(n11424), .A2(n11423), .A3(n11422), .A4(n11421), .ZN(
        n11430) );
  AOI22_X1 U14328 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14329 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14330 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14331 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11425) );
  NAND4_X1 U14332 ( .A1(n11428), .A2(n11427), .A3(n11426), .A4(n11425), .ZN(
        n11429) );
  AOI22_X1 U14333 ( .A1(n11999), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11990), .B2(n14008), .ZN(n11436) );
  NAND2_X1 U14334 ( .A1(n11435), .A2(n11436), .ZN(n13996) );
  INV_X1 U14335 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11433) );
  XNOR2_X1 U14336 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B(n11441), .ZN(
        n20319) );
  AOI22_X1 U14337 ( .A1(n11928), .A2(n20319), .B1(n12142), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11432) );
  OAI21_X1 U14338 ( .B1(n11902), .B2(n11433), .A(n11432), .ZN(n11434) );
  INV_X1 U14339 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11439) );
  NAND2_X1 U14340 ( .A1(n11990), .A2(n14010), .ZN(n11438) );
  OAI21_X1 U14341 ( .B1(n11995), .B2(n11439), .A(n11438), .ZN(n11440) );
  NAND2_X1 U14342 ( .A1(n14006), .A2(n11590), .ZN(n11450) );
  INV_X1 U14343 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13805) );
  INV_X1 U14344 ( .A(n11462), .ZN(n11446) );
  INV_X1 U14345 ( .A(n11442), .ZN(n11444) );
  INV_X1 U14346 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11443) );
  NAND2_X1 U14347 ( .A1(n11444), .A2(n11443), .ZN(n11445) );
  NAND2_X1 U14348 ( .A1(n11446), .A2(n11445), .ZN(n20307) );
  AOI22_X1 U14349 ( .A1(n20307), .A2(n11928), .B1(n12142), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11447) );
  INV_X1 U14350 ( .A(n11448), .ZN(n11449) );
  NAND2_X1 U14351 ( .A1(n11450), .A2(n11449), .ZN(n13803) );
  NAND2_X1 U14352 ( .A1(n13802), .A2(n13803), .ZN(n13801) );
  AOI22_X1 U14353 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14354 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9698), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14355 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14356 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11451) );
  AND4_X1 U14357 ( .A1(n11454), .A2(n11453), .A3(n11452), .A4(n11451), .ZN(
        n11461) );
  AOI22_X1 U14358 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9699), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14359 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11457) );
  AOI22_X1 U14360 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11456) );
  NAND2_X1 U14361 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11455) );
  AND3_X1 U14362 ( .A1(n11457), .A2(n11456), .A3(n11455), .ZN(n11459) );
  NAND2_X1 U14363 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11458) );
  NAND4_X1 U14364 ( .A1(n11461), .A2(n11460), .A3(n11459), .A4(n11458), .ZN(
        n11465) );
  NOR2_X1 U14365 ( .A1(n11462), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11463) );
  NOR2_X1 U14366 ( .A1(n11498), .A2(n11463), .ZN(n20289) );
  INV_X1 U14367 ( .A(n12142), .ZN(n13631) );
  INV_X1 U14368 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21209) );
  OAI22_X1 U14369 ( .A1(n20289), .A2(n10196), .B1(n13631), .B2(n21209), .ZN(
        n11464) );
  AOI21_X1 U14370 ( .B1(n11590), .B2(n11465), .A(n11464), .ZN(n11467) );
  NAND2_X1 U14371 ( .A1(n12143), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11466) );
  NAND2_X1 U14372 ( .A1(n12143), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14373 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14374 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14375 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14376 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11468) );
  AND4_X1 U14377 ( .A1(n11471), .A2(n11470), .A3(n11469), .A4(n11468), .ZN(
        n11478) );
  AOI22_X1 U14378 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11891), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14379 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14380 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11473) );
  NAND2_X1 U14381 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11472) );
  AND3_X1 U14382 ( .A1(n11474), .A2(n11473), .A3(n11472), .ZN(n11476) );
  NAND2_X1 U14383 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11475) );
  NAND4_X1 U14384 ( .A1(n11478), .A2(n11477), .A3(n11476), .A4(n11475), .ZN(
        n11479) );
  NAND2_X1 U14385 ( .A1(n11590), .A2(n11479), .ZN(n11482) );
  XOR2_X1 U14386 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11498), .Z(n20273) );
  INV_X1 U14387 ( .A(n20273), .ZN(n11480) );
  AOI22_X1 U14388 ( .A1(n12142), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n11928), .B2(n11480), .ZN(n11481) );
  INV_X1 U14389 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11486) );
  NAND2_X1 U14390 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11485) );
  NAND2_X1 U14391 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11484) );
  OAI211_X1 U14392 ( .C1(n11934), .C2(n11486), .A(n11485), .B(n11484), .ZN(
        n11487) );
  INV_X1 U14393 ( .A(n11487), .ZN(n11491) );
  AOI22_X1 U14394 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14395 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11489) );
  NAND2_X1 U14396 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11488) );
  NAND4_X1 U14397 ( .A1(n11491), .A2(n11490), .A3(n11489), .A4(n11488), .ZN(
        n11497) );
  AOI22_X1 U14398 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14399 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11494) );
  AOI22_X1 U14400 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14401 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11492) );
  NAND4_X1 U14402 ( .A1(n11495), .A2(n11494), .A3(n11493), .A4(n11492), .ZN(
        n11496) );
  NOR2_X1 U14403 ( .A1(n11497), .A2(n11496), .ZN(n11502) );
  NAND2_X1 U14404 ( .A1(n12143), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11501) );
  INV_X1 U14405 ( .A(n11504), .ZN(n11499) );
  XNOR2_X1 U14406 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B(n11499), .ZN(
        n14034) );
  AOI22_X1 U14407 ( .A1(n11928), .A2(n14034), .B1(n12142), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11500) );
  OAI211_X1 U14408 ( .C1(n11503), .C2(n11502), .A(n11501), .B(n11500), .ZN(
        n14028) );
  NAND2_X1 U14409 ( .A1(n12143), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11507) );
  OAI21_X1 U14410 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11505), .A(
        n11538), .ZN(n16331) );
  AOI22_X1 U14411 ( .A1(n11928), .A2(n16331), .B1(n12142), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11506) );
  NAND2_X1 U14412 ( .A1(n11507), .A2(n11506), .ZN(n14843) );
  AOI22_X1 U14413 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11891), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14414 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14415 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U14416 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11508) );
  AND4_X1 U14417 ( .A1(n11511), .A2(n11510), .A3(n11509), .A4(n11508), .ZN(
        n11519) );
  AOI22_X1 U14418 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11518) );
  NAND2_X1 U14419 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11515) );
  AOI22_X1 U14420 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11514) );
  NAND2_X1 U14421 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11513) );
  NAND2_X1 U14422 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11512) );
  AND4_X1 U14423 ( .A1(n11515), .A2(n11514), .A3(n11513), .A4(n11512), .ZN(
        n11517) );
  NAND2_X1 U14424 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11516) );
  NAND4_X1 U14425 ( .A1(n11519), .A2(n11518), .A3(n11517), .A4(n11516), .ZN(
        n11520) );
  AND2_X1 U14426 ( .A1(n11590), .A2(n11520), .ZN(n14891) );
  NAND2_X1 U14427 ( .A1(n14027), .A2(n14891), .ZN(n11521) );
  XOR2_X1 U14428 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11556), .Z(
        n15193) );
  INV_X1 U14429 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11884) );
  NAND2_X1 U14430 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11523) );
  NAND2_X1 U14431 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11522) );
  OAI211_X1 U14432 ( .C1(n11934), .C2(n11884), .A(n11523), .B(n11522), .ZN(
        n11524) );
  INV_X1 U14433 ( .A(n11524), .ZN(n11528) );
  AOI22_X1 U14434 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14435 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11526) );
  NAND2_X1 U14436 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11525) );
  NAND4_X1 U14437 ( .A1(n11528), .A2(n11527), .A3(n11526), .A4(n11525), .ZN(
        n11534) );
  AOI22_X1 U14438 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14439 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14440 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14441 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11529) );
  NAND4_X1 U14442 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(
        n11533) );
  OR2_X1 U14443 ( .A1(n11534), .A2(n11533), .ZN(n11535) );
  AOI22_X1 U14444 ( .A1(n11590), .A2(n11535), .B1(n12142), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11537) );
  NAND2_X1 U14445 ( .A1(n12143), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11536) );
  OAI211_X1 U14446 ( .C1(n15193), .C2(n10196), .A(n11537), .B(n11536), .ZN(
        n14846) );
  INV_X1 U14447 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14989) );
  XOR2_X1 U14448 ( .A(n16293), .B(n11538), .Z(n16320) );
  INV_X1 U14449 ( .A(n16320), .ZN(n11539) );
  AOI22_X1 U14450 ( .A1(n12142), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n11928), .B2(n11539), .ZN(n11553) );
  AOI22_X1 U14451 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14452 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11270), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14453 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9698), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14454 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n9690), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11540) );
  AND4_X1 U14455 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(
        n11550) );
  AOI22_X1 U14456 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11891), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14457 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14458 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11545) );
  NAND2_X1 U14459 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11544) );
  AND3_X1 U14460 ( .A1(n11546), .A2(n11545), .A3(n11544), .ZN(n11548) );
  NAND2_X1 U14461 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11547) );
  NAND4_X1 U14462 ( .A1(n11550), .A2(n11549), .A3(n11548), .A4(n11547), .ZN(
        n11551) );
  NAND2_X1 U14463 ( .A1(n11590), .A2(n11551), .ZN(n11552) );
  OAI211_X1 U14464 ( .C1(n11902), .C2(n14989), .A(n11553), .B(n11552), .ZN(
        n14981) );
  AND2_X1 U14465 ( .A1(n14846), .A2(n14981), .ZN(n11554) );
  NAND2_X1 U14466 ( .A1(n11557), .A2(n21218), .ZN(n11559) );
  INV_X1 U14467 ( .A(n11613), .ZN(n11558) );
  NAND2_X1 U14468 ( .A1(n11559), .A2(n11558), .ZN(n14835) );
  AOI22_X1 U14469 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11891), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14470 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14471 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14472 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11560) );
  NAND4_X1 U14473 ( .A1(n11563), .A2(n11562), .A3(n11561), .A4(n11560), .ZN(
        n11573) );
  INV_X1 U14474 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11566) );
  NAND2_X1 U14475 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11565) );
  NAND2_X1 U14476 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11564) );
  OAI211_X1 U14477 ( .C1(n11934), .C2(n11566), .A(n11565), .B(n11564), .ZN(
        n11567) );
  INV_X1 U14478 ( .A(n11567), .ZN(n11571) );
  AOI22_X1 U14479 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14480 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11569) );
  NAND2_X1 U14481 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11568) );
  NAND4_X1 U14482 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n11572) );
  OAI21_X1 U14483 ( .B1(n11573), .B2(n11572), .A(n11590), .ZN(n11576) );
  NAND2_X1 U14484 ( .A1(n12143), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11575) );
  NAND2_X1 U14485 ( .A1(n12142), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11574) );
  NAND3_X1 U14486 ( .A1(n11576), .A2(n11575), .A3(n11574), .ZN(n11577) );
  AOI21_X1 U14487 ( .B1(n14835), .B2(n11928), .A(n11577), .ZN(n14831) );
  NAND2_X1 U14488 ( .A1(n12143), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14489 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14490 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14491 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11891), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14492 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n9698), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11578) );
  AND4_X1 U14493 ( .A1(n11581), .A2(n11580), .A3(n11579), .A4(n11578), .ZN(
        n11588) );
  AOI22_X1 U14494 ( .A1(n11941), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U14495 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14496 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11583) );
  NAND2_X1 U14497 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11582) );
  AND3_X1 U14498 ( .A1(n11584), .A2(n11583), .A3(n11582), .ZN(n11586) );
  NAND2_X1 U14499 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11585) );
  NAND4_X1 U14500 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n11589) );
  NAND2_X1 U14501 ( .A1(n11590), .A2(n11589), .ZN(n11593) );
  XOR2_X1 U14502 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11613), .Z(
        n16315) );
  INV_X1 U14503 ( .A(n16315), .ZN(n11591) );
  AOI22_X1 U14504 ( .A1(n12142), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n11928), .B2(n11591), .ZN(n11592) );
  NAND2_X1 U14505 ( .A1(n14829), .A2(n11595), .ZN(n14811) );
  AOI22_X1 U14506 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14507 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14508 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11891), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14509 ( .A1(n9700), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11596) );
  NAND4_X1 U14510 ( .A1(n11599), .A2(n11598), .A3(n11597), .A4(n11596), .ZN(
        n11609) );
  NAND2_X1 U14511 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11603) );
  NAND2_X1 U14512 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11602) );
  NAND2_X1 U14513 ( .A1(n11339), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11601) );
  NAND2_X1 U14514 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11600) );
  AND4_X1 U14515 ( .A1(n11603), .A2(n11602), .A3(n11601), .A4(n11600), .ZN(
        n11607) );
  AOI22_X1 U14516 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11606) );
  NAND2_X1 U14517 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11605) );
  NAND2_X1 U14518 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11604) );
  NAND4_X1 U14519 ( .A1(n11607), .A2(n11606), .A3(n11605), .A4(n11604), .ZN(
        n11608) );
  NOR2_X1 U14520 ( .A1(n11609), .A2(n11608), .ZN(n11612) );
  AOI21_X1 U14521 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15167), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11610) );
  AOI21_X1 U14522 ( .B1(n12143), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11610), .ZN(
        n11611) );
  OAI21_X1 U14523 ( .B1(n11953), .B2(n11612), .A(n11611), .ZN(n11615) );
  XNOR2_X1 U14524 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B(n11629), .ZN(
        n15169) );
  NAND2_X1 U14525 ( .A1(n11928), .A2(n15169), .ZN(n11614) );
  NAND2_X1 U14526 ( .A1(n11615), .A2(n11614), .ZN(n14813) );
  INV_X1 U14527 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11781) );
  NAND2_X1 U14528 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11617) );
  NAND2_X1 U14529 ( .A1(n9700), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11616) );
  OAI211_X1 U14530 ( .C1(n11934), .C2(n11781), .A(n11617), .B(n11616), .ZN(
        n11618) );
  INV_X1 U14531 ( .A(n11618), .ZN(n11622) );
  AOI22_X1 U14532 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14533 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11620) );
  NAND2_X1 U14534 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11619) );
  NAND4_X1 U14535 ( .A1(n11622), .A2(n11621), .A3(n11620), .A4(n11619), .ZN(
        n11628) );
  AOI22_X1 U14536 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11891), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14537 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14538 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14539 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11623) );
  NAND4_X1 U14540 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11627) );
  NOR2_X1 U14541 ( .A1(n11628), .A2(n11627), .ZN(n11632) );
  XNOR2_X1 U14542 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11649), .ZN(
        n16279) );
  OAI22_X1 U14543 ( .A1(n16279), .A2(n10196), .B1(n13631), .B2(n16277), .ZN(
        n11630) );
  AOI21_X1 U14544 ( .B1(n12143), .B2(P1_EAX_REG_17__SCAN_IN), .A(n11630), .ZN(
        n11631) );
  OAI21_X1 U14545 ( .B1(n11953), .B2(n11632), .A(n11631), .ZN(n14956) );
  NAND2_X1 U14546 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11636) );
  NAND2_X1 U14547 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11635) );
  NAND2_X1 U14548 ( .A1(n11339), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11634) );
  NAND2_X1 U14549 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11633) );
  AND4_X1 U14550 ( .A1(n11636), .A2(n11635), .A3(n11634), .A4(n11633), .ZN(
        n11640) );
  AOI22_X1 U14551 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11639) );
  NAND2_X1 U14552 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11638) );
  NAND2_X1 U14553 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11637) );
  NAND4_X1 U14554 ( .A1(n11640), .A2(n11639), .A3(n11638), .A4(n11637), .ZN(
        n11646) );
  AOI22_X1 U14555 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14556 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14557 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14558 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11118), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11641) );
  NAND4_X1 U14559 ( .A1(n11644), .A2(n11643), .A3(n11642), .A4(n11641), .ZN(
        n11645) );
  NOR2_X1 U14560 ( .A1(n11646), .A2(n11645), .ZN(n11648) );
  AOI22_X1 U14561 ( .A1(n12143), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20966), .ZN(n11647) );
  OAI21_X1 U14562 ( .B1(n11953), .B2(n11648), .A(n11647), .ZN(n11651) );
  XNOR2_X1 U14563 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B(n11670), .ZN(
        n15145) );
  AOI21_X1 U14564 ( .B1(n11651), .B2(n10196), .A(n11650), .ZN(n14796) );
  AOI22_X1 U14565 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14566 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14567 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11118), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14568 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11652) );
  NAND4_X1 U14569 ( .A1(n11655), .A2(n11654), .A3(n11653), .A4(n11652), .ZN(
        n11665) );
  NAND2_X1 U14570 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11659) );
  NAND2_X1 U14571 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11658) );
  NAND2_X1 U14572 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11657) );
  NAND2_X1 U14573 ( .A1(n11339), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11656) );
  AND4_X1 U14574 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(
        n11663) );
  AOI22_X1 U14575 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11662) );
  NAND2_X1 U14576 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11661) );
  NAND2_X1 U14577 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11660) );
  NAND4_X1 U14578 ( .A1(n11663), .A2(n11662), .A3(n11661), .A4(n11660), .ZN(
        n11664) );
  NOR2_X1 U14579 ( .A1(n11665), .A2(n11664), .ZN(n11669) );
  NAND2_X1 U14580 ( .A1(n20966), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11666) );
  NAND2_X1 U14581 ( .A1(n10196), .A2(n11666), .ZN(n11667) );
  AOI21_X1 U14582 ( .B1(n12143), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11667), .ZN(
        n11668) );
  OAI21_X1 U14583 ( .B1(n11953), .B2(n11669), .A(n11668), .ZN(n11676) );
  INV_X1 U14584 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11673) );
  INV_X1 U14585 ( .A(n11671), .ZN(n11672) );
  NAND2_X1 U14586 ( .A1(n11673), .A2(n11672), .ZN(n11674) );
  AND2_X1 U14587 ( .A1(n11694), .A2(n11674), .ZN(n14790) );
  NAND2_X1 U14588 ( .A1(n14790), .A2(n11928), .ZN(n11675) );
  NAND2_X1 U14589 ( .A1(n11676), .A2(n11675), .ZN(n14783) );
  INV_X1 U14590 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11679) );
  NAND2_X1 U14591 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11678) );
  NAND2_X1 U14592 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11677) );
  OAI211_X1 U14593 ( .C1(n11934), .C2(n11679), .A(n11678), .B(n11677), .ZN(
        n11680) );
  INV_X1 U14594 ( .A(n11680), .ZN(n11684) );
  AOI22_X1 U14595 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14596 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11270), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11682) );
  NAND2_X1 U14597 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11681) );
  NAND4_X1 U14598 ( .A1(n11684), .A2(n11683), .A3(n11682), .A4(n11681), .ZN(
        n11690) );
  AOI22_X1 U14599 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11940), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14600 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n9690), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14601 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14602 ( .A1(n9700), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11685) );
  NAND4_X1 U14603 ( .A1(n11688), .A2(n11687), .A3(n11686), .A4(n11685), .ZN(
        n11689) );
  NOR2_X1 U14604 ( .A1(n11690), .A2(n11689), .ZN(n11693) );
  OAI21_X1 U14605 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21227), .A(n10196), 
        .ZN(n11691) );
  AOI21_X1 U14606 ( .B1(n12143), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11691), .ZN(
        n11692) );
  OAI21_X1 U14607 ( .B1(n11953), .B2(n11693), .A(n11692), .ZN(n11697) );
  INV_X1 U14608 ( .A(n11716), .ZN(n11717) );
  NAND2_X1 U14609 ( .A1(n11694), .A2(n21227), .ZN(n11695) );
  NAND2_X1 U14610 ( .A1(n15130), .A2(n11928), .ZN(n11696) );
  AOI22_X1 U14611 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U14612 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11891), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14613 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14614 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11698) );
  NAND4_X1 U14615 ( .A1(n11701), .A2(n11700), .A3(n11699), .A4(n11698), .ZN(
        n11711) );
  AOI22_X1 U14616 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11709) );
  NAND2_X1 U14617 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11705) );
  NAND2_X1 U14618 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11704) );
  NAND2_X1 U14619 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11703) );
  NAND2_X1 U14620 ( .A1(n11339), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11702) );
  AND4_X1 U14621 ( .A1(n11705), .A2(n11704), .A3(n11703), .A4(n11702), .ZN(
        n11708) );
  NAND2_X1 U14622 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11707) );
  NAND2_X1 U14623 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11706) );
  NAND4_X1 U14624 ( .A1(n11709), .A2(n11708), .A3(n11707), .A4(n11706), .ZN(
        n11710) );
  NOR2_X1 U14625 ( .A1(n11711), .A2(n11710), .ZN(n11715) );
  NAND2_X1 U14626 ( .A1(n20966), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11712) );
  NAND2_X1 U14627 ( .A1(n10196), .A2(n11712), .ZN(n11713) );
  AOI21_X1 U14628 ( .B1(n12143), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11713), .ZN(
        n11714) );
  OAI21_X1 U14629 ( .B1(n11953), .B2(n11715), .A(n11714), .ZN(n11720) );
  INV_X1 U14630 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14762) );
  NAND2_X1 U14631 ( .A1(n11717), .A2(n14762), .ZN(n11718) );
  NAND2_X1 U14632 ( .A1(n11741), .A2(n11718), .ZN(n15121) );
  INV_X1 U14633 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11723) );
  NAND2_X1 U14634 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11722) );
  NAND2_X1 U14635 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11721) );
  OAI211_X1 U14636 ( .C1(n11934), .C2(n11723), .A(n11722), .B(n11721), .ZN(
        n11724) );
  INV_X1 U14637 ( .A(n11724), .ZN(n11728) );
  AOI22_X1 U14638 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U14639 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11726) );
  NAND2_X1 U14640 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11725) );
  NAND4_X1 U14641 ( .A1(n11728), .A2(n11727), .A3(n11726), .A4(n11725), .ZN(
        n11734) );
  AOI22_X1 U14642 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14643 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14644 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U14645 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11729) );
  NAND4_X1 U14646 ( .A1(n11732), .A2(n11731), .A3(n11730), .A4(n11729), .ZN(
        n11733) );
  NOR2_X1 U14647 ( .A1(n11734), .A2(n11733), .ZN(n11737) );
  INV_X1 U14648 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11740) );
  AOI21_X1 U14649 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n11740), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11735) );
  AOI21_X1 U14650 ( .B1(n12143), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11735), .ZN(
        n11736) );
  OAI21_X1 U14651 ( .B1(n11953), .B2(n11737), .A(n11736), .ZN(n11739) );
  XNOR2_X1 U14652 ( .A(n11741), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15110) );
  NAND2_X1 U14653 ( .A1(n15110), .A2(n11928), .ZN(n11738) );
  NAND2_X1 U14654 ( .A1(n11739), .A2(n11738), .ZN(n14743) );
  INV_X1 U14655 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14731) );
  NAND2_X1 U14656 ( .A1(n11742), .A2(n14731), .ZN(n11743) );
  NAND2_X1 U14657 ( .A1(n11776), .A2(n11743), .ZN(n15103) );
  INV_X1 U14658 ( .A(n15103), .ZN(n11775) );
  OAI21_X1 U14659 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14731), .A(n10196), 
        .ZN(n11773) );
  INV_X1 U14660 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11745) );
  INV_X1 U14661 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11744) );
  OAI22_X1 U14662 ( .A1(n11830), .A2(n11745), .B1(n11880), .B2(n11744), .ZN(
        n11749) );
  INV_X1 U14663 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11746) );
  OAI22_X1 U14664 ( .A1(n9674), .A2(n11747), .B1(n11123), .B2(n11746), .ZN(
        n11748) );
  AOI211_X1 U14665 ( .C1(n11236), .C2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n11749), .B(n11748), .ZN(n11757) );
  AOI22_X1 U14666 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U14667 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U14668 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14669 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11750) );
  AND4_X1 U14670 ( .A1(n11753), .A2(n11752), .A3(n11751), .A4(n11750), .ZN(
        n11756) );
  AOI22_X1 U14671 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11755) );
  NAND2_X1 U14672 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11754) );
  NAND4_X1 U14673 ( .A1(n11757), .A2(n11756), .A3(n11755), .A4(n11754), .ZN(
        n11778) );
  INV_X1 U14674 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11759) );
  INV_X1 U14675 ( .A(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11758) );
  OAI22_X1 U14676 ( .A1(n11830), .A2(n11759), .B1(n11880), .B2(n11758), .ZN(
        n11762) );
  INV_X1 U14677 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n21203) );
  OAI22_X1 U14678 ( .A1(n9674), .A2(n11760), .B1(n11123), .B2(n21203), .ZN(
        n11761) );
  AOI211_X1 U14679 ( .C1(n11236), .C2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n11762), .B(n11761), .ZN(n11770) );
  AOI22_X1 U14680 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U14681 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U14682 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14683 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9700), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11763) );
  AND4_X1 U14684 ( .A1(n11766), .A2(n11765), .A3(n11764), .A4(n11763), .ZN(
        n11769) );
  AOI22_X1 U14685 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11768) );
  NAND2_X1 U14686 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11767) );
  NAND4_X1 U14687 ( .A1(n11770), .A2(n11769), .A3(n11768), .A4(n11767), .ZN(
        n11779) );
  XNOR2_X1 U14688 ( .A(n11778), .B(n11779), .ZN(n11771) );
  NOR2_X1 U14689 ( .A1(n11771), .A2(n11953), .ZN(n11772) );
  AOI211_X1 U14690 ( .C1(n12143), .C2(P1_EAX_REG_23__SCAN_IN), .A(n11773), .B(
        n11772), .ZN(n11774) );
  AOI21_X1 U14691 ( .B1(n11928), .B2(n11775), .A(n11774), .ZN(n14730) );
  INV_X1 U14692 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14721) );
  INV_X1 U14693 ( .A(n11803), .ZN(n11804) );
  NAND2_X1 U14694 ( .A1(n11776), .A2(n14721), .ZN(n11777) );
  NAND2_X1 U14695 ( .A1(n11804), .A2(n11777), .ZN(n15096) );
  INV_X1 U14696 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n11801) );
  NAND2_X1 U14697 ( .A1(n11779), .A2(n11778), .ZN(n11806) );
  INV_X1 U14698 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11790) );
  INV_X1 U14699 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11782) );
  OAI22_X1 U14700 ( .A1(n11885), .A2(n11782), .B1(n11880), .B2(n11781), .ZN(
        n11786) );
  INV_X1 U14701 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11784) );
  INV_X1 U14702 ( .A(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11783) );
  OAI22_X1 U14703 ( .A1(n11882), .A2(n11784), .B1(n9682), .B2(n11783), .ZN(
        n11785) );
  AOI211_X1 U14704 ( .C1(n11787), .C2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n11786), .B(n11785), .ZN(n11789) );
  AOI22_X1 U14705 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11788) );
  OAI211_X1 U14706 ( .C1(n11086), .C2(n11790), .A(n11789), .B(n11788), .ZN(
        n11797) );
  AOI22_X1 U14707 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11215), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U14708 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14709 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U14710 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11792) );
  NAND4_X1 U14711 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(
        n11796) );
  NOR2_X1 U14712 ( .A1(n11797), .A2(n11796), .ZN(n11807) );
  XOR2_X1 U14713 ( .A(n11806), .B(n11807), .Z(n11798) );
  INV_X1 U14714 ( .A(n11953), .ZN(n11920) );
  NAND2_X1 U14715 ( .A1(n11798), .A2(n11920), .ZN(n11800) );
  AOI21_X1 U14716 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20966), .A(
        n11928), .ZN(n11799) );
  OAI211_X1 U14717 ( .C1(n11902), .C2(n11801), .A(n11800), .B(n11799), .ZN(
        n11802) );
  INV_X1 U14718 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14707) );
  NAND2_X1 U14719 ( .A1(n11804), .A2(n14707), .ZN(n11805) );
  AND2_X1 U14720 ( .A1(n11851), .A2(n11805), .ZN(n14706) );
  OAI21_X1 U14721 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14707), .A(n10196), 
        .ZN(n11824) );
  NOR2_X1 U14722 ( .A1(n11807), .A2(n11806), .ZN(n11827) );
  INV_X1 U14723 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11810) );
  NAND2_X1 U14724 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11809) );
  NAND2_X1 U14725 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11808) );
  OAI211_X1 U14726 ( .C1(n11934), .C2(n11810), .A(n11809), .B(n11808), .ZN(
        n11811) );
  INV_X1 U14727 ( .A(n11811), .ZN(n11815) );
  AOI22_X1 U14728 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14729 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11813) );
  NAND2_X1 U14730 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11812) );
  NAND4_X1 U14731 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n11812), .ZN(
        n11821) );
  AOI22_X1 U14732 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U14733 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U14734 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11817) );
  AOI22_X1 U14735 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11816) );
  NAND4_X1 U14736 ( .A1(n11819), .A2(n11818), .A3(n11817), .A4(n11816), .ZN(
        n11820) );
  OR2_X1 U14737 ( .A1(n11821), .A2(n11820), .ZN(n11826) );
  XNOR2_X1 U14738 ( .A(n11827), .B(n11826), .ZN(n11822) );
  NOR2_X1 U14739 ( .A1(n11822), .A2(n11953), .ZN(n11823) );
  AOI211_X1 U14740 ( .C1(n12143), .C2(P1_EAX_REG_25__SCAN_IN), .A(n11824), .B(
        n11823), .ZN(n11825) );
  AOI21_X1 U14741 ( .B1(n11928), .B2(n14706), .A(n11825), .ZN(n14702) );
  NAND2_X1 U14742 ( .A1(n14701), .A2(n14702), .ZN(n14691) );
  INV_X1 U14743 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14693) );
  XNOR2_X1 U14744 ( .A(n11851), .B(n14693), .ZN(n15076) );
  INV_X1 U14745 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U14746 ( .A1(n11827), .A2(n11826), .ZN(n11855) );
  INV_X1 U14747 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11837) );
  INV_X1 U14748 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11829) );
  INV_X1 U14749 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11828) );
  OAI22_X1 U14750 ( .A1(n11830), .A2(n11829), .B1(n11880), .B2(n11828), .ZN(
        n11834) );
  INV_X1 U14751 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11831) );
  OAI22_X1 U14752 ( .A1(n9674), .A2(n11832), .B1(n11123), .B2(n11831), .ZN(
        n11833) );
  AOI211_X1 U14753 ( .C1(n11236), .C2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n11834), .B(n11833), .ZN(n11836) );
  AOI22_X1 U14754 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11891), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11835) );
  OAI211_X1 U14755 ( .C1(n11934), .C2(n11837), .A(n11836), .B(n11835), .ZN(
        n11845) );
  AOI22_X1 U14756 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11270), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U14757 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U14758 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9700), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U14759 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11840) );
  NAND4_X1 U14760 ( .A1(n11843), .A2(n11842), .A3(n11841), .A4(n11840), .ZN(
        n11844) );
  NOR2_X1 U14761 ( .A1(n11845), .A2(n11844), .ZN(n11856) );
  XOR2_X1 U14762 ( .A(n11855), .B(n11856), .Z(n11846) );
  NAND2_X1 U14763 ( .A1(n11846), .A2(n11920), .ZN(n11848) );
  INV_X1 U14764 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20852) );
  OAI21_X1 U14765 ( .B1(n20852), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n20966), .ZN(n11847) );
  OAI211_X1 U14766 ( .C1(n11902), .C2(n11849), .A(n11848), .B(n11847), .ZN(
        n11850) );
  INV_X1 U14767 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11854) );
  INV_X1 U14768 ( .A(n11924), .ZN(n11876) );
  NAND2_X1 U14769 ( .A1(n11852), .A2(n11854), .ZN(n11853) );
  OAI21_X1 U14770 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n11854), .A(n10196), 
        .ZN(n11874) );
  NOR2_X1 U14771 ( .A1(n11856), .A2(n11855), .ZN(n11878) );
  INV_X1 U14772 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11859) );
  NAND2_X1 U14773 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11858) );
  NAND2_X1 U14774 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11857) );
  OAI211_X1 U14775 ( .C1(n11934), .C2(n11859), .A(n11858), .B(n11857), .ZN(
        n11860) );
  INV_X1 U14776 ( .A(n11860), .ZN(n11865) );
  AOI22_X1 U14777 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14778 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11863) );
  NAND2_X1 U14779 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11862) );
  NAND4_X1 U14780 ( .A1(n11865), .A2(n11864), .A3(n11863), .A4(n11862), .ZN(
        n11871) );
  AOI22_X1 U14781 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11270), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14782 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11940), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U14783 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U14784 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11866) );
  NAND4_X1 U14785 ( .A1(n11869), .A2(n11868), .A3(n11867), .A4(n11866), .ZN(
        n11870) );
  OR2_X1 U14786 ( .A1(n11871), .A2(n11870), .ZN(n11877) );
  XNOR2_X1 U14787 ( .A(n11878), .B(n11877), .ZN(n11872) );
  NOR2_X1 U14788 ( .A1(n11872), .A2(n11953), .ZN(n11873) );
  AOI211_X1 U14789 ( .C1(n12143), .C2(P1_EAX_REG_27__SCAN_IN), .A(n11874), .B(
        n11873), .ZN(n11875) );
  INV_X1 U14790 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14670) );
  XNOR2_X1 U14791 ( .A(n11876), .B(n14670), .ZN(n15058) );
  INV_X1 U14792 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n11901) );
  NAND2_X1 U14793 ( .A1(n11878), .A2(n11877), .ZN(n11904) );
  INV_X1 U14794 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11890) );
  INV_X1 U14795 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11881) );
  INV_X1 U14796 ( .A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11879) );
  OAI22_X1 U14797 ( .A1(n11882), .A2(n11881), .B1(n11880), .B2(n11879), .ZN(
        n11887) );
  OAI22_X1 U14798 ( .A1(n11885), .A2(n11884), .B1(n9674), .B2(n11883), .ZN(
        n11886) );
  AOI211_X1 U14799 ( .C1(n11236), .C2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n11887), .B(n11886), .ZN(n11889) );
  AOI22_X1 U14800 ( .A1(n9698), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11839), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11888) );
  OAI211_X1 U14801 ( .C1(n11934), .C2(n11890), .A(n11889), .B(n11888), .ZN(
        n11897) );
  AOI22_X1 U14802 ( .A1(n9690), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11791), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U14803 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11891), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U14804 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11213), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U14805 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11892) );
  NAND4_X1 U14806 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11896) );
  NOR2_X1 U14807 ( .A1(n11897), .A2(n11896), .ZN(n11905) );
  XOR2_X1 U14808 ( .A(n11904), .B(n11905), .Z(n11898) );
  NAND2_X1 U14809 ( .A1(n11898), .A2(n11920), .ZN(n11900) );
  AOI21_X1 U14810 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20966), .A(
        n11928), .ZN(n11899) );
  OAI211_X1 U14811 ( .C1(n11902), .C2(n11901), .A(n11900), .B(n11899), .ZN(
        n11903) );
  NOR2_X1 U14812 ( .A1(n11905), .A2(n11904), .ZN(n11922) );
  INV_X1 U14813 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11908) );
  NAND2_X1 U14814 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11907) );
  NAND2_X1 U14815 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11906) );
  OAI211_X1 U14816 ( .C1(n11934), .C2(n11908), .A(n11907), .B(n11906), .ZN(
        n11909) );
  INV_X1 U14817 ( .A(n11909), .ZN(n11913) );
  AOI22_X1 U14818 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U14819 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11911) );
  NAND2_X1 U14820 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11910) );
  NAND4_X1 U14821 ( .A1(n11913), .A2(n11912), .A3(n11911), .A4(n11910), .ZN(
        n11919) );
  AOI22_X1 U14822 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11917) );
  AOI22_X1 U14823 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11916) );
  AOI22_X1 U14824 ( .A1(n9704), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U14825 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11914) );
  NAND4_X1 U14826 ( .A1(n11917), .A2(n11916), .A3(n11915), .A4(n11914), .ZN(
        n11918) );
  OR2_X1 U14827 ( .A1(n11919), .A2(n11918), .ZN(n11921) );
  NAND2_X1 U14828 ( .A1(n11922), .A2(n11921), .ZN(n11949) );
  OAI211_X1 U14829 ( .C1(n11922), .C2(n11921), .A(n11949), .B(n11920), .ZN(
        n11930) );
  INV_X1 U14830 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14321) );
  NOR2_X1 U14831 ( .A1(n14321), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11923) );
  AOI211_X1 U14832 ( .C1(n12143), .C2(P1_EAX_REG_29__SCAN_IN), .A(n11928), .B(
        n11923), .ZN(n11929) );
  INV_X1 U14833 ( .A(n11925), .ZN(n11926) );
  NAND2_X1 U14834 ( .A1(n11926), .A2(n14321), .ZN(n11927) );
  AOI22_X1 U14835 ( .A1(n11930), .A2(n11929), .B1(n11928), .B2(n14320), .ZN(
        n14317) );
  INV_X1 U14836 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11933) );
  NAND2_X1 U14837 ( .A1(n11118), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11932) );
  NAND2_X1 U14838 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11931) );
  OAI211_X1 U14839 ( .C1(n11934), .C2(n11933), .A(n11932), .B(n11931), .ZN(
        n11935) );
  INV_X1 U14840 ( .A(n11935), .ZN(n11939) );
  AOI22_X1 U14841 ( .A1(n11213), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11339), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U14842 ( .A1(n11215), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11937) );
  NAND2_X1 U14843 ( .A1(n11236), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11936) );
  NAND4_X1 U14844 ( .A1(n11939), .A2(n11938), .A3(n11937), .A4(n11936), .ZN(
        n11947) );
  AOI22_X1 U14845 ( .A1(n11270), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9690), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U14846 ( .A1(n11940), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U14847 ( .A1(n9703), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9698), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U14848 ( .A1(n11791), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11941), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11942) );
  NAND4_X1 U14849 ( .A1(n11945), .A2(n11944), .A3(n11943), .A4(n11942), .ZN(
        n11946) );
  NOR2_X1 U14850 ( .A1(n11947), .A2(n11946), .ZN(n11948) );
  XNOR2_X1 U14851 ( .A(n11949), .B(n11948), .ZN(n11954) );
  NAND2_X1 U14852 ( .A1(n20966), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11950) );
  NAND2_X1 U14853 ( .A1(n10196), .A2(n11950), .ZN(n11951) );
  AOI21_X1 U14854 ( .B1(n12143), .B2(P1_EAX_REG_30__SCAN_IN), .A(n11951), .ZN(
        n11952) );
  OAI21_X1 U14855 ( .B1(n11954), .B2(n11953), .A(n11952), .ZN(n11957) );
  XNOR2_X1 U14856 ( .A(n11955), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15036) );
  NAND2_X1 U14857 ( .A1(n15036), .A2(n11928), .ZN(n11956) );
  NAND2_X1 U14858 ( .A1(n11957), .A2(n11956), .ZN(n12140) );
  XNOR2_X2 U14859 ( .A(n12141), .B(n12140), .ZN(n15040) );
  XNOR2_X1 U14860 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11974) );
  NAND2_X1 U14861 ( .A1(n11973), .A2(n11974), .ZN(n11959) );
  NAND2_X1 U14862 ( .A1(n20722), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11958) );
  XNOR2_X1 U14863 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11985) );
  XNOR2_X1 U14864 ( .A(n13581), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11964) );
  INV_X1 U14865 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20418) );
  NOR2_X1 U14866 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20418), .ZN(
        n11960) );
  NAND2_X1 U14867 ( .A1(n12015), .A2(n11998), .ZN(n12007) );
  NAND2_X1 U14868 ( .A1(n12015), .A2(n11990), .ZN(n12005) );
  NAND3_X1 U14869 ( .A1(n16422), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n11961), .ZN(n12013) );
  INV_X1 U14870 ( .A(n11998), .ZN(n12002) );
  AOI21_X1 U14871 ( .B1(n11964), .B2(n11963), .A(n11962), .ZN(n11965) );
  INV_X1 U14872 ( .A(n11965), .ZN(n12010) );
  INV_X1 U14873 ( .A(n11973), .ZN(n11966) );
  OAI21_X1 U14874 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20820), .A(
        n11966), .ZN(n11967) );
  NOR2_X1 U14875 ( .A1(n11987), .A2(n11967), .ZN(n11972) );
  INV_X1 U14876 ( .A(n11967), .ZN(n11969) );
  OAI21_X1 U14877 ( .B1(n11170), .B2(n13642), .A(n11968), .ZN(n11989) );
  OAI211_X1 U14878 ( .C1(n13030), .C2(n11970), .A(n11969), .B(n11989), .ZN(
        n11971) );
  OAI21_X1 U14879 ( .B1(n11998), .B2(n11972), .A(n11971), .ZN(n11979) );
  INV_X1 U14880 ( .A(n11979), .ZN(n11984) );
  XNOR2_X1 U14881 ( .A(n11974), .B(n11973), .ZN(n12012) );
  NOR2_X1 U14882 ( .A1(n13642), .A2(n20963), .ZN(n11976) );
  NOR2_X1 U14883 ( .A1(n11987), .A2(n11968), .ZN(n11975) );
  AOI211_X1 U14884 ( .C1(n11999), .C2(n12012), .A(n11976), .B(n11975), .ZN(
        n11980) );
  INV_X1 U14885 ( .A(n11980), .ZN(n11983) );
  INV_X1 U14886 ( .A(n11976), .ZN(n11977) );
  NAND2_X1 U14887 ( .A1(n11977), .A2(n13637), .ZN(n11978) );
  OR2_X1 U14888 ( .A1(n11978), .A2(n11990), .ZN(n11981) );
  AOI22_X1 U14889 ( .A1(n12012), .A2(n11981), .B1(n11980), .B2(n11979), .ZN(
        n11982) );
  AOI21_X1 U14890 ( .B1(n11984), .B2(n11983), .A(n11982), .ZN(n11994) );
  XNOR2_X1 U14891 ( .A(n11986), .B(n11985), .ZN(n12011) );
  OAI21_X1 U14892 ( .B1(n11987), .B2(n12011), .A(n11989), .ZN(n11988) );
  AOI21_X1 U14893 ( .B1(n11999), .B2(n12011), .A(n11988), .ZN(n11993) );
  INV_X1 U14894 ( .A(n11989), .ZN(n11991) );
  NAND2_X1 U14895 ( .A1(n11991), .A2(n11990), .ZN(n11992) );
  OAI22_X1 U14896 ( .A1(n11994), .A2(n11993), .B1(n12011), .B2(n11992), .ZN(
        n11997) );
  NAND2_X1 U14897 ( .A1(n11995), .A2(n12010), .ZN(n11996) );
  AOI22_X1 U14898 ( .A1(n11998), .A2(n12010), .B1(n11997), .B2(n11996), .ZN(
        n12001) );
  NOR2_X1 U14899 ( .A1(n11999), .A2(n12013), .ZN(n12000) );
  OAI22_X1 U14900 ( .A1(n12013), .A2(n12002), .B1(n12001), .B2(n12000), .ZN(
        n12003) );
  AOI21_X1 U14901 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20963), .A(
        n12003), .ZN(n12004) );
  NAND2_X1 U14902 ( .A1(n12005), .A2(n12004), .ZN(n12006) );
  NAND2_X1 U14903 ( .A1(n16243), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20238) );
  INV_X1 U14904 ( .A(n12008), .ZN(n13028) );
  NOR2_X1 U14905 ( .A1(n12009), .A2(n20238), .ZN(n12016) );
  NOR3_X1 U14906 ( .A1(n12012), .A2(n12011), .A3(n12010), .ZN(n12014) );
  OAI21_X1 U14907 ( .B1(n12015), .B2(n12014), .A(n12013), .ZN(n13281) );
  NAND2_X1 U14908 ( .A1(n12016), .A2(n13281), .ZN(n12943) );
  AND2_X1 U14909 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20963), .ZN(n12018) );
  NAND2_X1 U14910 ( .A1(n20966), .A2(n20962), .ZN(n16429) );
  INV_X1 U14911 ( .A(n16429), .ZN(n21054) );
  NAND2_X1 U14912 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21054), .ZN(n16244) );
  INV_X1 U14913 ( .A(n16244), .ZN(n12017) );
  AOI22_X1 U14914 ( .A1(n11928), .A2(n12018), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n12017), .ZN(n12019) );
  AND2_X1 U14915 ( .A1(n20393), .A2(n12019), .ZN(n12020) );
  NAND2_X1 U14916 ( .A1(n12021), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12022) );
  XNOR2_X1 U14917 ( .A(n12022), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15030) );
  AND2_X1 U14918 ( .A1(n15030), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12023) );
  NAND2_X1 U14919 ( .A1(n12033), .A2(n9656), .ZN(n12024) );
  INV_X1 U14920 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13920) );
  OAI22_X1 U14921 ( .A1(n12105), .A2(n13920), .B1(n12472), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13326) );
  XNOR2_X1 U14922 ( .A(n12026), .B(n13326), .ZN(n13108) );
  NAND2_X1 U14923 ( .A1(n13108), .A2(n13107), .ZN(n12028) );
  INV_X1 U14924 ( .A(n12026), .ZN(n12027) );
  NAND2_X1 U14925 ( .A1(n12028), .A2(n12027), .ZN(n13430) );
  INV_X1 U14926 ( .A(n13430), .ZN(n12032) );
  MUX2_X1 U14927 ( .A(n9724), .B(n9656), .S(P1_EBX_REG_2__SCAN_IN), .Z(n12029)
         );
  INV_X1 U14928 ( .A(n12029), .ZN(n12030) );
  NAND2_X1 U14929 ( .A1(n12030), .A2(n10187), .ZN(n13429) );
  MUX2_X1 U14930 ( .A(n12112), .B(n12053), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12035) );
  INV_X1 U14931 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20387) );
  NAND2_X1 U14932 ( .A1(n12053), .A2(n12033), .ZN(n12055) );
  OAI21_X1 U14933 ( .B1(n13107), .B2(n20387), .A(n12055), .ZN(n12034) );
  NOR2_X1 U14934 ( .A1(n12035), .A2(n12034), .ZN(n13468) );
  INV_X1 U14935 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13969) );
  NAND2_X1 U14936 ( .A1(n9724), .A2(n13969), .ZN(n12038) );
  NAND2_X1 U14937 ( .A1(n12472), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12036) );
  OAI211_X1 U14938 ( .C1(n12033), .C2(P1_EBX_REG_4__SCAN_IN), .A(n12105), .B(
        n12036), .ZN(n12037) );
  AND2_X1 U14939 ( .A1(n12038), .A2(n12037), .ZN(n13448) );
  MUX2_X1 U14940 ( .A(n12112), .B(n12053), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n12041) );
  NAND2_X1 U14941 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12033), .ZN(
        n12039) );
  NAND2_X1 U14942 ( .A1(n12055), .A2(n12039), .ZN(n12040) );
  NOR2_X1 U14943 ( .A1(n12041), .A2(n12040), .ZN(n13736) );
  INV_X1 U14944 ( .A(n9724), .ZN(n12091) );
  NAND2_X1 U14945 ( .A1(n12472), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12044) );
  OAI211_X1 U14946 ( .C1(n12033), .C2(P1_EBX_REG_6__SCAN_IN), .A(n12105), .B(
        n12044), .ZN(n12045) );
  OAI21_X1 U14947 ( .B1(n12091), .B2(P1_EBX_REG_6__SCAN_IN), .A(n12045), .ZN(
        n16398) );
  MUX2_X1 U14948 ( .A(n12112), .B(n12053), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n12048) );
  NAND2_X1 U14949 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n12033), .ZN(
        n12046) );
  NAND2_X1 U14950 ( .A1(n12055), .A2(n12046), .ZN(n12047) );
  NOR2_X1 U14951 ( .A1(n12048), .A2(n12047), .ZN(n13825) );
  INV_X1 U14952 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n12049) );
  NAND2_X1 U14953 ( .A1(n9724), .A2(n12049), .ZN(n12052) );
  NAND2_X1 U14954 ( .A1(n12472), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12050) );
  OAI211_X1 U14955 ( .C1(n12033), .C2(P1_EBX_REG_8__SCAN_IN), .A(n12105), .B(
        n12050), .ZN(n12051) );
  MUX2_X1 U14956 ( .A(n12112), .B(n12053), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n12057) );
  NAND2_X1 U14957 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n12033), .ZN(
        n12054) );
  NAND2_X1 U14958 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  NOR2_X1 U14959 ( .A1(n12057), .A2(n12056), .ZN(n14024) );
  MUX2_X1 U14960 ( .A(n9724), .B(n9656), .S(P1_EBX_REG_10__SCAN_IN), .Z(n12058) );
  INV_X1 U14961 ( .A(n12058), .ZN(n12059) );
  NAND2_X1 U14962 ( .A1(n12059), .A2(n10180), .ZN(n14031) );
  INV_X1 U14963 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15005) );
  NAND2_X1 U14964 ( .A1(n12105), .A2(n15005), .ZN(n12061) );
  OAI211_X1 U14965 ( .C1(n12033), .C2(P1_EBX_REG_11__SCAN_IN), .A(n12472), .B(
        n12061), .ZN(n12062) );
  OAI21_X1 U14966 ( .B1(n12106), .B2(P1_EBX_REG_11__SCAN_IN), .A(n12062), .ZN(
        n14893) );
  INV_X1 U14967 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n16311) );
  NAND2_X1 U14968 ( .A1(n9724), .A2(n16311), .ZN(n12065) );
  NAND2_X1 U14969 ( .A1(n12472), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12063) );
  OAI211_X1 U14970 ( .C1(n12033), .C2(P1_EBX_REG_12__SCAN_IN), .A(n12105), .B(
        n12063), .ZN(n12064) );
  INV_X1 U14971 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14887) );
  NAND2_X1 U14972 ( .A1(n12112), .A2(n14887), .ZN(n12068) );
  INV_X1 U14973 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15008) );
  NAND2_X1 U14974 ( .A1(n12105), .A2(n15008), .ZN(n12066) );
  OAI211_X1 U14975 ( .C1(n12033), .C2(P1_EBX_REG_13__SCAN_IN), .A(n12472), .B(
        n12066), .ZN(n12067) );
  MUX2_X1 U14976 ( .A(n9724), .B(n9656), .S(P1_EBX_REG_14__SCAN_IN), .Z(n12069) );
  INV_X1 U14977 ( .A(n12069), .ZN(n12071) );
  INV_X1 U14978 ( .A(n13325), .ZN(n13206) );
  INV_X1 U14979 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15376) );
  NAND2_X1 U14980 ( .A1(n13206), .A2(n15376), .ZN(n12070) );
  NAND2_X1 U14981 ( .A1(n12071), .A2(n12070), .ZN(n14836) );
  INV_X1 U14982 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15368) );
  NAND2_X1 U14983 ( .A1(n12105), .A2(n15368), .ZN(n12072) );
  OAI211_X1 U14984 ( .C1(n12033), .C2(P1_EBX_REG_15__SCAN_IN), .A(n12472), .B(
        n12072), .ZN(n12073) );
  OAI21_X1 U14985 ( .B1(n12106), .B2(P1_EBX_REG_15__SCAN_IN), .A(n12073), .ZN(
        n14878) );
  MUX2_X1 U14986 ( .A(n9724), .B(n9656), .S(P1_EBX_REG_16__SCAN_IN), .Z(n12075) );
  NOR2_X1 U14987 ( .A1(n13325), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12074) );
  NOR2_X1 U14988 ( .A1(n12075), .A2(n12074), .ZN(n14823) );
  INV_X1 U14989 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n21212) );
  NAND2_X1 U14990 ( .A1(n12112), .A2(n21212), .ZN(n12078) );
  INV_X1 U14991 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15208) );
  NAND2_X1 U14992 ( .A1(n12105), .A2(n15208), .ZN(n12076) );
  OAI211_X1 U14993 ( .C1(n12033), .C2(P1_EBX_REG_17__SCAN_IN), .A(n12472), .B(
        n12076), .ZN(n12077) );
  NAND2_X1 U14994 ( .A1(n12472), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12079) );
  OAI211_X1 U14995 ( .C1(n12033), .C2(P1_EBX_REG_18__SCAN_IN), .A(n12105), .B(
        n12079), .ZN(n12080) );
  OAI21_X1 U14996 ( .B1(n12091), .B2(P1_EBX_REG_18__SCAN_IN), .A(n12080), .ZN(
        n14800) );
  INV_X1 U14997 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14791) );
  NAND2_X1 U14998 ( .A1(n12112), .A2(n14791), .ZN(n12083) );
  INV_X1 U14999 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15352) );
  NAND2_X1 U15000 ( .A1(n12105), .A2(n15352), .ZN(n12081) );
  OAI211_X1 U15001 ( .C1(n12033), .C2(P1_EBX_REG_19__SCAN_IN), .A(n12472), .B(
        n12081), .ZN(n12082) );
  INV_X1 U15002 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14874) );
  NAND2_X1 U15003 ( .A1(n9724), .A2(n14874), .ZN(n12086) );
  NAND2_X1 U15004 ( .A1(n12472), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12084) );
  OAI211_X1 U15005 ( .C1(n12033), .C2(P1_EBX_REG_20__SCAN_IN), .A(n12105), .B(
        n12084), .ZN(n12085) );
  MUX2_X1 U15006 ( .A(n12106), .B(n12105), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12088) );
  NAND2_X1 U15007 ( .A1(n12033), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12087) );
  AND2_X1 U15008 ( .A1(n12088), .A2(n12087), .ZN(n14759) );
  NAND2_X1 U15009 ( .A1(n12472), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12089) );
  OAI211_X1 U15010 ( .C1(n12033), .C2(P1_EBX_REG_22__SCAN_IN), .A(n12105), .B(
        n12089), .ZN(n12090) );
  OAI21_X1 U15011 ( .B1(n12091), .B2(P1_EBX_REG_22__SCAN_IN), .A(n12090), .ZN(
        n14744) );
  INV_X1 U15012 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15300) );
  NAND2_X1 U15013 ( .A1(n12105), .A2(n15300), .ZN(n12092) );
  OAI211_X1 U15014 ( .C1(n12033), .C2(P1_EBX_REG_23__SCAN_IN), .A(n12472), .B(
        n12092), .ZN(n12093) );
  OAI21_X1 U15015 ( .B1(n12106), .B2(P1_EBX_REG_23__SCAN_IN), .A(n12093), .ZN(
        n14729) );
  MUX2_X1 U15016 ( .A(n9724), .B(n9656), .S(P1_EBX_REG_24__SCAN_IN), .Z(n12094) );
  INV_X1 U15017 ( .A(n12094), .ZN(n12096) );
  INV_X1 U15018 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15221) );
  NAND2_X1 U15019 ( .A1(n13206), .A2(n15221), .ZN(n12095) );
  NAND2_X1 U15020 ( .A1(n12096), .A2(n12095), .ZN(n14718) );
  INV_X1 U15021 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n12097) );
  NAND2_X1 U15022 ( .A1(n12112), .A2(n12097), .ZN(n12100) );
  INV_X1 U15023 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15273) );
  NAND2_X1 U15024 ( .A1(n12105), .A2(n15273), .ZN(n12098) );
  OAI211_X1 U15025 ( .C1(n12033), .C2(P1_EBX_REG_25__SCAN_IN), .A(n12472), .B(
        n12098), .ZN(n12099) );
  AND2_X1 U15026 ( .A1(n12100), .A2(n12099), .ZN(n14704) );
  MUX2_X1 U15027 ( .A(n9724), .B(n9656), .S(P1_EBX_REG_26__SCAN_IN), .Z(n12102) );
  NOR2_X1 U15028 ( .A1(n13325), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12101) );
  NOR2_X1 U15029 ( .A1(n12102), .A2(n12101), .ZN(n14688) );
  MUX2_X1 U15030 ( .A(n9724), .B(n9656), .S(P1_EBX_REG_28__SCAN_IN), .Z(n12104) );
  NOR2_X1 U15031 ( .A1(n13325), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12103) );
  NOR2_X1 U15032 ( .A1(n12104), .A2(n12103), .ZN(n14666) );
  MUX2_X1 U15033 ( .A(n12106), .B(n12105), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12108) );
  NAND2_X1 U15034 ( .A1(n12033), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12107) );
  NAND2_X1 U15035 ( .A1(n12108), .A2(n12107), .ZN(n14678) );
  AND2_X1 U15036 ( .A1(n14666), .A2(n14678), .ZN(n12109) );
  OR2_X1 U15037 ( .A1(n12033), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12110) );
  OAI21_X1 U15038 ( .B1(n13325), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12110), .ZN(n12115) );
  OR2_X1 U15039 ( .A1(n12115), .A2(n9656), .ZN(n12114) );
  INV_X1 U15040 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n12111) );
  NAND2_X1 U15041 ( .A1(n12112), .A2(n12111), .ZN(n12113) );
  AND2_X1 U15042 ( .A1(n12114), .A2(n12113), .ZN(n14319) );
  OAI22_X1 U15043 ( .A1(n14318), .A2(n12472), .B1(n9730), .B2(n12115), .ZN(
        n12118) );
  NAND2_X1 U15044 ( .A1(n13325), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n12117) );
  NAND2_X1 U15045 ( .A1(n12033), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12116) );
  NAND2_X1 U15046 ( .A1(n12117), .A2(n12116), .ZN(n12471) );
  OR2_X1 U15047 ( .A1(n13854), .A2(n11170), .ZN(n12128) );
  AND2_X1 U15048 ( .A1(n13637), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12129) );
  NAND2_X1 U15049 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21050) );
  NAND2_X1 U15050 ( .A1(n21050), .A2(n20852), .ZN(n12121) );
  NAND2_X1 U15051 ( .A1(n12129), .A2(n12121), .ZN(n12119) );
  INV_X1 U15052 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20969) );
  NAND2_X1 U15053 ( .A1(n12120), .A2(n20969), .ZN(n16262) );
  NAND2_X1 U15054 ( .A1(n11968), .A2(n16262), .ZN(n13292) );
  INV_X1 U15055 ( .A(n12121), .ZN(n12122) );
  NAND2_X1 U15056 ( .A1(n13292), .A2(n12122), .ZN(n12131) );
  INV_X1 U15057 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15085) );
  INV_X1 U15058 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21037) );
  INV_X1 U15059 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20987) );
  INV_X1 U15060 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20986) );
  INV_X1 U15061 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20392) );
  NOR4_X1 U15062 ( .A1(n21037), .A2(n20987), .A3(n20986), .A4(n20392), .ZN(
        n20262) );
  NAND4_X1 U15063 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n20263)
         );
  NAND2_X1 U15064 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14833) );
  NOR2_X1 U15065 ( .A1(n20263), .A2(n14833), .ZN(n14036) );
  INV_X1 U15066 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21001) );
  NAND2_X1 U15067 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14853) );
  NOR2_X1 U15068 ( .A1(n21001), .A2(n14853), .ZN(n14834) );
  NAND4_X1 U15069 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n20262), .A3(n14036), 
        .A4(n14834), .ZN(n14815) );
  NAND3_X1 U15070 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14732) );
  NOR2_X1 U15071 ( .A1(n14815), .A2(n14732), .ZN(n14784) );
  NAND3_X1 U15072 ( .A1(n14784), .A2(P1_REIP_REG_19__SCAN_IN), .A3(
        P1_REIP_REG_18__SCAN_IN), .ZN(n14763) );
  AND2_X1 U15073 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14752) );
  AND2_X1 U15074 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n14752), .ZN(n14735) );
  NAND2_X1 U15075 ( .A1(n14735), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n12123) );
  NOR2_X1 U15076 ( .A1(n14763), .A2(n12123), .ZN(n14705) );
  NAND2_X1 U15077 ( .A1(n14705), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14708) );
  NOR2_X1 U15078 ( .A1(n15085), .A2(n14708), .ZN(n14694) );
  NAND2_X1 U15079 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n14694), .ZN(n14682) );
  INV_X1 U15080 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21021) );
  NOR3_X1 U15081 ( .A1(n14817), .A2(n14682), .A3(n21021), .ZN(n14671) );
  NAND2_X1 U15082 ( .A1(n14671), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14322) );
  INV_X1 U15083 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21025) );
  INV_X1 U15084 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n15033) );
  OAI21_X1 U15085 ( .B1(n14322), .B2(n21025), .A(n15033), .ZN(n12127) );
  NAND2_X1 U15086 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n12477) );
  INV_X1 U15087 ( .A(n12477), .ZN(n12126) );
  INV_X1 U15088 ( .A(n20261), .ZN(n20332) );
  AOI21_X1 U15089 ( .B1(n20333), .B2(n14682), .A(n20332), .ZN(n14696) );
  NAND2_X1 U15090 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n12124) );
  NAND2_X1 U15091 ( .A1(n20333), .A2(n12124), .ZN(n12125) );
  AND2_X1 U15092 ( .A1(n14696), .A2(n12125), .ZN(n14672) );
  OAI21_X1 U15093 ( .B1(n12126), .B2(n14817), .A(n14672), .ZN(n12480) );
  NAND2_X1 U15094 ( .A1(n12127), .A2(n12480), .ZN(n12138) );
  INV_X1 U15095 ( .A(n12128), .ZN(n12133) );
  INV_X1 U15096 ( .A(n12129), .ZN(n12130) );
  AND2_X1 U15097 ( .A1(n12131), .A2(n12130), .ZN(n12132) );
  INV_X1 U15098 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n21239) );
  NOR2_X1 U15099 ( .A1(n15030), .A2(n20962), .ZN(n12134) );
  AOI22_X1 U15100 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n15036), .ZN(n12135) );
  OAI21_X1 U15101 ( .B1(n20308), .B2(n21239), .A(n12135), .ZN(n12136) );
  AOI22_X1 U15102 ( .A1(n12143), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12142), .ZN(n12144) );
  INV_X1 U15103 ( .A(n12146), .ZN(n13205) );
  NAND2_X1 U15104 ( .A1(n15412), .A2(n11170), .ZN(n12147) );
  NAND3_X1 U15105 ( .A1(n12148), .A2(n13205), .A3(n12147), .ZN(n13194) );
  NAND2_X1 U15106 ( .A1(n13107), .A2(n21050), .ZN(n12150) );
  OR2_X1 U15107 ( .A1(n12149), .A2(n12150), .ZN(n12151) );
  NAND2_X1 U15108 ( .A1(n11968), .A2(n21050), .ZN(n12153) );
  NOR2_X1 U15109 ( .A1(n12009), .A2(n12153), .ZN(n12154) );
  NAND2_X1 U15110 ( .A1(n12154), .A2(n13281), .ZN(n13195) );
  AND3_X1 U15111 ( .A1(n20457), .A2(n20446), .A3(n12155), .ZN(n13104) );
  INV_X1 U15112 ( .A(n20238), .ZN(n13290) );
  AND2_X1 U15113 ( .A1(n14988), .A2(n20457), .ZN(n12159) );
  NAND2_X1 U15114 ( .A1(n15026), .A2(n12159), .ZN(n12175) );
  NOR4_X1 U15115 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n12163) );
  NOR4_X1 U15116 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n12162) );
  NOR4_X1 U15117 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_6__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n12161) );
  NOR4_X1 U15118 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_11__SCAN_IN), .A3(P1_ADDRESS_REG_10__SCAN_IN), .A4(
        P1_ADDRESS_REG_9__SCAN_IN), .ZN(n12160) );
  AND4_X1 U15119 ( .A1(n12163), .A2(n12162), .A3(n12161), .A4(n12160), .ZN(
        n12168) );
  NOR4_X1 U15120 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_0__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12166) );
  NOR4_X1 U15121 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n12165) );
  NOR4_X1 U15122 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(
        P1_ADDRESS_REG_28__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n12164) );
  INV_X1 U15123 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20988) );
  AND4_X1 U15124 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n20988), .ZN(
        n12167) );
  NAND2_X1 U15125 ( .A1(n12168), .A2(n12167), .ZN(n12169) );
  AND2_X2 U15126 ( .A1(n12169), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20419)
         );
  AOI22_X1 U15127 ( .A1(n14970), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14991), .ZN(n12170) );
  INV_X1 U15128 ( .A(n12170), .ZN(n12173) );
  INV_X1 U15129 ( .A(n20419), .ZN(n20421) );
  INV_X1 U15130 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16701) );
  NOR2_X1 U15131 ( .A1(n12173), .A2(n12172), .ZN(n12174) );
  NAND2_X1 U15132 ( .A1(n12175), .A2(n12174), .ZN(P1_U2873) );
  NOR2_X2 U15133 ( .A1(n12177), .A2(n12178), .ZN(n12239) );
  AOI22_X1 U15134 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15135 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12189) );
  INV_X1 U15136 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14178) );
  NOR2_X2 U15137 ( .A1(n14265), .A2(n17175), .ZN(n17392) );
  INV_X2 U15138 ( .A(n17208), .ZN(n17353) );
  AOI22_X1 U15139 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12176) );
  OAI21_X1 U15140 ( .B1(n14178), .B2(n9665), .A(n12176), .ZN(n12187) );
  AOI22_X1 U15141 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12185) );
  INV_X2 U15142 ( .A(n9721), .ZN(n17319) );
  AOI22_X1 U15143 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15144 ( .A1(n17423), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15145 ( .A1(n17406), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12182) );
  NAND4_X1 U15146 ( .A1(n12185), .A2(n12184), .A3(n12183), .A4(n12182), .ZN(
        n12186) );
  AOI211_X1 U15147 ( .C1(n9673), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n12187), .B(n12186), .ZN(n12188) );
  NAND3_X1 U15148 ( .A1(n12190), .A2(n12189), .A3(n12188), .ZN(n16681) );
  AOI22_X1 U15149 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12249), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15150 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15151 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12193) );
  INV_X1 U15152 ( .A(n12191), .ZN(n12237) );
  AOI22_X1 U15153 ( .A1(n17440), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12192) );
  NAND4_X1 U15154 ( .A1(n12195), .A2(n12194), .A3(n12193), .A4(n12192), .ZN(
        n12201) );
  AOI22_X1 U15155 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15156 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15157 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15158 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12196) );
  NAND4_X1 U15159 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12196), .ZN(
        n12200) );
  AOI22_X1 U15160 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15161 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15162 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15163 ( .A1(n17406), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12202) );
  NAND4_X1 U15164 ( .A1(n12205), .A2(n12204), .A3(n12203), .A4(n12202), .ZN(
        n12211) );
  AOI22_X1 U15165 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15166 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12249), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15167 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17440), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15168 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12206) );
  NAND4_X1 U15169 ( .A1(n12209), .A2(n12208), .A3(n12207), .A4(n12206), .ZN(
        n12210) );
  AOI22_X1 U15170 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17440), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15171 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14166), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15172 ( .A1(n12239), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12249), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15173 ( .A1(n17392), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12191), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15174 ( .A1(n12266), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12335), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15175 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12217) );
  INV_X1 U15176 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18482) );
  INV_X1 U15177 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12220) );
  INV_X1 U15178 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12219) );
  INV_X1 U15179 ( .A(n12221), .ZN(n12222) );
  OAI21_X1 U15180 ( .B1(n9721), .B2(n18482), .A(n12222), .ZN(n12223) );
  INV_X1 U15181 ( .A(n12223), .ZN(n12224) );
  AOI22_X1 U15182 ( .A1(n12307), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12249), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15183 ( .A1(n9688), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17440), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15184 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15185 ( .A1(n12239), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12191), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12226) );
  INV_X1 U15186 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18488) );
  AOI22_X1 U15187 ( .A1(n14166), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12335), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12230) );
  OAI21_X1 U15188 ( .B1(n9721), .B2(n18488), .A(n12230), .ZN(n12231) );
  INV_X4 U15189 ( .A(n17148), .ZN(n17441) );
  AOI22_X1 U15190 ( .A1(n17441), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15191 ( .A1(n12266), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12232) );
  INV_X1 U15192 ( .A(n12232), .ZN(n12233) );
  AOI21_X1 U15193 ( .B1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B2(n17196), .A(
        n12233), .ZN(n12234) );
  NAND4_X1 U15194 ( .A1(n10171), .A2(n12236), .A3(n12235), .A4(n12234), .ZN(
        n17628) );
  NAND2_X1 U15195 ( .A1(n17634), .A2(n17628), .ZN(n12277) );
  AOI22_X1 U15196 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15197 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17428), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15198 ( .A1(n17440), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12238) );
  OAI21_X1 U15199 ( .B1(n9721), .B2(n18500), .A(n12238), .ZN(n12245) );
  AOI22_X1 U15200 ( .A1(n17392), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15201 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15202 ( .A1(n12239), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12249), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15203 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12240) );
  NAND4_X1 U15204 ( .A1(n12243), .A2(n12242), .A3(n12241), .A4(n12240), .ZN(
        n12244) );
  AOI211_X1 U15205 ( .C1(n9687), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n12245), .B(n12244), .ZN(n12246) );
  NAND3_X1 U15206 ( .A1(n12248), .A2(n12247), .A3(n12246), .ZN(n17618) );
  NAND2_X1 U15207 ( .A1(n12261), .A2(n17618), .ZN(n12281) );
  AOI22_X1 U15208 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17440), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15209 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12258) );
  INV_X1 U15210 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18513) );
  AOI22_X1 U15211 ( .A1(n17406), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12250) );
  OAI21_X1 U15212 ( .B1(n9721), .B2(n18513), .A(n12250), .ZN(n12256) );
  AOI22_X1 U15213 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U15214 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9687), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15215 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15216 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12251) );
  NAND4_X1 U15217 ( .A1(n12254), .A2(n12253), .A3(n12252), .A4(n12251), .ZN(
        n12255) );
  AOI211_X1 U15218 ( .C1(n17348), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12256), .B(n12255), .ZN(n12257) );
  NAND3_X1 U15219 ( .A1(n12259), .A2(n12258), .A3(n12257), .ZN(n17609) );
  INV_X1 U15220 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21233) );
  XOR2_X1 U15221 ( .A(n12260), .B(n17609), .Z(n12285) );
  XOR2_X1 U15222 ( .A(n12261), .B(n17618), .Z(n12279) );
  XNOR2_X1 U15223 ( .A(n17628), .B(n17634), .ZN(n12275) );
  INV_X1 U15224 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19073) );
  NOR2_X1 U15225 ( .A1(n17634), .A2(n19073), .ZN(n12273) );
  AOI22_X1 U15226 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15227 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15228 ( .A1(n12239), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12265), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15229 ( .A1(n12249), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17440), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15230 ( .A1(n12307), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15231 ( .A1(n12266), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14166), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12267) );
  NAND2_X1 U15232 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18124), .ZN(
        n18123) );
  NOR2_X1 U15233 ( .A1(n12273), .A2(n18116), .ZN(n18108) );
  XNOR2_X1 U15234 ( .A(n12275), .B(n12274), .ZN(n18107) );
  INV_X1 U15235 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18412) );
  NOR2_X1 U15236 ( .A1(n12276), .A2(n18412), .ZN(n12278) );
  XNOR2_X1 U15237 ( .A(n12277), .B(n17623), .ZN(n18095) );
  INV_X1 U15238 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18403) );
  XOR2_X1 U15239 ( .A(n18403), .B(n12279), .Z(n18088) );
  NOR2_X1 U15240 ( .A1(n18089), .A2(n18088), .ZN(n18087) );
  XNOR2_X1 U15241 ( .A(n12281), .B(n17613), .ZN(n12283) );
  NOR2_X1 U15242 ( .A1(n12282), .A2(n12283), .ZN(n12284) );
  INV_X1 U15243 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18072) );
  INV_X1 U15244 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21195) );
  XOR2_X1 U15245 ( .A(n21195), .B(n12285), .Z(n18059) );
  OAI21_X1 U15246 ( .B1(n12286), .B2(n16681), .A(n17933), .ZN(n12288) );
  NOR2_X1 U15247 ( .A1(n12287), .A2(n12288), .ZN(n12289) );
  INV_X1 U15248 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18378) );
  INV_X1 U15249 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18360) );
  INV_X1 U15250 ( .A(n12290), .ZN(n12292) );
  NAND2_X1 U15251 ( .A1(n18037), .A2(n12290), .ZN(n17935) );
  NAND2_X1 U15252 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18329) );
  INV_X1 U15253 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17991) );
  NOR2_X1 U15254 ( .A1(n18329), .A2(n17991), .ZN(n18300) );
  NAND2_X1 U15255 ( .A1(n18300), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18283) );
  INV_X1 U15256 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18286) );
  NOR2_X1 U15257 ( .A1(n18283), .A2(n18286), .ZN(n18285) );
  NAND2_X1 U15258 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18285), .ZN(
        n18267) );
  INV_X1 U15259 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18274) );
  NOR2_X1 U15260 ( .A1(n18267), .A2(n18274), .ZN(n18237) );
  INV_X1 U15261 ( .A(n18237), .ZN(n16189) );
  NOR2_X1 U15262 ( .A1(n17935), .A2(n16189), .ZN(n12295) );
  INV_X1 U15263 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18343) );
  INV_X1 U15264 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18339) );
  NAND2_X1 U15265 ( .A1(n18343), .A2(n18339), .ZN(n18005) );
  INV_X1 U15266 ( .A(n18005), .ZN(n17988) );
  NOR4_X1 U15267 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12291) );
  NAND4_X1 U15268 ( .A1(n12292), .A2(n17988), .A3(n12291), .A4(n18274), .ZN(
        n12293) );
  NAND2_X1 U15269 ( .A1(n17933), .A2(n12293), .ZN(n12294) );
  OAI221_X1 U15270 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17933), 
        .C1(n21233), .C2(n12295), .A(n12294), .ZN(n17901) );
  NOR2_X1 U15271 ( .A1(n17901), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17900) );
  INV_X1 U15272 ( .A(n12294), .ZN(n12296) );
  NAND2_X1 U15273 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18242) );
  INV_X1 U15274 ( .A(n18242), .ZN(n17893) );
  NAND2_X1 U15275 ( .A1(n17893), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18204) );
  INV_X1 U15276 ( .A(n18204), .ZN(n17868) );
  INV_X1 U15277 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18208) );
  NAND2_X1 U15278 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18207) );
  NOR2_X1 U15279 ( .A1(n18208), .A2(n18207), .ZN(n18184) );
  NAND2_X1 U15280 ( .A1(n17868), .A2(n18184), .ZN(n18190) );
  INV_X1 U15281 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18195) );
  NOR2_X1 U15282 ( .A1(n18190), .A2(n18195), .ZN(n18178) );
  NAND2_X1 U15283 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18178), .ZN(
        n17806) );
  INV_X1 U15284 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17895) );
  NAND2_X1 U15285 ( .A1(n17933), .A2(n17895), .ZN(n17894) );
  NOR2_X1 U15286 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17894), .ZN(
        n12297) );
  INV_X1 U15287 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18225) );
  NAND2_X1 U15288 ( .A1(n12297), .A2(n18225), .ZN(n17853) );
  NOR2_X1 U15289 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17853), .ZN(
        n17835) );
  INV_X1 U15290 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18171) );
  NAND3_X1 U15291 ( .A1(n17835), .A2(n18171), .A3(n18195), .ZN(n12298) );
  INV_X1 U15292 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17814) );
  INV_X1 U15293 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18155) );
  NOR2_X1 U15294 ( .A1(n17914), .A2(n18242), .ZN(n17851) );
  NOR2_X1 U15295 ( .A1(n17819), .A2(n17851), .ZN(n17852) );
  NAND2_X1 U15296 ( .A1(n18184), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16190) );
  NOR3_X2 U15297 ( .A1(n17852), .A2(n17895), .A3(n16190), .ZN(n17818) );
  NAND3_X1 U15298 ( .A1(n17818), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17813), .ZN(n12302) );
  NAND2_X1 U15299 ( .A1(n12302), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12300) );
  INV_X1 U15300 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17787) );
  NAND2_X1 U15301 ( .A1(n18038), .A2(n12302), .ZN(n17800) );
  NAND2_X1 U15302 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16203) );
  INV_X1 U15303 ( .A(n16203), .ZN(n18135) );
  INV_X1 U15304 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18140) );
  INV_X1 U15305 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17755) );
  NAND2_X1 U15306 ( .A1(n9705), .A2(n18038), .ZN(n16686) );
  NAND2_X1 U15307 ( .A1(n17755), .A2(n18038), .ZN(n16683) );
  INV_X1 U15308 ( .A(n16683), .ZN(n12304) );
  INV_X1 U15309 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16628) );
  AOI22_X1 U15310 ( .A1(n17392), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12311) );
  CLKBUF_X3 U15311 ( .A(n12307), .Z(n17428) );
  AOI22_X1 U15312 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15313 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15314 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12308) );
  NAND4_X1 U15315 ( .A1(n12311), .A2(n12310), .A3(n12309), .A4(n12308), .ZN(
        n12317) );
  AOI22_X1 U15316 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U15317 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12314) );
  BUF_X4 U15318 ( .A(n9658), .Z(n17422) );
  AOI22_X1 U15319 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15320 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17440), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12312) );
  NAND4_X1 U15321 ( .A1(n12315), .A2(n12314), .A3(n12313), .A4(n12312), .ZN(
        n12316) );
  NAND2_X1 U15322 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19075), .ZN(n18970) );
  NAND2_X1 U15323 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18940), .ZN(
        n12326) );
  AOI22_X1 U15324 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18947), .B2(n12320), .ZN(
        n12322) );
  XOR2_X1 U15325 ( .A(n12321), .B(n12322), .Z(n12334) );
  OAI22_X1 U15326 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18951), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12324), .ZN(n12329) );
  NOR2_X1 U15327 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18951), .ZN(
        n12325) );
  NAND2_X1 U15328 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12324), .ZN(
        n12328) );
  AOI22_X1 U15329 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12329), .B1(
        n12325), .B2(n12328), .ZN(n12327) );
  OAI211_X1 U15330 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18940), .A(
        n12327), .B(n12326), .ZN(n12428) );
  INV_X1 U15331 ( .A(n12428), .ZN(n12333) );
  XNOR2_X1 U15332 ( .A(n12326), .B(n12429), .ZN(n12332) );
  NAND2_X1 U15333 ( .A1(n12327), .A2(n12334), .ZN(n12426) );
  AND2_X1 U15334 ( .A1(n12328), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12330) );
  OAI22_X1 U15335 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18916), .B1(
        n12330), .B2(n12329), .ZN(n12331) );
  INV_X1 U15336 ( .A(n12331), .ZN(n12427) );
  AOI21_X1 U15337 ( .B1(n12334), .B2(n12333), .A(n16786), .ZN(n18911) );
  INV_X1 U15338 ( .A(n18911), .ZN(n12430) );
  AOI22_X1 U15339 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15340 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15341 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U15342 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12336) );
  NAND4_X1 U15343 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12345) );
  AOI22_X1 U15344 ( .A1(n17440), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U15345 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U15346 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U15347 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12340) );
  NAND4_X1 U15348 ( .A1(n12343), .A2(n12342), .A3(n12341), .A4(n12340), .ZN(
        n12344) );
  AOI22_X1 U15349 ( .A1(n17440), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15350 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12348) );
  AOI22_X1 U15351 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15352 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17428), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12346) );
  NAND4_X1 U15353 ( .A1(n12349), .A2(n12348), .A3(n12347), .A4(n12346), .ZN(
        n12355) );
  AOI22_X1 U15354 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15355 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15356 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15357 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14205), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12350) );
  NAND4_X1 U15358 ( .A1(n12353), .A2(n12352), .A3(n12351), .A4(n12350), .ZN(
        n12354) );
  AOI22_X1 U15359 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15360 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17411), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17440), .ZN(n12358) );
  AOI22_X1 U15361 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n16181), .ZN(n12357) );
  AOI22_X1 U15362 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17406), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17382), .ZN(n12356) );
  NAND4_X1 U15363 ( .A1(n12359), .A2(n12358), .A3(n12357), .A4(n12356), .ZN(
        n12365) );
  AOI22_X1 U15364 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17423), .ZN(n12363) );
  AOI22_X1 U15365 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12249), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15366 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17441), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15367 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17392), .B1(
        n9687), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12360) );
  NAND4_X1 U15368 ( .A1(n12363), .A2(n12362), .A3(n12361), .A4(n12360), .ZN(
        n12364) );
  AOI22_X1 U15369 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15370 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12373) );
  AOI22_X1 U15371 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12366) );
  OAI21_X1 U15372 ( .B1(n12367), .B2(n18478), .A(n12366), .ZN(n12372) );
  AOI22_X1 U15373 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15374 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12249), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15375 ( .A1(n17440), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U15376 ( .A1(n17406), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U15377 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U15378 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17440), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U15379 ( .A1(n17406), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15380 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12375) );
  NAND4_X1 U15381 ( .A1(n12378), .A2(n12377), .A3(n12376), .A4(n12375), .ZN(
        n12384) );
  AOI22_X1 U15382 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15383 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15384 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14205), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15385 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12379) );
  NAND4_X1 U15386 ( .A1(n12382), .A2(n12381), .A3(n12380), .A4(n12379), .ZN(
        n12383) );
  AOI22_X1 U15387 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U15388 ( .A1(n17440), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15389 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15390 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12385) );
  NAND4_X1 U15391 ( .A1(n12388), .A2(n12387), .A3(n12386), .A4(n12385), .ZN(
        n12394) );
  AOI22_X1 U15392 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12392) );
  AOI22_X1 U15393 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12391) );
  AOI22_X1 U15394 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12390) );
  AOI22_X1 U15395 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12389) );
  NAND4_X1 U15396 ( .A1(n12392), .A2(n12391), .A3(n12390), .A4(n12389), .ZN(
        n12393) );
  NOR2_X1 U15397 ( .A1(n18510), .A2(n18503), .ZN(n12407) );
  AOI22_X1 U15398 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15399 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U15400 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12249), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12396) );
  AOI22_X1 U15401 ( .A1(n17406), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12395) );
  NAND4_X1 U15402 ( .A1(n12398), .A2(n12397), .A3(n12396), .A4(n12395), .ZN(
        n12404) );
  AOI22_X1 U15403 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U15404 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15405 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U15406 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17440), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12399) );
  NAND4_X1 U15407 ( .A1(n12402), .A2(n12401), .A3(n12400), .A4(n12399), .ZN(
        n12403) );
  NAND2_X1 U15408 ( .A1(n18485), .A2(n17495), .ZN(n16200) );
  INV_X1 U15409 ( .A(n18497), .ZN(n14132) );
  NAND2_X1 U15410 ( .A1(n18510), .A2(n14132), .ZN(n18919) );
  INV_X1 U15411 ( .A(n18510), .ZN(n16194) );
  NAND2_X1 U15412 ( .A1(n18503), .A2(n16194), .ZN(n12415) );
  NAND3_X1 U15413 ( .A1(n18485), .A2(n18919), .A3(n12415), .ZN(n12405) );
  NOR2_X1 U15414 ( .A1(n18475), .A2(n16828), .ZN(n12420) );
  OAI21_X1 U15415 ( .B1(n18518), .B2(n18936), .A(n12420), .ZN(n14256) );
  INV_X1 U15416 ( .A(n12405), .ZN(n12414) );
  NOR2_X1 U15417 ( .A1(n17642), .A2(n19112), .ZN(n12421) );
  INV_X1 U15418 ( .A(n12421), .ZN(n12406) );
  AOI21_X1 U15419 ( .B1(n18485), .B2(n12406), .A(n12407), .ZN(n12413) );
  NOR2_X1 U15420 ( .A1(n18518), .A2(n12407), .ZN(n12411) );
  NAND2_X1 U15421 ( .A1(n18497), .A2(n18936), .ZN(n12409) );
  OAI211_X1 U15422 ( .C1(n18497), .C2(n12411), .A(n12410), .B(n12409), .ZN(
        n12412) );
  OAI211_X1 U15423 ( .C1(n18491), .C2(n12417), .A(n14256), .B(n9655), .ZN(
        n12424) );
  NAND2_X1 U15424 ( .A1(n18485), .A2(n18491), .ZN(n18918) );
  NAND3_X1 U15425 ( .A1(n12416), .A2(n14134), .A3(n19112), .ZN(n12419) );
  NOR2_X2 U15426 ( .A1(n14249), .A2(n14250), .ZN(n18937) );
  NOR2_X1 U15427 ( .A1(n12421), .A2(n12420), .ZN(n19125) );
  NOR2_X2 U15428 ( .A1(n18919), .A2(n14255), .ZN(n14259) );
  INV_X1 U15429 ( .A(n12422), .ZN(n16821) );
  NOR3_X1 U15430 ( .A1(n12423), .A2(n19112), .A3(n16821), .ZN(n12425) );
  XNOR2_X1 U15431 ( .A(n16828), .B(n18485), .ZN(n16193) );
  OAI211_X1 U15432 ( .C1(n12429), .C2(n12428), .A(n12427), .B(n12426), .ZN(
        n16198) );
  NAND2_X1 U15433 ( .A1(n9726), .A2(n18039), .ZN(n12468) );
  NOR2_X1 U15434 ( .A1(n18140), .A2(n17755), .ZN(n16252) );
  NOR2_X1 U15435 ( .A1(n12306), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16251) );
  NOR2_X1 U15436 ( .A1(n18171), .A2(n17814), .ZN(n18133) );
  NAND3_X1 U15437 ( .A1(n18178), .A2(n18135), .A3(n18133), .ZN(n16680) );
  AND2_X1 U15438 ( .A1(n17634), .A2(n18124), .ZN(n12438) );
  NOR2_X1 U15439 ( .A1(n12438), .A2(n17628), .ZN(n12436) );
  NOR2_X1 U15440 ( .A1(n17623), .A2(n12436), .ZN(n12435) );
  NAND2_X1 U15441 ( .A1(n12435), .A2(n17618), .ZN(n12433) );
  NOR2_X1 U15442 ( .A1(n17613), .A2(n12433), .ZN(n12432) );
  NAND2_X1 U15443 ( .A1(n12432), .A2(n17609), .ZN(n12431) );
  NOR2_X1 U15444 ( .A1(n17605), .A2(n12431), .ZN(n12453) );
  XOR2_X1 U15445 ( .A(n17605), .B(n12431), .Z(n18043) );
  XOR2_X1 U15446 ( .A(n17609), .B(n12432), .Z(n12446) );
  XOR2_X1 U15447 ( .A(n17613), .B(n12433), .Z(n12434) );
  NAND2_X1 U15448 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12434), .ZN(
        n12445) );
  XOR2_X1 U15449 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12434), .Z(
        n18069) );
  XOR2_X1 U15450 ( .A(n17618), .B(n12435), .Z(n18083) );
  XOR2_X1 U15451 ( .A(n17623), .B(n12436), .Z(n12437) );
  NAND2_X1 U15452 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12437), .ZN(
        n12443) );
  XOR2_X1 U15453 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n12437), .Z(
        n18099) );
  XOR2_X1 U15454 ( .A(n17628), .B(n12438), .Z(n12439) );
  OR2_X1 U15455 ( .A1(n12274), .A2(n12439), .ZN(n12442) );
  XOR2_X1 U15456 ( .A(n12274), .B(n12439), .Z(n18431) );
  AOI21_X1 U15457 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17634), .A(
        n18124), .ZN(n12441) );
  INV_X1 U15458 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19091) );
  NOR2_X1 U15459 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17634), .ZN(
        n12440) );
  AOI221_X1 U15460 ( .B1(n18124), .B2(n17634), .C1(n12441), .C2(n19091), .A(
        n12440), .ZN(n18430) );
  NAND2_X1 U15461 ( .A1(n18431), .A2(n18430), .ZN(n18429) );
  NAND2_X1 U15462 ( .A1(n12442), .A2(n18429), .ZN(n18098) );
  NAND2_X1 U15463 ( .A1(n18099), .A2(n18098), .ZN(n18097) );
  NAND2_X1 U15464 ( .A1(n12443), .A2(n18097), .ZN(n18082) );
  NAND2_X1 U15465 ( .A1(n18083), .A2(n18082), .ZN(n12444) );
  NOR2_X1 U15466 ( .A1(n18083), .A2(n18082), .ZN(n18081) );
  AOI21_X1 U15467 ( .B1(n18403), .B2(n12444), .A(n18081), .ZN(n18068) );
  NAND2_X1 U15468 ( .A1(n18069), .A2(n18068), .ZN(n18067) );
  NAND2_X1 U15469 ( .A1(n12445), .A2(n18067), .ZN(n12447) );
  NAND2_X1 U15470 ( .A1(n12446), .A2(n12447), .ZN(n12448) );
  XOR2_X1 U15471 ( .A(n12447), .B(n12446), .Z(n18056) );
  NAND2_X1 U15472 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18056), .ZN(
        n18055) );
  NAND2_X1 U15473 ( .A1(n12448), .A2(n18055), .ZN(n18044) );
  NOR2_X1 U15474 ( .A1(n18043), .A2(n18044), .ZN(n12449) );
  NOR2_X1 U15475 ( .A1(n12449), .A2(n18378), .ZN(n12450) );
  NAND2_X1 U15476 ( .A1(n12453), .A2(n12450), .ZN(n12454) );
  INV_X1 U15477 ( .A(n12450), .ZN(n12452) );
  NAND2_X1 U15478 ( .A1(n18043), .A2(n18044), .ZN(n18042) );
  NAND2_X1 U15479 ( .A1(n12453), .A2(n12452), .ZN(n12451) );
  OAI211_X1 U15480 ( .C1(n12453), .C2(n12452), .A(n18042), .B(n12451), .ZN(
        n18026) );
  NAND2_X1 U15481 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18026), .ZN(
        n18025) );
  NAND2_X1 U15482 ( .A1(n12455), .A2(n17933), .ZN(n17934) );
  NOR2_X1 U15483 ( .A1(n16680), .A2(n17927), .ZN(n17777) );
  NAND3_X1 U15484 ( .A1(n16252), .A2(n16251), .A3(n17777), .ZN(n12467) );
  INV_X1 U15485 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16844) );
  INV_X1 U15486 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16862) );
  INV_X1 U15487 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n21234) );
  INV_X1 U15488 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17863) );
  NAND2_X1 U15489 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17795) );
  INV_X1 U15490 ( .A(n12458), .ZN(n17783) );
  NOR2_X1 U15491 ( .A1(n21234), .A2(n17783), .ZN(n17772) );
  NAND3_X1 U15492 ( .A1(n17772), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16651) );
  NOR2_X1 U15493 ( .A1(n16862), .A2(n16651), .ZN(n12459) );
  INV_X1 U15494 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n21075) );
  NAND2_X1 U15495 ( .A1(n21075), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18126) );
  NAND2_X1 U15496 ( .A1(n19075), .A2(n19068), .ZN(n19078) );
  NAND2_X1 U15497 ( .A1(n19123), .A2(n19068), .ZN(n16789) );
  AND2_X1 U15498 ( .A1(n19078), .A2(n16789), .ZN(n19106) );
  NAND2_X1 U15499 ( .A1(n18916), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19077) );
  OAI221_X1 U15500 ( .B1(n19123), .B2(P3_STATE2_REG_1__SCAN_IN), .C1(
        P3_STATE2_REG_2__SCAN_IN), .C2(n19075), .A(n19077), .ZN(n18473) );
  NAND3_X1 U15501 ( .A1(n19123), .A2(n19068), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18823) );
  NOR2_X2 U15502 ( .A1(n18597), .A2(n18823), .ZN(n18854) );
  AOI21_X1 U15503 ( .B1(n17841), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n18854), .ZN(n17880) );
  NAND2_X1 U15504 ( .A1(n12459), .A2(n17976), .ZN(n16641) );
  INV_X1 U15505 ( .A(n17841), .ZN(n17781) );
  NOR2_X1 U15506 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17781), .ZN(
        n16661) );
  NOR2_X1 U15507 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16641), .ZN(
        n12462) );
  INV_X1 U15508 ( .A(n18126), .ZN(n17839) );
  INV_X2 U15509 ( .A(n18854), .ZN(n18507) );
  OAI21_X1 U15510 ( .B1(n18507), .B2(n12459), .A(n18125), .ZN(n12460) );
  AOI21_X1 U15511 ( .B1(n16810), .B2(n17839), .A(n12460), .ZN(n12461) );
  INV_X1 U15512 ( .A(n12461), .ZN(n16653) );
  NOR3_X1 U15513 ( .A1(n16661), .A2(n12462), .A3(n16653), .ZN(n16642) );
  AOI21_X1 U15514 ( .B1(n16844), .B2(n16641), .A(n16642), .ZN(n12464) );
  INV_X1 U15515 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19111) );
  NOR2_X1 U15516 ( .A1(n19075), .A2(n19111), .ZN(n18080) );
  NAND2_X1 U15517 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16660), .ZN(
        n16640) );
  OAI21_X1 U15518 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16660), .A(
        n16640), .ZN(n16841) );
  OR3_X2 U15519 ( .A1(n19078), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18384) );
  INV_X2 U15520 ( .A(n18384), .ZN(n18385) );
  NAND2_X1 U15521 ( .A1(n18385), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16256) );
  OAI21_X1 U15522 ( .B1(n17965), .B2(n16841), .A(n16256), .ZN(n12463) );
  NAND2_X1 U15523 ( .A1(n17828), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17799) );
  NAND2_X1 U15524 ( .A1(n18139), .A2(n16252), .ZN(n16655) );
  INV_X1 U15525 ( .A(n16655), .ZN(n16688) );
  NAND2_X1 U15526 ( .A1(n16688), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16646) );
  NAND2_X1 U15527 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18170), .ZN(
        n17792) );
  NAND2_X1 U15528 ( .A1(n16252), .A2(n18131), .ZN(n16691) );
  NOR2_X1 U15529 ( .A1(n12306), .A2(n16691), .ZN(n16656) );
  INV_X1 U15530 ( .A(n16656), .ZN(n16207) );
  AOI22_X1 U15531 ( .A1(n9802), .A2(n16646), .B1(n18115), .B2(n16207), .ZN(
        n12465) );
  NAND2_X1 U15532 ( .A1(n15026), .A2(n20317), .ZN(n12484) );
  NAND2_X1 U15533 ( .A1(n13325), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12470) );
  NAND2_X1 U15534 ( .A1(n12033), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12469) );
  NAND2_X1 U15535 ( .A1(n12470), .A2(n12469), .ZN(n12473) );
  XNOR2_X1 U15536 ( .A(n12473), .B(n12471), .ZN(n12476) );
  NAND2_X1 U15537 ( .A1(n12473), .A2(n12472), .ZN(n12475) );
  INV_X1 U15538 ( .A(n14318), .ZN(n12474) );
  MUX2_X1 U15539 ( .A(n12476), .B(n12475), .S(n12474), .Z(n15231) );
  INV_X1 U15540 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14857) );
  INV_X1 U15541 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15028) );
  OAI22_X1 U15542 ( .A1(n20308), .A2(n14857), .B1(n15028), .B2(n20279), .ZN(
        n12479) );
  NOR3_X1 U15543 ( .A1(n14322), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n12477), 
        .ZN(n12478) );
  AOI211_X1 U15544 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n12480), .A(n12479), 
        .B(n12478), .ZN(n12481) );
  NAND2_X1 U15545 ( .A1(n12484), .A2(n12483), .ZN(P1_U2809) );
  INV_X1 U15546 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14285) );
  AND2_X1 U15547 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n12504), .ZN(
        n12506) );
  OAI21_X1 U15548 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12506), .A(
        n12487), .ZN(n15794) );
  INV_X1 U15549 ( .A(n15794), .ZN(n19176) );
  AOI21_X1 U15550 ( .B1(n15817), .B2(n9707), .A(n12488), .ZN(n19222) );
  AOI21_X1 U15551 ( .B1(n15840), .B2(n12489), .A(n12490), .ZN(n12814) );
  INV_X1 U15552 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15854) );
  NAND2_X1 U15553 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n12491), .ZN(
        n12503) );
  AOI21_X1 U15554 ( .B1(n15854), .B2(n12503), .A(n12492), .ZN(n19246) );
  AOI21_X1 U15555 ( .B1(n15864), .B2(n12493), .A(n12491), .ZN(n13729) );
  AOI21_X1 U15556 ( .B1(n19262), .B2(n12494), .A(n12495), .ZN(n19268) );
  NAND2_X1 U15557 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n12496), .ZN(
        n12502) );
  AOI21_X1 U15558 ( .B1(n10727), .B2(n12502), .A(n12497), .ZN(n19274) );
  AOI21_X1 U15559 ( .B1(n10719), .B2(n12498), .A(n12496), .ZN(n19306) );
  AOI21_X1 U15560 ( .B1(n12501), .B2(n12499), .A(n12500), .ZN(n13611) );
  INV_X1 U15561 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14338) );
  AND2_X1 U15562 ( .A1(n19332), .A2(n13720), .ZN(n13677) );
  OAI21_X1 U15563 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12499), .ZN(n14648) );
  NAND2_X1 U15564 ( .A1(n13677), .A2(n14648), .ZN(n13451) );
  NOR2_X1 U15565 ( .A1(n13611), .A2(n13451), .ZN(n13549) );
  OAI21_X1 U15566 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12500), .A(
        n12498), .ZN(n19495) );
  NAND2_X1 U15567 ( .A1(n13549), .A2(n19495), .ZN(n19304) );
  NOR2_X1 U15568 ( .A1(n19306), .A2(n19304), .ZN(n19288) );
  OAI21_X1 U15569 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12496), .A(
        n12502), .ZN(n19291) );
  NAND2_X1 U15570 ( .A1(n19288), .A2(n19291), .ZN(n19273) );
  NOR2_X1 U15571 ( .A1(n19274), .A2(n19273), .ZN(n13596) );
  OAI21_X1 U15572 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12497), .A(
        n12494), .ZN(n16525) );
  NAND2_X1 U15573 ( .A1(n13596), .A2(n16525), .ZN(n19266) );
  NOR2_X1 U15574 ( .A1(n19268), .A2(n19266), .ZN(n15512) );
  OAI21_X1 U15575 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12495), .A(
        n12493), .ZN(n16514) );
  NAND2_X1 U15576 ( .A1(n15512), .A2(n16514), .ZN(n13726) );
  NOR2_X1 U15577 ( .A1(n13729), .A2(n13726), .ZN(n13725) );
  OAI21_X1 U15578 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12491), .A(
        n12503), .ZN(n19251) );
  NAND2_X1 U15579 ( .A1(n13725), .A2(n19251), .ZN(n19238) );
  NOR2_X1 U15580 ( .A1(n19246), .A2(n19238), .ZN(n19237) );
  OAI21_X1 U15581 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12492), .A(
        n12489), .ZN(n19225) );
  NAND2_X1 U15582 ( .A1(n19237), .A2(n19225), .ZN(n12812) );
  NOR2_X1 U15583 ( .A1(n12814), .A2(n12812), .ZN(n15498) );
  OAI21_X1 U15584 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12490), .A(
        n9707), .ZN(n15828) );
  NAND2_X1 U15585 ( .A1(n15498), .A2(n15828), .ZN(n19216) );
  NOR2_X1 U15586 ( .A1(n19222), .A2(n19216), .ZN(n19215) );
  OAI21_X1 U15587 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12488), .A(
        n12507), .ZN(n16496) );
  INV_X1 U15588 ( .A(n16496), .ZN(n19200) );
  INV_X1 U15589 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19187) );
  AOI21_X1 U15590 ( .B1(n19187), .B2(n12507), .A(n12506), .ZN(n19186) );
  NOR2_X1 U15591 ( .A1(n19176), .A2(n19175), .ZN(n19174) );
  NOR2_X1 U15592 ( .A1(n19289), .A2(n19174), .ZN(n19157) );
  NOR2_X1 U15593 ( .A1(n10763), .A2(n12487), .ZN(n12508) );
  AOI21_X1 U15594 ( .B1(n10763), .B2(n12487), .A(n12508), .ZN(n19159) );
  NOR2_X1 U15595 ( .A1(n19157), .A2(n19159), .ZN(n19158) );
  NOR2_X1 U15596 ( .A1(n19289), .A2(n19158), .ZN(n15491) );
  OAI21_X1 U15597 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12508), .A(
        n9778), .ZN(n16491) );
  INV_X1 U15598 ( .A(n16491), .ZN(n15493) );
  NOR2_X1 U15599 ( .A1(n15491), .A2(n15493), .ZN(n15492) );
  NOR2_X1 U15600 ( .A1(n19289), .A2(n15492), .ZN(n15466) );
  AOI21_X1 U15601 ( .B1(n15754), .B2(n9778), .A(n12509), .ZN(n15756) );
  NOR2_X1 U15602 ( .A1(n15467), .A2(n19289), .ZN(n16471) );
  OAI21_X1 U15603 ( .B1(n12509), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n9785), .ZN(n15747) );
  INV_X1 U15604 ( .A(n15747), .ZN(n16472) );
  NOR2_X1 U15605 ( .A1(n16471), .A2(n16472), .ZN(n16470) );
  NOR2_X1 U15606 ( .A1(n19289), .A2(n16470), .ZN(n15460) );
  AOI21_X1 U15607 ( .B1(n15736), .B2(n9785), .A(n12510), .ZN(n15739) );
  NOR2_X2 U15608 ( .A1(n15460), .A2(n15739), .ZN(n15459) );
  NOR2_X1 U15609 ( .A1(n19289), .A2(n15459), .ZN(n16449) );
  OAI21_X1 U15610 ( .B1(n12510), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n12511), .ZN(n15722) );
  INV_X1 U15611 ( .A(n15722), .ZN(n16451) );
  NOR2_X1 U15612 ( .A1(n16449), .A2(n16451), .ZN(n16450) );
  NOR2_X1 U15613 ( .A1(n19289), .A2(n16450), .ZN(n12824) );
  AND2_X1 U15614 ( .A1(n12511), .A2(n15714), .ZN(n12512) );
  NOR2_X1 U15615 ( .A1(n12513), .A2(n12512), .ZN(n15716) );
  NOR2_X1 U15616 ( .A1(n12824), .A2(n15716), .ZN(n12825) );
  NOR2_X1 U15617 ( .A1(n19289), .A2(n12825), .ZN(n15441) );
  OR2_X1 U15618 ( .A1(n12513), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12514) );
  AND2_X1 U15619 ( .A1(n12514), .A2(n9789), .ZN(n15704) );
  NOR2_X1 U15620 ( .A1(n15441), .A2(n15704), .ZN(n15440) );
  NOR2_X1 U15621 ( .A1(n19289), .A2(n15440), .ZN(n16435) );
  NOR2_X1 U15622 ( .A1(n16435), .A2(n16434), .ZN(n15427) );
  NOR2_X1 U15623 ( .A1(n19289), .A2(n15427), .ZN(n12516) );
  INV_X1 U15624 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15693) );
  XNOR2_X1 U15625 ( .A(n12515), .B(n15693), .ZN(n15692) );
  XNOR2_X1 U15626 ( .A(n12516), .B(n15692), .ZN(n12517) );
  INV_X1 U15627 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19953) );
  INV_X1 U15628 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20228) );
  NAND4_X1 U15629 ( .A1(n19953), .A2(n16267), .A3(n20228), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20099) );
  INV_X1 U15630 ( .A(n20099), .ZN(n19308) );
  NAND2_X1 U15631 ( .A1(n12517), .A2(n19308), .ZN(n12797) );
  NAND2_X1 U15632 ( .A1(n12519), .A2(n12518), .ZN(n14274) );
  NAND2_X1 U15633 ( .A1(n10812), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12520) );
  XNOR2_X1 U15634 ( .A(n14274), .B(n12520), .ZN(n14273) );
  AND2_X1 U15635 ( .A1(n12837), .A2(n16591), .ZN(n20221) );
  NAND2_X1 U15636 ( .A1(READY12_REG_SCAN_IN), .A2(READY21_REG_SCAN_IN), .ZN(
        n20226) );
  INV_X1 U15637 ( .A(n20226), .ZN(n20114) );
  OR2_X1 U15638 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20114), .ZN(n12791) );
  NAND2_X1 U15639 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12791), .ZN(n12521) );
  NOR2_X1 U15640 ( .A1(n12963), .A2(n12521), .ZN(n12522) );
  INV_X1 U15641 ( .A(n12531), .ZN(n12526) );
  NOR2_X1 U15642 ( .A1(n10305), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12543) );
  NAND2_X1 U15643 ( .A1(n14295), .A2(P2_EAX_REG_5__SCAN_IN), .ZN(n12524) );
  NAND2_X1 U15644 ( .A1(n9657), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12523) );
  OAI211_X1 U15645 ( .C1(n12526), .C2(n12525), .A(n12524), .B(n12523), .ZN(
        n12529) );
  INV_X1 U15646 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n12527) );
  NOR2_X1 U15647 ( .A1(n12766), .A2(n12527), .ZN(n12528) );
  INV_X1 U15648 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U15649 ( .A1(n14295), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12535) );
  INV_X1 U15650 ( .A(n12532), .ZN(n12533) );
  OR2_X1 U15651 ( .A1(n12740), .A2(n12533), .ZN(n12534) );
  OAI211_X1 U15652 ( .C1(n12766), .C2(n12536), .A(n12535), .B(n12534), .ZN(
        n13556) );
  MUX2_X1 U15653 ( .A(n10305), .B(n20208), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12538) );
  NAND2_X1 U15654 ( .A1(n10293), .A2(n12537), .ZN(n12553) );
  AND2_X1 U15655 ( .A1(n12538), .A2(n12553), .ZN(n12539) );
  INV_X1 U15656 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19315) );
  AOI21_X1 U15657 ( .B1(n9676), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12542) );
  NAND2_X1 U15658 ( .A1(n10322), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12541) );
  OAI211_X1 U15659 ( .C1(n12766), .C2(n19315), .A(n12542), .B(n12541), .ZN(
        n13001) );
  INV_X1 U15660 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20121) );
  AOI22_X1 U15661 ( .A1(n12543), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12537), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12544) );
  OAI21_X1 U15662 ( .B1(n12766), .B2(n20121), .A(n12544), .ZN(n12551) );
  INV_X1 U15663 ( .A(n12551), .ZN(n12545) );
  OR2_X1 U15664 ( .A1(n12546), .A2(n12740), .ZN(n12549) );
  NAND2_X1 U15665 ( .A1(n12984), .A2(n10305), .ZN(n12547) );
  MUX2_X1 U15666 ( .A(n12547), .B(n20199), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12548) );
  NAND2_X1 U15667 ( .A1(n12549), .A2(n12548), .ZN(n13713) );
  INV_X1 U15668 ( .A(n13713), .ZN(n12550) );
  NAND2_X1 U15669 ( .A1(n13712), .A2(n12550), .ZN(n13716) );
  OAI211_X1 U15670 ( .C1(n20041), .C2(n20190), .A(n12554), .B(n12553), .ZN(
        n12555) );
  AND3_X1 U15671 ( .A1(n13716), .A2(n10195), .A3(n12555), .ZN(n12556) );
  OR2_X1 U15672 ( .A1(n12556), .A2(n12558), .ZN(n13680) );
  INV_X1 U15673 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n21208) );
  AOI22_X1 U15674 ( .A1(n14295), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12557) );
  OAI21_X1 U15675 ( .B1(n12766), .B2(n21208), .A(n12557), .ZN(n13679) );
  NOR2_X1 U15676 ( .A1(n13680), .A2(n13679), .ZN(n13681) );
  INV_X1 U15677 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13609) );
  AOI22_X1 U15678 ( .A1(n9657), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12560) );
  NAND2_X1 U15679 ( .A1(n14295), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12559) );
  AND2_X1 U15680 ( .A1(n12560), .A2(n12559), .ZN(n12563) );
  OR2_X1 U15681 ( .A1(n12740), .A2(n12561), .ZN(n12562) );
  OAI211_X1 U15682 ( .C1(n12766), .C2(n13609), .A(n12563), .B(n12562), .ZN(
        n13455) );
  OR2_X1 U15683 ( .A1(n12740), .A2(n12564), .ZN(n12565) );
  INV_X1 U15684 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20127) );
  AOI22_X1 U15685 ( .A1(n14295), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12567) );
  OAI21_X1 U15686 ( .B1(n12766), .B2(n20127), .A(n12567), .ZN(n14073) );
  NAND2_X1 U15687 ( .A1(n14074), .A2(n14073), .ZN(n12569) );
  OR2_X1 U15688 ( .A1(n12740), .A2(n10869), .ZN(n12568) );
  INV_X1 U15689 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20129) );
  AOI22_X1 U15690 ( .A1(n14295), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12570) );
  OAI21_X1 U15691 ( .B1(n12766), .B2(n20129), .A(n12570), .ZN(n16563) );
  INV_X1 U15692 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12590) );
  AOI22_X1 U15693 ( .A1(n14295), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15694 ( .A1(n14432), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14431), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12574) );
  NAND2_X1 U15695 ( .A1(n10430), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12573) );
  NAND2_X1 U15696 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12572) );
  NAND2_X1 U15697 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12571) );
  AND4_X1 U15698 ( .A1(n12574), .A2(n12573), .A3(n12572), .A4(n12571), .ZN(
        n12587) );
  AOI22_X1 U15699 ( .A1(n14404), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12578) );
  NAND2_X1 U15700 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12577) );
  INV_X1 U15701 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n19728) );
  OR2_X1 U15702 ( .A1(n14417), .A2(n19728), .ZN(n12576) );
  INV_X1 U15703 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13900) );
  OR2_X1 U15704 ( .A1(n14416), .A2(n13900), .ZN(n12575) );
  AOI22_X1 U15705 ( .A1(n14430), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12586) );
  INV_X1 U15706 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12579) );
  OR2_X1 U15707 ( .A1(n14412), .A2(n12579), .ZN(n12584) );
  INV_X1 U15708 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12580) );
  OR2_X1 U15709 ( .A1(n14411), .A2(n12580), .ZN(n12583) );
  NAND2_X1 U15710 ( .A1(n10578), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12582) );
  NAND2_X1 U15711 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12581) );
  AND4_X1 U15712 ( .A1(n12584), .A2(n12583), .A3(n12582), .A4(n12581), .ZN(
        n12585) );
  NAND4_X1 U15713 ( .A1(n12587), .A2(n10166), .A3(n12586), .A4(n12585), .ZN(
        n13344) );
  INV_X1 U15714 ( .A(n13344), .ZN(n13531) );
  OR2_X1 U15715 ( .A1(n12740), .A2(n13531), .ZN(n12588) );
  OAI211_X1 U15716 ( .C1(n12766), .C2(n12590), .A(n12589), .B(n12588), .ZN(
        n13602) );
  INV_X1 U15717 ( .A(n13602), .ZN(n12591) );
  AOI22_X1 U15718 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14404), .B1(
        n14432), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12595) );
  NAND2_X1 U15719 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12594) );
  NAND2_X1 U15720 ( .A1(n10430), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12593) );
  NAND2_X1 U15721 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12592) );
  AND4_X1 U15722 ( .A1(n12595), .A2(n12594), .A3(n12593), .A4(n12592), .ZN(
        n12610) );
  AOI22_X1 U15723 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14431), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12601) );
  NAND2_X1 U15724 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12600) );
  INV_X1 U15725 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12596) );
  OR2_X1 U15726 ( .A1(n14417), .A2(n12596), .ZN(n12599) );
  OR2_X1 U15727 ( .A1(n14411), .A2(n12597), .ZN(n12598) );
  AND4_X1 U15728 ( .A1(n12601), .A2(n12600), .A3(n12599), .A4(n12598), .ZN(
        n12609) );
  AOI22_X1 U15729 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10578), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12608) );
  INV_X1 U15730 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12602) );
  OR2_X1 U15731 ( .A1(n14412), .A2(n12602), .ZN(n12606) );
  INV_X1 U15732 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13874) );
  OR2_X1 U15733 ( .A1(n14416), .A2(n13874), .ZN(n12605) );
  NAND2_X1 U15734 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12604) );
  NAND2_X1 U15735 ( .A1(n14430), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12603) );
  AND4_X1 U15736 ( .A1(n12606), .A2(n12605), .A3(n12604), .A4(n12603), .ZN(
        n12607) );
  NAND4_X1 U15737 ( .A1(n12610), .A2(n12609), .A3(n12608), .A4(n12607), .ZN(
        n13417) );
  INV_X1 U15738 ( .A(n13417), .ZN(n12613) );
  NAND2_X1 U15739 ( .A1(n14296), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12612) );
  AOI22_X1 U15740 ( .A1(n14295), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12611) );
  OAI211_X1 U15741 ( .C1(n12613), .C2(n12740), .A(n12612), .B(n12611), .ZN(
        n16167) );
  INV_X1 U15742 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U15743 ( .A1(n14295), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U15744 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10494), .B1(
        n14430), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15745 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10645), .B1(
        n14433), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U15746 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14431), .B1(
        n14432), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12615) );
  NAND2_X1 U15747 ( .A1(n10430), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12614) );
  AND4_X1 U15748 ( .A1(n12617), .A2(n12616), .A3(n12615), .A4(n12614), .ZN(
        n12632) );
  AOI22_X1 U15749 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n14404), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12623) );
  NAND2_X1 U15750 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12622) );
  OR2_X1 U15751 ( .A1(n14412), .A2(n12618), .ZN(n12621) );
  INV_X1 U15752 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12619) );
  OR2_X1 U15753 ( .A1(n14417), .A2(n12619), .ZN(n12620) );
  NAND4_X1 U15754 ( .A1(n12623), .A2(n12622), .A3(n12621), .A4(n12620), .ZN(
        n12630) );
  INV_X1 U15755 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14044) );
  OR2_X1 U15756 ( .A1(n14416), .A2(n14044), .ZN(n12628) );
  INV_X1 U15757 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12624) );
  OR2_X1 U15758 ( .A1(n14411), .A2(n12624), .ZN(n12627) );
  NAND2_X1 U15759 ( .A1(n10578), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12626) );
  NAND2_X1 U15760 ( .A1(n10468), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12625) );
  NAND4_X1 U15761 ( .A1(n12628), .A2(n12627), .A3(n12626), .A4(n12625), .ZN(
        n12629) );
  NOR2_X1 U15762 ( .A1(n12630), .A2(n12629), .ZN(n12631) );
  OR2_X1 U15763 ( .A1(n12740), .A2(n13349), .ZN(n12633) );
  OAI211_X1 U15764 ( .C1(n12766), .C2(n12635), .A(n12634), .B(n12633), .ZN(
        n12636) );
  INV_X1 U15765 ( .A(n12636), .ZN(n15521) );
  AOI22_X1 U15766 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n14404), .B1(
        n14432), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12640) );
  NAND2_X1 U15767 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12639) );
  NAND2_X1 U15768 ( .A1(n10430), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12638) );
  NAND2_X1 U15769 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12637) );
  AND4_X1 U15770 ( .A1(n12640), .A2(n12639), .A3(n12638), .A4(n12637), .ZN(
        n12655) );
  AOI22_X1 U15771 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14431), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12646) );
  NAND2_X1 U15772 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12645) );
  INV_X1 U15773 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12641) );
  OR2_X1 U15774 ( .A1(n14417), .A2(n12641), .ZN(n12644) );
  INV_X1 U15775 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12642) );
  OR2_X1 U15776 ( .A1(n14411), .A2(n12642), .ZN(n12643) );
  AND4_X1 U15777 ( .A1(n12646), .A2(n12645), .A3(n12644), .A4(n12643), .ZN(
        n12654) );
  AOI22_X1 U15778 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10578), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12653) );
  INV_X1 U15779 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12647) );
  OR2_X1 U15780 ( .A1(n14412), .A2(n12647), .ZN(n12651) );
  INV_X1 U15781 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14109) );
  OR2_X1 U15782 ( .A1(n14416), .A2(n14109), .ZN(n12650) );
  NAND2_X1 U15783 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12649) );
  NAND2_X1 U15784 ( .A1(n14430), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12648) );
  AND4_X1 U15785 ( .A1(n12651), .A2(n12650), .A3(n12649), .A4(n12648), .ZN(
        n12652) );
  NAND4_X1 U15786 ( .A1(n12655), .A2(n12654), .A3(n12653), .A4(n12652), .ZN(
        n13505) );
  AOI22_X1 U15787 ( .A1(n14296), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n9916), 
        .B2(n13505), .ZN(n12657) );
  AOI22_X1 U15788 ( .A1(n14295), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12656) );
  NAND2_X1 U15789 ( .A1(n12657), .A2(n12656), .ZN(n13724) );
  AOI22_X1 U15790 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14431), .B1(
        n14432), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12661) );
  NAND2_X1 U15791 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12660) );
  NAND2_X1 U15792 ( .A1(n10430), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12659) );
  NAND2_X1 U15793 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12658) );
  AND4_X1 U15794 ( .A1(n12661), .A2(n12660), .A3(n12659), .A4(n12658), .ZN(
        n12676) );
  AOI22_X1 U15795 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n14404), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12667) );
  NAND2_X1 U15796 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12666) );
  INV_X1 U15797 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12662) );
  OR2_X1 U15798 ( .A1(n14417), .A2(n12662), .ZN(n12665) );
  INV_X1 U15799 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12663) );
  OR2_X1 U15800 ( .A1(n14411), .A2(n12663), .ZN(n12664) );
  AND4_X1 U15801 ( .A1(n12667), .A2(n12666), .A3(n12665), .A4(n12664), .ZN(
        n12675) );
  AOI22_X1 U15802 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10578), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12674) );
  INV_X1 U15803 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12668) );
  OR2_X1 U15804 ( .A1(n14412), .A2(n12668), .ZN(n12672) );
  INV_X1 U15805 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14358) );
  OR2_X1 U15806 ( .A1(n14416), .A2(n14358), .ZN(n12671) );
  NAND2_X1 U15807 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12670) );
  NAND2_X1 U15808 ( .A1(n14430), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12669) );
  AND4_X1 U15809 ( .A1(n12672), .A2(n12671), .A3(n12670), .A4(n12669), .ZN(
        n12673) );
  NAND4_X1 U15810 ( .A1(n12676), .A2(n12675), .A3(n12674), .A4(n12673), .ZN(
        n13436) );
  INV_X1 U15811 ( .A(n13436), .ZN(n13438) );
  AOI22_X1 U15812 ( .A1(n14295), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12677) );
  OAI21_X1 U15813 ( .B1(n13438), .B2(n12740), .A(n12677), .ZN(n12678) );
  AOI21_X1 U15814 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n14296), .A(n12678), 
        .ZN(n16124) );
  AOI22_X1 U15815 ( .A1(n14295), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U15816 ( .A1(n14432), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14404), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12682) );
  NAND2_X1 U15817 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12681) );
  NAND2_X1 U15818 ( .A1(n10430), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12680) );
  NAND2_X1 U15819 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12679) );
  AND4_X1 U15820 ( .A1(n12682), .A2(n12681), .A3(n12680), .A4(n12679), .ZN(
        n12697) );
  AOI22_X1 U15821 ( .A1(n14431), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12688) );
  NAND2_X1 U15822 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12687) );
  INV_X1 U15823 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12683) );
  OR2_X1 U15824 ( .A1(n14417), .A2(n12683), .ZN(n12686) );
  INV_X1 U15825 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12684) );
  OR2_X1 U15826 ( .A1(n14411), .A2(n12684), .ZN(n12685) );
  AND4_X1 U15827 ( .A1(n12688), .A2(n12687), .A3(n12686), .A4(n12685), .ZN(
        n12696) );
  AOI22_X1 U15828 ( .A1(n10578), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12695) );
  INV_X1 U15829 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12689) );
  OR2_X1 U15830 ( .A1(n14412), .A2(n12689), .ZN(n12693) );
  INV_X1 U15831 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14379) );
  OR2_X1 U15832 ( .A1(n14416), .A2(n14379), .ZN(n12692) );
  NAND2_X1 U15833 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12691) );
  NAND2_X1 U15834 ( .A1(n14430), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12690) );
  AND4_X1 U15835 ( .A1(n12693), .A2(n12692), .A3(n12691), .A4(n12690), .ZN(
        n12694) );
  NAND4_X1 U15836 ( .A1(n12697), .A2(n12696), .A3(n12695), .A4(n12694), .ZN(
        n13477) );
  INV_X1 U15837 ( .A(n13477), .ZN(n12698) );
  OR2_X1 U15838 ( .A1(n12740), .A2(n12698), .ZN(n12699) );
  OAI211_X1 U15839 ( .C1(n12766), .C2(n16109), .A(n12700), .B(n12699), .ZN(
        n16108) );
  AOI22_X1 U15840 ( .A1(n14295), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U15841 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n14430), .B1(
        n10494), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12704) );
  AOI22_X1 U15842 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10645), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U15843 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14431), .B1(
        n14432), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12702) );
  NAND2_X1 U15844 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12701) );
  AND4_X1 U15845 ( .A1(n12704), .A2(n12703), .A3(n12702), .A4(n12701), .ZN(
        n12718) );
  AOI22_X1 U15846 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n14404), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12710) );
  NAND2_X1 U15847 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12709) );
  INV_X1 U15848 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12705) );
  OR2_X1 U15849 ( .A1(n14417), .A2(n12705), .ZN(n12708) );
  INV_X1 U15850 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12706) );
  OR2_X1 U15851 ( .A1(n14412), .A2(n12706), .ZN(n12707) );
  NAND4_X1 U15852 ( .A1(n12710), .A2(n12709), .A3(n12708), .A4(n12707), .ZN(
        n12716) );
  INV_X1 U15853 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14392) );
  OR2_X1 U15854 ( .A1(n14416), .A2(n14392), .ZN(n12714) );
  OR2_X1 U15855 ( .A1(n14411), .A2(n21187), .ZN(n12713) );
  NAND2_X1 U15856 ( .A1(n10578), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12712) );
  NAND2_X1 U15857 ( .A1(n10468), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12711) );
  NAND4_X1 U15858 ( .A1(n12714), .A2(n12713), .A3(n12712), .A4(n12711), .ZN(
        n12715) );
  NOR2_X1 U15859 ( .A1(n12716), .A2(n12715), .ZN(n12717) );
  OR2_X1 U15860 ( .A1(n12740), .A2(n13622), .ZN(n12719) );
  OAI211_X1 U15861 ( .C1(n12766), .C2(n12721), .A(n12720), .B(n12719), .ZN(
        n16098) );
  AOI22_X1 U15862 ( .A1(n14295), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U15863 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10578), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U15864 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10645), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U15865 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n14404), .B1(
        n14432), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12723) );
  NAND2_X1 U15866 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12722) );
  AND4_X1 U15867 ( .A1(n12725), .A2(n12724), .A3(n12723), .A4(n12722), .ZN(
        n12739) );
  AOI22_X1 U15868 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n14431), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12730) );
  NAND2_X1 U15869 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12729) );
  OR2_X1 U15870 ( .A1(n14417), .A2(n14424), .ZN(n12728) );
  OR2_X1 U15871 ( .A1(n14411), .A2(n12726), .ZN(n12727) );
  NAND4_X1 U15872 ( .A1(n12730), .A2(n12729), .A3(n12728), .A4(n12727), .ZN(
        n12737) );
  OR2_X1 U15873 ( .A1(n14412), .A2(n12731), .ZN(n12735) );
  OR2_X1 U15874 ( .A1(n14416), .A2(n14413), .ZN(n12734) );
  NAND2_X1 U15875 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12733) );
  NAND2_X1 U15876 ( .A1(n14430), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12732) );
  NAND4_X1 U15877 ( .A1(n12735), .A2(n12734), .A3(n12733), .A4(n12732), .ZN(
        n12736) );
  NOR2_X1 U15878 ( .A1(n12737), .A2(n12736), .ZN(n12738) );
  OR2_X1 U15879 ( .A1(n12740), .A2(n13831), .ZN(n12741) );
  OAI211_X1 U15880 ( .C1(n12766), .C2(n15841), .A(n12742), .B(n12741), .ZN(
        n12819) );
  INV_X1 U15881 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20141) );
  AOI22_X1 U15882 ( .A1(n14295), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12743) );
  OAI21_X1 U15883 ( .B1(n12766), .B2(n20141), .A(n12743), .ZN(n15501) );
  INV_X1 U15884 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20143) );
  AOI22_X1 U15885 ( .A1(n14295), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12744) );
  OAI21_X1 U15886 ( .B1(n12766), .B2(n20143), .A(n12744), .ZN(n15675) );
  NAND2_X1 U15887 ( .A1(n14296), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12746) );
  AOI22_X1 U15888 ( .A1(n14295), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12745) );
  AOI22_X1 U15889 ( .A1(n14295), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12747) );
  OAI21_X1 U15890 ( .B1(n12766), .B2(n10759), .A(n12747), .ZN(n15659) );
  AOI22_X1 U15891 ( .A1(n14295), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12748) );
  OAI21_X1 U15892 ( .B1(n12766), .B2(n12749), .A(n12748), .ZN(n15999) );
  INV_X1 U15893 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20148) );
  AOI22_X1 U15894 ( .A1(n14295), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12750) );
  OAI21_X1 U15895 ( .B1(n12766), .B2(n20148), .A(n12750), .ZN(n15645) );
  NAND2_X1 U15896 ( .A1(n14296), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U15897 ( .A1(n14295), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12751) );
  NAND2_X1 U15898 ( .A1(n12752), .A2(n12751), .ZN(n15486) );
  AOI22_X1 U15899 ( .A1(n14295), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12753) );
  OAI21_X1 U15900 ( .B1(n12766), .B2(n10770), .A(n12753), .ZN(n15471) );
  NAND2_X1 U15901 ( .A1(n14296), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U15902 ( .A1(n14295), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12755) );
  AND2_X1 U15903 ( .A1(n12756), .A2(n12755), .ZN(n15624) );
  NAND2_X1 U15904 ( .A1(n14296), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U15905 ( .A1(n14295), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12757) );
  AND2_X1 U15906 ( .A1(n12758), .A2(n12757), .ZN(n15454) );
  NAND2_X1 U15907 ( .A1(n14296), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U15908 ( .A1(n14295), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12759) );
  NAND2_X1 U15909 ( .A1(n12760), .A2(n12759), .ZN(n15612) );
  NAND2_X1 U15910 ( .A1(n14296), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U15911 ( .A1(n14295), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12761) );
  AND2_X1 U15912 ( .A1(n12762), .A2(n12761), .ZN(n12830) );
  NAND2_X1 U15913 ( .A1(n14296), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U15914 ( .A1(n14295), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12763) );
  AND2_X1 U15915 ( .A1(n12764), .A2(n12763), .ZN(n15444) );
  INV_X1 U15916 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20160) );
  AOI22_X1 U15917 ( .A1(n14295), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12765) );
  OAI21_X1 U15918 ( .B1(n12766), .B2(n20160), .A(n12765), .ZN(n14607) );
  NAND2_X1 U15919 ( .A1(n14296), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U15920 ( .A1(n14295), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n9657), .B2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12767) );
  NAND2_X1 U15921 ( .A1(n12768), .A2(n12767), .ZN(n12769) );
  NAND2_X1 U15922 ( .A1(n14609), .A2(n12769), .ZN(n14298) );
  INV_X1 U15923 ( .A(n14609), .ZN(n12771) );
  INV_X1 U15924 ( .A(n12769), .ZN(n12770) );
  NAND2_X1 U15925 ( .A1(n12771), .A2(n12770), .ZN(n12772) );
  NAND2_X1 U15926 ( .A1(n14298), .A2(n12772), .ZN(n15880) );
  INV_X1 U15927 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n21221) );
  INV_X1 U15928 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20120) );
  INV_X1 U15929 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20103) );
  NAND2_X1 U15930 ( .A1(n21221), .A2(n20120), .ZN(n19136) );
  OAI211_X1 U15931 ( .C1(n21221), .C2(n20120), .A(n20103), .B(n19136), .ZN(
        n20227) );
  NOR2_X1 U15932 ( .A1(n20227), .A2(n20114), .ZN(n13059) );
  INV_X1 U15933 ( .A(n13059), .ZN(n13016) );
  NOR2_X1 U15934 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13016), .ZN(n12777) );
  AND2_X1 U15935 ( .A1(n12837), .A2(n12775), .ZN(n12848) );
  AOI21_X1 U15936 ( .B1(n20228), .B2(n20226), .A(P2_EBX_REG_31__SCAN_IN), .ZN(
        n12776) );
  NAND2_X1 U15937 ( .A1(n12848), .A2(n12776), .ZN(n12779) );
  INV_X1 U15938 ( .A(n12777), .ZN(n16613) );
  NAND2_X1 U15939 ( .A1(n19480), .A2(n16613), .ZN(n12778) );
  NAND2_X1 U15940 ( .A1(n12779), .A2(n12778), .ZN(n19320) );
  NOR2_X1 U15941 ( .A1(n20041), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19758) );
  INV_X1 U15942 ( .A(n19758), .ZN(n12780) );
  NOR2_X1 U15943 ( .A1(n19133), .A2(n12780), .ZN(n16608) );
  INV_X1 U15944 ( .A(n16608), .ZN(n12781) );
  NAND3_X1 U15945 ( .A1(n12781), .A2(n19277), .A3(n20099), .ZN(n12782) );
  NOR2_X2 U15946 ( .A1(n20221), .A2(n12782), .ZN(n19318) );
  AOI22_X1 U15947 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19320), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19318), .ZN(n12784) );
  NAND2_X1 U15948 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19298), .ZN(
        n12783) );
  OAI211_X1 U15949 ( .C1(n15880), .C2(n19312), .A(n12784), .B(n12783), .ZN(
        n12785) );
  AOI21_X1 U15950 ( .B1(n14273), .B2(n19317), .A(n12785), .ZN(n12795) );
  INV_X1 U15951 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U15952 ( .A1(n9663), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12786) );
  OAI21_X1 U15953 ( .B1(n12788), .B2(n12787), .A(n12786), .ZN(n12789) );
  AOI21_X1 U15954 ( .B1(n12790), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12789), .ZN(n14281) );
  INV_X1 U15955 ( .A(n15888), .ZN(n12793) );
  NOR2_X1 U15956 ( .A1(n12963), .A2(n12791), .ZN(n12792) );
  NAND2_X1 U15957 ( .A1(n20221), .A2(n12792), .ZN(n19292) );
  NAND2_X1 U15958 ( .A1(n12797), .A2(n12796), .ZN(P2_U2825) );
  INV_X1 U15959 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21045) );
  NOR3_X1 U15960 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21045), .ZN(n12799) );
  NOR4_X1 U15961 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12798) );
  NAND4_X1 U15962 ( .A1(n20419), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12799), .A4(
        n12798), .ZN(U214) );
  NOR4_X1 U15963 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12803) );
  NOR4_X1 U15964 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12802) );
  NOR4_X1 U15965 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12801) );
  NOR4_X1 U15966 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12800) );
  NAND4_X1 U15967 ( .A1(n12803), .A2(n12802), .A3(n12801), .A4(n12800), .ZN(
        n12808) );
  NOR4_X1 U15968 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12806) );
  NOR4_X1 U15969 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12805) );
  NOR4_X1 U15970 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12804) );
  INV_X1 U15971 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20124) );
  NAND4_X1 U15972 ( .A1(n12806), .A2(n12805), .A3(n12804), .A4(n20124), .ZN(
        n12807) );
  NOR2_X1 U15973 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12810) );
  NOR4_X1 U15974 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12809) );
  NAND4_X1 U15975 ( .A1(n12810), .A2(P2_W_R_N_REG_SCAN_IN), .A3(
        P2_M_IO_N_REG_SCAN_IN), .A4(n12809), .ZN(n12836) );
  NOR2_X1 U15976 ( .A1(n19517), .A2(n12836), .ZN(n16700) );
  NAND2_X1 U15977 ( .A1(n16700), .A2(U214), .ZN(U212) );
  NAND2_X1 U15978 ( .A1(n19308), .A2(n12811), .ZN(n19331) );
  AOI211_X1 U15979 ( .C1(n12814), .C2(n12812), .A(n15498), .B(n19331), .ZN(
        n12823) );
  AOI22_X1 U15980 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n19320), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19298), .ZN(n12813) );
  OAI211_X1 U15981 ( .C1(n15841), .C2(n19260), .A(n12813), .B(n19277), .ZN(
        n12822) );
  NAND2_X1 U15982 ( .A1(n19308), .A2(n19289), .ZN(n19325) );
  INV_X1 U15983 ( .A(n12814), .ZN(n15839) );
  OAI22_X1 U15984 ( .A1(n12815), .A2(n19300), .B1(n19325), .B2(n15839), .ZN(
        n12821) );
  AND2_X1 U15985 ( .A1(n13620), .A2(n12816), .ZN(n12817) );
  OR2_X1 U15986 ( .A1(n12817), .A2(n13931), .ZN(n15842) );
  INV_X1 U15987 ( .A(n12818), .ZN(n15503) );
  OAI21_X1 U15988 ( .B1(n16099), .B2(n12819), .A(n15503), .ZN(n19349) );
  OAI22_X1 U15989 ( .A1(n15842), .A2(n19292), .B1(n19312), .B2(n19349), .ZN(
        n12820) );
  OR4_X1 U15990 ( .A1(n12823), .A2(n12822), .A3(n12821), .A4(n12820), .ZN(
        P2_U2840) );
  AOI211_X1 U15991 ( .C1(n15716), .C2(n12824), .A(n12825), .B(n20099), .ZN(
        n12835) );
  INV_X1 U15992 ( .A(n19320), .ZN(n19285) );
  INV_X1 U15993 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12826) );
  OAI22_X1 U15994 ( .A1(n12827), .A2(n19300), .B1(n19285), .B2(n12826), .ZN(
        n12834) );
  OAI22_X1 U15995 ( .A1(n15714), .A2(n19326), .B1(n20157), .B2(n19260), .ZN(
        n12833) );
  AND2_X1 U15996 ( .A1(n9722), .A2(n12828), .ZN(n12829) );
  OR2_X1 U15997 ( .A1(n12829), .A2(n15437), .ZN(n15914) );
  NAND2_X1 U15998 ( .A1(n15611), .A2(n12830), .ZN(n12831) );
  NAND2_X1 U15999 ( .A1(n9723), .A2(n12831), .ZN(n15909) );
  OAI22_X1 U16000 ( .A1(n15914), .A2(n19292), .B1(n15909), .B2(n19312), .ZN(
        n12832) );
  OR4_X1 U16001 ( .A1(n12835), .A2(n12834), .A3(n12833), .A4(n12832), .ZN(
        P2_U2828) );
  NOR2_X1 U16002 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12836), .ZN(n16778)
         );
  INV_X2 U16003 ( .A(n21255), .ZN(U215) );
  INV_X1 U16004 ( .A(n12987), .ZN(n19409) );
  AND2_X1 U16005 ( .A1(n12837), .A2(n19409), .ZN(n19329) );
  INV_X1 U16006 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12839) );
  INV_X1 U16007 ( .A(n12848), .ZN(n12838) );
  OAI211_X1 U16008 ( .C1(n19329), .C2(n12839), .A(n12838), .B(n12841), .ZN(
        P2_U2814) );
  INV_X1 U16009 ( .A(n12840), .ZN(n13070) );
  INV_X1 U16010 ( .A(n20221), .ZN(n12844) );
  INV_X1 U16011 ( .A(n12841), .ZN(n12842) );
  OAI21_X1 U16012 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n12842), .A(n12844), 
        .ZN(n12843) );
  OAI21_X1 U16013 ( .B1(n13070), .B2(n12844), .A(n12843), .ZN(P2_U3612) );
  AND2_X1 U16014 ( .A1(n12840), .A2(n20226), .ZN(n12996) );
  NOR2_X1 U16015 ( .A1(n12996), .A2(n13059), .ZN(n12845) );
  AND2_X1 U16016 ( .A1(n16591), .A2(n12845), .ZN(n12846) );
  NAND2_X1 U16017 ( .A1(n16590), .A2(n12846), .ZN(n16602) );
  AND2_X1 U16018 ( .A1(n16602), .A2(n20095), .ZN(n20218) );
  OAI21_X1 U16019 ( .B1(n10688), .B2(n20218), .A(n12847), .ZN(P2_U2819) );
  INV_X1 U16020 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19444) );
  NAND3_X1 U16021 ( .A1(n12848), .A2(n9675), .A3(n20226), .ZN(n12946) );
  AOI22_X1 U16022 ( .A1(n19519), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19517), .ZN(n19536) );
  INV_X1 U16023 ( .A(n19536), .ZN(n15677) );
  NAND2_X1 U16024 ( .A1(n12884), .A2(n15677), .ZN(n12894) );
  NAND2_X1 U16025 ( .A1(n12848), .A2(n20226), .ZN(n12849) );
  NAND2_X1 U16026 ( .A1(n19481), .A2(P2_UWORD_REG_1__SCAN_IN), .ZN(n12850) );
  OAI211_X1 U16027 ( .C1(n19444), .C2(n19410), .A(n12894), .B(n12850), .ZN(
        P2_U2953) );
  INV_X1 U16028 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n12856) );
  INV_X1 U16029 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n12851) );
  OR2_X1 U16030 ( .A1(n19517), .A2(n12851), .ZN(n12853) );
  NAND2_X1 U16031 ( .A1(n12872), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12852) );
  AND2_X1 U16032 ( .A1(n12853), .A2(n12852), .ZN(n19358) );
  INV_X1 U16033 ( .A(n19358), .ZN(n12854) );
  NAND2_X1 U16034 ( .A1(n12884), .A2(n12854), .ZN(n12880) );
  NAND2_X1 U16035 ( .A1(n19481), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n12855) );
  OAI211_X1 U16036 ( .C1(n19410), .C2(n12856), .A(n12880), .B(n12855), .ZN(
        P2_U2978) );
  INV_X1 U16037 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n21198) );
  NAND2_X1 U16038 ( .A1(n12872), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12858) );
  INV_X1 U16039 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16733) );
  OR2_X1 U16040 ( .A1(n19517), .A2(n16733), .ZN(n12857) );
  NAND2_X1 U16041 ( .A1(n12858), .A2(n12857), .ZN(n19355) );
  NAND2_X1 U16042 ( .A1(n12884), .A2(n19355), .ZN(n12878) );
  NAND2_X1 U16043 ( .A1(n19481), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12859) );
  OAI211_X1 U16044 ( .C1(n21198), .C2(n19410), .A(n12878), .B(n12859), .ZN(
        P2_U2964) );
  INV_X1 U16045 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19450) );
  NAND2_X1 U16046 ( .A1(n12872), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12862) );
  INV_X1 U16047 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n12860) );
  OR2_X1 U16048 ( .A1(n12872), .A2(n12860), .ZN(n12861) );
  NAND2_X1 U16049 ( .A1(n12862), .A2(n12861), .ZN(n19350) );
  NAND2_X1 U16050 ( .A1(n12884), .A2(n19350), .ZN(n12887) );
  NAND2_X1 U16051 ( .A1(n19481), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12863) );
  OAI211_X1 U16052 ( .C1(n19450), .C2(n19410), .A(n12887), .B(n12863), .ZN(
        P2_U2981) );
  INV_X1 U16053 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19462) );
  NAND2_X1 U16054 ( .A1(n12872), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12865) );
  INV_X1 U16055 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16738) );
  OR2_X1 U16056 ( .A1(n12872), .A2(n16738), .ZN(n12864) );
  NAND2_X1 U16057 ( .A1(n12865), .A2(n12864), .ZN(n19366) );
  NAND2_X1 U16058 ( .A1(n12884), .A2(n19366), .ZN(n12889) );
  NAND2_X1 U16059 ( .A1(n19481), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12866) );
  OAI211_X1 U16060 ( .C1(n19462), .C2(n19410), .A(n12889), .B(n12866), .ZN(
        P2_U2975) );
  INV_X1 U16061 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19427) );
  INV_X1 U16062 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n12867) );
  OR2_X1 U16063 ( .A1(n12872), .A2(n12867), .ZN(n12869) );
  NAND2_X1 U16064 ( .A1(n12872), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12868) );
  AND2_X1 U16065 ( .A1(n12869), .A2(n12868), .ZN(n19363) );
  INV_X1 U16066 ( .A(n19363), .ZN(n12870) );
  NAND2_X1 U16067 ( .A1(n12884), .A2(n12870), .ZN(n12891) );
  NAND2_X1 U16068 ( .A1(n19481), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12871) );
  OAI211_X1 U16069 ( .C1(n19410), .C2(n19427), .A(n12891), .B(n12871), .ZN(
        P2_U2961) );
  INV_X1 U16070 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19420) );
  INV_X1 U16071 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16731) );
  OR2_X1 U16072 ( .A1(n19517), .A2(n16731), .ZN(n12874) );
  NAND2_X1 U16073 ( .A1(n12872), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12873) );
  AND2_X1 U16074 ( .A1(n12874), .A2(n12873), .ZN(n19353) );
  INV_X1 U16075 ( .A(n19353), .ZN(n12875) );
  NAND2_X1 U16076 ( .A1(n12884), .A2(n12875), .ZN(n12940) );
  NAND2_X1 U16077 ( .A1(n19481), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n12876) );
  OAI211_X1 U16078 ( .C1(n19410), .C2(n19420), .A(n12940), .B(n12876), .ZN(
        P2_U2965) );
  INV_X1 U16079 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19454) );
  NAND2_X1 U16080 ( .A1(n19481), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12877) );
  OAI211_X1 U16081 ( .C1(n19454), .C2(n19410), .A(n12878), .B(n12877), .ZN(
        P2_U2979) );
  INV_X1 U16082 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19423) );
  NAND2_X1 U16083 ( .A1(n19481), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12879) );
  OAI211_X1 U16084 ( .C1(n19410), .C2(n19423), .A(n12880), .B(n12879), .ZN(
        P2_U2963) );
  INV_X1 U16085 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19425) );
  NAND2_X1 U16086 ( .A1(n19517), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12883) );
  INV_X1 U16087 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n12881) );
  OR2_X1 U16088 ( .A1(n19517), .A2(n12881), .ZN(n12882) );
  NAND2_X1 U16089 ( .A1(n12883), .A2(n12882), .ZN(n19360) );
  NAND2_X1 U16090 ( .A1(n12884), .A2(n19360), .ZN(n19482) );
  NAND2_X1 U16091 ( .A1(n19481), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12885) );
  OAI211_X1 U16092 ( .C1(n19425), .C2(n19410), .A(n19482), .B(n12885), .ZN(
        P2_U2962) );
  INV_X1 U16093 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n19418) );
  NAND2_X1 U16094 ( .A1(n19481), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12886) );
  OAI211_X1 U16095 ( .C1(n19418), .C2(n19410), .A(n12887), .B(n12886), .ZN(
        P2_U2966) );
  INV_X1 U16096 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19429) );
  NAND2_X1 U16097 ( .A1(n19481), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12888) );
  OAI211_X1 U16098 ( .C1(n19429), .C2(n19410), .A(n12889), .B(n12888), .ZN(
        P2_U2960) );
  INV_X1 U16099 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n12892) );
  NAND2_X1 U16100 ( .A1(n19481), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n12890) );
  OAI211_X1 U16101 ( .C1(n12892), .C2(n19410), .A(n12891), .B(n12890), .ZN(
        P2_U2976) );
  INV_X1 U16102 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n12895) );
  NAND2_X1 U16103 ( .A1(n19481), .A2(P2_LWORD_REG_1__SCAN_IN), .ZN(n12893) );
  OAI211_X1 U16104 ( .C1(n12895), .C2(n19410), .A(n12894), .B(n12893), .ZN(
        P2_U2968) );
  OAI21_X1 U16105 ( .B1(n19484), .B2(n13147), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12903) );
  OAI21_X1 U16106 ( .B1(n12897), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12896), .ZN(n13084) );
  INV_X1 U16107 ( .A(n13084), .ZN(n12901) );
  NAND2_X1 U16108 ( .A1(n19303), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13092) );
  NAND2_X1 U16109 ( .A1(n13092), .A2(n12898), .ZN(n12900) );
  OAI21_X1 U16110 ( .B1(n19316), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14336), .ZN(n13083) );
  NOR2_X1 U16111 ( .A1(n16537), .A2(n13083), .ZN(n12899) );
  AOI211_X1 U16112 ( .C1(n12901), .C2(n16529), .A(n12900), .B(n12899), .ZN(
        n12902) );
  NAND2_X1 U16113 ( .A1(n12903), .A2(n12902), .ZN(P2_U3014) );
  INV_X1 U16114 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U16115 ( .A1(n19519), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19517), .ZN(n19560) );
  NOR2_X1 U16116 ( .A1(n12946), .A2(n19560), .ZN(n12910) );
  AOI21_X1 U16117 ( .B1(n19480), .B2(P2_EAX_REG_6__SCAN_IN), .A(n12910), .ZN(
        n12904) );
  OAI21_X1 U16118 ( .B1(n12947), .B2(n12905), .A(n12904), .ZN(P2_U2973) );
  INV_X1 U16119 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U16120 ( .A1(n19519), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19517), .ZN(n19540) );
  NOR2_X1 U16121 ( .A1(n12946), .A2(n19540), .ZN(n12919) );
  AOI21_X1 U16122 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n19480), .A(n12919), .ZN(
        n12906) );
  OAI21_X1 U16123 ( .B1(n12947), .B2(n12907), .A(n12906), .ZN(P2_U2969) );
  INV_X1 U16124 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n12909) );
  OAI22_X1 U16125 ( .A1(n19517), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19519), .ZN(n19550) );
  NOR2_X1 U16126 ( .A1(n12946), .A2(n19550), .ZN(n12936) );
  AOI21_X1 U16127 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(n19480), .A(n12936), .ZN(
        n12908) );
  OAI21_X1 U16128 ( .B1(n12947), .B2(n12909), .A(n12908), .ZN(P2_U2971) );
  INV_X1 U16129 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n12912) );
  AOI21_X1 U16130 ( .B1(n19480), .B2(P2_EAX_REG_22__SCAN_IN), .A(n12910), .ZN(
        n12911) );
  OAI21_X1 U16131 ( .B1(n12947), .B2(n12912), .A(n12911), .ZN(P2_U2958) );
  INV_X1 U16132 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n12914) );
  AOI22_X1 U16133 ( .A1(n19519), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19517), .ZN(n19553) );
  NOR2_X1 U16134 ( .A1(n12946), .A2(n19553), .ZN(n12922) );
  AOI21_X1 U16135 ( .B1(n19480), .B2(P2_EAX_REG_21__SCAN_IN), .A(n12922), .ZN(
        n12913) );
  OAI21_X1 U16136 ( .B1(n12947), .B2(n12914), .A(n12913), .ZN(P2_U2957) );
  INV_X1 U16137 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n12916) );
  AOI22_X1 U16138 ( .A1(n19519), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19517), .ZN(n19546) );
  NOR2_X1 U16139 ( .A1(n12946), .A2(n19546), .ZN(n12925) );
  AOI21_X1 U16140 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n19480), .A(n12925), .ZN(
        n12915) );
  OAI21_X1 U16141 ( .B1(n12947), .B2(n12916), .A(n12915), .ZN(P2_U2970) );
  INV_X1 U16142 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U16143 ( .A1(n19519), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19517), .ZN(n19567) );
  NOR2_X1 U16144 ( .A1(n12946), .A2(n19567), .ZN(n12928) );
  AOI21_X1 U16145 ( .B1(n19480), .B2(P2_EAX_REG_7__SCAN_IN), .A(n12928), .ZN(
        n12917) );
  OAI21_X1 U16146 ( .B1(n12947), .B2(n12918), .A(n12917), .ZN(P2_U2974) );
  INV_X1 U16147 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n12921) );
  AOI21_X1 U16148 ( .B1(P2_EAX_REG_18__SCAN_IN), .B2(n19480), .A(n12919), .ZN(
        n12920) );
  OAI21_X1 U16149 ( .B1(n12947), .B2(n12921), .A(n12920), .ZN(P2_U2954) );
  INV_X1 U16150 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n12924) );
  AOI21_X1 U16151 ( .B1(P2_EAX_REG_5__SCAN_IN), .B2(n19480), .A(n12922), .ZN(
        n12923) );
  OAI21_X1 U16152 ( .B1(n12947), .B2(n12924), .A(n12923), .ZN(P2_U2972) );
  INV_X1 U16153 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n12927) );
  AOI21_X1 U16154 ( .B1(n19480), .B2(P2_EAX_REG_19__SCAN_IN), .A(n12925), .ZN(
        n12926) );
  OAI21_X1 U16155 ( .B1(n12947), .B2(n12927), .A(n12926), .ZN(P2_U2955) );
  INV_X1 U16156 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n12930) );
  AOI21_X1 U16157 ( .B1(n19480), .B2(P2_EAX_REG_23__SCAN_IN), .A(n12928), .ZN(
        n12929) );
  OAI21_X1 U16158 ( .B1(n12947), .B2(n12930), .A(n12929), .ZN(P2_U2959) );
  INV_X1 U16159 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12932) );
  OAI22_X1 U16160 ( .A1(n19517), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19519), .ZN(n19527) );
  NOR2_X1 U16161 ( .A1(n12946), .A2(n19527), .ZN(n12933) );
  AOI21_X1 U16162 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n19480), .A(n12933), .ZN(
        n12931) );
  OAI21_X1 U16163 ( .B1(n12947), .B2(n12932), .A(n12931), .ZN(P2_U2967) );
  INV_X1 U16164 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12935) );
  AOI21_X1 U16165 ( .B1(P2_EAX_REG_16__SCAN_IN), .B2(n19480), .A(n12933), .ZN(
        n12934) );
  OAI21_X1 U16166 ( .B1(n12947), .B2(n12935), .A(n12934), .ZN(P2_U2952) );
  INV_X1 U16167 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n12938) );
  AOI21_X1 U16168 ( .B1(P2_EAX_REG_20__SCAN_IN), .B2(n19480), .A(n12936), .ZN(
        n12937) );
  OAI21_X1 U16169 ( .B1(n12947), .B2(n12938), .A(n12937), .ZN(P2_U2956) );
  INV_X1 U16170 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n12941) );
  NAND2_X1 U16171 ( .A1(n19480), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n12939) );
  OAI211_X1 U16172 ( .C1(n12947), .C2(n12941), .A(n12940), .B(n12939), .ZN(
        P2_U2980) );
  NOR2_X2 U16173 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20909) );
  NAND2_X1 U16174 ( .A1(n20909), .A2(n20962), .ZN(n20241) );
  INV_X1 U16175 ( .A(n20241), .ZN(n13964) );
  AOI21_X1 U16176 ( .B1(n12943), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13964), 
        .ZN(n12944) );
  NAND2_X1 U16177 ( .A1(n13098), .A2(n12944), .ZN(P1_U2801) );
  INV_X1 U16178 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12948) );
  AOI22_X1 U16179 ( .A1(n19519), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19517), .ZN(n19348) );
  INV_X1 U16180 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12945) );
  OAI222_X1 U16181 ( .A1(n12948), .A2(n12947), .B1(n12946), .B2(n19348), .C1(
        n19410), .C2(n12945), .ZN(P2_U2982) );
  OAI21_X1 U16182 ( .B1(n10300), .B2(n16267), .A(n20041), .ZN(n13160) );
  AOI22_X1 U16183 ( .A1(n13160), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19989), .B2(n20208), .ZN(n12949) );
  NAND2_X1 U16184 ( .A1(n9675), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12951) );
  AND4_X1 U16185 ( .A1(n10300), .A2(n12951), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20041), .ZN(n12952) );
  NAND2_X1 U16186 ( .A1(n10297), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12977) );
  NAND2_X1 U16187 ( .A1(n12977), .A2(n9675), .ZN(n12953) );
  MUX2_X1 U16188 ( .A(n12953), .B(n12963), .S(n12954), .Z(n12966) );
  INV_X1 U16189 ( .A(n12954), .ZN(n12960) );
  INV_X1 U16190 ( .A(n12955), .ZN(n12958) );
  INV_X1 U16191 ( .A(n12956), .ZN(n12957) );
  OAI21_X1 U16192 ( .B1(n9676), .B2(n12958), .A(n12957), .ZN(n12959) );
  OAI21_X1 U16193 ( .B1(n9675), .B2(n12960), .A(n12959), .ZN(n12961) );
  NAND2_X1 U16194 ( .A1(n12961), .A2(n13056), .ZN(n12962) );
  OAI21_X1 U16195 ( .B1(n12964), .B2(n12963), .A(n12962), .ZN(n12965) );
  NAND2_X1 U16196 ( .A1(n12966), .A2(n12965), .ZN(n12969) );
  INV_X1 U16197 ( .A(n12967), .ZN(n12968) );
  NAND2_X1 U16198 ( .A1(n12969), .A2(n12968), .ZN(n12970) );
  OAI21_X1 U16199 ( .B1(n12971), .B2(n13082), .A(n12970), .ZN(n12975) );
  NAND2_X1 U16200 ( .A1(n12972), .A2(n13082), .ZN(n12973) );
  NAND3_X1 U16201 ( .A1(n12975), .A2(n12974), .A3(n12973), .ZN(n12976) );
  MUX2_X1 U16202 ( .A(n12976), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n16267), .Z(n13057) );
  NAND2_X1 U16203 ( .A1(n12978), .A2(n19416), .ZN(n12979) );
  OR2_X1 U16204 ( .A1(n12988), .A2(n10322), .ZN(n12983) );
  INV_X1 U16205 ( .A(n12981), .ZN(n12982) );
  NAND2_X1 U16206 ( .A1(n12983), .A2(n12982), .ZN(n13067) );
  NAND2_X1 U16207 ( .A1(n12984), .A2(n12989), .ZN(n12985) );
  NAND2_X1 U16208 ( .A1(n12985), .A2(n19539), .ZN(n12986) );
  NAND2_X1 U16209 ( .A1(n12987), .A2(n12986), .ZN(n12994) );
  AOI21_X1 U16210 ( .B1(n12988), .B2(n19549), .A(n13073), .ZN(n12993) );
  NAND2_X1 U16211 ( .A1(n12989), .A2(n10452), .ZN(n12995) );
  NAND2_X1 U16212 ( .A1(n12995), .A2(n13056), .ZN(n12990) );
  NAND2_X1 U16213 ( .A1(n12990), .A2(n10305), .ZN(n12991) );
  NAND2_X1 U16214 ( .A1(n12991), .A2(n19539), .ZN(n12992) );
  NAND4_X1 U16215 ( .A1(n13067), .A2(n12994), .A3(n12993), .A4(n12992), .ZN(
        n13017) );
  NOR2_X1 U16216 ( .A1(n13017), .A2(n12995), .ZN(n13404) );
  AND3_X1 U16217 ( .A1(n16590), .A2(n12996), .A3(n16591), .ZN(n12997) );
  AOI21_X1 U16218 ( .B1(n16597), .B2(n13404), .A(n12997), .ZN(n13020) );
  NAND2_X1 U16219 ( .A1(n12999), .A2(n12998), .ZN(n13076) );
  NAND2_X1 U16220 ( .A1(n13020), .A2(n13076), .ZN(n13000) );
  AOI21_X1 U16221 ( .B1(n20203), .B2(n19404), .A(n19400), .ZN(n13010) );
  INV_X1 U16222 ( .A(n13001), .ZN(n13002) );
  XNOR2_X1 U16223 ( .A(n13003), .B(n13002), .ZN(n19373) );
  INV_X1 U16224 ( .A(n19373), .ZN(n13009) );
  NOR2_X1 U16225 ( .A1(n10322), .A2(n10300), .ZN(n13005) );
  NAND2_X1 U16226 ( .A1(n19371), .A2(n13005), .ZN(n14624) );
  INV_X1 U16227 ( .A(n14624), .ZN(n13006) );
  INV_X1 U16228 ( .A(n19527), .ZN(n19337) );
  AOI22_X1 U16229 ( .A1(n19365), .A2(n19337), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19399), .ZN(n13008) );
  NAND3_X1 U16230 ( .A1(n19784), .A2(n19404), .A3(n13009), .ZN(n13007) );
  OAI211_X1 U16231 ( .C1(n13010), .C2(n13009), .A(n13008), .B(n13007), .ZN(
        P2_U2919) );
  NAND2_X1 U16232 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20200) );
  NOR2_X1 U16233 ( .A1(n16267), .A2(n20200), .ZN(n16610) );
  INV_X1 U16234 ( .A(n16597), .ZN(n13015) );
  INV_X1 U16235 ( .A(n13013), .ZN(n13014) );
  NAND2_X1 U16236 ( .A1(n13693), .A2(n13014), .ZN(n13405) );
  INV_X1 U16237 ( .A(n13405), .ZN(n16593) );
  NAND2_X1 U16238 ( .A1(n13015), .A2(n16593), .ZN(n13048) );
  NOR2_X1 U16239 ( .A1(n10330), .A2(n13016), .ZN(n13018) );
  AOI21_X1 U16240 ( .B1(n16590), .B2(n13018), .A(n13017), .ZN(n13055) );
  AND2_X1 U16241 ( .A1(n13048), .A2(n13055), .ZN(n13021) );
  NAND2_X1 U16242 ( .A1(n16597), .A2(n9675), .ZN(n19412) );
  INV_X1 U16243 ( .A(n19412), .ZN(n13060) );
  NAND3_X1 U16244 ( .A1(n13060), .A2(n19409), .A3(n13059), .ZN(n13019) );
  OAI22_X1 U16245 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20041), .B1(n16589), 
        .B2(n16622), .ZN(n13022) );
  AOI21_X1 U16246 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16610), .A(n13022), .ZN(
        n13850) );
  INV_X1 U16247 ( .A(n13850), .ZN(n13027) );
  NOR2_X1 U16248 ( .A1(n9676), .A2(n13023), .ZN(n13024) );
  NAND2_X1 U16249 ( .A1(n19409), .A2(n13024), .ZN(n16600) );
  OR3_X1 U16250 ( .A1(n13850), .A2(n13403), .A3(n16600), .ZN(n13025) );
  OAI21_X1 U16251 ( .B1(n13027), .B2(n13026), .A(n13025), .ZN(P2_U3595) );
  NAND2_X1 U16252 ( .A1(n12008), .A2(n13281), .ZN(n20239) );
  INV_X1 U16253 ( .A(n21050), .ZN(n20976) );
  AOI21_X1 U16254 ( .B1(n13029), .B2(n16262), .A(n20976), .ZN(n21053) );
  NOR2_X1 U16255 ( .A1(n20239), .A2(n21053), .ZN(n16226) );
  NOR2_X1 U16256 ( .A1(n16226), .A2(n20238), .ZN(n20245) );
  INV_X1 U16257 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13039) );
  NAND2_X1 U16258 ( .A1(n13248), .A2(n13637), .ZN(n13283) );
  OR2_X1 U16259 ( .A1(n13194), .A2(n13030), .ZN(n16229) );
  AND2_X1 U16260 ( .A1(n13224), .A2(n16229), .ZN(n13300) );
  NAND3_X1 U16261 ( .A1(n13031), .A2(n13205), .A3(n13310), .ZN(n13032) );
  NAND2_X1 U16262 ( .A1(n13300), .A2(n13032), .ZN(n13033) );
  MUX2_X1 U16263 ( .A(n13308), .B(n13033), .S(n13285), .Z(n13035) );
  NOR2_X1 U16264 ( .A1(n13281), .A2(n12009), .ZN(n13034) );
  OR2_X1 U16265 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  NAND2_X1 U16266 ( .A1(n13036), .A2(n11165), .ZN(n16228) );
  INV_X1 U16267 ( .A(n16228), .ZN(n13037) );
  NAND2_X1 U16268 ( .A1(n20245), .A2(n13037), .ZN(n13038) );
  OAI21_X1 U16269 ( .B1(n20245), .B2(n13039), .A(n13038), .ZN(P1_U3484) );
  NOR2_X1 U16270 ( .A1(n13209), .A2(n9656), .ZN(n13041) );
  OAI21_X1 U16271 ( .B1(n13964), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n21047), 
        .ZN(n13040) );
  OAI21_X1 U16272 ( .B1(n21047), .B2(n13041), .A(n13040), .ZN(P1_U3487) );
  NAND2_X1 U16273 ( .A1(n19506), .A2(n13147), .ZN(n13043) );
  NAND2_X1 U16274 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19888) );
  OAI21_X1 U16275 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n19888), .ZN(n19659) );
  NOR2_X1 U16276 ( .A1(n19659), .A2(n20183), .ZN(n19857) );
  AOI21_X1 U16277 ( .B1(n13160), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19857), .ZN(n13042) );
  NAND2_X1 U16278 ( .A1(n13043), .A2(n13042), .ZN(n13045) );
  NOR2_X1 U16279 ( .A1(n14477), .A2(n10442), .ZN(n13156) );
  NAND2_X1 U16280 ( .A1(n13045), .A2(n13044), .ZN(n13046) );
  NAND2_X1 U16281 ( .A1(n10315), .A2(n13047), .ZN(n13808) );
  NAND2_X1 U16282 ( .A1(n13048), .A2(n13808), .ZN(n13049) );
  NAND2_X1 U16283 ( .A1(n15572), .A2(n10305), .ZN(n15594) );
  MUX2_X1 U16284 ( .A(n13708), .B(n13845), .S(n15572), .Z(n13050) );
  OAI21_X1 U16285 ( .B1(n19657), .B2(n15594), .A(n13050), .ZN(P2_U2886) );
  INV_X1 U16286 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19497) );
  INV_X1 U16287 ( .A(n13051), .ZN(n13064) );
  MUX2_X1 U16288 ( .A(n19539), .B(n10330), .S(n9675), .Z(n13052) );
  NOR2_X1 U16289 ( .A1(n13052), .A2(n20114), .ZN(n13053) );
  NAND2_X1 U16290 ( .A1(n16590), .A2(n13053), .ZN(n13054) );
  AND2_X1 U16291 ( .A1(n13055), .A2(n13054), .ZN(n13063) );
  AOI21_X1 U16292 ( .B1(n13057), .B2(n13056), .A(n19549), .ZN(n13058) );
  NAND2_X1 U16293 ( .A1(n19412), .A2(n13058), .ZN(n13062) );
  NAND3_X1 U16294 ( .A1(n13060), .A2(n13069), .A3(n13059), .ZN(n13061) );
  NAND4_X1 U16295 ( .A1(n13064), .A2(n13063), .A3(n13062), .A4(n13061), .ZN(
        n13065) );
  OR2_X1 U16296 ( .A1(n13066), .A2(n10452), .ZN(n13695) );
  NAND2_X1 U16297 ( .A1(n13695), .A2(n13067), .ZN(n13079) );
  NAND2_X1 U16298 ( .A1(n10308), .A2(n19549), .ZN(n13071) );
  AOI22_X1 U16299 ( .A1(n13071), .A2(n13070), .B1(n10297), .B2(n13069), .ZN(
        n13075) );
  NAND3_X1 U16300 ( .A1(n10318), .A2(n13073), .A3(n13072), .ZN(n13074) );
  NAND4_X1 U16301 ( .A1(n13068), .A2(n13076), .A3(n13075), .A4(n13074), .ZN(
        n13077) );
  AOI21_X1 U16302 ( .B1(n13079), .B2(n13078), .A(n13077), .ZN(n13844) );
  NAND2_X1 U16303 ( .A1(n13844), .A2(n13808), .ZN(n13080) );
  INV_X1 U16304 ( .A(n13081), .ZN(n20212) );
  AND2_X1 U16305 ( .A1(n16598), .A2(n13082), .ZN(n20210) );
  OAI22_X1 U16306 ( .A1(n19515), .A2(n13084), .B1(n19502), .B2(n13083), .ZN(
        n13095) );
  OR2_X1 U16307 ( .A1(n13091), .A2(n19303), .ZN(n19501) );
  NAND2_X1 U16308 ( .A1(n16591), .A2(n9676), .ZN(n13085) );
  NAND2_X1 U16309 ( .A1(n13405), .A2(n13085), .ZN(n13086) );
  NAND2_X2 U16310 ( .A1(n13091), .A2(n13086), .ZN(n19508) );
  INV_X1 U16311 ( .A(n19508), .ZN(n16544) );
  NAND2_X1 U16312 ( .A1(n13087), .A2(n10452), .ZN(n13089) );
  NAND2_X1 U16313 ( .A1(n13089), .A2(n13809), .ZN(n13090) );
  AOI22_X1 U16314 ( .A1(n16544), .A2(n19373), .B1(n19505), .B2(n19314), .ZN(
        n13093) );
  OAI211_X1 U16315 ( .C1(n19497), .C2(n19501), .A(n13093), .B(n13092), .ZN(
        n13094) );
  AOI211_X1 U16316 ( .C1(n19497), .C2(n19499), .A(n13095), .B(n13094), .ZN(
        n13096) );
  INV_X1 U16317 ( .A(n13096), .ZN(P2_U3046) );
  AND2_X1 U16318 ( .A1(n14094), .A2(n20976), .ZN(n13097) );
  INV_X1 U16319 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14974) );
  NAND2_X1 U16320 ( .A1(n13114), .A2(n13637), .ZN(n13110) );
  INV_X1 U16321 ( .A(DATAI_15_), .ZN(n13100) );
  INV_X1 U16322 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13099) );
  MUX2_X1 U16323 ( .A(n13100), .B(n13099), .S(n20419), .Z(n14973) );
  INV_X1 U16324 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13101) );
  OAI222_X1 U16325 ( .A1(n13357), .A2(n14974), .B1(n13110), .B2(n14973), .C1(
        n13114), .C2(n13101), .ZN(P1_U2967) );
  OAI21_X1 U16326 ( .B1(n13103), .B2(n13102), .A(n13426), .ZN(n13943) );
  NAND2_X1 U16327 ( .A1(n13285), .A2(n13308), .ZN(n13198) );
  NAND4_X1 U16328 ( .A1(n13107), .A2(n13104), .A3(n20450), .A4(n11172), .ZN(
        n13105) );
  NAND2_X1 U16329 ( .A1(n13198), .A2(n13105), .ZN(n13106) );
  XNOR2_X1 U16330 ( .A(n13108), .B(n13107), .ZN(n20405) );
  AOI22_X1 U16331 ( .A1(n20351), .A2(n20405), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14885), .ZN(n13109) );
  OAI21_X1 U16332 ( .B1(n13943), .B2(n14890), .A(n13109), .ZN(P1_U2871) );
  INV_X1 U16333 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14966) );
  NAND2_X1 U16334 ( .A1(n20421), .A2(DATAI_0_), .ZN(n13112) );
  NAND2_X1 U16335 ( .A1(n20419), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13111) );
  AND2_X1 U16336 ( .A1(n13112), .A2(n13111), .ZN(n20428) );
  INV_X1 U16337 ( .A(n20428), .ZN(n13113) );
  NAND2_X1 U16338 ( .A1(n13388), .A2(n13113), .ZN(n13394) );
  NAND2_X1 U16339 ( .A1(n13366), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13115) );
  OAI211_X1 U16340 ( .C1(n14966), .C2(n13357), .A(n13394), .B(n13115), .ZN(
        P1_U2937) );
  INV_X1 U16341 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n13773) );
  INV_X1 U16342 ( .A(DATAI_14_), .ZN(n13117) );
  NAND2_X1 U16343 ( .A1(n20419), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13116) );
  OAI21_X1 U16344 ( .B1(n20419), .B2(n13117), .A(n13116), .ZN(n14976) );
  NAND2_X1 U16345 ( .A1(n13388), .A2(n14976), .ZN(n13123) );
  NAND2_X1 U16346 ( .A1(n13366), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n13118) );
  OAI211_X1 U16347 ( .C1(n13773), .C2(n13357), .A(n13123), .B(n13118), .ZN(
        P1_U2966) );
  INV_X1 U16348 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13490) );
  INV_X1 U16349 ( .A(DATAI_11_), .ZN(n13120) );
  NAND2_X1 U16350 ( .A1(n20419), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13119) );
  OAI21_X1 U16351 ( .B1(n20419), .B2(n13120), .A(n13119), .ZN(n14992) );
  NAND2_X1 U16352 ( .A1(n13388), .A2(n14992), .ZN(n13137) );
  NAND2_X1 U16353 ( .A1(n13366), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13121) );
  OAI211_X1 U16354 ( .C1(n13490), .C2(n13357), .A(n13137), .B(n13121), .ZN(
        P1_U2948) );
  INV_X1 U16355 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13498) );
  NAND2_X1 U16356 ( .A1(n13366), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13122) );
  OAI211_X1 U16357 ( .C1(n13498), .C2(n13357), .A(n13123), .B(n13122), .ZN(
        P1_U2951) );
  INV_X1 U16358 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13503) );
  INV_X1 U16359 ( .A(DATAI_13_), .ZN(n21085) );
  NAND2_X1 U16360 ( .A1(n20419), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13124) );
  OAI21_X1 U16361 ( .B1(n20419), .B2(n21085), .A(n13124), .ZN(n14978) );
  NAND2_X1 U16362 ( .A1(n13388), .A2(n14978), .ZN(n13130) );
  NAND2_X1 U16363 ( .A1(n13366), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13125) );
  OAI211_X1 U16364 ( .C1(n13503), .C2(n13357), .A(n13130), .B(n13125), .ZN(
        P1_U2950) );
  INV_X1 U16365 ( .A(DATAI_12_), .ZN(n13127) );
  NAND2_X1 U16366 ( .A1(n20419), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13126) );
  OAI21_X1 U16367 ( .B1(n20419), .B2(n13127), .A(n13126), .ZN(n14985) );
  NAND2_X1 U16368 ( .A1(n13388), .A2(n14985), .ZN(n13142) );
  NAND2_X1 U16369 ( .A1(n13366), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n13128) );
  OAI211_X1 U16370 ( .C1(n14989), .C2(n13357), .A(n13142), .B(n13128), .ZN(
        P1_U2964) );
  INV_X1 U16371 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n13767) );
  NAND2_X1 U16372 ( .A1(n13366), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n13129) );
  OAI211_X1 U16373 ( .C1(n13767), .C2(n13357), .A(n13130), .B(n13129), .ZN(
        P1_U2965) );
  INV_X1 U16374 ( .A(DATAI_10_), .ZN(n13132) );
  NAND2_X1 U16375 ( .A1(n20419), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13131) );
  OAI21_X1 U16376 ( .B1(n20419), .B2(n13132), .A(n13131), .ZN(n14911) );
  NAND2_X1 U16377 ( .A1(n13388), .A2(n14911), .ZN(n13135) );
  NAND2_X1 U16378 ( .A1(n13366), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13133) );
  OAI211_X1 U16379 ( .C1(n11849), .C2(n13357), .A(n13135), .B(n13133), .ZN(
        P1_U2947) );
  INV_X1 U16380 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13776) );
  NAND2_X1 U16381 ( .A1(n13366), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n13134) );
  OAI211_X1 U16382 ( .C1(n13776), .C2(n13357), .A(n13135), .B(n13134), .ZN(
        P1_U2962) );
  INV_X1 U16383 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13764) );
  NAND2_X1 U16384 ( .A1(n13366), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n13136) );
  OAI211_X1 U16385 ( .C1(n13764), .C2(n13357), .A(n13137), .B(n13136), .ZN(
        P1_U2963) );
  INV_X1 U16386 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13761) );
  INV_X1 U16387 ( .A(DATAI_9_), .ZN(n13139) );
  NAND2_X1 U16388 ( .A1(n20419), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13138) );
  OAI21_X1 U16389 ( .B1(n20419), .B2(n13139), .A(n13138), .ZN(n14917) );
  NAND2_X1 U16390 ( .A1(n13388), .A2(n14917), .ZN(n13144) );
  NAND2_X1 U16391 ( .A1(n13366), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n13140) );
  OAI211_X1 U16392 ( .C1(n13761), .C2(n13357), .A(n13144), .B(n13140), .ZN(
        P1_U2961) );
  NAND2_X1 U16393 ( .A1(n13366), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13141) );
  OAI211_X1 U16394 ( .C1(n11901), .C2(n13357), .A(n13142), .B(n13141), .ZN(
        P1_U2949) );
  INV_X1 U16395 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13487) );
  NAND2_X1 U16396 ( .A1(n13366), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13143) );
  OAI211_X1 U16397 ( .C1(n13487), .C2(n13357), .A(n13144), .B(n13143), .ZN(
        P1_U2946) );
  NAND2_X1 U16398 ( .A1(n13454), .A2(n13147), .ZN(n13151) );
  NOR2_X1 U16399 ( .A1(n20190), .A2(n20199), .ZN(n19987) );
  INV_X1 U16400 ( .A(n20085), .ZN(n20029) );
  NOR2_X1 U16401 ( .A1(n13161), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13148) );
  NOR2_X1 U16402 ( .A1(n13148), .A2(n20183), .ZN(n13149) );
  AND2_X1 U16403 ( .A1(n20029), .A2(n13149), .ZN(n19921) );
  AOI21_X1 U16404 ( .B1(n13160), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19921), .ZN(n13150) );
  NAND2_X1 U16405 ( .A1(n13151), .A2(n13150), .ZN(n13152) );
  NAND2_X1 U16406 ( .A1(n13152), .A2(n13153), .ZN(n13176) );
  OAI21_X1 U16407 ( .B1(n13153), .B2(n13152), .A(n13176), .ZN(n13154) );
  INV_X1 U16408 ( .A(n13155), .ZN(n13701) );
  INV_X1 U16409 ( .A(n13156), .ZN(n13157) );
  NAND2_X1 U16410 ( .A1(n13701), .A2(n13157), .ZN(n13158) );
  NAND2_X1 U16411 ( .A1(n13160), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13170) );
  NAND2_X1 U16412 ( .A1(n19888), .A2(n20190), .ZN(n13163) );
  INV_X1 U16413 ( .A(n13161), .ZN(n13162) );
  NAND2_X1 U16414 ( .A1(n13163), .A2(n13162), .ZN(n19660) );
  OR2_X1 U16415 ( .A1(n19660), .A2(n20183), .ZN(n13169) );
  NAND2_X1 U16416 ( .A1(n13170), .A2(n13169), .ZN(n13166) );
  NAND4_X1 U16417 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A3(
        P2_STATE2_REG_0__SCAN_IN), .A4(n9676), .ZN(n13164) );
  OR2_X1 U16418 ( .A1(n13166), .A2(n13167), .ZN(n13165) );
  NAND2_X1 U16419 ( .A1(n13166), .A2(n13167), .ZN(n13174) );
  NAND4_X1 U16420 ( .A1(n13164), .A2(n13170), .A3(n13169), .A4(n13168), .ZN(
        n13171) );
  AND2_X1 U16421 ( .A1(n13174), .A2(n13171), .ZN(n13172) );
  NAND2_X1 U16422 ( .A1(n13259), .A2(n13260), .ZN(n13261) );
  NAND2_X1 U16423 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10306), .ZN(
        n13175) );
  NOR2_X1 U16424 ( .A1(n14477), .A2(n13178), .ZN(n13179) );
  NAND2_X1 U16425 ( .A1(n13347), .A2(n13179), .ZN(n13272) );
  OR2_X1 U16426 ( .A1(n13347), .A2(n13179), .ZN(n13180) );
  NAND2_X1 U16427 ( .A1(n13272), .A2(n13180), .ZN(n19382) );
  NAND2_X1 U16428 ( .A1(n13183), .A2(n13182), .ZN(n13184) );
  AND2_X1 U16429 ( .A1(n13181), .A2(n13184), .ZN(n19487) );
  NOR2_X1 U16430 ( .A1(n15572), .A2(n13185), .ZN(n13186) );
  AOI21_X1 U16431 ( .B1(n19487), .B2(n15572), .A(n13186), .ZN(n13187) );
  OAI21_X1 U16432 ( .B1(n19382), .B2(n15594), .A(n13187), .ZN(P2_U2883) );
  OR3_X1 U16433 ( .A1(n13285), .A2(n20976), .A3(n16262), .ZN(n16236) );
  NAND2_X1 U16434 ( .A1(n13188), .A2(n16236), .ZN(n13191) );
  NOR2_X1 U16435 ( .A1(n12009), .A2(n11968), .ZN(n16211) );
  NAND2_X1 U16436 ( .A1(n13224), .A2(n12149), .ZN(n13189) );
  OR2_X1 U16437 ( .A1(n16211), .A2(n13189), .ZN(n13190) );
  NAND2_X1 U16438 ( .A1(n13191), .A2(n13190), .ZN(n13200) );
  AND2_X1 U16439 ( .A1(n13283), .A2(n13310), .ZN(n13192) );
  AND2_X1 U16440 ( .A1(n13193), .A2(n13192), .ZN(n13208) );
  AOI21_X1 U16441 ( .B1(n12009), .B2(n13194), .A(n13208), .ZN(n13286) );
  OAI211_X1 U16442 ( .C1(n13852), .C2(n9954), .A(n13195), .B(n13286), .ZN(
        n13196) );
  INV_X1 U16443 ( .A(n13196), .ZN(n13197) );
  AND2_X1 U16444 ( .A1(n13198), .A2(n13197), .ZN(n13199) );
  INV_X1 U16445 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21176) );
  NAND2_X1 U16446 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16432) );
  INV_X1 U16447 ( .A(n16432), .ZN(n16427) );
  NAND2_X1 U16448 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16427), .ZN(n13590) );
  OR2_X1 U16449 ( .A1(n21176), .A2(n13590), .ZN(n13201) );
  OAI21_X1 U16450 ( .B1(n13583), .B2(n20238), .A(n13201), .ZN(n16418) );
  AOI21_X1 U16451 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20963), .A(n16418), 
        .ZN(n16417) );
  OAI211_X1 U16452 ( .C1(n13206), .C2(n13205), .A(n13204), .B(n13203), .ZN(
        n13207) );
  NOR2_X1 U16453 ( .A1(n13208), .A2(n13207), .ZN(n13212) );
  NAND2_X1 U16454 ( .A1(n13210), .A2(n13209), .ZN(n13211) );
  AND2_X1 U16455 ( .A1(n13212), .A2(n13211), .ZN(n13315) );
  AND3_X1 U16456 ( .A1(n13213), .A2(n12149), .A3(n13311), .ZN(n13214) );
  AND2_X1 U16457 ( .A1(n13315), .A2(n13214), .ZN(n13218) );
  NAND2_X1 U16458 ( .A1(n9954), .A2(n13293), .ZN(n13215) );
  OAI21_X1 U16459 ( .B1(n9731), .B2(n13310), .A(n13215), .ZN(n13313) );
  NOR2_X1 U16460 ( .A1(n13313), .A2(n11172), .ZN(n13216) );
  MUX2_X1 U16461 ( .A(n12009), .B(n13216), .S(n13637), .Z(n13217) );
  NAND2_X1 U16462 ( .A1(n13218), .A2(n13217), .ZN(n13580) );
  INV_X1 U16463 ( .A(n13219), .ZN(n13222) );
  INV_X1 U16464 ( .A(n11008), .ZN(n13220) );
  NAND2_X1 U16465 ( .A1(n13220), .A2(n11302), .ZN(n13221) );
  NAND2_X1 U16466 ( .A1(n13222), .A2(n13221), .ZN(n13227) );
  INV_X1 U16467 ( .A(n13227), .ZN(n13231) );
  NAND2_X1 U16468 ( .A1(n11172), .A2(n13231), .ZN(n13230) );
  INV_X1 U16469 ( .A(n13580), .ZN(n15413) );
  OR2_X1 U16470 ( .A1(n13223), .A2(n15413), .ZN(n13229) );
  INV_X1 U16471 ( .A(n13224), .ZN(n13225) );
  OR2_X1 U16472 ( .A1(n13308), .A2(n13225), .ZN(n13573) );
  XNOR2_X1 U16473 ( .A(n10996), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13226) );
  AOI22_X1 U16474 ( .A1(n13573), .A2(n13227), .B1(n16211), .B2(n13226), .ZN(
        n13228) );
  OAI211_X1 U16475 ( .C1(n13580), .C2(n13230), .A(n13229), .B(n13228), .ZN(
        n13582) );
  INV_X1 U16476 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14018) );
  NOR2_X1 U16477 ( .A1(n20962), .A2(n14018), .ZN(n15417) );
  INV_X1 U16478 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21205) );
  OAI22_X1 U16479 ( .A1(n21205), .A2(n9877), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15418) );
  INV_X1 U16480 ( .A(n15418), .ZN(n13232) );
  INV_X1 U16481 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20674) );
  AOI222_X1 U16482 ( .A1(n13582), .A2(n16419), .B1(n15417), .B2(n13232), .C1(
        n13231), .C2(n16247), .ZN(n13234) );
  NAND2_X1 U16483 ( .A1(n16417), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13233) );
  OAI21_X1 U16484 ( .B1(n16417), .B2(n13234), .A(n13233), .ZN(P1_U3472) );
  MUX2_X1 U16485 ( .A(n13699), .B(n13235), .S(n15592), .Z(n13236) );
  OAI21_X1 U16486 ( .B1(n20203), .B2(n15594), .A(n13236), .ZN(P2_U2887) );
  INV_X1 U16487 ( .A(n13237), .ZN(n13238) );
  NAND2_X1 U16488 ( .A1(n13239), .A2(n13238), .ZN(n13241) );
  MUX2_X1 U16489 ( .A(n14655), .B(n10358), .S(n15592), .Z(n13242) );
  OAI21_X1 U16490 ( .B1(n19520), .B2(n15594), .A(n13242), .ZN(P2_U2885) );
  XOR2_X1 U16491 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13272), .Z(n13247)
         );
  AND2_X1 U16492 ( .A1(n13181), .A2(n13243), .ZN(n13244) );
  OR2_X1 U16493 ( .A1(n13276), .A2(n13244), .ZN(n16534) );
  MUX2_X1 U16494 ( .A(n16534), .B(n13245), .S(n15592), .Z(n13246) );
  OAI21_X1 U16495 ( .B1(n13247), .B2(n15594), .A(n13246), .ZN(P2_U2882) );
  OR2_X1 U16496 ( .A1(n13248), .A2(n20457), .ZN(n13249) );
  INV_X1 U16497 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n13524) );
  NAND2_X1 U16498 ( .A1(n20421), .A2(DATAI_1_), .ZN(n13251) );
  NAND2_X1 U16499 ( .A1(n20419), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13250) );
  AND2_X1 U16500 ( .A1(n13251), .A2(n13250), .ZN(n20435) );
  OAI222_X1 U16501 ( .A1(n14995), .A2(n13943), .B1(n14988), .B2(n13524), .C1(
        n14987), .C2(n20435), .ZN(P1_U2903) );
  INV_X1 U16502 ( .A(n13252), .ZN(n13255) );
  OAI21_X1 U16503 ( .B1(n13255), .B2(n13254), .A(n13253), .ZN(n13927) );
  INV_X1 U16504 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n13784) );
  OAI222_X1 U16505 ( .A1(n14995), .A2(n13927), .B1(n14988), .B2(n13784), .C1(
        n14987), .C2(n20428), .ZN(P1_U2904) );
  NAND2_X1 U16506 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13342) );
  NOR2_X1 U16507 ( .A1(n13272), .A2(n13342), .ZN(n13416) );
  XNOR2_X1 U16508 ( .A(n13416), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13258) );
  AOI21_X1 U16509 ( .B1(n13256), .B2(n13277), .A(n13527), .ZN(n16559) );
  INV_X1 U16510 ( .A(n16559), .ZN(n19279) );
  MUX2_X1 U16511 ( .A(n19279), .B(n10813), .S(n15592), .Z(n13257) );
  OAI21_X1 U16512 ( .B1(n13258), .B2(n15594), .A(n13257), .ZN(P2_U2880) );
  NOR2_X1 U16513 ( .A1(n13263), .A2(n15592), .ZN(n13264) );
  AOI21_X1 U16514 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n15592), .A(n13264), .ZN(
        n13265) );
  OAI21_X1 U16515 ( .B1(n20177), .B2(n15594), .A(n13265), .ZN(P2_U2884) );
  INV_X1 U16516 ( .A(n13852), .ZN(n13266) );
  INV_X1 U16517 ( .A(n16262), .ZN(n13282) );
  NAND2_X1 U16518 ( .A1(n13266), .A2(n13282), .ZN(n13269) );
  NOR2_X1 U16519 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16432), .ZN(n21051) );
  AOI222_X1 U16520 ( .A1(n13512), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n16264), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .C1(n21051), .C2(P1_LWORD_REG_4__SCAN_IN), .ZN(n13270) );
  INV_X1 U16521 ( .A(n13270), .ZN(P1_U2932) );
  NOR2_X1 U16522 ( .A1(n13272), .A2(n13271), .ZN(n13274) );
  INV_X1 U16523 ( .A(n13416), .ZN(n13273) );
  OAI211_X1 U16524 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13274), .A(
        n13273), .B(n15575), .ZN(n13280) );
  OR2_X1 U16525 ( .A1(n13276), .A2(n13275), .ZN(n13278) );
  NAND2_X1 U16526 ( .A1(n13278), .A2(n13277), .ZN(n19293) );
  INV_X1 U16527 ( .A(n19293), .ZN(n14084) );
  NAND2_X1 U16528 ( .A1(n14084), .A2(n15572), .ZN(n13279) );
  OAI211_X1 U16529 ( .C1(n15572), .C2(n19284), .A(n13280), .B(n13279), .ZN(
        P2_U2881) );
  INV_X1 U16530 ( .A(n13281), .ZN(n13289) );
  OAI211_X1 U16531 ( .C1(n11968), .C2(n13282), .A(n9954), .B(n21050), .ZN(
        n13288) );
  INV_X1 U16532 ( .A(n13283), .ZN(n13284) );
  NAND2_X1 U16533 ( .A1(n13285), .A2(n13284), .ZN(n13287) );
  OAI211_X1 U16534 ( .C1(n13289), .C2(n13288), .A(n13287), .B(n13286), .ZN(
        n13291) );
  NAND2_X1 U16535 ( .A1(n13291), .A2(n13290), .ZN(n13298) );
  NAND2_X1 U16536 ( .A1(n13292), .A2(n21050), .ZN(n13294) );
  OAI211_X1 U16537 ( .C1(n12149), .C2(n13294), .A(n13310), .B(n13293), .ZN(
        n13295) );
  NAND2_X1 U16538 ( .A1(n13295), .A2(n20438), .ZN(n13296) );
  OAI211_X1 U16539 ( .C1(n20446), .C2(n13322), .A(n9670), .B(n13300), .ZN(
        n13301) );
  NAND2_X1 U16540 ( .A1(n11170), .A2(n13303), .ZN(n13657) );
  OAI21_X1 U16541 ( .B1(n14094), .B2(n13641), .A(n13657), .ZN(n13304) );
  INV_X1 U16542 ( .A(n13304), .ZN(n13305) );
  NAND2_X1 U16543 ( .A1(n13306), .A2(n13305), .ZN(n13307) );
  OAI21_X1 U16544 ( .B1(n13307), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13646), .ZN(n13331) );
  NAND2_X1 U16545 ( .A1(n13324), .A2(n13308), .ZN(n20370) );
  OR2_X1 U16546 ( .A1(n13324), .A2(n20407), .ZN(n13318) );
  OAI21_X1 U16547 ( .B1(n10038), .B2(n13637), .A(n11172), .ZN(n13309) );
  OAI21_X1 U16548 ( .B1(n13311), .B2(n13310), .A(n13309), .ZN(n13312) );
  AOI21_X1 U16549 ( .B1(n13637), .B2(n13313), .A(n13312), .ZN(n13314) );
  NAND2_X1 U16550 ( .A1(n13315), .A2(n13314), .ZN(n13316) );
  NAND2_X1 U16551 ( .A1(n13324), .A2(n13316), .ZN(n14016) );
  NOR2_X1 U16552 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14016), .ZN(
        n13319) );
  INV_X1 U16553 ( .A(n13319), .ZN(n13317) );
  INV_X1 U16554 ( .A(n20371), .ZN(n14019) );
  AOI21_X1 U16555 ( .B1(n20390), .B2(n14018), .A(n14019), .ZN(n20416) );
  NAND2_X1 U16556 ( .A1(n13324), .A2(n16211), .ZN(n16364) );
  NOR3_X1 U16557 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20390), .A3(
        n13319), .ZN(n13320) );
  AOI21_X1 U16558 ( .B1(n20416), .B2(n16364), .A(n13320), .ZN(n13321) );
  INV_X1 U16559 ( .A(n13321), .ZN(n13329) );
  OAI22_X1 U16560 ( .A1(n13322), .A2(n11168), .B1(n12149), .B2(n14094), .ZN(
        n13323) );
  NOR2_X1 U16561 ( .A1(n13325), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13327) );
  OR2_X1 U16562 ( .A1(n13327), .A2(n13326), .ZN(n13356) );
  INV_X1 U16563 ( .A(n13356), .ZN(n13925) );
  INV_X1 U16564 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13921) );
  NOR2_X1 U16565 ( .A1(n20393), .A2(n13921), .ZN(n13338) );
  AOI21_X1 U16566 ( .B1(n20406), .B2(n13925), .A(n13338), .ZN(n13328) );
  OAI211_X1 U16567 ( .C1(n20408), .C2(n13331), .A(n13329), .B(n13328), .ZN(
        P1_U3031) );
  NAND3_X1 U16568 ( .A1(n20963), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16425) );
  INV_X1 U16569 ( .A(n16425), .ZN(n13330) );
  INV_X1 U16570 ( .A(n13331), .ZN(n13339) );
  INV_X1 U16571 ( .A(n20909), .ZN(n20903) );
  NAND2_X1 U16572 ( .A1(n20903), .A2(n13333), .ZN(n21049) );
  NAND2_X1 U16573 ( .A1(n21049), .A2(n20963), .ZN(n13334) );
  NAND2_X1 U16574 ( .A1(n20963), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16237) );
  NAND2_X1 U16575 ( .A1(n20852), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13335) );
  AND2_X1 U16576 ( .A1(n16237), .A2(n13335), .ZN(n13648) );
  INV_X1 U16577 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13336) );
  AOI21_X1 U16578 ( .B1(n15201), .B2(n13648), .A(n13336), .ZN(n13337) );
  AOI211_X1 U16579 ( .C1(n13339), .C2(n16345), .A(n13338), .B(n13337), .ZN(
        n13340) );
  OAI21_X1 U16580 ( .B1(n20422), .B2(n13927), .A(n13340), .ZN(P1_U2999) );
  NAND2_X1 U16581 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13341) );
  NOR2_X1 U16582 ( .A1(n13342), .A2(n13341), .ZN(n13343) );
  NAND3_X1 U16583 ( .A1(n13344), .A2(n13417), .A3(n13343), .ZN(n13345) );
  NOR2_X1 U16584 ( .A1(n14477), .A2(n13345), .ZN(n13346) );
  INV_X1 U16585 ( .A(n13348), .ZN(n13351) );
  INV_X1 U16586 ( .A(n13349), .ZN(n13350) );
  OAI211_X1 U16587 ( .C1(n13351), .C2(n13350), .A(n15575), .B(n13437), .ZN(
        n13355) );
  OR2_X1 U16588 ( .A1(n13352), .A2(n13419), .ZN(n13353) );
  AND2_X1 U16589 ( .A1(n13353), .A2(n13507), .ZN(n16510) );
  NAND2_X1 U16590 ( .A1(n15572), .A2(n16510), .ZN(n13354) );
  OAI211_X1 U16591 ( .C1(n15572), .C2(n10704), .A(n13355), .B(n13354), .ZN(
        P2_U2877) );
  OAI222_X1 U16592 ( .A1(n13927), .A2(n14890), .B1(n13920), .B2(n20356), .C1(
        n13356), .C2(n14896), .ZN(P1_U2872) );
  AOI22_X1 U16593 ( .A1(n13400), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n13366), .ZN(n13358) );
  INV_X1 U16594 ( .A(n20435), .ZN(n14958) );
  NAND2_X1 U16595 ( .A1(n13388), .A2(n14958), .ZN(n13372) );
  NAND2_X1 U16596 ( .A1(n13358), .A2(n13372), .ZN(P1_U2953) );
  AOI22_X1 U16597 ( .A1(n13400), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n13366), .ZN(n13361) );
  NAND2_X1 U16598 ( .A1(n20421), .A2(DATAI_2_), .ZN(n13360) );
  NAND2_X1 U16599 ( .A1(n20419), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13359) );
  AND2_X1 U16600 ( .A1(n13360), .A2(n13359), .ZN(n20439) );
  INV_X1 U16601 ( .A(n20439), .ZN(n14951) );
  NAND2_X1 U16602 ( .A1(n13388), .A2(n14951), .ZN(n13384) );
  NAND2_X1 U16603 ( .A1(n13361), .A2(n13384), .ZN(P1_U2954) );
  AOI22_X1 U16604 ( .A1(n13400), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n13366), .ZN(n13365) );
  NAND2_X1 U16605 ( .A1(n20421), .A2(DATAI_4_), .ZN(n13363) );
  NAND2_X1 U16606 ( .A1(n20419), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13362) );
  AND2_X1 U16607 ( .A1(n13363), .A2(n13362), .ZN(n20447) );
  INV_X1 U16608 ( .A(n20447), .ZN(n13364) );
  NAND2_X1 U16609 ( .A1(n13388), .A2(n13364), .ZN(n13367) );
  NAND2_X1 U16610 ( .A1(n13365), .A2(n13367), .ZN(P1_U2956) );
  AOI22_X1 U16611 ( .A1(n13400), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n13366), .ZN(n13368) );
  NAND2_X1 U16612 ( .A1(n13368), .A2(n13367), .ZN(P1_U2941) );
  AOI22_X1 U16613 ( .A1(n13400), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n13366), .ZN(n13371) );
  INV_X1 U16614 ( .A(DATAI_6_), .ZN(n13370) );
  NAND2_X1 U16615 ( .A1(n20419), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13369) );
  OAI21_X1 U16616 ( .B1(n20419), .B2(n13370), .A(n13369), .ZN(n14932) );
  NAND2_X1 U16617 ( .A1(n13388), .A2(n14932), .ZN(n13401) );
  NAND2_X1 U16618 ( .A1(n13371), .A2(n13401), .ZN(P1_U2943) );
  AOI22_X1 U16619 ( .A1(n13400), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n13366), .ZN(n13373) );
  NAND2_X1 U16620 ( .A1(n13373), .A2(n13372), .ZN(P1_U2938) );
  AOI22_X1 U16621 ( .A1(n13400), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n13366), .ZN(n13377) );
  NAND2_X1 U16622 ( .A1(n20421), .A2(DATAI_3_), .ZN(n13375) );
  NAND2_X1 U16623 ( .A1(n20419), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13374) );
  AND2_X1 U16624 ( .A1(n13375), .A2(n13374), .ZN(n20443) );
  INV_X1 U16625 ( .A(n20443), .ZN(n13376) );
  NAND2_X1 U16626 ( .A1(n13388), .A2(n13376), .ZN(n13392) );
  NAND2_X1 U16627 ( .A1(n13377), .A2(n13392), .ZN(P1_U2955) );
  AOI22_X1 U16628 ( .A1(n13400), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n13366), .ZN(n13380) );
  INV_X1 U16629 ( .A(DATAI_5_), .ZN(n13379) );
  NAND2_X1 U16630 ( .A1(n20419), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13378) );
  OAI21_X1 U16631 ( .B1(n20419), .B2(n13379), .A(n13378), .ZN(n14937) );
  NAND2_X1 U16632 ( .A1(n13388), .A2(n14937), .ZN(n13398) );
  NAND2_X1 U16633 ( .A1(n13380), .A2(n13398), .ZN(P1_U2942) );
  AOI22_X1 U16634 ( .A1(n13400), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n13366), .ZN(n13383) );
  INV_X1 U16635 ( .A(DATAI_8_), .ZN(n13382) );
  NAND2_X1 U16636 ( .A1(n20419), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13381) );
  OAI21_X1 U16637 ( .B1(n20419), .B2(n13382), .A(n13381), .ZN(n14922) );
  NAND2_X1 U16638 ( .A1(n13388), .A2(n14922), .ZN(n13390) );
  NAND2_X1 U16639 ( .A1(n13383), .A2(n13390), .ZN(P1_U2945) );
  AOI22_X1 U16640 ( .A1(n13400), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n13366), .ZN(n13385) );
  NAND2_X1 U16641 ( .A1(n13385), .A2(n13384), .ZN(P1_U2939) );
  AOI22_X1 U16642 ( .A1(n13400), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n13366), .ZN(n13389) );
  INV_X1 U16643 ( .A(DATAI_7_), .ZN(n13387) );
  NAND2_X1 U16644 ( .A1(n20419), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13386) );
  OAI21_X1 U16645 ( .B1(n20419), .B2(n13387), .A(n13386), .ZN(n14927) );
  NAND2_X1 U16646 ( .A1(n13388), .A2(n14927), .ZN(n13396) );
  NAND2_X1 U16647 ( .A1(n13389), .A2(n13396), .ZN(P1_U2959) );
  AOI22_X1 U16648 ( .A1(n13400), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n13366), .ZN(n13391) );
  NAND2_X1 U16649 ( .A1(n13391), .A2(n13390), .ZN(P1_U2960) );
  AOI22_X1 U16650 ( .A1(n13400), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n13366), .ZN(n13393) );
  NAND2_X1 U16651 ( .A1(n13393), .A2(n13392), .ZN(P1_U2940) );
  AOI22_X1 U16652 ( .A1(n13400), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n13366), .ZN(n13395) );
  NAND2_X1 U16653 ( .A1(n13395), .A2(n13394), .ZN(P1_U2952) );
  AOI22_X1 U16654 ( .A1(n13400), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n13366), .ZN(n13397) );
  NAND2_X1 U16655 ( .A1(n13397), .A2(n13396), .ZN(P1_U2944) );
  AOI22_X1 U16656 ( .A1(n13400), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n13366), .ZN(n13399) );
  NAND2_X1 U16657 ( .A1(n13399), .A2(n13398), .ZN(P1_U2957) );
  AOI22_X1 U16658 ( .A1(n13400), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n13366), .ZN(n13402) );
  NAND2_X1 U16659 ( .A1(n13402), .A2(n13401), .ZN(P1_U2958) );
  INV_X1 U16660 ( .A(n13403), .ZN(n20176) );
  INV_X1 U16661 ( .A(n13404), .ZN(n16596) );
  NAND2_X1 U16662 ( .A1(n16596), .A2(n13405), .ZN(n13815) );
  INV_X1 U16663 ( .A(n10431), .ZN(n13406) );
  NAND2_X1 U16664 ( .A1(n13406), .A2(n16575), .ZN(n13806) );
  INV_X1 U16665 ( .A(n13087), .ZN(n13811) );
  INV_X1 U16666 ( .A(n10417), .ZN(n13407) );
  OAI211_X1 U16667 ( .C1(n13811), .C2(n13407), .A(n10261), .B(n13807), .ZN(
        n13408) );
  AOI21_X1 U16668 ( .B1(n13815), .B2(n13806), .A(n13408), .ZN(n13413) );
  NAND3_X1 U16669 ( .A1(n13809), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n13808), .ZN(n13410) );
  OAI21_X1 U16670 ( .B1(n13811), .B2(n10417), .A(n13806), .ZN(n13409) );
  AOI21_X1 U16671 ( .B1(n13411), .B2(n13410), .A(n13409), .ZN(n13412) );
  OAI22_X1 U16672 ( .A1(n13263), .A2(n13844), .B1(n13413), .B2(n13412), .ZN(
        n16574) );
  AOI22_X1 U16673 ( .A1(n19521), .A2(n16616), .B1(n20176), .B2(n16574), .ZN(
        n13415) );
  NAND2_X1 U16674 ( .A1(n13850), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13414) );
  OAI21_X1 U16675 ( .B1(n13415), .B2(n13850), .A(n13414), .ZN(P2_U3596) );
  NAND2_X1 U16676 ( .A1(n13416), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13530) );
  NOR2_X1 U16677 ( .A1(n13530), .A2(n13531), .ZN(n13529) );
  OAI211_X1 U16678 ( .C1(n13529), .C2(n13417), .A(n15575), .B(n13348), .ZN(
        n13422) );
  NAND2_X1 U16679 ( .A1(n13418), .A2(n13526), .ZN(n13420) );
  NAND2_X1 U16680 ( .A1(n13420), .A2(n10121), .ZN(n15876) );
  INV_X1 U16681 ( .A(n15876), .ZN(n19269) );
  NAND2_X1 U16682 ( .A1(n15572), .A2(n19269), .ZN(n13421) );
  OAI211_X1 U16683 ( .C1(n15572), .C2(n13423), .A(n13422), .B(n13421), .ZN(
        P2_U2878) );
  INV_X1 U16684 ( .A(n13424), .ZN(n13425) );
  AOI21_X1 U16685 ( .B1(n13427), .B2(n13426), .A(n13425), .ZN(n20346) );
  INV_X1 U16686 ( .A(n20346), .ZN(n13432) );
  INV_X1 U16687 ( .A(n13469), .ZN(n13428) );
  AOI21_X1 U16688 ( .B1(n13430), .B2(n13429), .A(n13428), .ZN(n20396) );
  AOI22_X1 U16689 ( .A1(n20351), .A2(n20396), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14885), .ZN(n13431) );
  OAI21_X1 U16690 ( .B1(n13432), .B2(n14890), .A(n13431), .ZN(P1_U2870) );
  INV_X1 U16691 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13516) );
  OAI222_X1 U16692 ( .A1(n14995), .A2(n13432), .B1(n14988), .B2(n13516), .C1(
        n14987), .C2(n20439), .ZN(P1_U2902) );
  OR2_X1 U16693 ( .A1(n13509), .A2(n13434), .ZN(n13435) );
  AND2_X1 U16694 ( .A1(n13433), .A2(n13435), .ZN(n16504) );
  INV_X1 U16695 ( .A(n16504), .ZN(n19255) );
  INV_X1 U16696 ( .A(n13476), .ZN(n13441) );
  INV_X1 U16697 ( .A(n13505), .ZN(n13439) );
  OAI21_X1 U16698 ( .B1(n13437), .B2(n13439), .A(n13438), .ZN(n13440) );
  NAND3_X1 U16699 ( .A1(n13441), .A2(n15575), .A3(n13440), .ZN(n13443) );
  NAND2_X1 U16700 ( .A1(n15578), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13442) );
  OAI211_X1 U16701 ( .C1(n19255), .C2(n15578), .A(n13443), .B(n13442), .ZN(
        P2_U2875) );
  NAND2_X1 U16702 ( .A1(n13446), .A2(n13445), .ZN(n13447) );
  NAND2_X1 U16703 ( .A1(n13444), .A2(n13447), .ZN(n20362) );
  OR2_X1 U16704 ( .A1(n13471), .A2(n13448), .ZN(n13449) );
  AND2_X1 U16705 ( .A1(n13737), .A2(n13449), .ZN(n20374) );
  AOI22_X1 U16706 ( .A1(n20351), .A2(n20374), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n14885), .ZN(n13450) );
  OAI21_X1 U16707 ( .B1(n20362), .B2(n14890), .A(n13450), .ZN(P1_U2868) );
  INV_X1 U16708 ( .A(n19329), .ZN(n13692) );
  NAND2_X1 U16709 ( .A1(n12811), .A2(n13451), .ZN(n13452) );
  XNOR2_X1 U16710 ( .A(n13611), .B(n13452), .ZN(n13453) );
  NAND2_X1 U16711 ( .A1(n13453), .A2(n19308), .ZN(n13464) );
  NAND2_X1 U16712 ( .A1(n10100), .A2(n10098), .ZN(n13456) );
  AND2_X1 U16713 ( .A1(n13553), .A2(n13456), .ZN(n20180) );
  OAI22_X1 U16714 ( .A1(n19285), .A2(n13457), .B1(n13609), .B2(n19260), .ZN(
        n13459) );
  NOR2_X1 U16715 ( .A1(n19326), .A2(n12501), .ZN(n13458) );
  AOI211_X1 U16716 ( .C1(n19319), .C2(n20180), .A(n13459), .B(n13458), .ZN(
        n13460) );
  OAI21_X1 U16717 ( .B1(n13461), .B2(n19300), .A(n13460), .ZN(n13462) );
  AOI21_X1 U16718 ( .B1(n13454), .B2(n19313), .A(n13462), .ZN(n13463) );
  OAI211_X1 U16719 ( .C1(n13692), .C2(n20177), .A(n13464), .B(n13463), .ZN(
        P2_U2852) );
  INV_X1 U16720 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n13465) );
  OAI222_X1 U16721 ( .A1(n20362), .A2(n14995), .B1(n13465), .B2(n14988), .C1(
        n14987), .C2(n20447), .ZN(P1_U2900) );
  XOR2_X1 U16722 ( .A(n13466), .B(n13467), .Z(n13856) );
  INV_X1 U16723 ( .A(n13856), .ZN(n13480) );
  INV_X1 U16724 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13473) );
  AND2_X1 U16725 ( .A1(n13469), .A2(n13468), .ZN(n13470) );
  NOR2_X1 U16726 ( .A1(n13471), .A2(n13470), .ZN(n20384) );
  INV_X1 U16727 ( .A(n20384), .ZN(n13472) );
  OAI222_X1 U16728 ( .A1(n13480), .A2(n14890), .B1(n20356), .B2(n13473), .C1(
        n13472), .C2(n14896), .ZN(P1_U2869) );
  NAND2_X1 U16729 ( .A1(n13433), .A2(n13474), .ZN(n13475) );
  NAND2_X1 U16730 ( .A1(n13618), .A2(n13475), .ZN(n16111) );
  OAI211_X1 U16731 ( .C1(n13476), .C2(n13477), .A(n13621), .B(n15575), .ZN(
        n13479) );
  NAND2_X1 U16732 ( .A1(n15578), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13478) );
  OAI211_X1 U16733 ( .C1(n16111), .C2(n15592), .A(n13479), .B(n13478), .ZN(
        P2_U2874) );
  INV_X1 U16734 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n13521) );
  OAI222_X1 U16735 ( .A1(n14995), .A2(n13480), .B1(n14988), .B2(n13521), .C1(
        n14987), .C2(n20443), .ZN(P1_U2901) );
  INV_X1 U16736 ( .A(P1_UWORD_REG_12__SCAN_IN), .ZN(n13482) );
  INV_X2 U16737 ( .A(n21051), .ZN(n13785) );
  INV_X1 U16738 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13481) );
  OAI222_X1 U16739 ( .A1(n13482), .A2(n13785), .B1(n13758), .B2(n11901), .C1(
        n13741), .C2(n13481), .ZN(P1_U2908) );
  INV_X1 U16740 ( .A(P1_UWORD_REG_7__SCAN_IN), .ZN(n13485) );
  INV_X1 U16741 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13484) );
  INV_X1 U16742 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n13483) );
  OAI222_X1 U16743 ( .A1(n13485), .A2(n13785), .B1(n13758), .B2(n13484), .C1(
        n13741), .C2(n13483), .ZN(P1_U2913) );
  INV_X1 U16744 ( .A(P1_UWORD_REG_9__SCAN_IN), .ZN(n13488) );
  INV_X1 U16745 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13486) );
  OAI222_X1 U16746 ( .A1(n13488), .A2(n13785), .B1(n13758), .B2(n13487), .C1(
        n13741), .C2(n13486), .ZN(P1_U2911) );
  INV_X1 U16747 ( .A(P1_UWORD_REG_11__SCAN_IN), .ZN(n13491) );
  INV_X1 U16748 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13489) );
  OAI222_X1 U16749 ( .A1(n13491), .A2(n13785), .B1(n13758), .B2(n13490), .C1(
        n13741), .C2(n13489), .ZN(P1_U2909) );
  INV_X1 U16750 ( .A(P1_UWORD_REG_8__SCAN_IN), .ZN(n13493) );
  INV_X1 U16751 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13492) );
  OAI222_X1 U16752 ( .A1(n13493), .A2(n13785), .B1(n13758), .B2(n11801), .C1(
        n13741), .C2(n13492), .ZN(P1_U2912) );
  INV_X1 U16753 ( .A(P1_UWORD_REG_5__SCAN_IN), .ZN(n13496) );
  INV_X1 U16754 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13495) );
  INV_X1 U16755 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n13494) );
  OAI222_X1 U16756 ( .A1(n13496), .A2(n13785), .B1(n13758), .B2(n13495), .C1(
        n13741), .C2(n13494), .ZN(P1_U2915) );
  INV_X1 U16757 ( .A(P1_UWORD_REG_14__SCAN_IN), .ZN(n13499) );
  INV_X1 U16758 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13497) );
  OAI222_X1 U16759 ( .A1(n13499), .A2(n13785), .B1(n13758), .B2(n13498), .C1(
        n13741), .C2(n13497), .ZN(P1_U2906) );
  INV_X1 U16760 ( .A(P1_UWORD_REG_10__SCAN_IN), .ZN(n13501) );
  INV_X1 U16761 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13500) );
  OAI222_X1 U16762 ( .A1(n13501), .A2(n13785), .B1(n13758), .B2(n11849), .C1(
        n13741), .C2(n13500), .ZN(P1_U2910) );
  INV_X1 U16763 ( .A(P1_UWORD_REG_13__SCAN_IN), .ZN(n13504) );
  INV_X1 U16764 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13502) );
  OAI222_X1 U16765 ( .A1(n13504), .A2(n13785), .B1(n13758), .B2(n13503), .C1(
        n13741), .C2(n13502), .ZN(P1_U2907) );
  XOR2_X1 U16766 ( .A(n13437), .B(n13505), .Z(n13511) );
  AND2_X1 U16767 ( .A1(n13507), .A2(n13506), .ZN(n13508) );
  OR2_X1 U16768 ( .A1(n13509), .A2(n13508), .ZN(n16135) );
  MUX2_X1 U16769 ( .A(n16135), .B(n21083), .S(n15592), .Z(n13510) );
  OAI21_X1 U16770 ( .B1(n13511), .B2(n15594), .A(n13510), .ZN(P2_U2876) );
  INV_X1 U16771 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n13514) );
  INV_X1 U16772 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n13513) );
  OAI222_X1 U16773 ( .A1(n13514), .A2(n13785), .B1(n13783), .B2(n13707), .C1(
        n13513), .C2(n13741), .ZN(P1_U2931) );
  INV_X1 U16774 ( .A(P1_LWORD_REG_2__SCAN_IN), .ZN(n13517) );
  INV_X1 U16775 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n13515) );
  OAI222_X1 U16776 ( .A1(n13517), .A2(n13785), .B1(n13516), .B2(n13783), .C1(
        n13515), .C2(n13741), .ZN(P1_U2934) );
  INV_X1 U16777 ( .A(P1_LWORD_REG_6__SCAN_IN), .ZN(n13519) );
  INV_X1 U16778 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n13518) );
  OAI222_X1 U16779 ( .A1(n13519), .A2(n13785), .B1(n11433), .B2(n13783), .C1(
        n13518), .C2(n13741), .ZN(P1_U2930) );
  INV_X1 U16780 ( .A(P1_LWORD_REG_3__SCAN_IN), .ZN(n13522) );
  INV_X1 U16781 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n13520) );
  OAI222_X1 U16782 ( .A1(n13522), .A2(n13785), .B1(n13521), .B2(n13783), .C1(
        n13520), .C2(n13741), .ZN(P1_U2933) );
  INV_X1 U16783 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n13525) );
  INV_X1 U16784 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n13523) );
  OAI222_X1 U16785 ( .A1(n13525), .A2(n13785), .B1(n13524), .B2(n13783), .C1(
        n13523), .C2(n13741), .ZN(P1_U2935) );
  OAI21_X1 U16786 ( .B1(n13528), .B2(n13527), .A(n13526), .ZN(n16548) );
  NOR2_X1 U16787 ( .A1(n16548), .A2(n15592), .ZN(n13533) );
  AOI211_X1 U16788 ( .C1(n13531), .C2(n13530), .A(n15594), .B(n13529), .ZN(
        n13532) );
  AOI211_X1 U16789 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n15592), .A(n13533), .B(
        n13532), .ZN(n13534) );
  INV_X1 U16790 ( .A(n13534), .ZN(P2_U2879) );
  XNOR2_X1 U16791 ( .A(n13535), .B(n14291), .ZN(n13536) );
  XNOR2_X1 U16792 ( .A(n13537), .B(n13536), .ZN(n13616) );
  XOR2_X1 U16793 ( .A(n13538), .B(n13539), .Z(n13614) );
  NAND2_X1 U16794 ( .A1(n13614), .A2(n16550), .ZN(n13548) );
  INV_X1 U16795 ( .A(n20180), .ZN(n13540) );
  OAI22_X1 U16796 ( .A1(n19508), .A2(n13540), .B1(n13609), .B2(n19277), .ZN(
        n13546) );
  AOI21_X1 U16797 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14638) );
  INV_X1 U16798 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19500) );
  NOR3_X1 U16799 ( .A1(n19497), .A2(n19500), .A3(n14633), .ZN(n14639) );
  OAI21_X1 U16800 ( .B1(n16045), .B2(n14639), .A(n19499), .ZN(n14292) );
  NOR2_X1 U16801 ( .A1(n14638), .A2(n14292), .ZN(n13793) );
  INV_X1 U16802 ( .A(n14639), .ZN(n13541) );
  NAND2_X1 U16803 ( .A1(n16046), .A2(n13541), .ZN(n13542) );
  AND2_X1 U16804 ( .A1(n13542), .A2(n19501), .ZN(n14301) );
  NAND2_X1 U16805 ( .A1(n16045), .A2(n14638), .ZN(n13543) );
  AND2_X1 U16806 ( .A1(n14301), .A2(n13543), .ZN(n13794) );
  INV_X1 U16807 ( .A(n13794), .ZN(n13544) );
  MUX2_X1 U16808 ( .A(n13793), .B(n13544), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n13545) );
  AOI211_X1 U16809 ( .C1(n19505), .C2(n13454), .A(n13546), .B(n13545), .ZN(
        n13547) );
  OAI211_X1 U16810 ( .C1(n13616), .C2(n19502), .A(n13548), .B(n13547), .ZN(
        P2_U3043) );
  INV_X1 U16811 ( .A(n19495), .ZN(n13552) );
  NOR2_X1 U16812 ( .A1(n19289), .A2(n13549), .ZN(n13551) );
  AOI21_X1 U16813 ( .B1(n13552), .B2(n13551), .A(n20099), .ZN(n13550) );
  OAI21_X1 U16814 ( .B1(n13552), .B2(n13551), .A(n13550), .ZN(n13563) );
  INV_X1 U16815 ( .A(n13553), .ZN(n13555) );
  INV_X1 U16816 ( .A(n13956), .ZN(n13554) );
  OAI21_X1 U16817 ( .B1(n13556), .B2(n13555), .A(n13554), .ZN(n19380) );
  AOI22_X1 U16818 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19298), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n19320), .ZN(n13557) );
  OAI211_X1 U16819 ( .C1(n19312), .C2(n19380), .A(n13557), .B(n19277), .ZN(
        n13558) );
  AOI21_X1 U16820 ( .B1(n19318), .B2(P2_REIP_REG_4__SCAN_IN), .A(n13558), .ZN(
        n13559) );
  OAI21_X1 U16821 ( .B1(n13560), .B2(n19300), .A(n13559), .ZN(n13561) );
  AOI21_X1 U16822 ( .B1(n19487), .B2(n19313), .A(n13561), .ZN(n13562) );
  OAI211_X1 U16823 ( .C1(n19382), .C2(n13692), .A(n13563), .B(n13562), .ZN(
        P2_U2851) );
  INV_X1 U16824 ( .A(n20552), .ZN(n20791) );
  NOR2_X1 U16825 ( .A1(n11328), .A2(n20791), .ZN(n13564) );
  XNOR2_X1 U16826 ( .A(n13564), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13970) );
  NOR3_X1 U16827 ( .A1(n13970), .A2(n12009), .A3(n13637), .ZN(n16420) );
  OR2_X1 U16828 ( .A1(n16420), .A2(n13583), .ZN(n13565) );
  OAI21_X1 U16829 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n16217), .A(
        n13565), .ZN(n13566) );
  NAND2_X1 U16830 ( .A1(n21176), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13587) );
  OAI22_X1 U16831 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n13566), .B1(n13587), 
        .B2(n16422), .ZN(n16232) );
  NOR2_X1 U16832 ( .A1(n13219), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13567) );
  NOR2_X1 U16833 ( .A1(n11236), .A2(n13567), .ZN(n15421) );
  NAND2_X1 U16834 ( .A1(n11172), .A2(n15421), .ZN(n13578) );
  MUX2_X1 U16835 ( .A(n13569), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n11008), .Z(n13571) );
  NOR2_X1 U16836 ( .A1(n13571), .A2(n13570), .ZN(n13572) );
  NAND2_X1 U16837 ( .A1(n13573), .A2(n13572), .ZN(n13577) );
  XNOR2_X1 U16838 ( .A(n13574), .B(n13581), .ZN(n13575) );
  NAND2_X1 U16839 ( .A1(n16211), .A2(n13575), .ZN(n13576) );
  OAI211_X1 U16840 ( .C1(n13580), .C2(n13578), .A(n13577), .B(n13576), .ZN(
        n13579) );
  AOI21_X1 U16841 ( .B1(n20426), .B2(n13580), .A(n13579), .ZN(n15425) );
  MUX2_X1 U16842 ( .A(n13581), .B(n15425), .S(n16217), .Z(n16225) );
  OAI22_X1 U16843 ( .A1(n16225), .A2(P1_STATE2_REG_1__SCAN_IN), .B1(n13587), 
        .B2(n13581), .ZN(n13589) );
  NAND2_X1 U16844 ( .A1(n13582), .A2(n16217), .ZN(n13585) );
  NAND2_X1 U16845 ( .A1(n13583), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13584) );
  NAND2_X1 U16846 ( .A1(n13585), .A2(n13584), .ZN(n16223) );
  NAND2_X1 U16847 ( .A1(n16223), .A2(n20962), .ZN(n13586) );
  OAI21_X1 U16848 ( .B1(n13587), .B2(n11302), .A(n13586), .ZN(n13588) );
  NAND2_X1 U16849 ( .A1(n13589), .A2(n13588), .ZN(n16230) );
  NOR2_X1 U16850 ( .A1(n16230), .A2(n11010), .ZN(n13592) );
  NOR3_X1 U16851 ( .A1(n16232), .A2(n13592), .A3(P1_FLUSH_REG_SCAN_IN), .ZN(
        n13591) );
  OAI21_X1 U16852 ( .B1(n13591), .B2(n13590), .A(n20557), .ZN(n20417) );
  OR2_X1 U16853 ( .A1(n13592), .A2(n16432), .ZN(n13593) );
  NOR2_X1 U16854 ( .A1(n16232), .A2(n13593), .ZN(n16241) );
  INV_X1 U16855 ( .A(n11320), .ZN(n20523) );
  AND2_X1 U16856 ( .A1(n20674), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15410) );
  OAI22_X1 U16857 ( .A1(n13302), .A2(n20903), .B1(n20523), .B2(n15410), .ZN(
        n13594) );
  OAI21_X1 U16858 ( .B1(n16241), .B2(n13594), .A(n20417), .ZN(n13595) );
  OAI21_X1 U16859 ( .B1(n20417), .B2(n20820), .A(n13595), .ZN(P1_U3478) );
  NOR2_X1 U16860 ( .A1(n19289), .A2(n13596), .ZN(n13597) );
  XNOR2_X1 U16861 ( .A(n13597), .B(n16525), .ZN(n13598) );
  NAND2_X1 U16862 ( .A1(n13598), .A2(n19308), .ZN(n13607) );
  INV_X1 U16863 ( .A(n13599), .ZN(n13601) );
  INV_X1 U16864 ( .A(n16166), .ZN(n13600) );
  OAI21_X1 U16865 ( .B1(n13602), .B2(n13601), .A(n13600), .ZN(n19368) );
  AOI22_X1 U16866 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19318), .ZN(n13603) );
  OAI211_X1 U16867 ( .C1(n19312), .C2(n19368), .A(n13603), .B(n19277), .ZN(
        n13605) );
  NOR2_X1 U16868 ( .A1(n16548), .A2(n19292), .ZN(n13604) );
  AOI211_X1 U16869 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n19320), .A(n13605), .B(
        n13604), .ZN(n13606) );
  OAI211_X1 U16870 ( .C1(n19300), .C2(n13608), .A(n13607), .B(n13606), .ZN(
        P2_U2847) );
  OAI22_X1 U16871 ( .A1(n16541), .A2(n12501), .B1(n13609), .B2(n19277), .ZN(
        n13610) );
  AOI21_X1 U16872 ( .B1(n16533), .B2(n13611), .A(n13610), .ZN(n13612) );
  OAI21_X1 U16873 ( .B1(n13263), .B2(n16526), .A(n13612), .ZN(n13613) );
  AOI21_X1 U16874 ( .B1(n13614), .B2(n16529), .A(n13613), .ZN(n13615) );
  OAI21_X1 U16875 ( .B1(n16537), .B2(n13616), .A(n13615), .ZN(P2_U3011) );
  NAND2_X1 U16876 ( .A1(n13618), .A2(n13617), .ZN(n13619) );
  NAND2_X1 U16877 ( .A1(n13620), .A2(n13619), .ZN(n19232) );
  OAI211_X1 U16878 ( .C1(n9994), .C2(n13623), .A(n15575), .B(n13830), .ZN(
        n13625) );
  NAND2_X1 U16879 ( .A1(n15578), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13624) );
  OAI211_X1 U16880 ( .C1(n19232), .C2(n15592), .A(n13625), .B(n13624), .ZN(
        P2_U2873) );
  INV_X1 U16881 ( .A(n20417), .ZN(n13636) );
  INV_X1 U16882 ( .A(n13627), .ZN(n13628) );
  OR2_X1 U16883 ( .A1(n20851), .A2(n9702), .ZN(n20785) );
  AOI211_X1 U16884 ( .C1(n20697), .C2(n20785), .A(P1_STATE2_REG_3__SCAN_IN), 
        .B(n13631), .ZN(n13633) );
  NAND3_X1 U16885 ( .A1(n9702), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n20909), 
        .ZN(n15408) );
  NOR2_X1 U16886 ( .A1(n20641), .A2(n15408), .ZN(n20640) );
  NAND2_X1 U16887 ( .A1(n20909), .A2(n20852), .ZN(n20789) );
  INV_X1 U16888 ( .A(n20426), .ZN(n20667) );
  OAI22_X1 U16889 ( .A1(n13626), .A2(n20789), .B1(n20667), .B2(n15410), .ZN(
        n13632) );
  NOR3_X1 U16890 ( .A1(n13633), .A2(n20640), .A3(n13632), .ZN(n13635) );
  NAND2_X1 U16891 ( .A1(n13636), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13634) );
  OAI21_X1 U16892 ( .B1(n13636), .B2(n13635), .A(n13634), .ZN(P1_U3475) );
  NAND2_X1 U16893 ( .A1(n13638), .A2(n13637), .ZN(n13645) );
  INV_X1 U16894 ( .A(n13639), .ZN(n13640) );
  NAND2_X1 U16895 ( .A1(n13640), .A2(n13641), .ZN(n13670) );
  OAI211_X1 U16896 ( .C1(n13641), .C2(n13640), .A(n16235), .B(n13670), .ZN(
        n13643) );
  AND3_X1 U16897 ( .A1(n13643), .A2(n20438), .A3(n13642), .ZN(n13644) );
  NOR2_X1 U16898 ( .A1(n13647), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20409) );
  NOR2_X1 U16899 ( .A1(n20409), .A2(n20363), .ZN(n13651) );
  AOI22_X1 U16900 ( .A1(n20357), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20407), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13649) );
  OAI21_X1 U16901 ( .B1(n20368), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13649), .ZN(n13650) );
  AOI21_X1 U16902 ( .B1(n13651), .B2(n13656), .A(n13650), .ZN(n13652) );
  OAI21_X1 U16903 ( .B1(n20422), .B2(n13943), .A(n13652), .ZN(P1_U2998) );
  INV_X1 U16904 ( .A(n13646), .ZN(n13654) );
  NAND2_X1 U16905 ( .A1(n13654), .A2(n13653), .ZN(n13655) );
  INV_X1 U16906 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20403) );
  XNOR2_X1 U16907 ( .A(n13666), .B(n20403), .ZN(n13662) );
  XNOR2_X1 U16908 ( .A(n13670), .B(n13669), .ZN(n13659) );
  INV_X1 U16909 ( .A(n13657), .ZN(n13658) );
  AOI21_X1 U16910 ( .B1(n13659), .B2(n16235), .A(n13658), .ZN(n13660) );
  OAI21_X1 U16911 ( .B1(n13662), .B2(n13661), .A(n13668), .ZN(n20397) );
  AOI22_X1 U16912 ( .A1(n20357), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20407), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13663) );
  OAI21_X1 U16913 ( .B1(n20368), .B2(n20337), .A(n13663), .ZN(n13664) );
  AOI21_X1 U16914 ( .B1(n20346), .B2(n16332), .A(n13664), .ZN(n13665) );
  OAI21_X1 U16915 ( .B1(n20363), .B2(n20397), .A(n13665), .ZN(P1_U2997) );
  NAND2_X1 U16916 ( .A1(n13666), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13667) );
  NAND2_X1 U16917 ( .A1(n13670), .A2(n13669), .ZN(n13990) );
  XNOR2_X1 U16918 ( .A(n13990), .B(n13988), .ZN(n13671) );
  OAI22_X1 U16919 ( .A1(n13626), .A2(n9971), .B1(n14094), .B2(n13671), .ZN(
        n13672) );
  OAI21_X1 U16920 ( .B1(n13673), .B2(n13672), .A(n9671), .ZN(n20382) );
  AOI22_X1 U16921 ( .A1(n20357), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20407), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13674) );
  OAI21_X1 U16922 ( .B1(n20368), .B2(n13858), .A(n13674), .ZN(n13675) );
  AOI21_X1 U16923 ( .B1(n13856), .B2(n16332), .A(n13675), .ZN(n13676) );
  OAI21_X1 U16924 ( .B1(n20382), .B2(n20363), .A(n13676), .ZN(P1_U2996) );
  NOR2_X1 U16925 ( .A1(n19289), .A2(n13677), .ZN(n13719) );
  XNOR2_X1 U16926 ( .A(n13719), .B(n14648), .ZN(n13678) );
  NAND2_X1 U16927 ( .A1(n13678), .A2(n19308), .ZN(n13691) );
  NAND2_X1 U16928 ( .A1(n13680), .A2(n13679), .ZN(n13683) );
  INV_X1 U16929 ( .A(n13681), .ZN(n13682) );
  NAND2_X1 U16930 ( .A1(n13683), .A2(n13682), .ZN(n20188) );
  NAND2_X1 U16931 ( .A1(n20188), .A2(n19319), .ZN(n13686) );
  OAI22_X1 U16932 ( .A1(n19285), .A2(n10358), .B1(n21208), .B2(n19260), .ZN(
        n13684) );
  AOI21_X1 U16933 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19298), .A(
        n13684), .ZN(n13685) );
  OAI211_X1 U16934 ( .C1(n19300), .C2(n13687), .A(n13686), .B(n13685), .ZN(
        n13688) );
  AOI21_X1 U16935 ( .B1(n13689), .B2(n19313), .A(n13688), .ZN(n13690) );
  OAI211_X1 U16936 ( .C1(n13692), .C2(n19520), .A(n13691), .B(n13690), .ZN(
        P2_U2853) );
  INV_X1 U16937 ( .A(n13693), .ZN(n13694) );
  NAND2_X1 U16938 ( .A1(n13695), .A2(n13694), .ZN(n13842) );
  INV_X1 U16939 ( .A(n13842), .ZN(n13697) );
  MUX2_X1 U16940 ( .A(n13811), .B(n13697), .S(n13696), .Z(n13698) );
  OAI21_X1 U16941 ( .B1(n13699), .B2(n13844), .A(n13698), .ZN(n16578) );
  INV_X1 U16942 ( .A(n19332), .ZN(n13700) );
  AOI22_X1 U16943 ( .A1(n19289), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n13700), .B2(n12811), .ZN(n13818) );
  AOI222_X1 U16944 ( .A1(n16578), .A2(n20176), .B1(n13701), .B2(n16616), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n13818), .ZN(n13703) );
  NAND2_X1 U16945 ( .A1(n13850), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13702) );
  OAI21_X1 U16946 ( .B1(n13703), .B2(n13850), .A(n13702), .ZN(P2_U3601) );
  INV_X1 U16947 ( .A(n13704), .ZN(n13705) );
  AOI21_X1 U16948 ( .B1(n13706), .B2(n13444), .A(n13705), .ZN(n20327) );
  INV_X1 U16949 ( .A(n20327), .ZN(n13739) );
  INV_X1 U16950 ( .A(n14937), .ZN(n20451) );
  OAI222_X1 U16951 ( .A1(n13739), .A2(n14995), .B1(n13707), .B2(n14988), .C1(
        n14987), .C2(n20451), .ZN(P1_U2899) );
  INV_X1 U16952 ( .A(n14335), .ZN(n13711) );
  OAI22_X1 U16953 ( .A1(n19285), .A2(n13708), .B1(n20121), .B2(n19260), .ZN(
        n13710) );
  NOR2_X1 U16954 ( .A1(n19326), .A2(n14338), .ZN(n13709) );
  AOI211_X1 U16955 ( .C1(n19317), .C2(n13711), .A(n13710), .B(n13709), .ZN(
        n13718) );
  INV_X1 U16956 ( .A(n13712), .ZN(n13714) );
  NAND2_X1 U16957 ( .A1(n13714), .A2(n13713), .ZN(n13715) );
  NAND2_X1 U16958 ( .A1(n13716), .A2(n13715), .ZN(n20197) );
  NAND2_X1 U16959 ( .A1(n19319), .A2(n20197), .ZN(n13717) );
  OAI211_X1 U16960 ( .C1(n13845), .C2(n19292), .A(n13718), .B(n13717), .ZN(
        n13722) );
  OAI21_X1 U16961 ( .B1(n19332), .B2(n13720), .A(n13719), .ZN(n13817) );
  OAI22_X1 U16962 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19325), .B1(
        n13817), .B2(n20099), .ZN(n13721) );
  AOI211_X1 U16963 ( .C1(n19329), .C2(n20193), .A(n13722), .B(n13721), .ZN(
        n13723) );
  INV_X1 U16964 ( .A(n13723), .ZN(P2_U2854) );
  OAI21_X1 U16965 ( .B1(n15520), .B2(n13724), .A(n16125), .ZN(n19359) );
  OR2_X1 U16966 ( .A1(n19289), .A2(n13725), .ZN(n19250) );
  AOI211_X1 U16967 ( .C1(n13726), .C2(n13729), .A(n20099), .B(n19250), .ZN(
        n13727) );
  INV_X1 U16968 ( .A(n13727), .ZN(n13735) );
  INV_X1 U16969 ( .A(n13728), .ZN(n13733) );
  INV_X1 U16970 ( .A(n13729), .ZN(n15865) );
  OAI22_X1 U16971 ( .A1(n16135), .A2(n19292), .B1(n19325), .B2(n15865), .ZN(
        n13732) );
  AOI22_X1 U16972 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19318), .ZN(n13730) );
  OAI211_X1 U16973 ( .C1(n19285), .C2(n21083), .A(n13730), .B(n19277), .ZN(
        n13731) );
  AOI211_X1 U16974 ( .C1(n19317), .C2(n13733), .A(n13732), .B(n13731), .ZN(
        n13734) );
  OAI211_X1 U16975 ( .C1(n19359), .C2(n19312), .A(n13735), .B(n13734), .ZN(
        P2_U2844) );
  NAND2_X1 U16976 ( .A1(n13737), .A2(n13736), .ZN(n13738) );
  NAND2_X1 U16977 ( .A1(n16399), .A2(n13738), .ZN(n20324) );
  INV_X1 U16978 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13740) );
  OAI222_X1 U16979 ( .A1(n20324), .A2(n14896), .B1(n13740), .B2(n20356), .C1(
        n13739), .C2(n14890), .ZN(P1_U2867) );
  INV_X1 U16980 ( .A(P1_UWORD_REG_3__SCAN_IN), .ZN(n13744) );
  INV_X1 U16981 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13743) );
  INV_X1 U16982 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n13742) );
  OAI222_X1 U16983 ( .A1(n13744), .A2(n13785), .B1(n13758), .B2(n13743), .C1(
        n13741), .C2(n13742), .ZN(P1_U2917) );
  INV_X1 U16984 ( .A(P1_UWORD_REG_1__SCAN_IN), .ZN(n13747) );
  INV_X1 U16985 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13746) );
  INV_X1 U16986 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n13745) );
  OAI222_X1 U16987 ( .A1(n13747), .A2(n13785), .B1(n13758), .B2(n13746), .C1(
        n13741), .C2(n13745), .ZN(P1_U2919) );
  INV_X1 U16988 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n13750) );
  INV_X1 U16989 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13749) );
  INV_X1 U16990 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n13748) );
  OAI222_X1 U16991 ( .A1(n13750), .A2(n13785), .B1(n13758), .B2(n13749), .C1(
        n13741), .C2(n13748), .ZN(P1_U2914) );
  INV_X1 U16992 ( .A(P1_UWORD_REG_0__SCAN_IN), .ZN(n13752) );
  INV_X1 U16993 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n13751) );
  OAI222_X1 U16994 ( .A1(n13752), .A2(n13785), .B1(n13758), .B2(n14966), .C1(
        n13741), .C2(n13751), .ZN(P1_U2920) );
  INV_X1 U16995 ( .A(P1_UWORD_REG_2__SCAN_IN), .ZN(n13755) );
  INV_X1 U16996 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13754) );
  INV_X1 U16997 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n13753) );
  OAI222_X1 U16998 ( .A1(n13755), .A2(n13785), .B1(n13758), .B2(n13754), .C1(
        n13741), .C2(n13753), .ZN(P1_U2918) );
  INV_X1 U16999 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n13759) );
  INV_X1 U17000 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13757) );
  INV_X1 U17001 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n13756) );
  OAI222_X1 U17002 ( .A1(n13759), .A2(n13785), .B1(n13758), .B2(n13757), .C1(
        n13741), .C2(n13756), .ZN(P1_U2916) );
  INV_X1 U17003 ( .A(P1_LWORD_REG_9__SCAN_IN), .ZN(n13762) );
  INV_X1 U17004 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n13760) );
  OAI222_X1 U17005 ( .A1(n13762), .A2(n13785), .B1(n13783), .B2(n13761), .C1(
        n13760), .C2(n13741), .ZN(P1_U2927) );
  INV_X1 U17006 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n13765) );
  INV_X1 U17007 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n13763) );
  OAI222_X1 U17008 ( .A1(n13765), .A2(n13785), .B1(n13783), .B2(n13764), .C1(
        n13763), .C2(n13741), .ZN(P1_U2925) );
  INV_X1 U17009 ( .A(P1_LWORD_REG_13__SCAN_IN), .ZN(n13768) );
  INV_X1 U17010 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n13766) );
  OAI222_X1 U17011 ( .A1(n13768), .A2(n13785), .B1(n13783), .B2(n13767), .C1(
        n13766), .C2(n13741), .ZN(P1_U2923) );
  INV_X1 U17012 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n13769) );
  OAI222_X1 U17013 ( .A1(n13101), .A2(n13785), .B1(n14974), .B2(n13783), .C1(
        n13769), .C2(n13741), .ZN(P1_U2921) );
  INV_X1 U17014 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n13771) );
  INV_X1 U17015 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n13770) );
  OAI222_X1 U17016 ( .A1(n13771), .A2(n13785), .B1(n13783), .B2(n13805), .C1(
        n13770), .C2(n13741), .ZN(P1_U2929) );
  INV_X1 U17017 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n13774) );
  INV_X1 U17018 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n13772) );
  OAI222_X1 U17019 ( .A1(n13774), .A2(n13785), .B1(n13783), .B2(n13773), .C1(
        n13772), .C2(n13741), .ZN(P1_U2922) );
  INV_X1 U17020 ( .A(P1_LWORD_REG_10__SCAN_IN), .ZN(n13777) );
  INV_X1 U17021 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n13775) );
  OAI222_X1 U17022 ( .A1(n13777), .A2(n13785), .B1(n13783), .B2(n13776), .C1(
        n13775), .C2(n13741), .ZN(P1_U2926) );
  INV_X1 U17023 ( .A(P1_LWORD_REG_8__SCAN_IN), .ZN(n13779) );
  INV_X1 U17024 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13836) );
  INV_X1 U17025 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n13778) );
  OAI222_X1 U17026 ( .A1(n13779), .A2(n13785), .B1(n13836), .B2(n13783), .C1(
        n13778), .C2(n13741), .ZN(P1_U2928) );
  INV_X1 U17027 ( .A(P1_LWORD_REG_12__SCAN_IN), .ZN(n13781) );
  INV_X1 U17028 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n13780) );
  OAI222_X1 U17029 ( .A1(n13781), .A2(n13785), .B1(n13783), .B2(n14989), .C1(
        n13780), .C2(n13741), .ZN(P1_U2924) );
  INV_X1 U17030 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n13786) );
  INV_X1 U17031 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n13782) );
  OAI222_X1 U17032 ( .A1(n13786), .A2(n13785), .B1(n13784), .B2(n13783), .C1(
        n13782), .C2(n13741), .ZN(P1_U2936) );
  NAND2_X1 U17033 ( .A1(n13788), .A2(n13787), .ZN(n13789) );
  XNOR2_X1 U17034 ( .A(n13789), .B(n13954), .ZN(n19491) );
  INV_X1 U17035 ( .A(n13790), .ZN(n13791) );
  XNOR2_X1 U17036 ( .A(n13792), .B(n13791), .ZN(n19485) );
  NAND2_X1 U17037 ( .A1(n19485), .A2(n16568), .ZN(n13800) );
  NAND2_X1 U17038 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13793), .ZN(
        n16552) );
  INV_X1 U17039 ( .A(n16552), .ZN(n13798) );
  NAND2_X1 U17040 ( .A1(n19487), .A2(n19505), .ZN(n13796) );
  INV_X1 U17041 ( .A(n19499), .ZN(n16093) );
  OAI21_X1 U17042 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16093), .A(
        n13794), .ZN(n14076) );
  AOI22_X1 U17043 ( .A1(n19303), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n14076), .ZN(n13795) );
  OAI211_X1 U17044 ( .C1(n19508), .C2(n19380), .A(n13796), .B(n13795), .ZN(
        n13797) );
  AOI21_X1 U17045 ( .B1(n13798), .B2(n13954), .A(n13797), .ZN(n13799) );
  OAI211_X1 U17046 ( .C1(n19491), .C2(n19515), .A(n13800), .B(n13799), .ZN(
        P2_U3042) );
  OR2_X1 U17047 ( .A1(n13802), .A2(n13803), .ZN(n13804) );
  AND2_X1 U17048 ( .A1(n13801), .A2(n13804), .ZN(n20297) );
  INV_X1 U17049 ( .A(n20297), .ZN(n13827) );
  INV_X1 U17050 ( .A(n14927), .ZN(n20462) );
  OAI222_X1 U17051 ( .A1(n13827), .A2(n14995), .B1(n13805), .B2(n14988), .C1(
        n14987), .C2(n20462), .ZN(P1_U2897) );
  NAND2_X1 U17052 ( .A1(n13807), .A2(n13806), .ZN(n13814) );
  AOI21_X1 U17053 ( .B1(n13809), .B2(n13808), .A(n13814), .ZN(n13813) );
  NOR3_X1 U17054 ( .A1(n13811), .A2(n13810), .A3(n10417), .ZN(n13812) );
  AOI211_X1 U17055 ( .C1(n13815), .C2(n13814), .A(n13813), .B(n13812), .ZN(
        n13816) );
  OAI21_X1 U17056 ( .B1(n14655), .B2(n13844), .A(n13816), .ZN(n16577) );
  OAI21_X1 U17057 ( .B1(n12811), .B2(n19500), .A(n13817), .ZN(n13846) );
  NOR2_X1 U17058 ( .A1(n13818), .A2(n10785), .ZN(n13847) );
  AOI222_X1 U17059 ( .A1(n16577), .A2(n20176), .B1(n16616), .B2(n20184), .C1(
        n13846), .C2(n13847), .ZN(n13820) );
  NAND2_X1 U17060 ( .A1(n13850), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13819) );
  OAI21_X1 U17061 ( .B1(n13820), .B2(n13850), .A(n13819), .ZN(P2_U3599) );
  OAI21_X1 U17062 ( .B1(n10037), .B2(n10176), .A(n13821), .ZN(n20286) );
  OAI21_X1 U17063 ( .B1(n9728), .B2(n13822), .A(n14025), .ZN(n13823) );
  INV_X1 U17064 ( .A(n13823), .ZN(n20284) );
  AOI22_X1 U17065 ( .A1(n20284), .A2(n20351), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14885), .ZN(n13824) );
  OAI21_X1 U17066 ( .B1(n20286), .B2(n14890), .A(n13824), .ZN(P1_U2864) );
  AND2_X1 U17067 ( .A1(n16401), .A2(n13825), .ZN(n13826) );
  OR2_X1 U17068 ( .A1(n13826), .A2(n9728), .ZN(n20298) );
  INV_X1 U17069 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13828) );
  OAI222_X1 U17070 ( .A1(n20298), .A2(n14896), .B1(n13828), .B2(n20356), .C1(
        n13827), .C2(n14890), .ZN(P1_U2865) );
  INV_X1 U17071 ( .A(n15842), .ZN(n16074) );
  INV_X1 U17072 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13829) );
  NOR2_X1 U17073 ( .A1(n15572), .A2(n13829), .ZN(n13833) );
  AOI211_X1 U17074 ( .C1(n13831), .C2(n13830), .A(n15594), .B(n13910), .ZN(
        n13832) );
  AOI211_X1 U17075 ( .C1(n16074), .C2(n15572), .A(n13833), .B(n13832), .ZN(
        n13834) );
  INV_X1 U17076 ( .A(n13834), .ZN(P2_U2872) );
  INV_X1 U17077 ( .A(n14922), .ZN(n13835) );
  OAI222_X1 U17078 ( .A1(n14995), .A2(n20286), .B1(n14988), .B2(n13836), .C1(
        n14987), .C2(n13835), .ZN(P1_U2896) );
  AND2_X1 U17079 ( .A1(n13704), .A2(n13837), .ZN(n13838) );
  NOR2_X1 U17080 ( .A1(n13802), .A2(n13838), .ZN(n20353) );
  INV_X1 U17081 ( .A(n20353), .ZN(n13839) );
  INV_X1 U17082 ( .A(n14932), .ZN(n20454) );
  OAI222_X1 U17083 ( .A1(n14995), .A2(n13839), .B1(n14988), .B2(n11433), .C1(
        n14987), .C2(n20454), .ZN(P1_U2898) );
  NOR2_X1 U17084 ( .A1(n10418), .A2(n10431), .ZN(n13841) );
  AOI22_X1 U17085 ( .A1(n13842), .A2(n13841), .B1(n13840), .B2(n13087), .ZN(
        n13843) );
  OAI21_X1 U17086 ( .B1(n13845), .B2(n13844), .A(n13843), .ZN(n16580) );
  INV_X1 U17087 ( .A(n13846), .ZN(n13848) );
  AOI222_X1 U17088 ( .A1(n16580), .A2(n20176), .B1(n13848), .B2(n13847), .C1(
        n20193), .C2(n16616), .ZN(n13851) );
  NAND2_X1 U17089 ( .A1(n13850), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13849) );
  OAI21_X1 U17090 ( .B1(n13851), .B2(n13850), .A(n13849), .ZN(P2_U3600) );
  OR2_X1 U17091 ( .A1(n13854), .A2(n13852), .ZN(n20342) );
  OR2_X1 U17092 ( .A1(n13854), .A2(n13853), .ZN(n13855) );
  INV_X1 U17093 ( .A(n13975), .ZN(n20345) );
  NAND2_X1 U17094 ( .A1(n13856), .A2(n20345), .ZN(n13868) );
  NAND2_X1 U17095 ( .A1(n20333), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20336) );
  NAND2_X1 U17096 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n20986), .ZN(n13865) );
  OAI221_X1 U17097 ( .B1(n14817), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n14817), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n20261), .ZN(n13857) );
  AOI22_X1 U17098 ( .A1(n20340), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n13857), .ZN(n13861) );
  INV_X1 U17099 ( .A(n13858), .ZN(n13859) );
  NAND2_X1 U17100 ( .A1(n20339), .A2(n13859), .ZN(n13860) );
  OAI211_X1 U17101 ( .C1(n20308), .C2(n13473), .A(n13861), .B(n13860), .ZN(
        n13862) );
  INV_X1 U17102 ( .A(n13862), .ZN(n13864) );
  NAND2_X1 U17103 ( .A1(n20334), .A2(n20384), .ZN(n13863) );
  OAI211_X1 U17104 ( .C1(n20336), .C2(n13865), .A(n13864), .B(n13863), .ZN(
        n13866) );
  INV_X1 U17105 ( .A(n13866), .ZN(n13867) );
  OAI211_X1 U17106 ( .C1(n20667), .C2(n20342), .A(n13868), .B(n13867), .ZN(
        P1_U2837) );
  OR2_X1 U17107 ( .A1(n13933), .A2(n13870), .ZN(n13871) );
  NAND2_X1 U17108 ( .A1(n13869), .A2(n13871), .ZN(n19213) );
  INV_X1 U17109 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13872) );
  OAI22_X1 U17110 ( .A1(n21236), .A2(n14417), .B1(n14411), .B2(n13872), .ZN(
        n13873) );
  INV_X1 U17111 ( .A(n13873), .ZN(n13884) );
  INV_X1 U17112 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13875) );
  OAI22_X1 U17113 ( .A1(n13875), .A2(n14416), .B1(n14412), .B2(n13874), .ZN(
        n13876) );
  INV_X1 U17114 ( .A(n13876), .ZN(n13883) );
  INV_X1 U17115 ( .A(n14431), .ZN(n14398) );
  NAND2_X1 U17116 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13878) );
  NAND2_X1 U17117 ( .A1(n14421), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13877) );
  OAI211_X1 U17118 ( .C1(n14398), .C2(n13879), .A(n13878), .B(n13877), .ZN(
        n13880) );
  INV_X1 U17119 ( .A(n13880), .ZN(n13882) );
  AOI22_X1 U17120 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10494), .B1(
        n14430), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13881) );
  NAND4_X1 U17121 ( .A1(n13884), .A2(n13883), .A3(n13882), .A4(n13881), .ZN(
        n13890) );
  AOI22_X1 U17122 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10578), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13888) );
  AOI22_X1 U17123 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10645), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13887) );
  AOI22_X1 U17124 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14432), .B1(
        n14404), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13886) );
  NAND2_X1 U17125 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13885) );
  NAND4_X1 U17126 ( .A1(n13888), .A2(n13887), .A3(n13886), .A4(n13885), .ZN(
        n13889) );
  NOR2_X1 U17127 ( .A1(n13890), .A2(n13889), .ZN(n13914) );
  AOI22_X1 U17128 ( .A1(n10578), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13894) );
  AOI22_X1 U17129 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U17130 ( .A1(n14432), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14404), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13892) );
  NAND2_X1 U17131 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13891) );
  AND4_X1 U17132 ( .A1(n13894), .A2(n13893), .A3(n13892), .A4(n13891), .ZN(
        n13909) );
  AOI22_X1 U17133 ( .A1(n14431), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13899) );
  NAND2_X1 U17134 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13898) );
  INV_X1 U17135 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n19764) );
  OR2_X1 U17136 ( .A1(n14417), .A2(n19764), .ZN(n13897) );
  INV_X1 U17137 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13895) );
  OR2_X1 U17138 ( .A1(n14411), .A2(n13895), .ZN(n13896) );
  NAND4_X1 U17139 ( .A1(n13899), .A2(n13898), .A3(n13897), .A4(n13896), .ZN(
        n13907) );
  OR2_X1 U17140 ( .A1(n14412), .A2(n13900), .ZN(n13905) );
  INV_X1 U17141 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13901) );
  OR2_X1 U17142 ( .A1(n14416), .A2(n13901), .ZN(n13904) );
  NAND2_X1 U17143 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13903) );
  NAND2_X1 U17144 ( .A1(n14430), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13902) );
  NAND4_X1 U17145 ( .A1(n13905), .A2(n13904), .A3(n13903), .A4(n13902), .ZN(
        n13906) );
  NOR2_X1 U17146 ( .A1(n13907), .A2(n13906), .ZN(n13908) );
  NAND2_X1 U17147 ( .A1(n13909), .A2(n13908), .ZN(n13928) );
  INV_X1 U17148 ( .A(n13912), .ZN(n13913) );
  AOI21_X1 U17149 ( .B1(n13914), .B2(n13911), .A(n13912), .ZN(n15681) );
  NAND2_X1 U17150 ( .A1(n15681), .A2(n15575), .ZN(n13916) );
  NAND2_X1 U17151 ( .A1(n15578), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13915) );
  OAI211_X1 U17152 ( .C1(n19213), .C2(n15578), .A(n13916), .B(n13915), .ZN(
        P2_U2870) );
  INV_X1 U17153 ( .A(n20342), .ZN(n13917) );
  NAND2_X1 U17154 ( .A1(n13917), .A2(n11320), .ZN(n13919) );
  OAI21_X1 U17155 ( .B1(n20340), .B2(n20339), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13918) );
  OAI211_X1 U17156 ( .C1(n20308), .C2(n13920), .A(n13919), .B(n13918), .ZN(
        n13924) );
  INV_X1 U17157 ( .A(n20292), .ZN(n13922) );
  NOR2_X1 U17158 ( .A1(n13922), .A2(n13921), .ZN(n13923) );
  AOI211_X1 U17159 ( .C1(n13925), .C2(n20334), .A(n13924), .B(n13923), .ZN(
        n13926) );
  OAI21_X1 U17160 ( .B1(n13975), .B2(n13927), .A(n13926), .ZN(P1_U2840) );
  OR2_X1 U17161 ( .A1(n13910), .A2(n13928), .ZN(n13929) );
  AND2_X1 U17162 ( .A1(n13911), .A2(n13929), .ZN(n19344) );
  NAND2_X1 U17163 ( .A1(n19344), .A2(n15575), .ZN(n13935) );
  NOR2_X1 U17164 ( .A1(n13931), .A2(n13930), .ZN(n13932) );
  OR2_X1 U17165 ( .A1(n13933), .A2(n13932), .ZN(n15827) );
  NAND2_X1 U17166 ( .A1(n16062), .A2(n15572), .ZN(n13934) );
  OAI211_X1 U17167 ( .C1(n15572), .C2(n13936), .A(n13935), .B(n13934), .ZN(
        P2_U2871) );
  AOI22_X1 U17168 ( .A1(n20335), .A2(P1_EBX_REG_1__SCAN_IN), .B1(n20333), .B2(
        n21037), .ZN(n13942) );
  NOR2_X1 U17169 ( .A1(n20342), .A2(n9697), .ZN(n13940) );
  AOI22_X1 U17170 ( .A1(n20340), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20332), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13938) );
  OAI21_X1 U17171 ( .B1(n20330), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13938), .ZN(n13939) );
  AOI211_X1 U17172 ( .C1(n20405), .C2(n20334), .A(n13940), .B(n13939), .ZN(
        n13941) );
  OAI211_X1 U17173 ( .C1(n13943), .C2(n13975), .A(n13942), .B(n13941), .ZN(
        P1_U2839) );
  AND2_X1 U17174 ( .A1(n13821), .A2(n13944), .ZN(n13945) );
  OR2_X1 U17175 ( .A1(n13945), .A2(n9763), .ZN(n20272) );
  AOI22_X1 U17176 ( .A1(n14993), .A2(n14917), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14991), .ZN(n13946) );
  OAI21_X1 U17177 ( .B1(n20272), .B2(n14995), .A(n13946), .ZN(P1_U2895) );
  XNOR2_X1 U17178 ( .A(n13947), .B(n13948), .ZN(n16536) );
  AND2_X1 U17179 ( .A1(n13950), .A2(n10636), .ZN(n13951) );
  OAI22_X1 U17180 ( .A1(n13953), .A2(n13952), .B1(n13949), .B2(n13951), .ZN(
        n16535) );
  NOR2_X1 U17181 ( .A1(n16535), .A2(n19515), .ZN(n13962) );
  NAND2_X1 U17182 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14075) );
  INV_X1 U17183 ( .A(n14075), .ZN(n14290) );
  AOI211_X1 U17184 ( .C1(n13955), .C2(n13954), .A(n14290), .B(n16552), .ZN(
        n13961) );
  NOR2_X1 U17185 ( .A1(n16534), .A2(n16547), .ZN(n13960) );
  XNOR2_X1 U17186 ( .A(n13957), .B(n13956), .ZN(n19378) );
  AOI22_X1 U17187 ( .A1(n19303), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n14076), .ZN(n13958) );
  OAI21_X1 U17188 ( .B1(n19508), .B2(n19378), .A(n13958), .ZN(n13959) );
  NOR4_X1 U17189 ( .A1(n13962), .A2(n13961), .A3(n13960), .A4(n13959), .ZN(
        n13963) );
  OAI21_X1 U17190 ( .B1(n19502), .B2(n16536), .A(n13963), .ZN(P2_U3041) );
  OR4_X1 U17191 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20986), .A3(n20392), .A4(
        n20336), .ZN(n13974) );
  NAND2_X1 U17192 ( .A1(n20261), .A2(n13964), .ZN(n20322) );
  OAI21_X1 U17193 ( .B1(n20262), .B2(n14817), .A(n20261), .ZN(n20321) );
  NAND2_X1 U17194 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20321), .ZN(n13965) );
  AND2_X1 U17195 ( .A1(n20322), .A2(n13965), .ZN(n13968) );
  INV_X1 U17196 ( .A(n20367), .ZN(n13966) );
  AOI22_X1 U17197 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n13966), .ZN(n13967) );
  OAI211_X1 U17198 ( .C1(n20308), .C2(n13969), .A(n13968), .B(n13967), .ZN(
        n13972) );
  NOR2_X1 U17199 ( .A1(n13970), .A2(n20342), .ZN(n13971) );
  AOI211_X1 U17200 ( .C1(n20334), .C2(n20374), .A(n13972), .B(n13971), .ZN(
        n13973) );
  OAI211_X1 U17201 ( .C1(n13975), .C2(n20362), .A(n13974), .B(n13973), .ZN(
        P1_U2836) );
  NAND2_X1 U17202 ( .A1(n13976), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13977) );
  NAND2_X1 U17203 ( .A1(n13978), .A2(n13977), .ZN(n20359) );
  NAND2_X1 U17204 ( .A1(n13979), .A2(n14005), .ZN(n13983) );
  NAND2_X1 U17205 ( .A1(n13990), .A2(n13988), .ZN(n13980) );
  XNOR2_X1 U17206 ( .A(n13980), .B(n13987), .ZN(n13981) );
  NAND2_X1 U17207 ( .A1(n13981), .A2(n16235), .ZN(n13982) );
  NAND2_X1 U17208 ( .A1(n13983), .A2(n13982), .ZN(n13984) );
  INV_X1 U17209 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20381) );
  XNOR2_X1 U17210 ( .A(n13984), .B(n20381), .ZN(n20358) );
  NAND2_X1 U17211 ( .A1(n13984), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13985) );
  NAND2_X1 U17212 ( .A1(n13986), .A2(n14005), .ZN(n13993) );
  AND2_X1 U17213 ( .A1(n13988), .A2(n13987), .ZN(n13989) );
  NAND2_X1 U17214 ( .A1(n13990), .A2(n13989), .ZN(n13999) );
  XNOR2_X1 U17215 ( .A(n13999), .B(n13997), .ZN(n13991) );
  NAND2_X1 U17216 ( .A1(n13991), .A2(n16235), .ZN(n13992) );
  INV_X1 U17217 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16409) );
  NAND2_X1 U17218 ( .A1(n13994), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13995) );
  NAND3_X1 U17219 ( .A1(n14093), .A2(n13996), .A3(n14005), .ZN(n14002) );
  INV_X1 U17220 ( .A(n13997), .ZN(n13998) );
  OR2_X1 U17221 ( .A1(n13999), .A2(n13998), .ZN(n14007) );
  XNOR2_X1 U17222 ( .A(n14007), .B(n14008), .ZN(n14000) );
  NAND2_X1 U17223 ( .A1(n14000), .A2(n16235), .ZN(n14001) );
  NAND2_X1 U17224 ( .A1(n14002), .A2(n14001), .ZN(n16337) );
  OR2_X1 U17225 ( .A1(n16337), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14003) );
  NAND2_X1 U17226 ( .A1(n16337), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14004) );
  NAND2_X1 U17227 ( .A1(n14006), .A2(n14005), .ZN(n14013) );
  INV_X1 U17228 ( .A(n14007), .ZN(n14009) );
  NAND2_X1 U17229 ( .A1(n14009), .A2(n14008), .ZN(n14096) );
  XNOR2_X1 U17230 ( .A(n14096), .B(n14010), .ZN(n14011) );
  NAND2_X1 U17231 ( .A1(n14011), .A2(n16235), .ZN(n14012) );
  NAND2_X1 U17232 ( .A1(n14013), .A2(n14012), .ZN(n14014) );
  OR2_X1 U17233 ( .A1(n14014), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14087) );
  NAND2_X1 U17234 ( .A1(n14014), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14089) );
  NAND2_X1 U17235 ( .A1(n14087), .A2(n14089), .ZN(n14015) );
  XNOR2_X1 U17236 ( .A(n14088), .B(n14015), .ZN(n16333) );
  INV_X1 U17237 ( .A(n16333), .ZN(n14022) );
  NOR2_X1 U17238 ( .A1(n20381), .A2(n20387), .ZN(n20375) );
  INV_X1 U17239 ( .A(n20375), .ZN(n14017) );
  NOR2_X1 U17240 ( .A1(n14018), .A2(n14016), .ZN(n15309) );
  INV_X1 U17241 ( .A(n16364), .ZN(n15314) );
  NOR2_X1 U17242 ( .A1(n20411), .A2(n9877), .ZN(n20398) );
  NAND2_X1 U17243 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n20398), .ZN(
        n15394) );
  NOR3_X1 U17244 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14017), .A3(
        n15394), .ZN(n16414) );
  INV_X1 U17245 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16397) );
  NOR3_X1 U17246 ( .A1(n20403), .A2(n9877), .A3(n14017), .ZN(n14219) );
  NOR2_X1 U17247 ( .A1(n16409), .A2(n14017), .ZN(n15390) );
  OAI21_X1 U17248 ( .B1(n14018), .B2(n9877), .A(n20403), .ZN(n20369) );
  NAND2_X1 U17249 ( .A1(n15390), .A2(n20369), .ZN(n15307) );
  AOI21_X1 U17250 ( .B1(n15307), .B2(n20390), .A(n14019), .ZN(n14220) );
  OAI21_X1 U17251 ( .B1(n20372), .B2(n14219), .A(n14220), .ZN(n16407) );
  NOR3_X1 U17252 ( .A1(n16414), .A2(n16397), .A3(n16407), .ZN(n16406) );
  NAND2_X1 U17253 ( .A1(n20372), .A2(n20370), .ZN(n15377) );
  INV_X1 U17254 ( .A(n15377), .ZN(n15361) );
  NAND2_X1 U17255 ( .A1(n15361), .A2(n20371), .ZN(n15217) );
  INV_X1 U17256 ( .A(n15217), .ZN(n14221) );
  NOR2_X1 U17257 ( .A1(n16406), .A2(n14221), .ZN(n16388) );
  NAND2_X1 U17258 ( .A1(n20390), .A2(n20369), .ZN(n16411) );
  NAND2_X1 U17259 ( .A1(n16411), .A2(n15394), .ZN(n16372) );
  NAND2_X1 U17260 ( .A1(n15390), .A2(n16372), .ZN(n16396) );
  NOR2_X1 U17261 ( .A1(n16397), .A2(n16396), .ZN(n16390) );
  INV_X1 U17262 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16391) );
  INV_X1 U17263 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20991) );
  OAI22_X1 U17264 ( .A1(n20393), .A2(n20991), .B1(n16412), .B2(n20298), .ZN(
        n14020) );
  AOI221_X1 U17265 ( .B1(n16388), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(
        n16390), .C2(n16391), .A(n14020), .ZN(n14021) );
  OAI21_X1 U17266 ( .B1(n14022), .B2(n20408), .A(n14021), .ZN(P1_U3024) );
  INV_X1 U17267 ( .A(n14023), .ZN(n14030) );
  NAND2_X1 U17268 ( .A1(n14025), .A2(n14024), .ZN(n14026) );
  NAND2_X1 U17269 ( .A1(n14030), .A2(n14026), .ZN(n20264) );
  INV_X1 U17270 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20266) );
  OAI222_X1 U17271 ( .A1(n20264), .A2(n14896), .B1(n20266), .B2(n20356), .C1(
        n20272), .C2(n14890), .ZN(P1_U2863) );
  NOR2_X1 U17272 ( .A1(n9763), .A2(n14028), .ZN(n14029) );
  OR2_X1 U17273 ( .A1(n14027), .A2(n14029), .ZN(n15206) );
  AOI21_X1 U17274 ( .B1(n14031), .B2(n14030), .A(n10175), .ZN(n16380) );
  AOI22_X1 U17275 ( .A1(n16380), .A2(n20351), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14885), .ZN(n14032) );
  OAI21_X1 U17276 ( .B1(n15206), .B2(n14890), .A(n14032), .ZN(P1_U2862) );
  AOI22_X1 U17277 ( .A1(n14993), .A2(n14911), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14991), .ZN(n14033) );
  OAI21_X1 U17278 ( .B1(n15206), .B2(n14995), .A(n14033), .ZN(P1_U2894) );
  INV_X1 U17279 ( .A(n14034), .ZN(n15203) );
  AOI22_X1 U17280 ( .A1(n20334), .A2(n16380), .B1(n20335), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n14035) );
  OAI211_X1 U17281 ( .C1(n20279), .C2(n15200), .A(n14035), .B(n20322), .ZN(
        n14039) );
  INV_X1 U17282 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20277) );
  INV_X1 U17283 ( .A(n20320), .ZN(n20280) );
  NOR2_X1 U17284 ( .A1(n20277), .A2(n20270), .ZN(n14037) );
  NAND3_X1 U17285 ( .A1(n20262), .A2(n14036), .A3(n20261), .ZN(n14847) );
  AND2_X1 U17286 ( .A1(n20292), .A2(n14847), .ZN(n16302) );
  MUX2_X1 U17287 ( .A(n14037), .B(n16302), .S(P1_REIP_REG_10__SCAN_IN), .Z(
        n14038) );
  AOI211_X1 U17288 ( .C1(n20339), .C2(n15203), .A(n14039), .B(n14038), .ZN(
        n14040) );
  OAI21_X1 U17289 ( .B1(n20287), .B2(n15206), .A(n14040), .ZN(P1_U2830) );
  INV_X1 U17290 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14042) );
  INV_X1 U17291 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14041) );
  OAI22_X1 U17292 ( .A1(n14042), .A2(n14417), .B1(n14411), .B2(n14041), .ZN(
        n14043) );
  INV_X1 U17293 ( .A(n14043), .ZN(n14054) );
  INV_X1 U17294 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14045) );
  OAI22_X1 U17295 ( .A1(n14045), .A2(n14416), .B1(n14412), .B2(n14044), .ZN(
        n14046) );
  INV_X1 U17296 ( .A(n14046), .ZN(n14053) );
  NAND2_X1 U17297 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14048) );
  NAND2_X1 U17298 ( .A1(n14421), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14047) );
  OAI211_X1 U17299 ( .C1(n14398), .C2(n14049), .A(n14048), .B(n14047), .ZN(
        n14050) );
  INV_X1 U17300 ( .A(n14050), .ZN(n14052) );
  AOI22_X1 U17301 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n14430), .B1(
        n10494), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14051) );
  NAND4_X1 U17302 ( .A1(n14054), .A2(n14053), .A3(n14052), .A4(n14051), .ZN(
        n14060) );
  AOI22_X1 U17303 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10578), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14058) );
  AOI22_X1 U17304 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10645), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14057) );
  AOI22_X1 U17305 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n14404), .B1(
        n14432), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14056) );
  NAND2_X1 U17306 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14055) );
  NAND4_X1 U17307 ( .A1(n14058), .A2(n14057), .A3(n14056), .A4(n14055), .ZN(
        n14059) );
  NOR2_X1 U17308 ( .A1(n14060), .A2(n14059), .ZN(n14126) );
  OR2_X1 U17309 ( .A1(n13913), .A2(n14126), .ZN(n14128) );
  INV_X1 U17310 ( .A(n14128), .ZN(n14061) );
  AOI21_X1 U17311 ( .B1(n14126), .B2(n13913), .A(n14061), .ZN(n15672) );
  NAND2_X1 U17312 ( .A1(n15672), .A2(n15575), .ZN(n14065) );
  NAND2_X1 U17313 ( .A1(n13869), .A2(n14062), .ZN(n14063) );
  AND2_X1 U17314 ( .A1(n14104), .A2(n14063), .ZN(n19205) );
  NAND2_X1 U17315 ( .A1(n19205), .A2(n15572), .ZN(n14064) );
  OAI211_X1 U17316 ( .C1(n15572), .C2(n14066), .A(n14065), .B(n14064), .ZN(
        P2_U2869) );
  XNOR2_X1 U17317 ( .A(n14068), .B(n14067), .ZN(n16527) );
  OAI21_X1 U17318 ( .B1(n14070), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14071), .ZN(n14072) );
  INV_X1 U17319 ( .A(n14072), .ZN(n16530) );
  NAND2_X1 U17320 ( .A1(n16530), .A2(n16550), .ZN(n14086) );
  XNOR2_X1 U17321 ( .A(n14074), .B(n14073), .ZN(n19370) );
  NOR2_X1 U17322 ( .A1(n19508), .A2(n19370), .ZN(n14083) );
  NOR3_X1 U17323 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14075), .A3(
        n16552), .ZN(n14080) );
  NAND2_X1 U17324 ( .A1(n19499), .A2(n14075), .ZN(n14078) );
  INV_X1 U17325 ( .A(n14076), .ZN(n14077) );
  NAND2_X1 U17326 ( .A1(n14078), .A2(n14077), .ZN(n14079) );
  OR2_X1 U17327 ( .A1(n14080), .A2(n14079), .ZN(n16560) );
  OAI21_X1 U17328 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14080), .A(
        n16560), .ZN(n14081) );
  OAI21_X1 U17329 ( .B1(n19277), .B2(n20127), .A(n14081), .ZN(n14082) );
  AOI211_X1 U17330 ( .C1(n14084), .C2(n19505), .A(n14083), .B(n14082), .ZN(
        n14085) );
  OAI211_X1 U17331 ( .C1(n16527), .C2(n19502), .A(n14086), .B(n14085), .ZN(
        P2_U3040) );
  NAND2_X1 U17332 ( .A1(n14088), .A2(n14087), .ZN(n14090) );
  NAND2_X1 U17333 ( .A1(n14090), .A2(n14089), .ZN(n14214) );
  NOR2_X1 U17334 ( .A1(n14091), .A2(n9971), .ZN(n14092) );
  OR3_X1 U17335 ( .A1(n14096), .A2(n14095), .A3(n14094), .ZN(n14097) );
  NAND2_X1 U17336 ( .A1(n15011), .A2(n14097), .ZN(n14215) );
  XNOR2_X1 U17337 ( .A(n14215), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14098) );
  XNOR2_X1 U17338 ( .A(n14214), .B(n14098), .ZN(n16389) );
  NAND2_X1 U17339 ( .A1(n16389), .A2(n16345), .ZN(n14102) );
  INV_X1 U17340 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n14099) );
  OAI22_X1 U17341 ( .A1(n15201), .A2(n21209), .B1(n20393), .B2(n14099), .ZN(
        n14100) );
  AOI21_X1 U17342 ( .B1(n20289), .B2(n16321), .A(n14100), .ZN(n14101) );
  OAI211_X1 U17343 ( .C1(n20422), .C2(n20286), .A(n14102), .B(n14101), .ZN(
        P1_U2991) );
  NAND2_X1 U17344 ( .A1(n14104), .A2(n14103), .ZN(n14105) );
  NAND2_X1 U17345 ( .A1(n15588), .A2(n14105), .ZN(n19193) );
  INV_X1 U17346 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14106) );
  OAI22_X1 U17347 ( .A1(n14107), .A2(n14417), .B1(n14411), .B2(n14106), .ZN(
        n14108) );
  INV_X1 U17348 ( .A(n14108), .ZN(n14119) );
  INV_X1 U17349 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14110) );
  OAI22_X1 U17350 ( .A1(n14110), .A2(n14416), .B1(n14412), .B2(n14109), .ZN(
        n14111) );
  INV_X1 U17351 ( .A(n14111), .ZN(n14118) );
  NAND2_X1 U17352 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14113) );
  NAND2_X1 U17353 ( .A1(n14421), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n14112) );
  OAI211_X1 U17354 ( .C1(n14398), .C2(n14114), .A(n14113), .B(n14112), .ZN(
        n14115) );
  INV_X1 U17355 ( .A(n14115), .ZN(n14117) );
  AOI22_X1 U17356 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10494), .B1(
        n14430), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14116) );
  NAND4_X1 U17357 ( .A1(n14119), .A2(n14118), .A3(n14117), .A4(n14116), .ZN(
        n14125) );
  AOI22_X1 U17358 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10578), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14123) );
  AOI22_X1 U17359 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10645), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U17360 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14432), .B1(
        n14404), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14121) );
  NAND2_X1 U17361 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14120) );
  NAND4_X1 U17362 ( .A1(n14123), .A2(n14122), .A3(n14121), .A4(n14120), .ZN(
        n14124) );
  NOR2_X1 U17363 ( .A1(n14125), .A2(n14124), .ZN(n14129) );
  AOI21_X1 U17364 ( .B1(n14129), .B2(n14128), .A(n14368), .ZN(n15665) );
  NAND2_X1 U17365 ( .A1(n15665), .A2(n15575), .ZN(n14131) );
  NAND2_X1 U17366 ( .A1(n15578), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14130) );
  OAI211_X1 U17367 ( .C1(n19193), .C2(n15578), .A(n14131), .B(n14130), .ZN(
        P2_U2868) );
  AND2_X1 U17368 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17227) );
  INV_X1 U17369 ( .A(n16198), .ZN(n18907) );
  NOR2_X1 U17370 ( .A1(n14132), .A2(n17597), .ZN(n14133) );
  NOR4_X2 U17371 ( .A1(n19112), .A2(n18475), .A3(n16269), .A4(n18967), .ZN(
        n17478) );
  INV_X1 U17372 ( .A(n17478), .ZN(n17481) );
  NOR2_X1 U17373 ( .A1(n17597), .A2(n17481), .ZN(n17464) );
  INV_X1 U17374 ( .A(n17464), .ZN(n17484) );
  INV_X1 U17375 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16902) );
  INV_X1 U17376 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17305) );
  INV_X1 U17377 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n14135) );
  INV_X1 U17378 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17419) );
  INV_X1 U17379 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17078) );
  INV_X1 U17380 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17451) );
  INV_X1 U17381 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17136) );
  INV_X1 U17382 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17466) );
  NAND3_X1 U17383 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17469) );
  NOR3_X1 U17384 ( .A1(n17136), .A2(n17466), .A3(n17469), .ZN(n17465) );
  AND2_X1 U17385 ( .A1(n17478), .A2(n17465), .ZN(n17462) );
  NAND4_X1 U17386 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(n17462), .ZN(n17452) );
  NAND4_X1 U17387 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .A4(P3_EBX_REG_12__SCAN_IN), .ZN(n17333)
         );
  NAND2_X1 U17388 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17331), .ZN(n17330) );
  NAND3_X1 U17389 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .ZN(n14245) );
  NOR2_X2 U17390 ( .A1(n17262), .A2(n14245), .ZN(n17251) );
  NAND2_X1 U17391 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17251), .ZN(n17238) );
  NAND2_X1 U17392 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17243), .ZN(n17234) );
  NAND2_X1 U17393 ( .A1(n17470), .A2(n17234), .ZN(n17232) );
  OAI21_X1 U17394 ( .B1(n17227), .B2(n17484), .A(n17232), .ZN(n17228) );
  AOI22_X1 U17395 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14139) );
  AOI22_X1 U17396 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14138) );
  AOI22_X1 U17397 ( .A1(n12239), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14137) );
  AOI22_X1 U17398 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14136) );
  NAND4_X1 U17399 ( .A1(n14139), .A2(n14138), .A3(n14137), .A4(n14136), .ZN(
        n14145) );
  AOI22_X1 U17400 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14143) );
  AOI22_X1 U17401 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14142) );
  AOI22_X1 U17402 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14141) );
  AOI22_X1 U17403 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14140) );
  NAND4_X1 U17404 ( .A1(n14143), .A2(n14142), .A3(n14141), .A4(n14140), .ZN(
        n14144) );
  NOR2_X1 U17405 ( .A1(n14145), .A2(n14144), .ZN(n14209) );
  AOI22_X1 U17406 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14149) );
  AOI22_X1 U17407 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14148) );
  AOI22_X1 U17408 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17440), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14147) );
  AOI22_X1 U17409 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14146) );
  NAND4_X1 U17410 ( .A1(n14149), .A2(n14148), .A3(n14147), .A4(n14146), .ZN(
        n14155) );
  AOI22_X1 U17411 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14153) );
  AOI22_X1 U17412 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14152) );
  AOI22_X1 U17413 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14151) );
  AOI22_X1 U17414 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14150) );
  NAND4_X1 U17415 ( .A1(n14153), .A2(n14152), .A3(n14151), .A4(n14150), .ZN(
        n14154) );
  NOR2_X1 U17416 ( .A1(n14155), .A2(n14154), .ZN(n17235) );
  AOI22_X1 U17417 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14159) );
  AOI22_X1 U17418 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9673), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14158) );
  AOI22_X1 U17419 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14157) );
  AOI22_X1 U17420 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14156) );
  NAND4_X1 U17421 ( .A1(n14159), .A2(n14158), .A3(n14157), .A4(n14156), .ZN(
        n14165) );
  AOI22_X1 U17422 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14163) );
  AOI22_X1 U17423 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14162) );
  AOI22_X1 U17424 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14161) );
  AOI22_X1 U17425 ( .A1(n17440), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14160) );
  NAND4_X1 U17426 ( .A1(n14163), .A2(n14162), .A3(n14161), .A4(n14160), .ZN(
        n14164) );
  NOR2_X1 U17427 ( .A1(n14165), .A2(n14164), .ZN(n17244) );
  AOI22_X1 U17428 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14176) );
  AOI22_X1 U17429 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14175) );
  AOI22_X1 U17430 ( .A1(n17423), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14167) );
  OAI21_X1 U17431 ( .B1(n17208), .B2(n18478), .A(n14167), .ZN(n14173) );
  AOI22_X1 U17432 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17440), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14171) );
  AOI22_X1 U17433 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14170) );
  AOI22_X1 U17434 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14169) );
  AOI22_X1 U17435 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14168) );
  NAND4_X1 U17436 ( .A1(n14171), .A2(n14170), .A3(n14169), .A4(n14168), .ZN(
        n14172) );
  AOI211_X1 U17437 ( .C1(n17411), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n14173), .B(n14172), .ZN(n14174) );
  NAND3_X1 U17438 ( .A1(n14176), .A2(n14175), .A3(n14174), .ZN(n17248) );
  AOI22_X1 U17439 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14187) );
  AOI22_X1 U17440 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17411), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14186) );
  AOI22_X1 U17441 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17441), .ZN(n14177) );
  OAI21_X1 U17442 ( .B1(n17209), .B2(n14178), .A(n14177), .ZN(n14184) );
  AOI22_X1 U17443 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17440), .ZN(n14182) );
  AOI22_X1 U17444 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n14205), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14181) );
  AOI22_X1 U17445 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n16181), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17423), .ZN(n14180) );
  AOI22_X1 U17446 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14179) );
  NAND4_X1 U17447 ( .A1(n14182), .A2(n14181), .A3(n14180), .A4(n14179), .ZN(
        n14183) );
  AOI211_X1 U17448 ( .C1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .C2(n17319), .A(
        n14184), .B(n14183), .ZN(n14185) );
  NAND3_X1 U17449 ( .A1(n14187), .A2(n14186), .A3(n14185), .ZN(n17249) );
  NAND2_X1 U17450 ( .A1(n17248), .A2(n17249), .ZN(n17247) );
  NOR2_X1 U17451 ( .A1(n17244), .A2(n17247), .ZN(n17241) );
  AOI22_X1 U17452 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14197) );
  AOI22_X1 U17453 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14196) );
  AOI22_X1 U17454 ( .A1(n17440), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14188) );
  OAI21_X1 U17455 ( .B1(n17208), .B2(n18488), .A(n14188), .ZN(n14194) );
  AOI22_X1 U17456 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14192) );
  AOI22_X1 U17457 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14191) );
  AOI22_X1 U17458 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9687), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14190) );
  AOI22_X1 U17459 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14189) );
  NAND4_X1 U17460 ( .A1(n14192), .A2(n14191), .A3(n14190), .A4(n14189), .ZN(
        n14193) );
  AOI211_X1 U17461 ( .C1(n14205), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n14194), .B(n14193), .ZN(n14195) );
  NAND3_X1 U17462 ( .A1(n14197), .A2(n14196), .A3(n14195), .ZN(n17240) );
  NAND2_X1 U17463 ( .A1(n17241), .A2(n17240), .ZN(n17239) );
  NOR2_X1 U17464 ( .A1(n17235), .A2(n17239), .ZN(n17511) );
  AOI22_X1 U17465 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14208) );
  AOI22_X1 U17466 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14207) );
  AOI22_X1 U17467 ( .A1(n17440), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14198) );
  OAI21_X1 U17468 ( .B1(n17208), .B2(n18500), .A(n14198), .ZN(n14204) );
  AOI22_X1 U17469 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14202) );
  AOI22_X1 U17470 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14201) );
  AOI22_X1 U17471 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14200) );
  AOI22_X1 U17472 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14199) );
  NAND4_X1 U17473 ( .A1(n14202), .A2(n14201), .A3(n14200), .A4(n14199), .ZN(
        n14203) );
  AOI211_X1 U17474 ( .C1(n14205), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n14204), .B(n14203), .ZN(n14206) );
  NAND3_X1 U17475 ( .A1(n14208), .A2(n14207), .A3(n14206), .ZN(n17510) );
  NAND2_X1 U17476 ( .A1(n17511), .A2(n17510), .ZN(n17509) );
  NOR2_X1 U17477 ( .A1(n14209), .A2(n17509), .ZN(n17225) );
  AOI21_X1 U17478 ( .B1(n14209), .B2(n17509), .A(n17225), .ZN(n17505) );
  AOI22_X1 U17479 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17228), .B1(n17482), 
        .B2(n17505), .ZN(n14212) );
  INV_X1 U17480 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14210) );
  INV_X1 U17481 ( .A(n17234), .ZN(n17237) );
  NAND3_X1 U17482 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14210), .A3(n17237), 
        .ZN(n14211) );
  NAND2_X1 U17483 ( .A1(n14212), .A2(n14211), .ZN(P3_U2675) );
  INV_X1 U17484 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16384) );
  MUX2_X1 U17485 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n16384), .S(
        n16312), .Z(n14218) );
  OR2_X1 U17486 ( .A1(n14215), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14213) );
  NAND2_X1 U17487 ( .A1(n14215), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14216) );
  XOR2_X1 U17488 ( .A(n14218), .B(n14997), .Z(n14229) );
  INV_X1 U17489 ( .A(n20372), .ZN(n20373) );
  NAND2_X1 U17490 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14219), .ZN(
        n15308) );
  NAND3_X1 U17491 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15207) );
  INV_X1 U17492 ( .A(n14220), .ZN(n15392) );
  AOI211_X1 U17493 ( .C1(n20373), .C2(n15308), .A(n15207), .B(n15392), .ZN(
        n14222) );
  NOR2_X1 U17494 ( .A1(n14222), .A2(n14221), .ZN(n16381) );
  NOR2_X1 U17495 ( .A1(n15207), .A2(n16396), .ZN(n16383) );
  OAI22_X1 U17496 ( .A1(n20393), .A2(n20277), .B1(n16412), .B2(n20264), .ZN(
        n14223) );
  AOI221_X1 U17497 ( .B1(n16381), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n16383), .C2(n16384), .A(n14223), .ZN(n14224) );
  OAI21_X1 U17498 ( .B1(n14229), .B2(n20408), .A(n14224), .ZN(P1_U3022) );
  AOI22_X1 U17499 ( .A1(n20357), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20407), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14226) );
  NAND2_X1 U17500 ( .A1(n16321), .A2(n20273), .ZN(n14225) );
  OAI211_X1 U17501 ( .C1(n20272), .C2(n20422), .A(n14226), .B(n14225), .ZN(
        n14227) );
  INV_X1 U17502 ( .A(n14227), .ZN(n14228) );
  OAI21_X1 U17503 ( .B1(n14229), .B2(n20363), .A(n14228), .ZN(P1_U2990) );
  XNOR2_X1 U17504 ( .A(n14231), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14232) );
  XNOR2_X1 U17505 ( .A(n14230), .B(n14232), .ZN(n16572) );
  INV_X1 U17506 ( .A(n14235), .ZN(n16517) );
  AND2_X1 U17507 ( .A1(n14235), .A2(n14234), .ZN(n14236) );
  OAI22_X1 U17508 ( .A1(n9864), .A2(n16517), .B1(n14237), .B2(n14236), .ZN(
        n16569) );
  OAI22_X1 U17509 ( .A1(n16541), .A2(n10727), .B1(n20129), .B2(n19277), .ZN(
        n14240) );
  INV_X1 U17510 ( .A(n19274), .ZN(n14238) );
  OAI22_X1 U17511 ( .A1(n16526), .A2(n19279), .B1(n19496), .B2(n14238), .ZN(
        n14239) );
  AOI211_X1 U17512 ( .C1(n16569), .C2(n10990), .A(n14240), .B(n14239), .ZN(
        n14241) );
  OAI21_X1 U17513 ( .B1(n19490), .B2(n16572), .A(n14241), .ZN(P2_U3007) );
  NAND2_X1 U17514 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17227), .ZN(n14244) );
  INV_X1 U17515 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n14242) );
  NOR2_X1 U17516 ( .A1(n14242), .A2(n17303), .ZN(n17276) );
  NAND4_X1 U17517 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(n17276), .ZN(n14243) );
  NOR3_X1 U17518 ( .A1(n14245), .A2(n14244), .A3(n14243), .ZN(n17220) );
  NAND2_X1 U17519 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17220), .ZN(n14246) );
  NOR2_X1 U17520 ( .A1(n17597), .A2(n14246), .ZN(n14248) );
  NAND2_X1 U17521 ( .A1(n17470), .A2(n14246), .ZN(n17221) );
  INV_X1 U17522 ( .A(n17221), .ZN(n14247) );
  MUX2_X1 U17523 ( .A(n14248), .B(n14247), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  OAI21_X1 U17524 ( .B1(n14265), .B2(n12318), .A(n18916), .ZN(n14251) );
  NAND2_X1 U17525 ( .A1(n16822), .A2(n14251), .ZN(n18914) );
  NOR2_X1 U17526 ( .A1(n19078), .A2(n18914), .ZN(n14263) );
  INV_X1 U17527 ( .A(n16786), .ZN(n18910) );
  NAND2_X1 U17528 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19113) );
  NAND2_X1 U17529 ( .A1(n18910), .A2(n19113), .ZN(n14261) );
  NAND2_X1 U17530 ( .A1(n19112), .A2(n17706), .ZN(n18960) );
  INV_X1 U17531 ( .A(n18960), .ZN(n14252) );
  INV_X2 U17532 ( .A(n19120), .ZN(n19121) );
  AND2_X1 U17533 ( .A1(n19121), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19002) );
  NOR2_X1 U17534 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18980) );
  NOR3_X1 U17535 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19002), .A3(n18980), 
        .ZN(n16824) );
  OAI21_X1 U17536 ( .B1(n14253), .B2(n14252), .A(n16824), .ZN(n17640) );
  INV_X1 U17537 ( .A(n19113), .ZN(n18988) );
  INV_X1 U17538 ( .A(n14255), .ZN(n14258) );
  OAI211_X1 U17539 ( .C1(n16792), .C2(n14258), .A(n9655), .B(n14256), .ZN(
        n16195) );
  AOI211_X1 U17540 ( .C1(n18907), .C2(n14259), .A(n16271), .B(n16195), .ZN(
        n14260) );
  OAI21_X1 U17541 ( .B1(n14261), .B2(n17640), .A(n14260), .ZN(n18934) );
  NOR2_X1 U17542 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19068), .ZN(n18474) );
  INV_X1 U17543 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18460) );
  NAND3_X1 U17544 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19066)
         );
  NOR2_X1 U17545 ( .A1(n18460), .A2(n19066), .ZN(n14262) );
  AOI211_X1 U17546 ( .C1(n19107), .C2(n18934), .A(n18474), .B(n14262), .ZN(
        n19094) );
  MUX2_X1 U17547 ( .A(n14263), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19094), .Z(P3_U3284) );
  OAI211_X1 U17548 ( .C1(n14265), .C2(n12318), .A(n14264), .B(n18916), .ZN(
        n18459) );
  NOR2_X1 U17549 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18459), .ZN(n14266) );
  OAI21_X1 U17550 ( .B1(n14266), .B2(n19066), .A(n18597), .ZN(n18470) );
  INV_X1 U17551 ( .A(n18470), .ZN(n14267) );
  NOR2_X1 U17552 ( .A1(n19106), .A2(n18080), .ZN(n18463) );
  AOI21_X1 U17553 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18463), .ZN(n18464) );
  NOR2_X1 U17554 ( .A1(n14267), .A2(n18464), .ZN(n14269) );
  INV_X1 U17555 ( .A(n18823), .ZN(n18465) );
  NOR2_X1 U17556 ( .A1(n19068), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18524) );
  OR2_X1 U17557 ( .A1(n18524), .A2(n14267), .ZN(n18462) );
  OR2_X1 U17558 ( .A1(n18465), .A2(n18462), .ZN(n14268) );
  MUX2_X1 U17559 ( .A(n14269), .B(n14268), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NAND2_X1 U17560 ( .A1(n14271), .A2(n14270), .ZN(n15684) );
  AOI21_X1 U17561 ( .B1(n14273), .B2(n14277), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15687) );
  AND2_X1 U17562 ( .A1(n14277), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14272) );
  NAND2_X1 U17563 ( .A1(n14273), .A2(n14272), .ZN(n15685) );
  NOR2_X1 U17564 ( .A1(n14274), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14275) );
  MUX2_X1 U17565 ( .A(n14276), .B(n14275), .S(n10812), .Z(n15432) );
  NAND2_X1 U17566 ( .A1(n15432), .A2(n14277), .ZN(n14278) );
  XNOR2_X1 U17567 ( .A(n14278), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14279) );
  XNOR2_X1 U17568 ( .A(n14280), .B(n14279), .ZN(n14665) );
  AOI22_X1 U17569 ( .A1(n9663), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14284) );
  NAND2_X1 U17570 ( .A1(n10736), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14283) );
  OAI211_X1 U17571 ( .C1(n14286), .C2(n14285), .A(n14284), .B(n14283), .ZN(
        n14287) );
  XNOR2_X1 U17572 ( .A(n14288), .B(n14287), .ZN(n15435) );
  INV_X1 U17573 ( .A(n15435), .ZN(n15525) );
  NAND2_X1 U17574 ( .A1(n16002), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16005) );
  NOR2_X1 U17575 ( .A1(n16008), .A2(n16005), .ZN(n14289) );
  NAND3_X1 U17576 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n14289), .ZN(n15989) );
  NOR2_X1 U17577 ( .A1(n15781), .A2(n15989), .ZN(n15968) );
  NAND3_X1 U17578 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n15968), .ZN(n14303) );
  NAND2_X1 U17579 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14290), .ZN(
        n16553) );
  NAND2_X1 U17580 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16554) );
  OR4_X1 U17581 ( .A1(n14638), .A2(n14291), .A3(n16553), .A4(n16554), .ZN(
        n14299) );
  NOR2_X1 U17582 ( .A1(n14299), .A2(n14292), .ZN(n16164) );
  INV_X1 U17583 ( .A(n16164), .ZN(n15959) );
  OR2_X1 U17584 ( .A1(n14303), .A2(n15959), .ZN(n15953) );
  AND2_X1 U17585 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15923) );
  NAND2_X1 U17586 ( .A1(n15923), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14293) );
  NOR2_X1 U17587 ( .A1(n15953), .A2(n14293), .ZN(n15893) );
  AND2_X1 U17588 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14294) );
  NAND2_X1 U17589 ( .A1(n15893), .A2(n14294), .ZN(n15883) );
  NOR4_X1 U17590 ( .A1(n15883), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15882), .A4(n15690), .ZN(n14312) );
  AOI222_X1 U17591 ( .A1(n14296), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n14295), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n9657), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14297) );
  NAND2_X1 U17592 ( .A1(n16093), .A2(n14301), .ZN(n14309) );
  INV_X1 U17593 ( .A(n14299), .ZN(n14300) );
  NAND2_X1 U17594 ( .A1(n14301), .A2(n14300), .ZN(n14302) );
  NAND2_X1 U17595 ( .A1(n14309), .A2(n14302), .ZN(n16172) );
  NAND2_X1 U17596 ( .A1(n19499), .A2(n14303), .ZN(n14304) );
  AND2_X1 U17597 ( .A1(n16172), .A2(n14304), .ZN(n15948) );
  NAND2_X1 U17598 ( .A1(n19499), .A2(n15947), .ZN(n14305) );
  AND2_X1 U17599 ( .A1(n15948), .A2(n14305), .ZN(n15938) );
  OAI21_X1 U17600 ( .B1(n15937), .B2(n15922), .A(n14309), .ZN(n14306) );
  AND2_X1 U17601 ( .A1(n15938), .A2(n14306), .ZN(n15907) );
  OR3_X1 U17602 ( .A1(n15882), .A2(n14612), .A3(n15894), .ZN(n14307) );
  AOI21_X1 U17603 ( .B1(n19499), .B2(n14307), .A(n15690), .ZN(n14308) );
  NAND2_X1 U17604 ( .A1(n15907), .A2(n14308), .ZN(n15884) );
  NAND3_X1 U17605 ( .A1(n15884), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14309), .ZN(n14310) );
  NAND2_X1 U17606 ( .A1(n19303), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14657) );
  OAI211_X1 U17607 ( .C1(n19333), .C2(n19508), .A(n14310), .B(n14657), .ZN(
        n14311) );
  NAND2_X1 U17608 ( .A1(n14663), .A2(n16550), .ZN(n14314) );
  OAI211_X1 U17609 ( .C1(n14665), .C2(n19502), .A(n14315), .B(n14314), .ZN(
        P2_U3015) );
  AOI21_X1 U17610 ( .B1(n14319), .B2(n9730), .A(n14318), .ZN(n15244) );
  INV_X1 U17611 ( .A(n14320), .ZN(n15044) );
  OAI22_X1 U17612 ( .A1(n14321), .A2(n20279), .B1(n20330), .B2(n15044), .ZN(
        n14324) );
  NOR2_X1 U17613 ( .A1(n14322), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14323) );
  AOI211_X1 U17614 ( .C1(P1_EBX_REG_29__SCAN_IN), .C2(n20335), .A(n14324), .B(
        n14323), .ZN(n14325) );
  OAI21_X1 U17615 ( .B1(n14672), .B2(n21025), .A(n14325), .ZN(n14326) );
  AOI21_X1 U17616 ( .B1(n15244), .B2(n20334), .A(n14326), .ZN(n14327) );
  OAI21_X1 U17617 ( .B1(n15047), .B2(n20287), .A(n14327), .ZN(P1_U2811) );
  AOI22_X1 U17618 ( .A1(n15244), .A2(n20351), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14885), .ZN(n14328) );
  OAI21_X1 U17619 ( .B1(n15047), .B2(n14890), .A(n14328), .ZN(P1_U2843) );
  INV_X1 U17620 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n14331) );
  AND2_X1 U17621 ( .A1(n20450), .A2(n11165), .ZN(n14329) );
  AOI22_X1 U17622 ( .A1(n14959), .A2(n14978), .B1(n14991), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n14330) );
  OAI21_X1 U17623 ( .B1(n14331), .B2(n14962), .A(n14330), .ZN(n14332) );
  AOI21_X1 U17624 ( .B1(n14970), .B2(DATAI_29_), .A(n14332), .ZN(n14333) );
  OAI21_X1 U17625 ( .B1(n15047), .B2(n14995), .A(n14333), .ZN(P1_U2875) );
  OAI21_X1 U17626 ( .B1(n14336), .B2(n14335), .A(n14334), .ZN(n14337) );
  XOR2_X1 U17627 ( .A(n14337), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n19503) );
  NOR2_X1 U17628 ( .A1(n16541), .A2(n14338), .ZN(n14342) );
  OAI21_X1 U17629 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14340), .A(
        n14339), .ZN(n19516) );
  NAND2_X1 U17630 ( .A1(n19303), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19513) );
  OAI21_X1 U17631 ( .B1(n19490), .B2(n19516), .A(n19513), .ZN(n14341) );
  AOI211_X1 U17632 ( .C1(n16533), .C2(n14338), .A(n14342), .B(n14341), .ZN(
        n14344) );
  NAND2_X1 U17633 ( .A1(n19506), .A2(n19486), .ZN(n14343) );
  OAI211_X1 U17634 ( .C1(n19503), .C2(n16537), .A(n14344), .B(n14343), .ZN(
        P2_U3013) );
  AOI21_X1 U17635 ( .B1(n16211), .B2(n16419), .A(n16417), .ZN(n14347) );
  OAI22_X1 U17636 ( .A1(n20523), .A2(n15413), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15412), .ZN(n16212) );
  OAI22_X1 U17637 ( .A1(n20962), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15422), .ZN(n14345) );
  AOI21_X1 U17638 ( .B1(n16212), .B2(n16419), .A(n14345), .ZN(n14346) );
  OAI22_X1 U17639 ( .A1(n14347), .A2(n16215), .B1(n16417), .B2(n14346), .ZN(
        P1_U3474) );
  AOI22_X1 U17640 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10578), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14351) );
  AOI22_X1 U17641 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10645), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14350) );
  AOI22_X1 U17642 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14432), .B1(
        n14404), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14349) );
  NAND2_X1 U17643 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14348) );
  AND4_X1 U17644 ( .A1(n14351), .A2(n14350), .A3(n14349), .A4(n14348), .ZN(
        n14367) );
  AOI22_X1 U17645 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n14431), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14357) );
  NAND2_X1 U17646 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14356) );
  INV_X1 U17647 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14352) );
  OR2_X1 U17648 ( .A1(n14417), .A2(n14352), .ZN(n14355) );
  INV_X1 U17649 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14353) );
  OR2_X1 U17650 ( .A1(n14411), .A2(n14353), .ZN(n14354) );
  NAND4_X1 U17651 ( .A1(n14357), .A2(n14356), .A3(n14355), .A4(n14354), .ZN(
        n14365) );
  OR2_X1 U17652 ( .A1(n14412), .A2(n14358), .ZN(n14363) );
  INV_X1 U17653 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14359) );
  OR2_X1 U17654 ( .A1(n14416), .A2(n14359), .ZN(n14362) );
  NAND2_X1 U17655 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14361) );
  NAND2_X1 U17656 ( .A1(n14430), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n14360) );
  NAND4_X1 U17657 ( .A1(n14363), .A2(n14362), .A3(n14361), .A4(n14360), .ZN(
        n14364) );
  NOR2_X1 U17658 ( .A1(n14365), .A2(n14364), .ZN(n14366) );
  NAND2_X1 U17659 ( .A1(n14367), .A2(n14366), .ZN(n15585) );
  AOI22_X1 U17660 ( .A1(n10578), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U17661 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14371) );
  AOI22_X1 U17662 ( .A1(n14432), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14404), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14370) );
  NAND2_X1 U17663 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14369) );
  AND4_X1 U17664 ( .A1(n14372), .A2(n14371), .A3(n14370), .A4(n14369), .ZN(
        n14388) );
  AOI22_X1 U17665 ( .A1(n14431), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14421), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14378) );
  NAND2_X1 U17666 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14377) );
  OR2_X1 U17667 ( .A1(n14417), .A2(n14373), .ZN(n14376) );
  INV_X1 U17668 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14374) );
  OR2_X1 U17669 ( .A1(n14411), .A2(n14374), .ZN(n14375) );
  NAND4_X1 U17670 ( .A1(n14378), .A2(n14377), .A3(n14376), .A4(n14375), .ZN(
        n14386) );
  OR2_X1 U17671 ( .A1(n14412), .A2(n14379), .ZN(n14384) );
  INV_X1 U17672 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14380) );
  OR2_X1 U17673 ( .A1(n14416), .A2(n14380), .ZN(n14383) );
  NAND2_X1 U17674 ( .A1(n10494), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n14382) );
  NAND2_X1 U17675 ( .A1(n14430), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n14381) );
  NAND4_X1 U17676 ( .A1(n14384), .A2(n14383), .A3(n14382), .A4(n14381), .ZN(
        n14385) );
  NOR2_X1 U17677 ( .A1(n14386), .A2(n14385), .ZN(n14387) );
  NAND2_X1 U17678 ( .A1(n14388), .A2(n14387), .ZN(n15580) );
  INV_X1 U17679 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14389) );
  OAI22_X1 U17680 ( .A1(n14390), .A2(n14417), .B1(n14411), .B2(n14389), .ZN(
        n14391) );
  INV_X1 U17681 ( .A(n14391), .ZN(n14403) );
  INV_X1 U17682 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14393) );
  OAI22_X1 U17683 ( .A1(n14393), .A2(n14416), .B1(n14412), .B2(n14392), .ZN(
        n14394) );
  INV_X1 U17684 ( .A(n14394), .ZN(n14402) );
  NAND2_X1 U17685 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n14396) );
  NAND2_X1 U17686 ( .A1(n14421), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n14395) );
  OAI211_X1 U17687 ( .C1(n14398), .C2(n14397), .A(n14396), .B(n14395), .ZN(
        n14399) );
  INV_X1 U17688 ( .A(n14399), .ZN(n14401) );
  AOI22_X1 U17689 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n14430), .B1(
        n10494), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14400) );
  NAND4_X1 U17690 ( .A1(n14403), .A2(n14402), .A3(n14401), .A4(n14400), .ZN(
        n14410) );
  AOI22_X1 U17691 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10578), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14408) );
  AOI22_X1 U17692 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10645), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U17693 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n14404), .B1(
        n14432), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14406) );
  NAND2_X1 U17694 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n14405) );
  NAND4_X1 U17695 ( .A1(n14408), .A2(n14407), .A3(n14406), .A4(n14405), .ZN(
        n14409) );
  NOR2_X1 U17696 ( .A1(n14410), .A2(n14409), .ZN(n15574) );
  INV_X1 U17697 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14587) );
  OAI22_X1 U17698 ( .A1(n14413), .A2(n14412), .B1(n14411), .B2(n14587), .ZN(
        n14414) );
  INV_X1 U17699 ( .A(n14414), .ZN(n14429) );
  INV_X1 U17700 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14418) );
  INV_X1 U17701 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14415) );
  OAI22_X1 U17702 ( .A1(n14418), .A2(n14417), .B1(n14416), .B2(n14415), .ZN(
        n14419) );
  INV_X1 U17703 ( .A(n14419), .ZN(n14428) );
  NAND2_X1 U17704 ( .A1(n14420), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14423) );
  NAND2_X1 U17705 ( .A1(n14421), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n14422) );
  OAI211_X1 U17706 ( .C1(n10164), .C2(n14424), .A(n14423), .B(n14422), .ZN(
        n14425) );
  INV_X1 U17707 ( .A(n14425), .ZN(n14427) );
  AOI22_X1 U17708 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10494), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14426) );
  NAND4_X1 U17709 ( .A1(n14429), .A2(n14428), .A3(n14427), .A4(n14426), .ZN(
        n14439) );
  AOI22_X1 U17710 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10578), .B1(
        n14430), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14437) );
  AOI22_X1 U17711 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10645), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14436) );
  AOI22_X1 U17712 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n14432), .B1(
        n14431), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14435) );
  NAND2_X1 U17713 ( .A1(n14433), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14434) );
  NAND4_X1 U17714 ( .A1(n14437), .A2(n14436), .A3(n14435), .A4(n14434), .ZN(
        n14438) );
  NOR2_X1 U17715 ( .A1(n14439), .A2(n14438), .ZN(n14459) );
  INV_X1 U17716 ( .A(n14459), .ZN(n14458) );
  AOI22_X1 U17717 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9692), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14449) );
  AND2_X1 U17718 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14441) );
  OR2_X1 U17719 ( .A1(n14441), .A2(n14440), .ZN(n14596) );
  INV_X1 U17720 ( .A(n14596), .ZN(n14564) );
  NAND2_X1 U17721 ( .A1(n14595), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14444) );
  NAND2_X1 U17722 ( .A1(n14589), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14443) );
  AND3_X1 U17723 ( .A1(n14564), .A2(n14444), .A3(n14443), .ZN(n14448) );
  AOI22_X1 U17724 ( .A1(n14590), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14447) );
  INV_X1 U17725 ( .A(n14588), .ZN(n14594) );
  AOI22_X1 U17726 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14446) );
  NAND4_X1 U17727 ( .A1(n14449), .A2(n14448), .A3(n14447), .A4(n14446), .ZN(
        n14457) );
  AOI22_X1 U17728 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9691), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14455) );
  AOI22_X1 U17729 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14589), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14454) );
  AOI22_X1 U17730 ( .A1(n14593), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14453) );
  NAND2_X1 U17731 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14451) );
  NAND2_X1 U17732 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n14450) );
  AND3_X1 U17733 ( .A1(n14451), .A2(n14596), .A3(n14450), .ZN(n14452) );
  NAND4_X1 U17734 ( .A1(n14455), .A2(n14454), .A3(n14453), .A4(n14452), .ZN(
        n14456) );
  NAND2_X1 U17735 ( .A1(n14457), .A2(n14456), .ZN(n14481) );
  INV_X1 U17736 ( .A(n14481), .ZN(n14462) );
  NAND2_X1 U17737 ( .A1(n14458), .A2(n14462), .ZN(n14483) );
  OAI21_X1 U17738 ( .B1(n10452), .B2(n14481), .A(n14459), .ZN(n14460) );
  OAI21_X1 U17739 ( .B1(n10452), .B2(n14483), .A(n14460), .ZN(n14482) );
  NAND2_X1 U17740 ( .A1(n10452), .A2(n14462), .ZN(n15567) );
  AOI22_X1 U17741 ( .A1(n9679), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n9691), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14468) );
  AOI22_X1 U17742 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14589), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14467) );
  AOI22_X1 U17743 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14466) );
  NAND2_X1 U17744 ( .A1(n14593), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14464) );
  NAND2_X1 U17745 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n14463) );
  AND3_X1 U17746 ( .A1(n14464), .A2(n14596), .A3(n14463), .ZN(n14465) );
  NAND4_X1 U17747 ( .A1(n14468), .A2(n14467), .A3(n14466), .A4(n14465), .ZN(
        n14476) );
  AOI22_X1 U17748 ( .A1(n10416), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14474) );
  NAND2_X1 U17749 ( .A1(n14593), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14470) );
  NAND2_X1 U17750 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n14469) );
  AND3_X1 U17751 ( .A1(n14564), .A2(n14470), .A3(n14469), .ZN(n14473) );
  AOI22_X1 U17752 ( .A1(n14590), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14589), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14472) );
  AOI22_X1 U17753 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14471) );
  NAND4_X1 U17754 ( .A1(n14474), .A2(n14473), .A3(n14472), .A4(n14471), .ZN(
        n14475) );
  NAND2_X1 U17755 ( .A1(n14476), .A2(n14475), .ZN(n14480) );
  XOR2_X1 U17756 ( .A(n14480), .B(n14483), .Z(n14478) );
  INV_X1 U17757 ( .A(n14477), .ZN(n14541) );
  NAND2_X1 U17758 ( .A1(n14478), .A2(n14541), .ZN(n15556) );
  INV_X1 U17759 ( .A(n15556), .ZN(n14479) );
  INV_X1 U17760 ( .A(n14480), .ZN(n14484) );
  NAND2_X1 U17761 ( .A1(n10292), .A2(n14484), .ZN(n15559) );
  INV_X1 U17762 ( .A(n14483), .ZN(n14485) );
  AND2_X1 U17763 ( .A1(n14485), .A2(n14484), .ZN(n14500) );
  AOI22_X1 U17764 ( .A1(n10416), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9691), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14491) );
  NAND2_X1 U17765 ( .A1(n14595), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14487) );
  NAND2_X1 U17766 ( .A1(n14589), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n14486) );
  AND3_X1 U17767 ( .A1(n14564), .A2(n14487), .A3(n14486), .ZN(n14490) );
  AOI22_X1 U17768 ( .A1(n14590), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14489) );
  AOI22_X1 U17769 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14488) );
  NAND4_X1 U17770 ( .A1(n14491), .A2(n14490), .A3(n14489), .A4(n14488), .ZN(
        n14499) );
  AOI22_X1 U17771 ( .A1(n9696), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9692), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14497) );
  AOI22_X1 U17772 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14589), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14496) );
  AOI22_X1 U17773 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14495) );
  NAND2_X1 U17774 ( .A1(n14595), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14493) );
  NAND2_X1 U17775 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n14492) );
  AND3_X1 U17776 ( .A1(n14493), .A2(n14596), .A3(n14492), .ZN(n14494) );
  NAND4_X1 U17777 ( .A1(n14497), .A2(n14496), .A3(n14495), .A4(n14494), .ZN(
        n14498) );
  AND2_X1 U17778 ( .A1(n14499), .A2(n14498), .ZN(n14501) );
  NAND2_X1 U17779 ( .A1(n14500), .A2(n14501), .ZN(n14537) );
  OAI211_X1 U17780 ( .C1(n14500), .C2(n14501), .A(n14541), .B(n14537), .ZN(
        n14504) );
  INV_X1 U17781 ( .A(n14501), .ZN(n14502) );
  NOR2_X1 U17782 ( .A1(n9675), .A2(n14502), .ZN(n15551) );
  NAND2_X1 U17783 ( .A1(n15552), .A2(n15551), .ZN(n15550) );
  INV_X1 U17784 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n19842) );
  NAND2_X1 U17785 ( .A1(n14593), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14507) );
  OAI211_X1 U17786 ( .C1(n14445), .C2(n19842), .A(n14564), .B(n14507), .ZN(
        n14508) );
  INV_X1 U17787 ( .A(n14508), .ZN(n14512) );
  AOI22_X1 U17788 ( .A1(n14590), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14589), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14511) );
  AOI22_X1 U17789 ( .A1(n9679), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9692), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14510) );
  AOI22_X1 U17790 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14509) );
  NAND4_X1 U17791 ( .A1(n14512), .A2(n14511), .A3(n14510), .A4(n14509), .ZN(
        n14520) );
  AOI22_X1 U17792 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n9691), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14518) );
  AOI22_X1 U17793 ( .A1(n9695), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14589), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14517) );
  AOI22_X1 U17794 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14516) );
  NAND2_X1 U17795 ( .A1(n14593), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14514) );
  NAND2_X1 U17796 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n14513) );
  AND3_X1 U17797 ( .A1(n14514), .A2(n14596), .A3(n14513), .ZN(n14515) );
  NAND4_X1 U17798 ( .A1(n14518), .A2(n14517), .A3(n14516), .A4(n14515), .ZN(
        n14519) );
  AND2_X1 U17799 ( .A1(n14520), .A2(n14519), .ZN(n14538) );
  XNOR2_X1 U17800 ( .A(n14537), .B(n14538), .ZN(n14521) );
  NAND2_X1 U17801 ( .A1(n10292), .A2(n14538), .ZN(n15543) );
  AOI22_X1 U17802 ( .A1(n9679), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n9691), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14528) );
  AOI22_X1 U17803 ( .A1(n10278), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14589), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14527) );
  AOI22_X1 U17804 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14526) );
  NAND2_X1 U17805 ( .A1(n14595), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n14524) );
  NAND2_X1 U17806 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n14523) );
  AND3_X1 U17807 ( .A1(n14524), .A2(n14596), .A3(n14523), .ZN(n14525) );
  NAND4_X1 U17808 ( .A1(n14528), .A2(n14527), .A3(n14526), .A4(n14525), .ZN(
        n14536) );
  INV_X1 U17809 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n19808) );
  AOI22_X1 U17810 ( .A1(n10416), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14534) );
  NAND2_X1 U17811 ( .A1(n14595), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14530) );
  NAND2_X1 U17812 ( .A1(n14589), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14529) );
  AND3_X1 U17813 ( .A1(n14564), .A2(n14530), .A3(n14529), .ZN(n14533) );
  INV_X1 U17814 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n21197) );
  AOI22_X1 U17815 ( .A1(n10278), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14532) );
  AOI22_X1 U17816 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14531) );
  NAND4_X1 U17817 ( .A1(n14534), .A2(n14533), .A3(n14532), .A4(n14531), .ZN(
        n14535) );
  NAND2_X1 U17818 ( .A1(n14536), .A2(n14535), .ZN(n14546) );
  INV_X1 U17819 ( .A(n14546), .ZN(n14543) );
  INV_X1 U17820 ( .A(n14537), .ZN(n14539) );
  NAND2_X1 U17821 ( .A1(n14539), .A2(n14538), .ZN(n14540) );
  INV_X1 U17822 ( .A(n14540), .ZN(n14542) );
  OR2_X1 U17823 ( .A1(n14540), .A2(n14546), .ZN(n15531) );
  OAI211_X1 U17824 ( .C1(n14543), .C2(n14542), .A(n14541), .B(n15531), .ZN(
        n14544) );
  AOI21_X1 U17825 ( .B1(n14545), .B2(n14544), .A(n14547), .ZN(n15537) );
  NOR2_X1 U17826 ( .A1(n9675), .A2(n14546), .ZN(n15539) );
  NAND2_X1 U17827 ( .A1(n15537), .A2(n15539), .ZN(n15538) );
  INV_X1 U17828 ( .A(n14547), .ZN(n15532) );
  AOI22_X1 U17829 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9691), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14553) );
  AOI22_X1 U17830 ( .A1(n10278), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14589), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14552) );
  AOI22_X1 U17831 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14551) );
  NAND2_X1 U17832 ( .A1(n14593), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14549) );
  NAND2_X1 U17833 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n14548) );
  AND3_X1 U17834 ( .A1(n14549), .A2(n14596), .A3(n14548), .ZN(n14550) );
  NAND4_X1 U17835 ( .A1(n14553), .A2(n14552), .A3(n14551), .A4(n14550), .ZN(
        n14561) );
  AOI22_X1 U17836 ( .A1(n10416), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14559) );
  NAND2_X1 U17837 ( .A1(n14593), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n14555) );
  NAND2_X1 U17838 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n14554) );
  AND3_X1 U17839 ( .A1(n14564), .A2(n14555), .A3(n14554), .ZN(n14558) );
  AOI22_X1 U17840 ( .A1(n10278), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14589), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14557) );
  AOI22_X1 U17841 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14556) );
  NAND4_X1 U17842 ( .A1(n14559), .A2(n14558), .A3(n14557), .A4(n14556), .ZN(
        n14560) );
  NAND2_X1 U17843 ( .A1(n14561), .A2(n14560), .ZN(n14577) );
  AOI21_X2 U17844 ( .B1(n15538), .B2(n15532), .A(n14577), .ZN(n15527) );
  AOI22_X1 U17845 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9691), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14568) );
  NAND2_X1 U17846 ( .A1(n14595), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14563) );
  NAND2_X1 U17847 ( .A1(n14589), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n14562) );
  AND3_X1 U17848 ( .A1(n14564), .A2(n14563), .A3(n14562), .ZN(n14567) );
  AOI22_X1 U17849 ( .A1(n10278), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14566) );
  AOI22_X1 U17850 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14565) );
  NAND4_X1 U17851 ( .A1(n14568), .A2(n14567), .A3(n14566), .A4(n14565), .ZN(
        n14576) );
  AOI22_X1 U17852 ( .A1(n10278), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9692), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14574) );
  AOI22_X1 U17853 ( .A1(n9679), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14589), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14573) );
  AOI22_X1 U17854 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14572) );
  NAND2_X1 U17855 ( .A1(n14595), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n14570) );
  NAND2_X1 U17856 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n14569) );
  AND3_X1 U17857 ( .A1(n14570), .A2(n14596), .A3(n14569), .ZN(n14571) );
  NAND4_X1 U17858 ( .A1(n14574), .A2(n14573), .A3(n14572), .A4(n14571), .ZN(
        n14575) );
  NAND2_X1 U17859 ( .A1(n14576), .A2(n14575), .ZN(n14580) );
  INV_X1 U17860 ( .A(n14577), .ZN(n15533) );
  NAND2_X1 U17861 ( .A1(n9676), .A2(n15533), .ZN(n14578) );
  OR2_X1 U17862 ( .A1(n15531), .A2(n14578), .ZN(n14579) );
  NOR2_X1 U17863 ( .A1(n14579), .A2(n14580), .ZN(n14581) );
  AOI21_X1 U17864 ( .B1(n14580), .B2(n14579), .A(n14581), .ZN(n15526) );
  INV_X1 U17865 ( .A(n14581), .ZN(n14582) );
  AOI22_X1 U17866 ( .A1(n10278), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14584) );
  AOI22_X1 U17867 ( .A1(n9691), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14589), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14583) );
  NAND2_X1 U17868 ( .A1(n14584), .A2(n14583), .ZN(n14603) );
  AOI21_X1 U17869 ( .B1(n10429), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n14596), .ZN(n14586) );
  AOI22_X1 U17870 ( .A1(n14593), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14585) );
  OAI211_X1 U17871 ( .C1(n14588), .C2(n14587), .A(n14586), .B(n14585), .ZN(
        n14602) );
  AOI22_X1 U17872 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9692), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14592) );
  AOI22_X1 U17873 ( .A1(n10278), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14589), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14591) );
  NAND2_X1 U17874 ( .A1(n14592), .A2(n14591), .ZN(n14601) );
  AOI22_X1 U17875 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14599) );
  NAND2_X1 U17876 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n14598) );
  NAND2_X1 U17877 ( .A1(n14595), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n14597) );
  NAND4_X1 U17878 ( .A1(n14599), .A2(n14598), .A3(n14597), .A4(n14596), .ZN(
        n14600) );
  OAI22_X1 U17879 ( .A1(n14603), .A2(n14602), .B1(n14601), .B2(n14600), .ZN(
        n14604) );
  NOR2_X1 U17880 ( .A1(n15888), .A2(n15592), .ZN(n14605) );
  AOI21_X1 U17881 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15592), .A(n14605), .ZN(
        n14606) );
  NOR2_X1 U17882 ( .A1(n15443), .A2(n14607), .ZN(n14608) );
  OAI21_X1 U17883 ( .B1(n19508), .B2(n16447), .A(n14610), .ZN(n14611) );
  INV_X1 U17884 ( .A(n14611), .ZN(n14619) );
  NOR2_X1 U17885 ( .A1(n15883), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14615) );
  NAND2_X1 U17886 ( .A1(n15893), .A2(n15894), .ZN(n15912) );
  NAND2_X1 U17887 ( .A1(n15912), .A2(n15907), .ZN(n15902) );
  AOI21_X1 U17888 ( .B1(n15893), .B2(n14612), .A(n15902), .ZN(n14613) );
  NOR2_X1 U17889 ( .A1(n14615), .A2(n14614), .ZN(n14618) );
  INV_X1 U17890 ( .A(n16441), .ZN(n14616) );
  NAND3_X1 U17891 ( .A1(n14619), .A2(n14618), .A3(n14617), .ZN(n14620) );
  AOI21_X1 U17892 ( .B1(n14621), .B2(n16550), .A(n14620), .ZN(n14622) );
  OAI21_X1 U17893 ( .B1(n14623), .B2(n19502), .A(n14622), .ZN(P2_U3017) );
  NOR2_X2 U17894 ( .A1(n14624), .A2(n19519), .ZN(n19340) );
  NOR2_X2 U17895 ( .A1(n14624), .A2(n19517), .ZN(n19339) );
  AOI22_X1 U17896 ( .A1(n19340), .A2(BUF2_REG_30__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n14626) );
  AOI22_X1 U17897 ( .A1(n19338), .A2(n19350), .B1(n19399), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14625) );
  OAI211_X1 U17898 ( .C1(n15880), .C2(n19342), .A(n14626), .B(n14625), .ZN(
        n14627) );
  INV_X1 U17899 ( .A(n14627), .ZN(n14628) );
  OAI21_X1 U17900 ( .B1(n14629), .B2(n16479), .A(n14628), .ZN(P2_U2889) );
  OAI21_X1 U17901 ( .B1(n14632), .B2(n14631), .A(n14630), .ZN(n14645) );
  OAI22_X1 U17902 ( .A1(n14633), .A2(n19501), .B1(n19515), .B2(n14645), .ZN(
        n14637) );
  NAND2_X1 U17903 ( .A1(n14635), .A2(n14634), .ZN(n14651) );
  AND3_X1 U17904 ( .A1(n16568), .A2(n14652), .A3(n14651), .ZN(n14636) );
  AOI211_X1 U17905 ( .C1(n16544), .C2(n20188), .A(n14637), .B(n14636), .ZN(
        n14644) );
  NOR2_X1 U17906 ( .A1(n14639), .A2(n14638), .ZN(n14640) );
  INV_X1 U17907 ( .A(n14640), .ZN(n14642) );
  AND2_X1 U17908 ( .A1(n19303), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14646) );
  AND2_X1 U17909 ( .A1(n16046), .A2(n14640), .ZN(n14641) );
  AOI211_X1 U17910 ( .C1(n16045), .C2(n14642), .A(n14646), .B(n14641), .ZN(
        n14643) );
  OAI211_X1 U17911 ( .C1(n14655), .C2(n16547), .A(n14644), .B(n14643), .ZN(
        P2_U3044) );
  INV_X1 U17912 ( .A(n14645), .ZN(n14650) );
  AOI21_X1 U17913 ( .B1(n19484), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14646), .ZN(n14647) );
  OAI21_X1 U17914 ( .B1(n19496), .B2(n14648), .A(n14647), .ZN(n14649) );
  AOI21_X1 U17915 ( .B1(n16529), .B2(n14650), .A(n14649), .ZN(n14654) );
  NAND3_X1 U17916 ( .A1(n14652), .A2(n10990), .A3(n14651), .ZN(n14653) );
  OAI211_X1 U17917 ( .C1(n16526), .C2(n14655), .A(n14654), .B(n14653), .ZN(
        P2_U3012) );
  NAND2_X1 U17918 ( .A1(n19484), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14656) );
  OAI211_X1 U17919 ( .C1(n14658), .C2(n19496), .A(n14657), .B(n14656), .ZN(
        n14659) );
  INV_X1 U17920 ( .A(n14659), .ZN(n14660) );
  OAI21_X1 U17921 ( .B1(n14665), .B2(n16537), .A(n14664), .ZN(P2_U2983) );
  AND2_X1 U17922 ( .A1(n14690), .A2(n14678), .ZN(n14667) );
  OAI21_X1 U17923 ( .B1(n14667), .B2(n14666), .A(n9730), .ZN(n15250) );
  NAND2_X1 U17924 ( .A1(n15060), .A2(n20317), .ZN(n14677) );
  OAI22_X1 U17925 ( .A1(n14670), .A2(n20279), .B1(n20330), .B2(n15058), .ZN(
        n14675) );
  INV_X1 U17926 ( .A(n14671), .ZN(n14673) );
  INV_X1 U17927 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n15056) );
  AOI21_X1 U17928 ( .B1(n14673), .B2(n15056), .A(n14672), .ZN(n14674) );
  AOI211_X1 U17929 ( .C1(n20335), .C2(P1_EBX_REG_28__SCAN_IN), .A(n14675), .B(
        n14674), .ZN(n14676) );
  OAI211_X1 U17930 ( .C1(n20325), .C2(n15250), .A(n14677), .B(n14676), .ZN(
        P1_U2812) );
  XNOR2_X1 U17931 ( .A(n14690), .B(n14678), .ZN(n15265) );
  OAI21_X1 U17932 ( .B1(n14679), .B2(n14680), .A(n14668), .ZN(n14861) );
  INV_X1 U17933 ( .A(n14861), .ZN(n15069) );
  NAND2_X1 U17934 ( .A1(n15069), .A2(n20317), .ZN(n14687) );
  INV_X1 U17935 ( .A(n14696), .ZN(n14685) );
  INV_X1 U17936 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14860) );
  AOI22_X1 U17937 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n15065), .ZN(n14681) );
  OAI21_X1 U17938 ( .B1(n20308), .B2(n14860), .A(n14681), .ZN(n14684) );
  NOR3_X1 U17939 ( .A1(n14817), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14682), 
        .ZN(n14683) );
  AOI211_X1 U17940 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14685), .A(n14684), 
        .B(n14683), .ZN(n14686) );
  OAI211_X1 U17941 ( .C1(n15265), .C2(n20325), .A(n14687), .B(n14686), .ZN(
        P1_U2813) );
  NOR2_X1 U17942 ( .A1(n14703), .A2(n14688), .ZN(n14689) );
  OR2_X1 U17943 ( .A1(n14690), .A2(n14689), .ZN(n15277) );
  AOI21_X1 U17944 ( .B1(n14692), .B2(n14691), .A(n14679), .ZN(n15078) );
  NAND2_X1 U17945 ( .A1(n15078), .A2(n20317), .ZN(n14700) );
  OAI22_X1 U17946 ( .A1(n14693), .A2(n20279), .B1(n20330), .B2(n15076), .ZN(
        n14698) );
  AOI21_X1 U17947 ( .B1(n20333), .B2(n14694), .A(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14695) );
  NOR2_X1 U17948 ( .A1(n14696), .A2(n14695), .ZN(n14697) );
  AOI211_X1 U17949 ( .C1(n20335), .C2(P1_EBX_REG_26__SCAN_IN), .A(n14698), .B(
        n14697), .ZN(n14699) );
  OAI211_X1 U17950 ( .C1(n20325), .C2(n15277), .A(n14700), .B(n14699), .ZN(
        P1_U2814) );
  OAI21_X1 U17951 ( .B1(n14701), .B2(n14702), .A(n14691), .ZN(n14916) );
  AOI21_X1 U17952 ( .B1(n14704), .B2(n14720), .A(n14703), .ZN(n15283) );
  INV_X1 U17953 ( .A(n14705), .ZN(n14722) );
  AOI21_X1 U17954 ( .B1(n20333), .B2(n14722), .A(n20332), .ZN(n14736) );
  INV_X1 U17955 ( .A(n14706), .ZN(n15087) );
  OAI22_X1 U17956 ( .A1(n14707), .A2(n20279), .B1(n20330), .B2(n15087), .ZN(
        n14712) );
  INV_X1 U17957 ( .A(n14708), .ZN(n14709) );
  NOR2_X1 U17958 ( .A1(n14709), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14710) );
  AOI211_X1 U17959 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(P1_REIP_REG_25__SCAN_IN), .A(n14710), .B(n14817), .ZN(n14711) );
  AOI211_X1 U17960 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n20335), .A(n14712), .B(
        n14711), .ZN(n14713) );
  OAI21_X1 U17961 ( .B1(n14736), .B2(n15085), .A(n14713), .ZN(n14714) );
  AOI21_X1 U17962 ( .B1(n15283), .B2(n20334), .A(n14714), .ZN(n14715) );
  OAI21_X1 U17963 ( .B1(n14916), .B2(n20287), .A(n14715), .ZN(P1_U2815) );
  AOI21_X1 U17964 ( .B1(n14717), .B2(n14716), .A(n14701), .ZN(n15098) );
  INV_X1 U17965 ( .A(n15098), .ZN(n14867) );
  NAND2_X1 U17966 ( .A1(n14728), .A2(n14718), .ZN(n14719) );
  NAND2_X1 U17967 ( .A1(n14720), .A2(n14719), .ZN(n14865) );
  INV_X1 U17968 ( .A(n14865), .ZN(n15291) );
  INV_X1 U17969 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n15094) );
  OAI22_X1 U17970 ( .A1(n14721), .A2(n20279), .B1(n20330), .B2(n15096), .ZN(
        n14724) );
  NOR3_X1 U17971 ( .A1(n14817), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n14722), 
        .ZN(n14723) );
  AOI211_X1 U17972 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n20335), .A(n14724), .B(
        n14723), .ZN(n14725) );
  OAI21_X1 U17973 ( .B1(n14736), .B2(n15094), .A(n14725), .ZN(n14726) );
  AOI21_X1 U17974 ( .B1(n15291), .B2(n20334), .A(n14726), .ZN(n14727) );
  OAI21_X1 U17975 ( .B1(n14867), .B2(n20287), .A(n14727), .ZN(P1_U2816) );
  OAI21_X1 U17976 ( .B1(n14745), .B2(n14729), .A(n14728), .ZN(n15297) );
  OAI21_X1 U17977 ( .B1(n9725), .B2(n14730), .A(n14716), .ZN(n14869) );
  INV_X1 U17978 ( .A(n14869), .ZN(n15105) );
  NAND2_X1 U17979 ( .A1(n15105), .A2(n20317), .ZN(n14741) );
  OAI22_X1 U17980 ( .A1(n14731), .A2(n20279), .B1(n20330), .B2(n15103), .ZN(
        n14739) );
  INV_X1 U17981 ( .A(n14815), .ZN(n14816) );
  AND2_X1 U17982 ( .A1(n20333), .A2(n14816), .ZN(n14818) );
  INV_X1 U17983 ( .A(n14732), .ZN(n14733) );
  AND2_X1 U17984 ( .A1(n14818), .A2(n14733), .ZN(n14807) );
  AND2_X1 U17985 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14734) );
  AND2_X1 U17986 ( .A1(n14807), .A2(n14734), .ZN(n14778) );
  AOI21_X1 U17987 ( .B1(n14778), .B2(n14735), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14737) );
  NOR2_X1 U17988 ( .A1(n14737), .A2(n14736), .ZN(n14738) );
  AOI211_X1 U17989 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n20335), .A(n14739), .B(
        n14738), .ZN(n14740) );
  OAI211_X1 U17990 ( .C1(n20325), .C2(n15297), .A(n14741), .B(n14740), .ZN(
        P1_U2817) );
  AOI21_X1 U17991 ( .B1(n14743), .B2(n14742), .A(n9725), .ZN(n15115) );
  AND2_X1 U17992 ( .A1(n14761), .A2(n14744), .ZN(n14746) );
  OR2_X1 U17993 ( .A1(n14746), .A2(n14745), .ZN(n15306) );
  INV_X1 U17994 ( .A(n14763), .ZN(n14747) );
  NAND3_X1 U17995 ( .A1(n20261), .A2(P1_REIP_REG_20__SCAN_IN), .A3(n14747), 
        .ZN(n14748) );
  NAND2_X1 U17996 ( .A1(n20292), .A2(n14748), .ZN(n14776) );
  OAI21_X1 U17997 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n14817), .A(n14776), 
        .ZN(n14751) );
  INV_X1 U17998 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14870) );
  AOI22_X1 U17999 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n15110), .ZN(n14749) );
  OAI21_X1 U18000 ( .B1(n20308), .B2(n14870), .A(n14749), .ZN(n14750) );
  AOI21_X1 U18001 ( .B1(n14751), .B2(P1_REIP_REG_22__SCAN_IN), .A(n14750), 
        .ZN(n14754) );
  INV_X1 U18002 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n15111) );
  NAND3_X1 U18003 ( .A1(n14778), .A2(n15111), .A3(n14752), .ZN(n14753) );
  OAI211_X1 U18004 ( .C1(n15306), .C2(n20325), .A(n14754), .B(n14753), .ZN(
        n14755) );
  AOI21_X1 U18005 ( .B1(n15115), .B2(n20317), .A(n14755), .ZN(n14756) );
  INV_X1 U18006 ( .A(n14756), .ZN(P1_U2818) );
  OAI21_X1 U18007 ( .B1(n14757), .B2(n14758), .A(n14742), .ZN(n15125) );
  NAND2_X1 U18008 ( .A1(n14774), .A2(n14759), .ZN(n14760) );
  AND2_X1 U18009 ( .A1(n14761), .A2(n14760), .ZN(n15330) );
  INV_X1 U18010 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15120) );
  OAI22_X1 U18011 ( .A1(n14762), .A2(n20279), .B1(n20330), .B2(n15121), .ZN(
        n14765) );
  INV_X1 U18012 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21012) );
  NOR4_X1 U18013 ( .A1(n14817), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n14763), 
        .A4(n21012), .ZN(n14764) );
  AOI211_X1 U18014 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n20335), .A(n14765), .B(
        n14764), .ZN(n14766) );
  OAI21_X1 U18015 ( .B1(n15120), .B2(n14776), .A(n14766), .ZN(n14767) );
  AOI21_X1 U18016 ( .B1(n15330), .B2(n20334), .A(n14767), .ZN(n14768) );
  OAI21_X1 U18017 ( .B1(n15125), .B2(n20287), .A(n14768), .ZN(P1_U2819) );
  INV_X1 U18018 ( .A(n14769), .ZN(n14773) );
  BUF_X1 U18019 ( .A(n14770), .Z(n14771) );
  INV_X1 U18020 ( .A(n14771), .ZN(n14772) );
  AOI21_X1 U18021 ( .B1(n14773), .B2(n14772), .A(n14757), .ZN(n15131) );
  INV_X1 U18022 ( .A(n15131), .ZN(n14945) );
  OAI21_X1 U18023 ( .B1(n14788), .B2(n14775), .A(n14774), .ZN(n14873) );
  INV_X1 U18024 ( .A(n14873), .ZN(n15336) );
  INV_X1 U18025 ( .A(n14776), .ZN(n14777) );
  OAI21_X1 U18026 ( .B1(n14778), .B2(P1_REIP_REG_20__SCAN_IN), .A(n14777), 
        .ZN(n14780) );
  AOI22_X1 U18027 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n15130), .ZN(n14779) );
  OAI211_X1 U18028 ( .C1(n14874), .C2(n20308), .A(n14780), .B(n14779), .ZN(
        n14781) );
  AOI21_X1 U18029 ( .B1(n15336), .B2(n20334), .A(n14781), .ZN(n14782) );
  OAI21_X1 U18030 ( .B1(n14945), .B2(n20287), .A(n14782), .ZN(P1_U2820) );
  AOI21_X1 U18031 ( .B1(n14783), .B2(n9741), .A(n14771), .ZN(n15140) );
  INV_X1 U18032 ( .A(n15140), .ZN(n14949) );
  OAI21_X1 U18033 ( .B1(n14784), .B2(n14817), .A(n20261), .ZN(n16276) );
  NAND2_X1 U18034 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14785) );
  OAI211_X1 U18035 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(P1_REIP_REG_18__SCAN_IN), .A(n14807), .B(n14785), .ZN(n14786) );
  OAI211_X1 U18036 ( .C1(n20279), .C2(n11673), .A(n14786), .B(n20322), .ZN(
        n14787) );
  AOI21_X1 U18037 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n16276), .A(n14787), 
        .ZN(n14794) );
  AOI21_X1 U18038 ( .B1(n14789), .B2(n14801), .A(n14788), .ZN(n15346) );
  INV_X1 U18039 ( .A(n14790), .ZN(n15138) );
  OAI22_X1 U18040 ( .A1(n20308), .A2(n14791), .B1(n20330), .B2(n15138), .ZN(
        n14792) );
  AOI21_X1 U18041 ( .B1(n15346), .B2(n20334), .A(n14792), .ZN(n14793) );
  OAI211_X1 U18042 ( .C1(n14949), .C2(n20287), .A(n14794), .B(n14793), .ZN(
        P1_U2821) );
  INV_X1 U18043 ( .A(n14795), .ZN(n14798) );
  INV_X1 U18044 ( .A(n14796), .ZN(n14797) );
  OAI21_X1 U18045 ( .B1(n14798), .B2(n14797), .A(n9741), .ZN(n14950) );
  OAI21_X1 U18046 ( .B1(n14799), .B2(n15365), .A(n14800), .ZN(n14802) );
  NAND2_X1 U18047 ( .A1(n14802), .A2(n14801), .ZN(n15355) );
  INV_X1 U18048 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21009) );
  INV_X1 U18049 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14805) );
  INV_X1 U18050 ( .A(n20322), .ZN(n20310) );
  NOR2_X1 U18051 ( .A1(n20330), .A2(n15145), .ZN(n14803) );
  AOI211_X1 U18052 ( .C1(n20340), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20310), .B(n14803), .ZN(n14804) );
  OAI21_X1 U18053 ( .B1(n14805), .B2(n20308), .A(n14804), .ZN(n14806) );
  AOI21_X1 U18054 ( .B1(n14807), .B2(n21009), .A(n14806), .ZN(n14808) );
  OAI21_X1 U18055 ( .B1(n15355), .B2(n20325), .A(n14808), .ZN(n14809) );
  AOI21_X1 U18056 ( .B1(n16276), .B2(P1_REIP_REG_18__SCAN_IN), .A(n14809), 
        .ZN(n14810) );
  OAI21_X1 U18057 ( .B1(n14950), .B2(n20287), .A(n14810), .ZN(P1_U2822) );
  AOI21_X1 U18058 ( .B1(n14813), .B2(n14811), .A(n14812), .ZN(n14814) );
  INV_X1 U18059 ( .A(n14814), .ZN(n15172) );
  INV_X1 U18060 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21003) );
  NOR3_X1 U18061 ( .A1(n14817), .A2(n14815), .A3(n21003), .ZN(n16275) );
  INV_X1 U18062 ( .A(n16275), .ZN(n14821) );
  OAI21_X1 U18063 ( .B1(n14817), .B2(n14816), .A(n20261), .ZN(n16284) );
  INV_X1 U18064 ( .A(n14818), .ZN(n14819) );
  NOR2_X1 U18065 ( .A1(n14819), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n16286) );
  NOR2_X1 U18066 ( .A1(n16284), .A2(n16286), .ZN(n14820) );
  MUX2_X1 U18067 ( .A(n14821), .B(n14820), .S(P1_REIP_REG_16__SCAN_IN), .Z(
        n14828) );
  NAND2_X1 U18068 ( .A1(n20339), .A2(n15169), .ZN(n14822) );
  OAI211_X1 U18069 ( .C1(n20279), .C2(n15167), .A(n20322), .B(n14822), .ZN(
        n14826) );
  OR2_X1 U18070 ( .A1(n14881), .A2(n14823), .ZN(n14824) );
  NAND2_X1 U18071 ( .A1(n14799), .A2(n14824), .ZN(n15381) );
  NOR2_X1 U18072 ( .A1(n15381), .A2(n20325), .ZN(n14825) );
  AOI211_X1 U18073 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n20335), .A(n14826), .B(
        n14825), .ZN(n14827) );
  OAI211_X1 U18074 ( .C1(n15172), .C2(n20287), .A(n14828), .B(n14827), .ZN(
        P1_U2824) );
  NAND2_X1 U18075 ( .A1(n14830), .A2(n14831), .ZN(n14832) );
  NAND2_X1 U18076 ( .A1(n9668), .A2(n14832), .ZN(n15183) );
  NOR2_X1 U18077 ( .A1(n14833), .A2(n20270), .ZN(n16303) );
  OAI221_X1 U18078 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n14834), .C1(
        P1_REIP_REG_14__SCAN_IN), .C2(n16303), .A(n16284), .ZN(n14841) );
  INV_X1 U18079 ( .A(n14835), .ZN(n15180) );
  AND2_X1 U18080 ( .A1(n14851), .A2(n14836), .ZN(n14837) );
  NOR2_X1 U18081 ( .A1(n14879), .A2(n14837), .ZN(n16356) );
  AOI22_X1 U18082 ( .A1(n16356), .A2(n20334), .B1(n20335), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14838) );
  OAI211_X1 U18083 ( .C1(n20279), .C2(n21218), .A(n14838), .B(n20322), .ZN(
        n14839) );
  AOI21_X1 U18084 ( .B1(n20339), .B2(n15180), .A(n14839), .ZN(n14840) );
  OAI211_X1 U18085 ( .C1(n15183), .C2(n20287), .A(n14841), .B(n14840), .ZN(
        P1_U2826) );
  OAI21_X1 U18086 ( .B1(n14027), .B2(n14843), .A(n14844), .ZN(n14892) );
  INV_X1 U18087 ( .A(n14891), .ZN(n14845) );
  OAI21_X1 U18088 ( .B1(n14892), .B2(n14845), .A(n14844), .ZN(n14980) );
  OAI21_X1 U18089 ( .B1(n14982), .B2(n14846), .A(n14830), .ZN(n15196) );
  OAI21_X1 U18090 ( .B1(n14853), .B2(n14847), .A(n20292), .ZN(n16297) );
  AOI22_X1 U18091 ( .A1(n20335), .A2(P1_EBX_REG_13__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n20340), .ZN(n14848) );
  OAI211_X1 U18092 ( .C1(n21001), .C2(n16297), .A(n14848), .B(n20322), .ZN(
        n14855) );
  NAND2_X1 U18093 ( .A1(n15399), .A2(n14849), .ZN(n14850) );
  NAND2_X1 U18094 ( .A1(n14851), .A2(n14850), .ZN(n16371) );
  NAND2_X1 U18095 ( .A1(n16303), .A2(n21001), .ZN(n14852) );
  OAI22_X1 U18096 ( .A1(n20325), .A2(n16371), .B1(n14853), .B2(n14852), .ZN(
        n14854) );
  AOI211_X1 U18097 ( .C1(n15193), .C2(n20339), .A(n14855), .B(n14854), .ZN(
        n14856) );
  OAI21_X1 U18098 ( .B1(n15196), .B2(n20287), .A(n14856), .ZN(P1_U2827) );
  OAI22_X1 U18099 ( .A1(n15231), .A2(n14896), .B1(n20356), .B2(n14857), .ZN(
        P1_U2841) );
  OAI222_X1 U18100 ( .A1(n14890), .A2(n15040), .B1(n21239), .B2(n20356), .C1(
        n15242), .C2(n14896), .ZN(P1_U2842) );
  INV_X1 U18101 ( .A(n15060), .ZN(n14859) );
  INV_X1 U18102 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14858) );
  OAI222_X1 U18103 ( .A1(n14890), .A2(n14859), .B1(n14858), .B2(n20356), .C1(
        n15250), .C2(n14896), .ZN(P1_U2844) );
  OAI222_X1 U18104 ( .A1(n14861), .A2(n14890), .B1(n14860), .B2(n20356), .C1(
        n14896), .C2(n15265), .ZN(P1_U2845) );
  INV_X1 U18105 ( .A(n15078), .ZN(n14863) );
  INV_X1 U18106 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14862) );
  OAI222_X1 U18107 ( .A1(n14890), .A2(n14863), .B1(n14862), .B2(n20356), .C1(
        n15277), .C2(n14896), .ZN(P1_U2846) );
  AOI22_X1 U18108 ( .A1(n15283), .A2(n20351), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n14885), .ZN(n14864) );
  OAI21_X1 U18109 ( .B1(n14916), .B2(n14890), .A(n14864), .ZN(P1_U2847) );
  INV_X1 U18110 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14866) );
  OAI222_X1 U18111 ( .A1(n14890), .A2(n14867), .B1(n14866), .B2(n20356), .C1(
        n14865), .C2(n14896), .ZN(P1_U2848) );
  INV_X1 U18112 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14868) );
  OAI222_X1 U18113 ( .A1(n14890), .A2(n14869), .B1(n14868), .B2(n20356), .C1(
        n15297), .C2(n14896), .ZN(P1_U2849) );
  INV_X1 U18114 ( .A(n15115), .ZN(n14871) );
  OAI222_X1 U18115 ( .A1(n14890), .A2(n14871), .B1(n14870), .B2(n20356), .C1(
        n15306), .C2(n14896), .ZN(P1_U2850) );
  AOI22_X1 U18116 ( .A1(n15330), .A2(n20351), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14885), .ZN(n14872) );
  OAI21_X1 U18117 ( .B1(n15125), .B2(n14890), .A(n14872), .ZN(P1_U2851) );
  OAI222_X1 U18118 ( .A1(n14945), .A2(n14890), .B1(n14874), .B2(n20356), .C1(
        n14873), .C2(n14896), .ZN(P1_U2852) );
  AOI22_X1 U18119 ( .A1(n15346), .A2(n20351), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14885), .ZN(n14875) );
  OAI21_X1 U18120 ( .B1(n14949), .B2(n14890), .A(n14875), .ZN(P1_U2853) );
  OAI222_X1 U18121 ( .A1(n14950), .A2(n14890), .B1(n14805), .B2(n20356), .C1(
        n15355), .C2(n14896), .ZN(P1_U2854) );
  INV_X1 U18122 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14876) );
  OAI222_X1 U18123 ( .A1(n15172), .A2(n14890), .B1(n14876), .B2(n20356), .C1(
        n15381), .C2(n14896), .ZN(P1_U2856) );
  AOI21_X1 U18124 ( .B1(n14877), .B2(n9668), .A(n10024), .ZN(n16316) );
  INV_X1 U18125 ( .A(n14890), .ZN(n20352) );
  NOR2_X1 U18126 ( .A1(n14879), .A2(n14878), .ZN(n14880) );
  OR2_X1 U18127 ( .A1(n14881), .A2(n14880), .ZN(n16348) );
  INV_X1 U18128 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14882) );
  OAI22_X1 U18129 ( .A1(n16348), .A2(n14896), .B1(n14882), .B2(n20356), .ZN(
        n14883) );
  AOI21_X1 U18130 ( .B1(n16316), .B2(n20352), .A(n14883), .ZN(n14884) );
  INV_X1 U18131 ( .A(n14884), .ZN(P1_U2857) );
  AOI22_X1 U18132 ( .A1(n16356), .A2(n20351), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14885), .ZN(n14886) );
  OAI21_X1 U18133 ( .B1(n15183), .B2(n14890), .A(n14886), .ZN(P1_U2858) );
  OAI22_X1 U18134 ( .A1(n16371), .A2(n14896), .B1(n14887), .B2(n20356), .ZN(
        n14888) );
  INV_X1 U18135 ( .A(n14888), .ZN(n14889) );
  OAI21_X1 U18136 ( .B1(n15196), .B2(n14890), .A(n14889), .ZN(P1_U2859) );
  XNOR2_X1 U18137 ( .A(n14892), .B(n14891), .ZN(n16328) );
  NOR2_X1 U18138 ( .A1(n10175), .A2(n14893), .ZN(n14894) );
  OR2_X1 U18139 ( .A1(n15401), .A2(n14894), .ZN(n16379) );
  INV_X1 U18140 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14895) );
  OAI22_X1 U18141 ( .A1(n16379), .A2(n14896), .B1(n14895), .B2(n20356), .ZN(
        n14897) );
  AOI21_X1 U18142 ( .B1(n16328), .B2(n20352), .A(n14897), .ZN(n14898) );
  INV_X1 U18143 ( .A(n14898), .ZN(P1_U2861) );
  INV_X1 U18144 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14900) );
  AOI22_X1 U18145 ( .A1(n14959), .A2(n14976), .B1(n14991), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n14899) );
  OAI21_X1 U18146 ( .B1(n14900), .B2(n14962), .A(n14899), .ZN(n14901) );
  AOI21_X1 U18147 ( .B1(n14970), .B2(DATAI_30_), .A(n14901), .ZN(n14902) );
  OAI21_X1 U18148 ( .B1(n15040), .B2(n14995), .A(n14902), .ZN(P1_U2874) );
  NAND2_X1 U18149 ( .A1(n15060), .A2(n14964), .ZN(n14906) );
  AOI22_X1 U18150 ( .A1(n14959), .A2(n14985), .B1(n14991), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n14905) );
  NAND2_X1 U18151 ( .A1(n14970), .A2(DATAI_28_), .ZN(n14904) );
  NAND2_X1 U18152 ( .A1(n14969), .A2(BUF1_REG_28__SCAN_IN), .ZN(n14903) );
  NAND4_X1 U18153 ( .A1(n14906), .A2(n14905), .A3(n14904), .A4(n14903), .ZN(
        P1_U2876) );
  NAND2_X1 U18154 ( .A1(n15069), .A2(n14964), .ZN(n14910) );
  AOI22_X1 U18155 ( .A1(n14959), .A2(n14992), .B1(n14991), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n14909) );
  NAND2_X1 U18156 ( .A1(n14970), .A2(DATAI_27_), .ZN(n14908) );
  NAND2_X1 U18157 ( .A1(n14969), .A2(BUF1_REG_27__SCAN_IN), .ZN(n14907) );
  NAND4_X1 U18158 ( .A1(n14910), .A2(n14909), .A3(n14908), .A4(n14907), .ZN(
        P1_U2877) );
  NAND2_X1 U18159 ( .A1(n15078), .A2(n14964), .ZN(n14915) );
  AOI22_X1 U18160 ( .A1(n14959), .A2(n14911), .B1(n14991), .B2(
        P1_EAX_REG_26__SCAN_IN), .ZN(n14914) );
  NAND2_X1 U18161 ( .A1(n14970), .A2(DATAI_26_), .ZN(n14913) );
  NAND2_X1 U18162 ( .A1(n14969), .A2(BUF1_REG_26__SCAN_IN), .ZN(n14912) );
  NAND4_X1 U18163 ( .A1(n14915), .A2(n14914), .A3(n14913), .A4(n14912), .ZN(
        P1_U2878) );
  INV_X1 U18164 ( .A(n14916), .ZN(n15089) );
  NAND2_X1 U18165 ( .A1(n15089), .A2(n14964), .ZN(n14921) );
  AOI22_X1 U18166 ( .A1(n14959), .A2(n14917), .B1(n14991), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n14920) );
  NAND2_X1 U18167 ( .A1(n14970), .A2(DATAI_25_), .ZN(n14919) );
  NAND2_X1 U18168 ( .A1(n14969), .A2(BUF1_REG_25__SCAN_IN), .ZN(n14918) );
  NAND4_X1 U18169 ( .A1(n14921), .A2(n14920), .A3(n14919), .A4(n14918), .ZN(
        P1_U2879) );
  NAND2_X1 U18170 ( .A1(n15098), .A2(n14964), .ZN(n14926) );
  AOI22_X1 U18171 ( .A1(n14959), .A2(n14922), .B1(n14991), .B2(
        P1_EAX_REG_24__SCAN_IN), .ZN(n14925) );
  NAND2_X1 U18172 ( .A1(n14970), .A2(DATAI_24_), .ZN(n14924) );
  NAND2_X1 U18173 ( .A1(n14969), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14923) );
  NAND4_X1 U18174 ( .A1(n14926), .A2(n14925), .A3(n14924), .A4(n14923), .ZN(
        P1_U2880) );
  NAND2_X1 U18175 ( .A1(n15105), .A2(n14964), .ZN(n14931) );
  AOI22_X1 U18176 ( .A1(n14959), .A2(n14927), .B1(n14991), .B2(
        P1_EAX_REG_23__SCAN_IN), .ZN(n14930) );
  NAND2_X1 U18177 ( .A1(n14970), .A2(DATAI_23_), .ZN(n14929) );
  NAND2_X1 U18178 ( .A1(n14969), .A2(BUF1_REG_23__SCAN_IN), .ZN(n14928) );
  NAND4_X1 U18179 ( .A1(n14931), .A2(n14930), .A3(n14929), .A4(n14928), .ZN(
        P1_U2881) );
  NAND2_X1 U18180 ( .A1(n15115), .A2(n14964), .ZN(n14936) );
  AOI22_X1 U18181 ( .A1(n14959), .A2(n14932), .B1(n14991), .B2(
        P1_EAX_REG_22__SCAN_IN), .ZN(n14935) );
  NAND2_X1 U18182 ( .A1(n14970), .A2(DATAI_22_), .ZN(n14934) );
  NAND2_X1 U18183 ( .A1(n14969), .A2(BUF1_REG_22__SCAN_IN), .ZN(n14933) );
  NAND4_X1 U18184 ( .A1(n14936), .A2(n14935), .A3(n14934), .A4(n14933), .ZN(
        P1_U2882) );
  INV_X1 U18185 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16717) );
  AOI22_X1 U18186 ( .A1(n14959), .A2(n14937), .B1(n14991), .B2(
        P1_EAX_REG_21__SCAN_IN), .ZN(n14939) );
  NAND2_X1 U18187 ( .A1(n14970), .A2(DATAI_21_), .ZN(n14938) );
  OAI211_X1 U18188 ( .C1(n14962), .C2(n16717), .A(n14939), .B(n14938), .ZN(
        n14940) );
  INV_X1 U18189 ( .A(n14940), .ZN(n14941) );
  OAI21_X1 U18190 ( .B1(n15125), .B2(n14995), .A(n14941), .ZN(P1_U2883) );
  INV_X1 U18191 ( .A(n14959), .ZN(n14967) );
  OAI22_X1 U18192 ( .A1(n14967), .A2(n20447), .B1(n14988), .B2(n13757), .ZN(
        n14942) );
  AOI21_X1 U18193 ( .B1(n14969), .B2(BUF1_REG_20__SCAN_IN), .A(n14942), .ZN(
        n14944) );
  NAND2_X1 U18194 ( .A1(n14970), .A2(DATAI_20_), .ZN(n14943) );
  OAI211_X1 U18195 ( .C1(n14945), .C2(n14995), .A(n14944), .B(n14943), .ZN(
        P1_U2884) );
  OAI22_X1 U18196 ( .A1(n14967), .A2(n20443), .B1(n14988), .B2(n13743), .ZN(
        n14946) );
  AOI21_X1 U18197 ( .B1(n14969), .B2(BUF1_REG_19__SCAN_IN), .A(n14946), .ZN(
        n14948) );
  NAND2_X1 U18198 ( .A1(n14970), .A2(DATAI_19_), .ZN(n14947) );
  OAI211_X1 U18199 ( .C1(n14949), .C2(n14995), .A(n14948), .B(n14947), .ZN(
        P1_U2885) );
  INV_X1 U18200 ( .A(n14950), .ZN(n15147) );
  NAND2_X1 U18201 ( .A1(n15147), .A2(n14964), .ZN(n14955) );
  AOI22_X1 U18202 ( .A1(n14959), .A2(n14951), .B1(n14991), .B2(
        P1_EAX_REG_18__SCAN_IN), .ZN(n14954) );
  NAND2_X1 U18203 ( .A1(n14970), .A2(DATAI_18_), .ZN(n14953) );
  NAND2_X1 U18204 ( .A1(n14969), .A2(BUF1_REG_18__SCAN_IN), .ZN(n14952) );
  NAND4_X1 U18205 ( .A1(n14955), .A2(n14954), .A3(n14953), .A4(n14952), .ZN(
        P1_U2886) );
  OR2_X1 U18206 ( .A1(n14812), .A2(n14956), .ZN(n14957) );
  AND2_X1 U18207 ( .A1(n14795), .A2(n14957), .ZN(n16307) );
  INV_X1 U18208 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16724) );
  AOI22_X1 U18209 ( .A1(n14959), .A2(n14958), .B1(n14991), .B2(
        P1_EAX_REG_17__SCAN_IN), .ZN(n14961) );
  NAND2_X1 U18210 ( .A1(n14970), .A2(DATAI_17_), .ZN(n14960) );
  OAI211_X1 U18211 ( .C1(n16724), .C2(n14962), .A(n14961), .B(n14960), .ZN(
        n14963) );
  AOI21_X1 U18212 ( .B1(n16307), .B2(n14964), .A(n14963), .ZN(n14965) );
  INV_X1 U18213 ( .A(n14965), .ZN(P1_U2887) );
  OAI22_X1 U18214 ( .A1(n14967), .A2(n20428), .B1(n14988), .B2(n14966), .ZN(
        n14968) );
  AOI21_X1 U18215 ( .B1(n14969), .B2(BUF1_REG_16__SCAN_IN), .A(n14968), .ZN(
        n14972) );
  NAND2_X1 U18216 ( .A1(n14970), .A2(DATAI_16_), .ZN(n14971) );
  OAI211_X1 U18217 ( .C1(n15172), .C2(n14995), .A(n14972), .B(n14971), .ZN(
        P1_U2888) );
  INV_X1 U18218 ( .A(n16316), .ZN(n14975) );
  OAI222_X1 U18219 ( .A1(n14995), .A2(n14975), .B1(n14988), .B2(n14974), .C1(
        n14987), .C2(n14973), .ZN(P1_U2889) );
  AOI22_X1 U18220 ( .A1(n14993), .A2(n14976), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14991), .ZN(n14977) );
  OAI21_X1 U18221 ( .B1(n15183), .B2(n14995), .A(n14977), .ZN(P1_U2890) );
  AOI22_X1 U18222 ( .A1(n14993), .A2(n14978), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14991), .ZN(n14979) );
  OAI21_X1 U18223 ( .B1(n15196), .B2(n14995), .A(n14979), .ZN(P1_U2891) );
  INV_X1 U18224 ( .A(n14980), .ZN(n14984) );
  INV_X1 U18225 ( .A(n14981), .ZN(n14983) );
  INV_X1 U18226 ( .A(n16319), .ZN(n14990) );
  INV_X1 U18227 ( .A(n14985), .ZN(n14986) );
  OAI222_X1 U18228 ( .A1(n14990), .A2(n14995), .B1(n14989), .B2(n14988), .C1(
        n14987), .C2(n14986), .ZN(P1_U2892) );
  INV_X1 U18229 ( .A(n16328), .ZN(n14996) );
  AOI22_X1 U18230 ( .A1(n14993), .A2(n14992), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14991), .ZN(n14994) );
  OAI21_X1 U18231 ( .B1(n14996), .B2(n14995), .A(n14994), .ZN(P1_U2893) );
  NAND2_X1 U18232 ( .A1(n15011), .A2(n16384), .ZN(n14998) );
  AND2_X1 U18233 ( .A1(n15011), .A2(n15208), .ZN(n15001) );
  OR2_X1 U18234 ( .A1(n9685), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15154) );
  NAND2_X1 U18235 ( .A1(n9685), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14999) );
  NAND2_X1 U18236 ( .A1(n15154), .A2(n14999), .ZN(n15162) );
  NAND2_X1 U18237 ( .A1(n9685), .A2(n15368), .ZN(n15000) );
  NAND2_X1 U18238 ( .A1(n15162), .A2(n15000), .ZN(n15153) );
  NAND2_X1 U18239 ( .A1(n15011), .A2(n15008), .ZN(n15002) );
  NAND2_X1 U18240 ( .A1(n15173), .A2(n15002), .ZN(n15190) );
  INV_X1 U18241 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15398) );
  NAND2_X1 U18242 ( .A1(n15011), .A2(n15398), .ZN(n15188) );
  NAND2_X1 U18243 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15003) );
  NAND2_X1 U18244 ( .A1(n15011), .A2(n15003), .ZN(n15185) );
  NAND2_X1 U18245 ( .A1(n15188), .A2(n15185), .ZN(n15004) );
  NOR2_X1 U18246 ( .A1(n15190), .A2(n15004), .ZN(n15150) );
  INV_X1 U18247 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15006) );
  NAND2_X1 U18248 ( .A1(n15006), .A2(n15005), .ZN(n15184) );
  NOR2_X1 U18249 ( .A1(n15184), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15007) );
  NOR2_X1 U18250 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15161) );
  AND4_X1 U18251 ( .A1(n15161), .A2(n15208), .A3(n15376), .A4(n15008), .ZN(
        n15009) );
  XNOR2_X1 U18252 ( .A(n15011), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15143) );
  AND2_X1 U18253 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15316) );
  NAND2_X1 U18254 ( .A1(n15012), .A2(n10184), .ZN(n15013) );
  INV_X1 U18255 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15356) );
  NAND2_X1 U18256 ( .A1(n15352), .A2(n15356), .ZN(n15015) );
  INV_X1 U18257 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15333) );
  INV_X1 U18258 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15337) );
  NAND2_X1 U18259 ( .A1(n15333), .A2(n15337), .ZN(n15016) );
  NAND3_X1 U18260 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15270) );
  NAND2_X1 U18261 ( .A1(n15050), .A2(n15270), .ZN(n15018) );
  NAND3_X1 U18262 ( .A1(n15018), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15081), .ZN(n15063) );
  NAND3_X1 U18263 ( .A1(n15300), .A2(n15273), .A3(n15221), .ZN(n15051) );
  AND2_X1 U18264 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15252) );
  NAND2_X1 U18265 ( .A1(n15252), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15211) );
  NAND2_X1 U18266 ( .A1(n15037), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15024) );
  NOR2_X1 U18267 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15251) );
  XNOR2_X1 U18268 ( .A(n15025), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15234) );
  NAND2_X1 U18269 ( .A1(n15026), .A2(n16332), .ZN(n15032) );
  INV_X1 U18270 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n15027) );
  NOR2_X1 U18271 ( .A1(n20393), .A2(n15027), .ZN(n15212) );
  NOR2_X1 U18272 ( .A1(n15201), .A2(n15028), .ZN(n15029) );
  AOI211_X1 U18273 ( .C1(n16321), .C2(n15030), .A(n15212), .B(n15029), .ZN(
        n15031) );
  OAI211_X1 U18274 ( .C1(n15234), .C2(n20363), .A(n15032), .B(n15031), .ZN(
        P1_U2968) );
  NOR2_X1 U18275 ( .A1(n20393), .A2(n15033), .ZN(n15237) );
  INV_X1 U18276 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15034) );
  NOR2_X1 U18277 ( .A1(n15201), .A2(n15034), .ZN(n15035) );
  AOI211_X1 U18278 ( .C1(n16321), .C2(n15036), .A(n15237), .B(n15035), .ZN(
        n15039) );
  NAND2_X1 U18279 ( .A1(n15235), .A2(n16345), .ZN(n15038) );
  OAI211_X1 U18280 ( .C1(n15040), .C2(n20422), .A(n15039), .B(n15038), .ZN(
        P1_U2969) );
  XNOR2_X1 U18281 ( .A(n16312), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15042) );
  XNOR2_X1 U18282 ( .A(n15041), .B(n15042), .ZN(n15249) );
  NOR2_X1 U18283 ( .A1(n20393), .A2(n21025), .ZN(n15243) );
  AOI21_X1 U18284 ( .B1(n20357), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15243), .ZN(n15043) );
  OAI21_X1 U18285 ( .B1(n20368), .B2(n15044), .A(n15043), .ZN(n15045) );
  INV_X1 U18286 ( .A(n15045), .ZN(n15046) );
  INV_X1 U18287 ( .A(n15048), .ZN(n15049) );
  OAI21_X1 U18288 ( .B1(n15249), .B2(n20363), .A(n15049), .ZN(P1_U2970) );
  NAND2_X1 U18289 ( .A1(n9685), .A2(n15270), .ZN(n15071) );
  NAND2_X1 U18290 ( .A1(n15050), .A2(n15071), .ZN(n15054) );
  OAI21_X1 U18291 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15051), .A(
        n15054), .ZN(n15053) );
  INV_X1 U18292 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15262) );
  MUX2_X1 U18293 ( .A(n15262), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n9685), .Z(n15052) );
  OAI211_X1 U18294 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15054), .A(
        n15053), .B(n15052), .ZN(n15055) );
  XOR2_X1 U18295 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n15055), .Z(
        n15259) );
  NOR2_X1 U18296 ( .A1(n20393), .A2(n15056), .ZN(n15254) );
  AOI21_X1 U18297 ( .B1(n20357), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15254), .ZN(n15057) );
  OAI21_X1 U18298 ( .B1(n20368), .B2(n15058), .A(n15057), .ZN(n15059) );
  AOI21_X1 U18299 ( .B1(n15060), .B2(n16332), .A(n15059), .ZN(n15061) );
  OAI21_X1 U18300 ( .B1(n20363), .B2(n15259), .A(n15061), .ZN(P1_U2971) );
  MUX2_X1 U18301 ( .A(n15063), .B(n15062), .S(n15135), .Z(n15064) );
  XNOR2_X1 U18302 ( .A(n15064), .B(n15262), .ZN(n15269) );
  INV_X1 U18303 ( .A(n15065), .ZN(n15067) );
  NOR2_X1 U18304 ( .A1(n20393), .A2(n21021), .ZN(n15261) );
  AOI21_X1 U18305 ( .B1(n20357), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15261), .ZN(n15066) );
  OAI21_X1 U18306 ( .B1(n20368), .B2(n15067), .A(n15066), .ZN(n15068) );
  AOI21_X1 U18307 ( .B1(n15069), .B2(n16332), .A(n15068), .ZN(n15070) );
  OAI21_X1 U18308 ( .B1(n20363), .B2(n15269), .A(n15070), .ZN(P1_U2972) );
  OAI211_X1 U18309 ( .C1(n15135), .C2(n15050), .A(n15072), .B(n15071), .ZN(
        n15073) );
  XOR2_X1 U18310 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15073), .Z(
        n15280) );
  INV_X1 U18311 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15074) );
  NOR2_X1 U18312 ( .A1(n20393), .A2(n15074), .ZN(n15271) );
  AOI21_X1 U18313 ( .B1(n20357), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15271), .ZN(n15075) );
  OAI21_X1 U18314 ( .B1(n20368), .B2(n15076), .A(n15075), .ZN(n15077) );
  AOI21_X1 U18315 ( .B1(n15078), .B2(n16332), .A(n15077), .ZN(n15079) );
  OAI21_X1 U18316 ( .B1(n20363), .B2(n15280), .A(n15079), .ZN(P1_U2973) );
  NAND2_X1 U18317 ( .A1(n15300), .A2(n15221), .ZN(n15080) );
  NOR2_X1 U18318 ( .A1(n15050), .A2(n15080), .ZN(n15083) );
  NAND2_X1 U18319 ( .A1(n15081), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15091) );
  NOR2_X1 U18320 ( .A1(n15091), .A2(n15221), .ZN(n15082) );
  MUX2_X1 U18321 ( .A(n15083), .B(n15082), .S(n16312), .Z(n15084) );
  XNOR2_X1 U18322 ( .A(n15084), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15287) );
  NOR2_X1 U18323 ( .A1(n20393), .A2(n15085), .ZN(n15282) );
  AOI21_X1 U18324 ( .B1(n20357), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15282), .ZN(n15086) );
  OAI21_X1 U18325 ( .B1(n20368), .B2(n15087), .A(n15086), .ZN(n15088) );
  AOI21_X1 U18326 ( .B1(n15089), .B2(n16332), .A(n15088), .ZN(n15090) );
  OAI21_X1 U18327 ( .B1(n20363), .B2(n15287), .A(n15090), .ZN(P1_U2974) );
  NOR2_X1 U18328 ( .A1(n15050), .A2(n16312), .ZN(n15092) );
  MUX2_X1 U18329 ( .A(n16312), .B(n15092), .S(n15091), .Z(n15093) );
  XNOR2_X1 U18330 ( .A(n15093), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15296) );
  NOR2_X1 U18331 ( .A1(n20393), .A2(n15094), .ZN(n15290) );
  AOI21_X1 U18332 ( .B1(n20357), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15290), .ZN(n15095) );
  OAI21_X1 U18333 ( .B1(n20368), .B2(n15096), .A(n15095), .ZN(n15097) );
  AOI21_X1 U18334 ( .B1(n15098), .B2(n16332), .A(n15097), .ZN(n15099) );
  OAI21_X1 U18335 ( .B1(n15296), .B2(n20363), .A(n15099), .ZN(P1_U2975) );
  XNOR2_X1 U18336 ( .A(n16312), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15100) );
  XNOR2_X1 U18337 ( .A(n15050), .B(n15100), .ZN(n15305) );
  INV_X1 U18338 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n15101) );
  NOR2_X1 U18339 ( .A1(n20393), .A2(n15101), .ZN(n15299) );
  AOI21_X1 U18340 ( .B1(n20357), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15299), .ZN(n15102) );
  OAI21_X1 U18341 ( .B1(n20368), .B2(n15103), .A(n15102), .ZN(n15104) );
  AOI21_X1 U18342 ( .B1(n15105), .B2(n16332), .A(n15104), .ZN(n15106) );
  OAI21_X1 U18343 ( .B1(n15305), .B2(n20363), .A(n15106), .ZN(P1_U2976) );
  NAND2_X1 U18344 ( .A1(n15108), .A2(n15107), .ZN(n15109) );
  XOR2_X1 U18345 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15109), .Z(
        n15325) );
  INV_X1 U18346 ( .A(n15110), .ZN(n15113) );
  NOR2_X1 U18347 ( .A1(n20393), .A2(n15111), .ZN(n15320) );
  AOI21_X1 U18348 ( .B1(n20357), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15320), .ZN(n15112) );
  OAI21_X1 U18349 ( .B1(n20368), .B2(n15113), .A(n15112), .ZN(n15114) );
  AOI21_X1 U18350 ( .B1(n15115), .B2(n16332), .A(n15114), .ZN(n15116) );
  OAI21_X1 U18351 ( .B1(n20363), .B2(n15325), .A(n15116), .ZN(P1_U2977) );
  NOR3_X1 U18352 ( .A1(n15142), .A2(n15135), .A3(n15352), .ZN(n15127) );
  NOR2_X1 U18353 ( .A1(n15118), .A2(n9685), .ZN(n15126) );
  AOI22_X1 U18354 ( .A1(n15127), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n15126), .B2(n15337), .ZN(n15119) );
  XNOR2_X1 U18355 ( .A(n15119), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15326) );
  NAND2_X1 U18356 ( .A1(n15326), .A2(n16345), .ZN(n15124) );
  NOR2_X1 U18357 ( .A1(n20393), .A2(n15120), .ZN(n15329) );
  NOR2_X1 U18358 ( .A1(n20368), .A2(n15121), .ZN(n15122) );
  AOI211_X1 U18359 ( .C1(n20357), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15329), .B(n15122), .ZN(n15123) );
  OAI211_X1 U18360 ( .C1(n20422), .C2(n15125), .A(n15124), .B(n15123), .ZN(
        P1_U2978) );
  NOR2_X1 U18361 ( .A1(n15127), .A2(n15126), .ZN(n15128) );
  XNOR2_X1 U18362 ( .A(n15128), .B(n15337), .ZN(n15345) );
  NOR2_X1 U18363 ( .A1(n20393), .A2(n21012), .ZN(n15335) );
  NOR2_X1 U18364 ( .A1(n15201), .A2(n21227), .ZN(n15129) );
  AOI211_X1 U18365 ( .C1(n16321), .C2(n15130), .A(n15335), .B(n15129), .ZN(
        n15133) );
  NAND2_X1 U18366 ( .A1(n15131), .A2(n16332), .ZN(n15132) );
  OAI211_X1 U18367 ( .C1(n15345), .C2(n20363), .A(n15133), .B(n15132), .ZN(
        P1_U2979) );
  NAND2_X1 U18368 ( .A1(n15135), .A2(n15356), .ZN(n15134) );
  MUX2_X1 U18369 ( .A(n15135), .B(n15134), .S(n15142), .Z(n15136) );
  XNOR2_X1 U18370 ( .A(n15136), .B(n15352), .ZN(n15354) );
  NAND2_X1 U18371 ( .A1(n20407), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15347) );
  NAND2_X1 U18372 ( .A1(n20357), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15137) );
  OAI211_X1 U18373 ( .C1(n20368), .C2(n15138), .A(n15347), .B(n15137), .ZN(
        n15139) );
  AOI21_X1 U18374 ( .B1(n15140), .B2(n16332), .A(n15139), .ZN(n15141) );
  OAI21_X1 U18375 ( .B1(n15354), .B2(n20363), .A(n15141), .ZN(P1_U2980) );
  OAI21_X1 U18376 ( .B1(n15014), .B2(n15143), .A(n15142), .ZN(n15364) );
  NOR2_X1 U18377 ( .A1(n20393), .A2(n21009), .ZN(n15358) );
  AOI21_X1 U18378 ( .B1(n20357), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15358), .ZN(n15144) );
  OAI21_X1 U18379 ( .B1(n20368), .B2(n15145), .A(n15144), .ZN(n15146) );
  AOI21_X1 U18380 ( .B1(n15147), .B2(n16332), .A(n15146), .ZN(n15148) );
  OAI21_X1 U18381 ( .B1(n20363), .B2(n15364), .A(n15148), .ZN(P1_U2981) );
  INV_X1 U18382 ( .A(n15150), .ZN(n15151) );
  AOI21_X1 U18383 ( .B1(n15149), .B2(n10172), .A(n15151), .ZN(n15175) );
  OAI21_X1 U18384 ( .B1(n15135), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15175), .ZN(n15152) );
  OAI211_X1 U18385 ( .C1(n15376), .C2(n9685), .A(n15152), .B(n15173), .ZN(
        n16314) );
  AOI21_X1 U18386 ( .B1(n15135), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16314), .ZN(n15160) );
  NOR2_X1 U18387 ( .A1(n15160), .A2(n15153), .ZN(n15165) );
  MUX2_X1 U18388 ( .A(n15160), .B(n15165), .S(n15154), .Z(n15155) );
  XNOR2_X1 U18389 ( .A(n15155), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15374) );
  INV_X1 U18390 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15156) );
  NOR2_X1 U18391 ( .A1(n20393), .A2(n15156), .ZN(n15367) );
  NOR2_X1 U18392 ( .A1(n15201), .A2(n16277), .ZN(n15157) );
  AOI211_X1 U18393 ( .C1(n16321), .C2(n16279), .A(n15367), .B(n15157), .ZN(
        n15159) );
  NAND2_X1 U18394 ( .A1(n16307), .A2(n16332), .ZN(n15158) );
  OAI211_X1 U18395 ( .C1(n15374), .C2(n20363), .A(n15159), .B(n15158), .ZN(
        P1_U2982) );
  INV_X1 U18396 ( .A(n15160), .ZN(n15164) );
  INV_X1 U18397 ( .A(n15161), .ZN(n15163) );
  AOI21_X1 U18398 ( .B1(n15164), .B2(n15163), .A(n15162), .ZN(n15166) );
  NOR2_X1 U18399 ( .A1(n15166), .A2(n15165), .ZN(n15375) );
  NAND2_X1 U18400 ( .A1(n15375), .A2(n16345), .ZN(n15171) );
  OR2_X1 U18401 ( .A1(n20393), .A2(n21006), .ZN(n15380) );
  OAI21_X1 U18402 ( .B1(n15201), .B2(n15167), .A(n15380), .ZN(n15168) );
  AOI21_X1 U18403 ( .B1(n16321), .B2(n15169), .A(n15168), .ZN(n15170) );
  OAI211_X1 U18404 ( .C1(n20422), .C2(n15172), .A(n15171), .B(n15170), .ZN(
        P1_U2983) );
  INV_X1 U18405 ( .A(n15173), .ZN(n15174) );
  NOR2_X1 U18406 ( .A1(n15175), .A2(n15174), .ZN(n15177) );
  XNOR2_X1 U18407 ( .A(n16312), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15176) );
  XNOR2_X1 U18408 ( .A(n15177), .B(n15176), .ZN(n16357) );
  NAND2_X1 U18409 ( .A1(n16357), .A2(n16345), .ZN(n15182) );
  INV_X1 U18410 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n15178) );
  OAI22_X1 U18411 ( .A1(n15201), .A2(n21218), .B1(n20393), .B2(n15178), .ZN(
        n15179) );
  AOI21_X1 U18412 ( .B1(n15180), .B2(n16321), .A(n15179), .ZN(n15181) );
  OAI211_X1 U18413 ( .C1(n20422), .C2(n15183), .A(n15182), .B(n15181), .ZN(
        P1_U2985) );
  INV_X1 U18414 ( .A(n15149), .ZN(n15186) );
  AOI22_X1 U18415 ( .A1(n15186), .A2(n15185), .B1(n15135), .B2(n15184), .ZN(
        n15388) );
  INV_X1 U18416 ( .A(n15188), .ZN(n15187) );
  AOI21_X1 U18417 ( .B1(n15135), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15187), .ZN(n15387) );
  NAND2_X1 U18418 ( .A1(n15388), .A2(n15387), .ZN(n15386) );
  NAND2_X1 U18419 ( .A1(n15386), .A2(n15188), .ZN(n15189) );
  XOR2_X1 U18420 ( .A(n15190), .B(n15189), .Z(n16368) );
  NAND2_X1 U18421 ( .A1(n16368), .A2(n16345), .ZN(n15195) );
  INV_X1 U18422 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15191) );
  OAI22_X1 U18423 ( .A1(n15201), .A2(n15191), .B1(n20393), .B2(n21001), .ZN(
        n15192) );
  AOI21_X1 U18424 ( .B1(n16321), .B2(n15193), .A(n15192), .ZN(n15194) );
  OAI211_X1 U18425 ( .C1(n20422), .C2(n15196), .A(n15195), .B(n15194), .ZN(
        P1_U2986) );
  MUX2_X1 U18426 ( .A(n15197), .B(n15149), .S(n16312), .Z(n15198) );
  XNOR2_X1 U18427 ( .A(n15198), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16382) );
  NAND2_X1 U18428 ( .A1(n16382), .A2(n16345), .ZN(n15205) );
  INV_X1 U18429 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15199) );
  OAI22_X1 U18430 ( .A1(n15201), .A2(n15200), .B1(n20393), .B2(n15199), .ZN(
        n15202) );
  AOI21_X1 U18431 ( .B1(n16321), .B2(n15203), .A(n15202), .ZN(n15204) );
  OAI211_X1 U18432 ( .C1(n20422), .C2(n15206), .A(n15205), .B(n15204), .ZN(
        P1_U2989) );
  NOR3_X1 U18433 ( .A1(n15006), .A2(n16384), .A3(n15207), .ZN(n15391) );
  NAND2_X1 U18434 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15391), .ZN(
        n15395) );
  NOR2_X1 U18435 ( .A1(n15398), .A2(n15395), .ZN(n16361) );
  NAND2_X1 U18436 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16361), .ZN(
        n15214) );
  NAND2_X1 U18437 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15218) );
  INV_X1 U18438 ( .A(n15218), .ZN(n15317) );
  INV_X1 U18439 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15369) );
  NOR4_X1 U18440 ( .A1(n15368), .A2(n15376), .A3(n15208), .A4(n15369), .ZN(
        n15360) );
  NAND2_X1 U18441 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15360), .ZN(
        n15311) );
  INV_X1 U18442 ( .A(n15311), .ZN(n15313) );
  AND3_X1 U18443 ( .A1(n15316), .A2(n15317), .A3(n15313), .ZN(n15209) );
  NAND2_X1 U18444 ( .A1(n16355), .A2(n15209), .ZN(n15288) );
  INV_X1 U18445 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15210) );
  NOR2_X1 U18446 ( .A1(n15260), .A2(n15211), .ZN(n15236) );
  NOR2_X1 U18447 ( .A1(n15023), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15213) );
  AOI21_X1 U18448 ( .B1(n15236), .B2(n15213), .A(n15212), .ZN(n15230) );
  NOR2_X1 U18449 ( .A1(n15308), .A2(n15214), .ZN(n15312) );
  OAI21_X1 U18450 ( .B1(n15214), .B2(n15307), .A(n20390), .ZN(n15215) );
  OAI211_X1 U18451 ( .C1(n20372), .C2(n15312), .A(n20371), .B(n15215), .ZN(
        n16367) );
  AND2_X1 U18452 ( .A1(n15377), .A2(n15311), .ZN(n15216) );
  NOR2_X1 U18453 ( .A1(n16367), .A2(n15216), .ZN(n15349) );
  NAND2_X1 U18454 ( .A1(n15349), .A2(n15316), .ZN(n15341) );
  NAND2_X1 U18455 ( .A1(n15341), .A2(n15217), .ZN(n15334) );
  NAND2_X1 U18456 ( .A1(n15377), .A2(n15218), .ZN(n15219) );
  NAND2_X1 U18457 ( .A1(n15334), .A2(n15219), .ZN(n15302) );
  NOR2_X1 U18458 ( .A1(n20370), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15220) );
  NAND2_X1 U18459 ( .A1(n15377), .A2(n15221), .ZN(n15222) );
  OAI21_X1 U18460 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n20372), .A(
        n15222), .ZN(n15223) );
  OR2_X1 U18461 ( .A1(n15293), .A2(n15223), .ZN(n15284) );
  NAND2_X1 U18462 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15224) );
  OR2_X1 U18463 ( .A1(n15293), .A2(n15377), .ZN(n15228) );
  OAI21_X1 U18464 ( .B1(n15284), .B2(n15224), .A(n15228), .ZN(n15256) );
  INV_X1 U18465 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15225) );
  AOI21_X1 U18466 ( .B1(n15228), .B2(n15019), .A(n15225), .ZN(n15226) );
  NAND2_X1 U18467 ( .A1(n15256), .A2(n15226), .ZN(n15245) );
  NAND2_X1 U18468 ( .A1(n15245), .A2(n15228), .ZN(n15227) );
  NAND2_X1 U18469 ( .A1(n15227), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15239) );
  NAND3_X1 U18470 ( .A1(n15239), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15228), .ZN(n15229) );
  OAI211_X1 U18471 ( .C1(n15231), .C2(n16412), .A(n15230), .B(n15229), .ZN(
        n15232) );
  INV_X1 U18472 ( .A(n15232), .ZN(n15233) );
  OAI21_X1 U18473 ( .B1(n15234), .B2(n20408), .A(n15233), .ZN(P1_U3000) );
  NAND2_X1 U18474 ( .A1(n15235), .A2(n20399), .ZN(n15241) );
  OR2_X1 U18475 ( .A1(n15236), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15238) );
  AOI21_X1 U18476 ( .B1(n15239), .B2(n15238), .A(n15237), .ZN(n15240) );
  OAI211_X1 U18477 ( .C1(n16412), .C2(n15242), .A(n15241), .B(n15240), .ZN(
        P1_U3001) );
  AOI21_X1 U18478 ( .B1(n15244), .B2(n20406), .A(n15243), .ZN(n15248) );
  NOR2_X1 U18479 ( .A1(n15260), .A2(n15019), .ZN(n15246) );
  OAI21_X1 U18480 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15246), .A(
        n15245), .ZN(n15247) );
  OAI211_X1 U18481 ( .C1(n15249), .C2(n20408), .A(n15248), .B(n15247), .ZN(
        P1_U3002) );
  INV_X1 U18482 ( .A(n15250), .ZN(n15255) );
  NOR3_X1 U18483 ( .A1(n15260), .A2(n15252), .A3(n15251), .ZN(n15253) );
  AOI211_X1 U18484 ( .C1(n15255), .C2(n20406), .A(n15254), .B(n15253), .ZN(
        n15258) );
  INV_X1 U18485 ( .A(n15256), .ZN(n15267) );
  NAND2_X1 U18486 ( .A1(n15267), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15257) );
  OAI211_X1 U18487 ( .C1(n15259), .C2(n20408), .A(n15258), .B(n15257), .ZN(
        P1_U3003) );
  INV_X1 U18488 ( .A(n15260), .ZN(n15263) );
  AOI21_X1 U18489 ( .B1(n15263), .B2(n15262), .A(n15261), .ZN(n15264) );
  OAI21_X1 U18490 ( .B1(n15265), .B2(n16412), .A(n15264), .ZN(n15266) );
  AOI21_X1 U18491 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15267), .A(
        n15266), .ZN(n15268) );
  OAI21_X1 U18492 ( .B1(n15269), .B2(n20408), .A(n15268), .ZN(P1_U3004) );
  INV_X1 U18493 ( .A(n15288), .ZN(n15301) );
  NOR2_X1 U18494 ( .A1(n15270), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15272) );
  AOI21_X1 U18495 ( .B1(n15301), .B2(n15272), .A(n15271), .ZN(n15276) );
  NAND3_X1 U18496 ( .A1(n15273), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15274) );
  NOR2_X1 U18497 ( .A1(n15288), .A2(n15274), .ZN(n15281) );
  OAI21_X1 U18498 ( .B1(n15284), .B2(n15281), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15275) );
  OAI211_X1 U18499 ( .C1(n15277), .C2(n16412), .A(n15276), .B(n15275), .ZN(
        n15278) );
  INV_X1 U18500 ( .A(n15278), .ZN(n15279) );
  OAI21_X1 U18501 ( .B1(n15280), .B2(n20408), .A(n15279), .ZN(P1_U3005) );
  AOI211_X1 U18502 ( .C1(n15283), .C2(n20406), .A(n15282), .B(n15281), .ZN(
        n15286) );
  NAND2_X1 U18503 ( .A1(n15284), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15285) );
  OAI211_X1 U18504 ( .C1(n15287), .C2(n20408), .A(n15286), .B(n15285), .ZN(
        P1_U3006) );
  NOR3_X1 U18505 ( .A1(n15288), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15300), .ZN(n15289) );
  AOI211_X1 U18506 ( .C1(n15291), .C2(n20406), .A(n15290), .B(n15289), .ZN(
        n15295) );
  NOR2_X1 U18507 ( .A1(n20411), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15292) );
  OAI21_X1 U18508 ( .B1(n15293), .B2(n15292), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15294) );
  OAI211_X1 U18509 ( .C1(n15296), .C2(n20408), .A(n15295), .B(n15294), .ZN(
        P1_U3007) );
  NOR2_X1 U18510 ( .A1(n15297), .A2(n16412), .ZN(n15298) );
  AOI211_X1 U18511 ( .C1(n15301), .C2(n15300), .A(n15299), .B(n15298), .ZN(
        n15304) );
  NAND2_X1 U18512 ( .A1(n15302), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15303) );
  OAI211_X1 U18513 ( .C1(n15305), .C2(n20408), .A(n15304), .B(n15303), .ZN(
        P1_U3008) );
  INV_X1 U18514 ( .A(n15306), .ZN(n15321) );
  INV_X1 U18515 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15318) );
  NOR2_X1 U18516 ( .A1(n20370), .A2(n15307), .ZN(n15310) );
  INV_X1 U18517 ( .A(n15308), .ZN(n16362) );
  OAI221_X1 U18518 ( .B1(n15310), .B2(n16362), .C1(n15310), .C2(n15309), .A(
        n16361), .ZN(n16363) );
  OR3_X1 U18519 ( .A1(n16363), .A2(n15008), .A3(n15311), .ZN(n15339) );
  NAND3_X1 U18520 ( .A1(n15314), .A2(n15313), .A3(n15312), .ZN(n15315) );
  NAND2_X1 U18521 ( .A1(n15339), .A2(n15315), .ZN(n15351) );
  NAND2_X1 U18522 ( .A1(n15351), .A2(n15316), .ZN(n15327) );
  AOI211_X1 U18523 ( .C1(n15333), .C2(n15318), .A(n15317), .B(n15327), .ZN(
        n15319) );
  AOI211_X1 U18524 ( .C1(n20406), .C2(n15321), .A(n15320), .B(n15319), .ZN(
        n15324) );
  INV_X1 U18525 ( .A(n15334), .ZN(n15322) );
  NAND2_X1 U18526 ( .A1(n15322), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15323) );
  OAI211_X1 U18527 ( .C1(n15325), .C2(n20408), .A(n15324), .B(n15323), .ZN(
        P1_U3009) );
  NAND2_X1 U18528 ( .A1(n15326), .A2(n20399), .ZN(n15332) );
  NOR2_X1 U18529 ( .A1(n15327), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15328) );
  AOI211_X1 U18530 ( .C1(n20406), .C2(n15330), .A(n15329), .B(n15328), .ZN(
        n15331) );
  OAI211_X1 U18531 ( .C1(n15334), .C2(n15333), .A(n15332), .B(n15331), .ZN(
        P1_U3010) );
  AOI21_X1 U18532 ( .B1(n15336), .B2(n20406), .A(n15335), .ZN(n15344) );
  INV_X1 U18533 ( .A(n15351), .ZN(n15338) );
  OAI21_X1 U18534 ( .B1(n15338), .B2(n15352), .A(n15337), .ZN(n15342) );
  NAND3_X1 U18535 ( .A1(n15349), .A2(n16364), .A3(n15339), .ZN(n15340) );
  NAND3_X1 U18536 ( .A1(n15342), .A2(n15341), .A3(n15340), .ZN(n15343) );
  OAI211_X1 U18537 ( .C1(n15345), .C2(n20408), .A(n15344), .B(n15343), .ZN(
        P1_U3011) );
  NAND2_X1 U18538 ( .A1(n15346), .A2(n20406), .ZN(n15348) );
  OAI211_X1 U18539 ( .C1(n15349), .C2(n15352), .A(n15348), .B(n15347), .ZN(
        n15350) );
  AOI21_X1 U18540 ( .B1(n15352), .B2(n15351), .A(n15350), .ZN(n15353) );
  OAI21_X1 U18541 ( .B1(n15354), .B2(n20408), .A(n15353), .ZN(P1_U3012) );
  INV_X1 U18542 ( .A(n15355), .ZN(n15359) );
  AND3_X1 U18543 ( .A1(n15356), .A2(n15360), .A3(n16355), .ZN(n15357) );
  AOI211_X1 U18544 ( .C1(n15359), .C2(n20406), .A(n15358), .B(n15357), .ZN(
        n15363) );
  INV_X1 U18545 ( .A(n16367), .ZN(n15379) );
  OAI21_X1 U18546 ( .B1(n15361), .B2(n15360), .A(n15379), .ZN(n15370) );
  NAND2_X1 U18547 ( .A1(n15370), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15362) );
  OAI211_X1 U18548 ( .C1(n15364), .C2(n20408), .A(n15363), .B(n15362), .ZN(
        P1_U3013) );
  INV_X1 U18549 ( .A(n15365), .ZN(n15366) );
  XNOR2_X1 U18550 ( .A(n14799), .B(n15366), .ZN(n16306) );
  AOI21_X1 U18551 ( .B1(n16306), .B2(n20406), .A(n15367), .ZN(n15373) );
  NAND2_X1 U18552 ( .A1(n16355), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16354) );
  NOR3_X1 U18553 ( .A1(n16354), .A2(n15369), .A3(n15368), .ZN(n15371) );
  OAI21_X1 U18554 ( .B1(n15371), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15370), .ZN(n15372) );
  OAI211_X1 U18555 ( .C1(n15374), .C2(n20408), .A(n15373), .B(n15372), .ZN(
        P1_U3014) );
  XNOR2_X1 U18556 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15385) );
  NAND2_X1 U18557 ( .A1(n15375), .A2(n20399), .ZN(n15384) );
  NAND2_X1 U18558 ( .A1(n15377), .A2(n15376), .ZN(n15378) );
  NAND2_X1 U18559 ( .A1(n15379), .A2(n15378), .ZN(n16352) );
  OAI21_X1 U18560 ( .B1(n15381), .B2(n16412), .A(n15380), .ZN(n15382) );
  AOI21_X1 U18561 ( .B1(n16352), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15382), .ZN(n15383) );
  OAI211_X1 U18562 ( .C1(n16354), .C2(n15385), .A(n15384), .B(n15383), .ZN(
        P1_U3015) );
  OAI21_X1 U18563 ( .B1(n15388), .B2(n15387), .A(n15386), .ZN(n15389) );
  INV_X1 U18564 ( .A(n15389), .ZN(n16324) );
  NAND3_X1 U18565 ( .A1(n15391), .A2(n15390), .A3(n15005), .ZN(n16374) );
  AOI21_X1 U18566 ( .B1(n16362), .B2(n15391), .A(n20372), .ZN(n15393) );
  AOI211_X1 U18567 ( .C1(n20390), .C2(n15395), .A(n15393), .B(n15392), .ZN(
        n16373) );
  OAI21_X1 U18568 ( .B1(n15394), .B2(n16374), .A(n16373), .ZN(n15397) );
  OAI21_X1 U18569 ( .B1(n15395), .B2(n16396), .A(n15398), .ZN(n15396) );
  OAI21_X1 U18570 ( .B1(n15398), .B2(n15397), .A(n15396), .ZN(n15404) );
  OAI21_X1 U18571 ( .B1(n15401), .B2(n15400), .A(n15399), .ZN(n15402) );
  INV_X1 U18572 ( .A(n15402), .ZN(n16309) );
  AOI22_X1 U18573 ( .A1(n16309), .A2(n20406), .B1(n20407), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15403) );
  OAI211_X1 U18574 ( .C1(n16324), .C2(n20408), .A(n15404), .B(n15403), .ZN(
        P1_U3019) );
  OR2_X1 U18575 ( .A1(n9702), .A2(n20903), .ZN(n15405) );
  NAND2_X1 U18576 ( .A1(n15405), .A2(n20789), .ZN(n20525) );
  OAI21_X1 U18577 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9702), .A(n20525), 
        .ZN(n15406) );
  OAI21_X1 U18578 ( .B1(n9697), .B2(n15410), .A(n15406), .ZN(n15407) );
  MUX2_X1 U18579 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15407), .S(
        n20417), .Z(P1_U3477) );
  INV_X1 U18580 ( .A(n20525), .ZN(n20902) );
  MUX2_X1 U18581 ( .A(n20902), .B(n15408), .S(n13627), .Z(n15409) );
  OAI21_X1 U18582 ( .B1(n15410), .B2(n13223), .A(n15409), .ZN(n15411) );
  MUX2_X1 U18583 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15411), .S(
        n20417), .Z(P1_U3476) );
  NOR3_X1 U18584 ( .A1(n15412), .A2(n11008), .A3(n11010), .ZN(n15415) );
  NOR2_X1 U18585 ( .A1(n9697), .A2(n15413), .ZN(n15414) );
  AOI211_X1 U18586 ( .C1(n16211), .C2(n10996), .A(n15415), .B(n15414), .ZN(
        n16216) );
  INV_X1 U18587 ( .A(n16419), .ZN(n15424) );
  NOR3_X1 U18588 ( .A1(n11010), .A2(n11008), .A3(n15422), .ZN(n15416) );
  AOI21_X1 U18589 ( .B1(n15418), .B2(n15417), .A(n15416), .ZN(n15419) );
  OAI21_X1 U18590 ( .B1(n16216), .B2(n15424), .A(n15419), .ZN(n15420) );
  MUX2_X1 U18591 ( .A(n15420), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n16417), .Z(P1_U3473) );
  INV_X1 U18592 ( .A(n15421), .ZN(n15423) );
  OAI22_X1 U18593 ( .A1(n15425), .A2(n15424), .B1(n15423), .B2(n15422), .ZN(
        n15426) );
  MUX2_X1 U18594 ( .A(n15426), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16417), .Z(P1_U3469) );
  NAND4_X1 U18595 ( .A1(n15427), .A2(n19308), .A3(n12811), .A4(n15692), .ZN(
        n15434) );
  INV_X1 U18596 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15428) );
  INV_X1 U18597 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20165) );
  OAI22_X1 U18598 ( .A1(n15428), .A2(n19326), .B1(n20165), .B2(n19260), .ZN(
        n15431) );
  NAND3_X1 U18599 ( .A1(n19480), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n16613), 
        .ZN(n15429) );
  OAI21_X1 U18600 ( .B1(n19333), .B2(n19312), .A(n15429), .ZN(n15430) );
  OAI211_X1 U18601 ( .C1(n15435), .C2(n19292), .A(n15434), .B(n15433), .ZN(
        P2_U2824) );
  NOR2_X1 U18602 ( .A1(n15437), .A2(n15436), .ZN(n15438) );
  AOI21_X1 U18603 ( .B1(n15441), .B2(n15704), .A(n15440), .ZN(n15442) );
  NAND2_X1 U18604 ( .A1(n15442), .A2(n19308), .ZN(n15452) );
  INV_X1 U18605 ( .A(n15443), .ZN(n15446) );
  NAND2_X1 U18606 ( .A1(n9723), .A2(n15444), .ZN(n15445) );
  NAND2_X1 U18607 ( .A1(n15446), .A2(n15445), .ZN(n15899) );
  AOI22_X1 U18608 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19320), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19318), .ZN(n15448) );
  NAND2_X1 U18609 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19298), .ZN(
        n15447) );
  OAI211_X1 U18610 ( .C1(n15899), .C2(n19312), .A(n15448), .B(n15447), .ZN(
        n15449) );
  AOI21_X1 U18611 ( .B1(n15450), .B2(n19317), .A(n15449), .ZN(n15451) );
  OAI211_X1 U18612 ( .C1(n19292), .C2(n15703), .A(n15452), .B(n15451), .ZN(
        P2_U2827) );
  OAI21_X1 U18613 ( .B1(n15563), .B2(n15453), .A(n9740), .ZN(n15933) );
  AND2_X1 U18614 ( .A1(n15627), .A2(n15454), .ZN(n15455) );
  OR2_X1 U18615 ( .A1(n15455), .A2(n9764), .ZN(n15618) );
  AOI22_X1 U18616 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19318), .ZN(n15456) );
  OAI21_X1 U18617 ( .B1(n19312), .B2(n15618), .A(n15456), .ZN(n15457) );
  AOI21_X1 U18618 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n19320), .A(n15457), .ZN(
        n15458) );
  OAI21_X1 U18619 ( .B1(n15933), .B2(n19292), .A(n15458), .ZN(n15462) );
  AOI211_X1 U18620 ( .C1(n15460), .C2(n15739), .A(n15459), .B(n20099), .ZN(
        n15461) );
  AOI211_X1 U18621 ( .C1(n19317), .C2(n15463), .A(n15462), .B(n15461), .ZN(
        n15464) );
  INV_X1 U18622 ( .A(n15464), .ZN(P2_U2830) );
  INV_X1 U18623 ( .A(n15465), .ZN(n15481) );
  AOI211_X1 U18624 ( .C1(n15756), .C2(n15466), .A(n15467), .B(n20099), .ZN(
        n15468) );
  INV_X1 U18625 ( .A(n15468), .ZN(n15480) );
  AND2_X1 U18626 ( .A1(n15485), .A2(n15469), .ZN(n15470) );
  NOR2_X1 U18627 ( .A1(n15561), .A2(n15470), .ZN(n15965) );
  INV_X1 U18628 ( .A(n15471), .ZN(n15474) );
  NAND2_X1 U18629 ( .A1(n15486), .A2(n15472), .ZN(n15473) );
  NAND2_X1 U18630 ( .A1(n15474), .A2(n15473), .ZN(n15475) );
  NAND2_X1 U18631 ( .A1(n15475), .A2(n15625), .ZN(n15963) );
  AOI22_X1 U18632 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n19320), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19318), .ZN(n15477) );
  NAND2_X1 U18633 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19298), .ZN(
        n15476) );
  OAI211_X1 U18634 ( .C1(n19312), .C2(n15963), .A(n15477), .B(n15476), .ZN(
        n15478) );
  AOI21_X1 U18635 ( .B1(n15965), .B2(n19313), .A(n15478), .ZN(n15479) );
  OAI211_X1 U18636 ( .C1(n15481), .C2(n19300), .A(n15480), .B(n15479), .ZN(
        P2_U2832) );
  NAND2_X1 U18637 ( .A1(n15482), .A2(n15483), .ZN(n15484) );
  NAND2_X1 U18638 ( .A1(n15485), .A2(n15484), .ZN(n16485) );
  XNOR2_X1 U18639 ( .A(n15486), .B(n15472), .ZN(n15978) );
  AOI22_X1 U18640 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n19320), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19318), .ZN(n15490) );
  OAI22_X1 U18641 ( .A1(n15487), .A2(n19300), .B1(n19326), .B2(n10795), .ZN(
        n15488) );
  INV_X1 U18642 ( .A(n15488), .ZN(n15489) );
  OAI211_X1 U18643 ( .C1(n15978), .C2(n19312), .A(n15490), .B(n15489), .ZN(
        n15495) );
  AOI211_X1 U18644 ( .C1(n15493), .C2(n15491), .A(n15492), .B(n20099), .ZN(
        n15494) );
  NOR2_X1 U18645 ( .A1(n15495), .A2(n15494), .ZN(n15496) );
  OAI21_X1 U18646 ( .B1(n19292), .B2(n16485), .A(n15496), .ZN(P2_U2833) );
  INV_X1 U18647 ( .A(n15497), .ZN(n15511) );
  NOR2_X1 U18648 ( .A1(n19289), .A2(n15498), .ZN(n15499) );
  XNOR2_X1 U18649 ( .A(n15499), .B(n15828), .ZN(n15500) );
  NAND2_X1 U18650 ( .A1(n15500), .A2(n19308), .ZN(n15510) );
  NOR2_X1 U18651 ( .A1(n19260), .A2(n20141), .ZN(n15508) );
  INV_X1 U18652 ( .A(n15676), .ZN(n15505) );
  INV_X1 U18653 ( .A(n15501), .ZN(n15502) );
  NAND2_X1 U18654 ( .A1(n15503), .A2(n15502), .ZN(n15504) );
  NAND2_X1 U18655 ( .A1(n15505), .A2(n15504), .ZN(n19341) );
  AOI22_X1 U18656 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(n19320), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19298), .ZN(n15506) );
  OAI211_X1 U18657 ( .C1(n19312), .C2(n19341), .A(n15506), .B(n19277), .ZN(
        n15507) );
  AOI211_X1 U18658 ( .C1(n16062), .C2(n19313), .A(n15508), .B(n15507), .ZN(
        n15509) );
  OAI211_X1 U18659 ( .C1(n19300), .C2(n15511), .A(n15510), .B(n15509), .ZN(
        P2_U2839) );
  NOR2_X1 U18660 ( .A1(n19289), .A2(n15512), .ZN(n15513) );
  XNOR2_X1 U18661 ( .A(n15513), .B(n16514), .ZN(n15514) );
  NAND2_X1 U18662 ( .A1(n15514), .A2(n19308), .ZN(n15524) );
  OAI22_X1 U18663 ( .A1(n15516), .A2(n19300), .B1(n19326), .B2(n15515), .ZN(
        n15517) );
  INV_X1 U18664 ( .A(n15517), .ZN(n15518) );
  OAI211_X1 U18665 ( .C1(n19285), .C2(n10704), .A(n15518), .B(n19277), .ZN(
        n15519) );
  AOI21_X1 U18666 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n19318), .A(n15519), 
        .ZN(n15523) );
  AOI21_X1 U18667 ( .B1(n15521), .B2(n16165), .A(n15520), .ZN(n16158) );
  AOI22_X1 U18668 ( .A1(n19313), .A2(n16510), .B1(n19319), .B2(n16158), .ZN(
        n15522) );
  NAND3_X1 U18669 ( .A1(n15524), .A2(n15523), .A3(n15522), .ZN(P2_U2845) );
  MUX2_X1 U18670 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n15525), .S(n15572), .Z(
        P2_U2856) );
  OR2_X1 U18671 ( .A1(n15527), .A2(n15526), .ZN(n15595) );
  NAND3_X1 U18672 ( .A1(n15595), .A2(n15528), .A3(n15575), .ZN(n15530) );
  NAND2_X1 U18673 ( .A1(n15578), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15529) );
  OAI211_X1 U18674 ( .C1(n15578), .C2(n16441), .A(n15530), .B(n15529), .ZN(
        P2_U2858) );
  NAND2_X1 U18675 ( .A1(n15532), .A2(n15531), .ZN(n15534) );
  XNOR2_X1 U18676 ( .A(n15534), .B(n15533), .ZN(n15605) );
  NOR2_X1 U18677 ( .A1(n15703), .A2(n15592), .ZN(n15535) );
  AOI21_X1 U18678 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15592), .A(n15535), .ZN(
        n15536) );
  OAI21_X1 U18679 ( .B1(n15605), .B2(n15594), .A(n15536), .ZN(P2_U2859) );
  OAI21_X1 U18680 ( .B1(n15537), .B2(n15539), .A(n15538), .ZN(n15610) );
  NOR2_X1 U18681 ( .A1(n15914), .A2(n15592), .ZN(n15540) );
  AOI21_X1 U18682 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n15592), .A(n15540), .ZN(
        n15541) );
  OAI21_X1 U18683 ( .B1(n15610), .B2(n15594), .A(n15541), .ZN(P2_U2860) );
  INV_X1 U18684 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n15549) );
  AOI21_X1 U18685 ( .B1(n15544), .B2(n15543), .A(n15542), .ZN(n15616) );
  NAND2_X1 U18686 ( .A1(n15616), .A2(n15575), .ZN(n15548) );
  INV_X1 U18687 ( .A(n9722), .ZN(n15545) );
  AOI21_X1 U18688 ( .B1(n15546), .B2(n9740), .A(n15545), .ZN(n16452) );
  NAND2_X1 U18689 ( .A1(n16452), .A2(n15572), .ZN(n15547) );
  OAI211_X1 U18690 ( .C1(n15572), .C2(n15549), .A(n15548), .B(n15547), .ZN(
        P2_U2861) );
  OAI21_X1 U18691 ( .B1(n15552), .B2(n15551), .A(n15550), .ZN(n15623) );
  MUX2_X1 U18692 ( .A(n15553), .B(n15933), .S(n15572), .Z(n15554) );
  OAI21_X1 U18693 ( .B1(n15623), .B2(n15594), .A(n15554), .ZN(P2_U2862) );
  INV_X1 U18694 ( .A(n15555), .ZN(n15557) );
  AOI21_X1 U18695 ( .B1(n15557), .B2(n15556), .A(n9772), .ZN(n15558) );
  XOR2_X1 U18696 ( .A(n15559), .B(n15558), .Z(n15632) );
  NOR2_X1 U18697 ( .A1(n15561), .A2(n15560), .ZN(n15562) );
  OR2_X1 U18698 ( .A1(n15563), .A2(n15562), .ZN(n15946) );
  NOR2_X1 U18699 ( .A1(n15946), .A2(n15592), .ZN(n15564) );
  AOI21_X1 U18700 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15578), .A(n15564), .ZN(
        n15565) );
  OAI21_X1 U18701 ( .B1(n15632), .B2(n15594), .A(n15565), .ZN(P2_U2863) );
  INV_X1 U18702 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n15571) );
  AOI21_X1 U18703 ( .B1(n15568), .B2(n15567), .A(n15566), .ZN(n15637) );
  NAND2_X1 U18704 ( .A1(n15637), .A2(n15575), .ZN(n15570) );
  NAND2_X1 U18705 ( .A1(n15965), .A2(n15572), .ZN(n15569) );
  OAI211_X1 U18706 ( .C1(n15572), .C2(n15571), .A(n15570), .B(n15569), .ZN(
        P2_U2864) );
  AOI21_X1 U18707 ( .B1(n15574), .B2(n15573), .A(n9738), .ZN(n15643) );
  NAND2_X1 U18708 ( .A1(n15643), .A2(n15575), .ZN(n15577) );
  NAND2_X1 U18709 ( .A1(n15578), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15576) );
  OAI211_X1 U18710 ( .C1(n16485), .C2(n15578), .A(n15577), .B(n15576), .ZN(
        P2_U2865) );
  OAI21_X1 U18711 ( .B1(n15579), .B2(n15580), .A(n15573), .ZN(n15656) );
  OR2_X1 U18712 ( .A1(n15590), .A2(n15581), .ZN(n15582) );
  NAND2_X1 U18713 ( .A1(n15482), .A2(n15582), .ZN(n19165) );
  MUX2_X1 U18714 ( .A(n19165), .B(n15583), .S(n15592), .Z(n15584) );
  OAI21_X1 U18715 ( .B1(n15656), .B2(n15594), .A(n15584), .ZN(P2_U2866) );
  NOR2_X1 U18716 ( .A1(n14368), .A2(n15585), .ZN(n15586) );
  OR2_X1 U18717 ( .A1(n15579), .A2(n15586), .ZN(n16480) );
  AND2_X1 U18718 ( .A1(n15588), .A2(n15587), .ZN(n15589) );
  NOR2_X1 U18719 ( .A1(n15590), .A2(n15589), .ZN(n19173) );
  INV_X1 U18720 ( .A(n19173), .ZN(n15797) );
  NOR2_X1 U18721 ( .A1(n15797), .A2(n15592), .ZN(n15591) );
  AOI21_X1 U18722 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n15592), .A(n15591), .ZN(
        n15593) );
  OAI21_X1 U18723 ( .B1(n16480), .B2(n15594), .A(n15593), .ZN(P2_U2867) );
  NAND3_X1 U18724 ( .A1(n15595), .A2(n15528), .A3(n19404), .ZN(n15600) );
  INV_X1 U18725 ( .A(n16447), .ZN(n15597) );
  INV_X1 U18726 ( .A(n19338), .ZN(n15619) );
  OAI22_X1 U18727 ( .A1(n15619), .A2(n19353), .B1(n19371), .B2(n19420), .ZN(
        n15596) );
  AOI21_X1 U18728 ( .B1(n19400), .B2(n15597), .A(n15596), .ZN(n15599) );
  AOI22_X1 U18729 ( .A1(n19340), .A2(BUF2_REG_29__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15598) );
  NAND3_X1 U18730 ( .A1(n15600), .A2(n15599), .A3(n15598), .ZN(P2_U2890) );
  AOI22_X1 U18731 ( .A1(n19340), .A2(BUF2_REG_28__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15602) );
  AOI22_X1 U18732 ( .A1(n19338), .A2(n19355), .B1(n19399), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15601) );
  OAI211_X1 U18733 ( .C1(n19342), .C2(n15899), .A(n15602), .B(n15601), .ZN(
        n15603) );
  INV_X1 U18734 ( .A(n15603), .ZN(n15604) );
  OAI21_X1 U18735 ( .B1(n15605), .B2(n16479), .A(n15604), .ZN(P2_U2891) );
  INV_X1 U18736 ( .A(n15909), .ZN(n15607) );
  OAI22_X1 U18737 ( .A1(n15619), .A2(n19358), .B1(n19371), .B2(n19423), .ZN(
        n15606) );
  AOI21_X1 U18738 ( .B1(n19400), .B2(n15607), .A(n15606), .ZN(n15609) );
  AOI22_X1 U18739 ( .A1(n19340), .A2(BUF2_REG_27__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15608) );
  OAI211_X1 U18740 ( .C1(n15610), .C2(n16479), .A(n15609), .B(n15608), .ZN(
        P2_U2892) );
  OAI21_X1 U18741 ( .B1(n9764), .B2(n15612), .A(n15611), .ZN(n16448) );
  AOI22_X1 U18742 ( .A1(n19340), .A2(BUF2_REG_26__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15614) );
  AOI22_X1 U18743 ( .A1(n19338), .A2(n19360), .B1(n19399), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15613) );
  OAI211_X1 U18744 ( .C1(n19342), .C2(n16448), .A(n15614), .B(n15613), .ZN(
        n15615) );
  AOI21_X1 U18745 ( .B1(n15616), .B2(n19404), .A(n15615), .ZN(n15617) );
  INV_X1 U18746 ( .A(n15617), .ZN(P2_U2893) );
  INV_X1 U18747 ( .A(n15618), .ZN(n15934) );
  OAI22_X1 U18748 ( .A1(n15619), .A2(n19363), .B1(n19371), .B2(n19427), .ZN(
        n15620) );
  AOI21_X1 U18749 ( .B1(n19400), .B2(n15934), .A(n15620), .ZN(n15622) );
  AOI22_X1 U18750 ( .A1(n19340), .A2(BUF2_REG_25__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15621) );
  OAI211_X1 U18751 ( .C1(n15623), .C2(n16479), .A(n15622), .B(n15621), .ZN(
        P2_U2894) );
  NAND2_X1 U18752 ( .A1(n15625), .A2(n15624), .ZN(n15626) );
  NAND2_X1 U18753 ( .A1(n15627), .A2(n15626), .ZN(n16467) );
  AOI22_X1 U18754 ( .A1(n19340), .A2(BUF2_REG_24__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15629) );
  AOI22_X1 U18755 ( .A1(n19338), .A2(n19366), .B1(n19399), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n15628) );
  OAI211_X1 U18756 ( .C1(n19342), .C2(n16467), .A(n15629), .B(n15628), .ZN(
        n15630) );
  INV_X1 U18757 ( .A(n15630), .ZN(n15631) );
  OAI21_X1 U18758 ( .B1(n15632), .B2(n16479), .A(n15631), .ZN(P2_U2895) );
  AOI22_X1 U18759 ( .A1(n19340), .A2(BUF2_REG_23__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15635) );
  INV_X1 U18760 ( .A(n19567), .ZN(n15633) );
  AOI22_X1 U18761 ( .A1(n19338), .A2(n15633), .B1(n19399), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15634) );
  OAI211_X1 U18762 ( .C1(n19342), .C2(n15963), .A(n15635), .B(n15634), .ZN(
        n15636) );
  AOI21_X1 U18763 ( .B1(n15637), .B2(n19404), .A(n15636), .ZN(n15638) );
  INV_X1 U18764 ( .A(n15638), .ZN(P2_U2896) );
  AOI22_X1 U18765 ( .A1(n19340), .A2(BUF2_REG_22__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15641) );
  INV_X1 U18766 ( .A(n19560), .ZN(n15639) );
  AOI22_X1 U18767 ( .A1(n19338), .A2(n15639), .B1(n19399), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15640) );
  OAI211_X1 U18768 ( .C1(n19342), .C2(n15978), .A(n15641), .B(n15640), .ZN(
        n15642) );
  AOI21_X1 U18769 ( .B1(n15643), .B2(n19404), .A(n15642), .ZN(n15644) );
  INV_X1 U18770 ( .A(n15644), .ZN(P2_U2897) );
  OR2_X1 U18771 ( .A1(n16001), .A2(n15645), .ZN(n15647) );
  AND2_X1 U18772 ( .A1(n15647), .A2(n15646), .ZN(n19163) );
  INV_X1 U18773 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19435) );
  INV_X1 U18774 ( .A(n19553), .ZN(n15648) );
  NAND2_X1 U18775 ( .A1(n19338), .A2(n15648), .ZN(n15649) );
  OAI21_X1 U18776 ( .B1(n19371), .B2(n19435), .A(n15649), .ZN(n15654) );
  INV_X1 U18777 ( .A(n19340), .ZN(n15652) );
  INV_X1 U18778 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15651) );
  INV_X1 U18779 ( .A(n19339), .ZN(n15650) );
  OAI22_X1 U18780 ( .A1(n15652), .A2(n15651), .B1(n15650), .B2(n16717), .ZN(
        n15653) );
  AOI211_X1 U18781 ( .C1(n19400), .C2(n19163), .A(n15654), .B(n15653), .ZN(
        n15655) );
  OAI21_X1 U18782 ( .B1(n15656), .B2(n16479), .A(n15655), .ZN(P2_U2898) );
  NOR2_X1 U18783 ( .A1(n15659), .A2(n15658), .ZN(n15660) );
  OR2_X1 U18784 ( .A1(n15657), .A2(n15660), .ZN(n19197) );
  AOI22_X1 U18785 ( .A1(n19340), .A2(BUF2_REG_19__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n15663) );
  INV_X1 U18786 ( .A(n19546), .ZN(n15661) );
  AOI22_X1 U18787 ( .A1(n19338), .A2(n15661), .B1(n19399), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15662) );
  OAI211_X1 U18788 ( .C1(n19342), .C2(n19197), .A(n15663), .B(n15662), .ZN(
        n15664) );
  AOI21_X1 U18789 ( .B1(n15665), .B2(n19404), .A(n15664), .ZN(n15666) );
  INV_X1 U18790 ( .A(n15666), .ZN(P2_U2900) );
  XNOR2_X1 U18791 ( .A(n15674), .B(n15667), .ZN(n19211) );
  AOI22_X1 U18792 ( .A1(n19340), .A2(BUF2_REG_18__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n15670) );
  INV_X1 U18793 ( .A(n19540), .ZN(n15668) );
  AOI22_X1 U18794 ( .A1(n19338), .A2(n15668), .B1(n19399), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15669) );
  OAI211_X1 U18795 ( .C1(n19211), .C2(n19342), .A(n15670), .B(n15669), .ZN(
        n15671) );
  AOI21_X1 U18796 ( .B1(n15672), .B2(n19404), .A(n15671), .ZN(n15673) );
  INV_X1 U18797 ( .A(n15673), .ZN(P2_U2901) );
  OAI21_X1 U18798 ( .B1(n15676), .B2(n15675), .A(n15674), .ZN(n19212) );
  AOI22_X1 U18799 ( .A1(n19340), .A2(BUF2_REG_17__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n15679) );
  AOI22_X1 U18800 ( .A1(n19338), .A2(n15677), .B1(n19399), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n15678) );
  OAI211_X1 U18801 ( .C1(n19342), .C2(n19212), .A(n15679), .B(n15678), .ZN(
        n15680) );
  AOI21_X1 U18802 ( .B1(n15681), .B2(n19404), .A(n15680), .ZN(n15682) );
  INV_X1 U18803 ( .A(n15682), .ZN(P2_U2902) );
  NAND2_X1 U18804 ( .A1(n15684), .A2(n15683), .ZN(n15689) );
  INV_X1 U18805 ( .A(n15685), .ZN(n15686) );
  NOR2_X1 U18806 ( .A1(n15687), .A2(n15686), .ZN(n15688) );
  XNOR2_X1 U18807 ( .A(n15689), .B(n15688), .ZN(n15892) );
  XNOR2_X1 U18808 ( .A(n15691), .B(n15690), .ZN(n15890) );
  INV_X1 U18809 ( .A(n15692), .ZN(n15695) );
  NAND2_X1 U18810 ( .A1(n19303), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15879) );
  OAI21_X1 U18811 ( .B1(n16541), .B2(n15693), .A(n15879), .ZN(n15694) );
  AOI21_X1 U18812 ( .B1(n15695), .B2(n16533), .A(n15694), .ZN(n15696) );
  OAI21_X1 U18813 ( .B1(n15888), .B2(n16526), .A(n15696), .ZN(n15697) );
  AOI21_X1 U18814 ( .B1(n15890), .B2(n16529), .A(n15697), .ZN(n15698) );
  OAI21_X1 U18815 ( .B1(n15892), .B2(n16537), .A(n15698), .ZN(P2_U2984) );
  INV_X1 U18816 ( .A(n15703), .ZN(n15896) );
  NAND2_X1 U18817 ( .A1(n15704), .A2(n16533), .ZN(n15705) );
  NAND2_X1 U18818 ( .A1(n19303), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15897) );
  OAI211_X1 U18819 ( .C1(n16541), .C2(n15706), .A(n15705), .B(n15897), .ZN(
        n15709) );
  OAI21_X1 U18820 ( .B1(n15713), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15707), .ZN(n15903) );
  NOR2_X1 U18821 ( .A1(n15903), .A2(n19490), .ZN(n15708) );
  AOI211_X2 U18822 ( .C1(n19486), .C2(n15896), .A(n15709), .B(n15708), .ZN(
        n15710) );
  OAI21_X1 U18823 ( .B1(n15906), .B2(n16537), .A(n15710), .ZN(P2_U2986) );
  XNOR2_X1 U18824 ( .A(n15711), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15918) );
  AOI21_X1 U18825 ( .B1(n15894), .B2(n15712), .A(n15713), .ZN(n15916) );
  NAND2_X1 U18826 ( .A1(n19303), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15908) );
  OAI21_X1 U18827 ( .B1(n16541), .B2(n15714), .A(n15908), .ZN(n15715) );
  AOI21_X1 U18828 ( .B1(n15716), .B2(n16533), .A(n15715), .ZN(n15717) );
  OAI21_X1 U18829 ( .B1(n15914), .B2(n16526), .A(n15717), .ZN(n15718) );
  AOI21_X1 U18830 ( .B1(n15916), .B2(n16529), .A(n15718), .ZN(n15719) );
  OAI21_X1 U18831 ( .B1(n15918), .B2(n16537), .A(n15719), .ZN(P2_U2987) );
  OAI21_X1 U18833 ( .B1(n9829), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15712), .ZN(n15931) );
  NOR2_X1 U18834 ( .A1(n15722), .A2(n19496), .ZN(n15725) );
  NAND2_X1 U18835 ( .A1(n19303), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15919) );
  OAI21_X1 U18836 ( .B1(n16541), .B2(n15723), .A(n15919), .ZN(n15724) );
  AOI211_X1 U18837 ( .C1(n16452), .C2(n19486), .A(n15725), .B(n15724), .ZN(
        n15730) );
  NAND2_X1 U18838 ( .A1(n15726), .A2(n15731), .ZN(n15728) );
  XNOR2_X1 U18839 ( .A(n15728), .B(n15727), .ZN(n15928) );
  NAND2_X1 U18840 ( .A1(n15928), .A2(n10990), .ZN(n15729) );
  OAI211_X1 U18841 ( .C1(n15931), .C2(n19490), .A(n15730), .B(n15729), .ZN(
        P2_U2988) );
  INV_X1 U18842 ( .A(n15731), .ZN(n15735) );
  AND2_X1 U18843 ( .A1(n15732), .A2(n15731), .ZN(n15733) );
  OAI22_X1 U18844 ( .A1(n15726), .A2(n15735), .B1(n15734), .B2(n15733), .ZN(
        n15945) );
  NAND2_X1 U18845 ( .A1(n9710), .A2(n15937), .ZN(n15932) );
  NAND3_X1 U18846 ( .A1(n15932), .A2(n16529), .A3(n15721), .ZN(n15741) );
  NAND2_X1 U18847 ( .A1(n19303), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15936) );
  OAI21_X1 U18848 ( .B1(n16541), .B2(n15736), .A(n15936), .ZN(n15738) );
  NOR2_X1 U18849 ( .A1(n15933), .A2(n16526), .ZN(n15737) );
  AOI211_X1 U18850 ( .C1(n16533), .C2(n15739), .A(n15738), .B(n15737), .ZN(
        n15740) );
  OAI211_X1 U18851 ( .C1(n15945), .C2(n16537), .A(n15741), .B(n15740), .ZN(
        P2_U2989) );
  OAI21_X1 U18852 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15742), .A(
        n9710), .ZN(n15957) );
  XNOR2_X1 U18853 ( .A(n15743), .B(n15947), .ZN(n15744) );
  XNOR2_X1 U18854 ( .A(n15745), .B(n15744), .ZN(n15955) );
  NOR2_X1 U18855 ( .A1(n15946), .A2(n16526), .ZN(n15749) );
  NAND2_X1 U18856 ( .A1(n19303), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15949) );
  NAND2_X1 U18857 ( .A1(n19484), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15746) );
  OAI211_X1 U18858 ( .C1(n15747), .C2(n19496), .A(n15949), .B(n15746), .ZN(
        n15748) );
  AOI211_X1 U18859 ( .C1(n15955), .C2(n10990), .A(n15749), .B(n15748), .ZN(
        n15750) );
  OAI21_X1 U18860 ( .B1(n15957), .B2(n19490), .A(n15750), .ZN(P2_U2990) );
  INV_X1 U18861 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15960) );
  INV_X1 U18863 ( .A(n15752), .ZN(n15753) );
  AOI21_X1 U18864 ( .B1(n15960), .B2(n15753), .A(n15742), .ZN(n15958) );
  NAND2_X1 U18865 ( .A1(n15958), .A2(n16529), .ZN(n15762) );
  OAI22_X1 U18866 ( .A1(n16541), .A2(n15754), .B1(n10770), .B2(n19277), .ZN(
        n15755) );
  AOI21_X1 U18867 ( .B1(n16533), .B2(n15756), .A(n15755), .ZN(n15761) );
  NOR2_X1 U18868 ( .A1(n15758), .A2(n15757), .ZN(n15966) );
  OR3_X1 U18869 ( .A1(n15967), .A2(n15966), .A3(n16537), .ZN(n15760) );
  NAND2_X1 U18870 ( .A1(n15965), .A2(n19486), .ZN(n15759) );
  NAND4_X1 U18871 ( .A1(n15762), .A2(n15761), .A3(n15760), .A4(n15759), .ZN(
        P2_U2991) );
  INV_X1 U18872 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16128) );
  INV_X1 U18873 ( .A(n16122), .ZN(n15764) );
  OAI21_X1 U18874 ( .B1(n15763), .B2(n16128), .A(n15764), .ZN(n15766) );
  NAND2_X1 U18875 ( .A1(n15763), .A2(n16128), .ZN(n15765) );
  AND2_X2 U18876 ( .A1(n15766), .A2(n15765), .ZN(n15848) );
  INV_X1 U18877 ( .A(n15846), .ZN(n15767) );
  AOI21_X2 U18878 ( .B1(n15848), .B2(n15847), .A(n15767), .ZN(n16086) );
  OR2_X2 U18879 ( .A1(n16086), .A2(n16084), .ZN(n15836) );
  INV_X1 U18880 ( .A(n15835), .ZN(n15768) );
  AOI21_X2 U18881 ( .B1(n15836), .B2(n15769), .A(n15768), .ZN(n15825) );
  NAND2_X1 U18882 ( .A1(n15825), .A2(n15824), .ZN(n15823) );
  INV_X1 U18883 ( .A(n15812), .ZN(n15770) );
  AOI21_X2 U18884 ( .B1(n15823), .B2(n15771), .A(n15770), .ZN(n16030) );
  AOI21_X1 U18885 ( .B1(n15788), .B2(n15773), .A(n15789), .ZN(n15777) );
  NAND2_X1 U18886 ( .A1(n15775), .A2(n15774), .ZN(n15776) );
  XNOR2_X1 U18887 ( .A(n15777), .B(n15776), .ZN(n15998) );
  NAND2_X1 U18888 ( .A1(n15780), .A2(n15781), .ZN(n15782) );
  AND2_X1 U18889 ( .A1(n15778), .A2(n15782), .ZN(n15996) );
  NOR2_X1 U18890 ( .A1(n20148), .A2(n19277), .ZN(n15992) );
  NOR2_X1 U18891 ( .A1(n16541), .A2(n10763), .ZN(n15783) );
  AOI211_X1 U18892 ( .C1(n19159), .C2(n16533), .A(n15992), .B(n15783), .ZN(
        n15784) );
  OAI21_X1 U18893 ( .B1(n19165), .B2(n16526), .A(n15784), .ZN(n15785) );
  AOI21_X1 U18894 ( .B1(n15996), .B2(n16529), .A(n15785), .ZN(n15786) );
  OAI21_X1 U18895 ( .B1(n15998), .B2(n16537), .A(n15786), .ZN(P2_U2993) );
  NAND2_X1 U18896 ( .A1(n15788), .A2(n15787), .ZN(n15792) );
  NAND2_X1 U18897 ( .A1(n10945), .A2(n15790), .ZN(n15791) );
  XNOR2_X1 U18898 ( .A(n15792), .B(n15791), .ZN(n16016) );
  AOI21_X1 U18899 ( .B1(n16010), .B2(n15793), .A(n10667), .ZN(n16013) );
  NAND2_X1 U18900 ( .A1(n19303), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n16003) );
  OAI21_X1 U18901 ( .B1(n19496), .B2(n15794), .A(n16003), .ZN(n15795) );
  AOI21_X1 U18902 ( .B1(n19484), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15795), .ZN(n15796) );
  OAI21_X1 U18903 ( .B1(n15797), .B2(n16526), .A(n15796), .ZN(n15798) );
  AOI21_X1 U18904 ( .B1(n16013), .B2(n16529), .A(n15798), .ZN(n15799) );
  OAI21_X1 U18905 ( .B1(n16016), .B2(n16537), .A(n15799), .ZN(P2_U2994) );
  OR2_X1 U18906 ( .A1(n15800), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15801) );
  NAND2_X1 U18907 ( .A1(n15793), .A2(n15801), .ZN(n16026) );
  NAND2_X1 U18908 ( .A1(n15803), .A2(n15802), .ZN(n15806) );
  INV_X1 U18909 ( .A(n16027), .ZN(n15804) );
  OAI21_X1 U18910 ( .B1(n16030), .B2(n15804), .A(n16028), .ZN(n15805) );
  XOR2_X1 U18911 ( .A(n15806), .B(n15805), .Z(n16017) );
  NAND2_X1 U18912 ( .A1(n16017), .A2(n10990), .ZN(n15810) );
  OAI22_X1 U18913 ( .A1(n16541), .A2(n19187), .B1(n10759), .B2(n19277), .ZN(
        n15808) );
  NOR2_X1 U18914 ( .A1(n19193), .A2(n16526), .ZN(n15807) );
  AOI211_X1 U18915 ( .C1(n16533), .C2(n19186), .A(n15808), .B(n15807), .ZN(
        n15809) );
  OAI211_X1 U18916 ( .C1(n19490), .C2(n16026), .A(n15810), .B(n15809), .ZN(
        P2_U2995) );
  NAND2_X1 U18917 ( .A1(n15812), .A2(n15811), .ZN(n15815) );
  NAND2_X1 U18918 ( .A1(n15823), .A2(n15813), .ZN(n15814) );
  XOR2_X1 U18919 ( .A(n15815), .B(n15814), .Z(n16060) );
  OR2_X1 U18920 ( .A1(n15816), .A2(n16055), .ZN(n16050) );
  XNOR2_X1 U18921 ( .A(n16050), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15821) );
  NAND2_X1 U18922 ( .A1(n19303), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16052) );
  OAI21_X1 U18923 ( .B1(n16541), .B2(n15817), .A(n16052), .ZN(n15818) );
  AOI21_X1 U18924 ( .B1(n19222), .B2(n16533), .A(n15818), .ZN(n15819) );
  OAI21_X1 U18925 ( .B1(n19213), .B2(n16526), .A(n15819), .ZN(n15820) );
  AOI21_X1 U18926 ( .B1(n15821), .B2(n16529), .A(n15820), .ZN(n15822) );
  OAI21_X1 U18927 ( .B1(n16060), .B2(n16537), .A(n15822), .ZN(P2_U2997) );
  OAI21_X1 U18928 ( .B1(n15825), .B2(n15824), .A(n15823), .ZN(n16070) );
  OAI22_X1 U18929 ( .A1(n15827), .A2(n16526), .B1(n15826), .B2(n16541), .ZN(
        n15830) );
  OAI22_X1 U18930 ( .A1(n20141), .A2(n19277), .B1(n19496), .B2(n15828), .ZN(
        n15829) );
  NOR2_X1 U18931 ( .A1(n15830), .A2(n15829), .ZN(n15833) );
  NOR2_X1 U18932 ( .A1(n15816), .A2(n16076), .ZN(n15831) );
  OAI211_X1 U18933 ( .C1(n15831), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16529), .B(n16050), .ZN(n15832) );
  OAI211_X1 U18934 ( .C1(n16070), .C2(n16537), .A(n15833), .B(n15832), .ZN(
        P2_U2998) );
  NAND2_X1 U18935 ( .A1(n15835), .A2(n15834), .ZN(n15838) );
  NAND2_X1 U18936 ( .A1(n15836), .A2(n16082), .ZN(n15837) );
  XOR2_X1 U18937 ( .A(n15838), .B(n15837), .Z(n16081) );
  XNOR2_X1 U18938 ( .A(n15816), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16079) );
  OAI22_X1 U18939 ( .A1(n16541), .A2(n15840), .B1(n19496), .B2(n15839), .ZN(
        n15844) );
  OAI22_X1 U18940 ( .A1(n15842), .A2(n16526), .B1(n15841), .B2(n19277), .ZN(
        n15843) );
  AOI211_X1 U18941 ( .C1(n16079), .C2(n16529), .A(n15844), .B(n15843), .ZN(
        n15845) );
  OAI21_X1 U18942 ( .B1(n16081), .B2(n16537), .A(n15845), .ZN(P2_U2999) );
  NAND2_X1 U18943 ( .A1(n15847), .A2(n15846), .ZN(n15849) );
  XOR2_X1 U18944 ( .A(n15849), .B(n15848), .Z(n16119) );
  NAND2_X1 U18945 ( .A1(n15850), .A2(n16138), .ZN(n16121) );
  INV_X1 U18946 ( .A(n16120), .ZN(n15852) );
  NAND2_X1 U18947 ( .A1(n16120), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16089) );
  INV_X1 U18948 ( .A(n16089), .ZN(n15851) );
  AOI21_X1 U18949 ( .B1(n15853), .B2(n15852), .A(n15851), .ZN(n16117) );
  OAI22_X1 U18950 ( .A1(n16541), .A2(n15854), .B1(n16109), .B2(n19277), .ZN(
        n15857) );
  INV_X1 U18951 ( .A(n19246), .ZN(n15855) );
  OAI22_X1 U18952 ( .A1(n16526), .A2(n16111), .B1(n19496), .B2(n15855), .ZN(
        n15856) );
  AOI211_X1 U18953 ( .C1(n16117), .C2(n16529), .A(n15857), .B(n15856), .ZN(
        n15858) );
  OAI21_X1 U18954 ( .B1(n16537), .B2(n16119), .A(n15858), .ZN(P2_U3001) );
  INV_X1 U18955 ( .A(n15850), .ZN(n15870) );
  OAI21_X1 U18956 ( .B1(n15870), .B2(n16156), .A(n16137), .ZN(n15859) );
  NAND2_X1 U18957 ( .A1(n15859), .A2(n16121), .ZN(n16145) );
  NAND2_X1 U18958 ( .A1(n15861), .A2(n15860), .ZN(n15863) );
  XOR2_X1 U18959 ( .A(n15863), .B(n15862), .Z(n16143) );
  OAI22_X1 U18960 ( .A1(n16541), .A2(n15864), .B1(n10738), .B2(n19277), .ZN(
        n15867) );
  OAI22_X1 U18961 ( .A1(n16526), .A2(n16135), .B1(n19496), .B2(n15865), .ZN(
        n15866) );
  AOI211_X1 U18962 ( .C1(n16143), .C2(n10990), .A(n15867), .B(n15866), .ZN(
        n15868) );
  OAI21_X1 U18963 ( .B1(n16145), .B2(n19490), .A(n15868), .ZN(P2_U3003) );
  OAI21_X1 U18964 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15869), .A(
        n15870), .ZN(n16176) );
  NAND2_X1 U18965 ( .A1(n16146), .A2(n16147), .ZN(n15873) );
  NAND2_X1 U18966 ( .A1(n15872), .A2(n15871), .ZN(n16149) );
  XOR2_X1 U18967 ( .A(n15873), .B(n16149), .Z(n16174) );
  INV_X1 U18968 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20132) );
  OAI22_X1 U18969 ( .A1(n16541), .A2(n19262), .B1(n20132), .B2(n19277), .ZN(
        n15874) );
  AOI21_X1 U18970 ( .B1(n16533), .B2(n19268), .A(n15874), .ZN(n15875) );
  OAI21_X1 U18971 ( .B1(n16526), .B2(n15876), .A(n15875), .ZN(n15877) );
  AOI21_X1 U18972 ( .B1(n16174), .B2(n10990), .A(n15877), .ZN(n15878) );
  OAI21_X1 U18973 ( .B1(n16176), .B2(n19490), .A(n15878), .ZN(P2_U3005) );
  OAI21_X1 U18974 ( .B1(n19508), .B2(n15880), .A(n15879), .ZN(n15881) );
  INV_X1 U18975 ( .A(n15881), .ZN(n15887) );
  OAI21_X1 U18976 ( .B1(n15883), .B2(n15882), .A(n15690), .ZN(n15885) );
  NAND2_X1 U18977 ( .A1(n15885), .A2(n15884), .ZN(n15886) );
  OAI211_X1 U18978 ( .C1(n15888), .C2(n16547), .A(n15887), .B(n15886), .ZN(
        n15889) );
  AOI21_X1 U18979 ( .B1(n15890), .B2(n16550), .A(n15889), .ZN(n15891) );
  OAI21_X1 U18980 ( .B1(n15892), .B2(n19502), .A(n15891), .ZN(P2_U3016) );
  INV_X1 U18981 ( .A(n15893), .ZN(n15895) );
  NOR3_X1 U18982 ( .A1(n15895), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15894), .ZN(n15901) );
  NAND2_X1 U18983 ( .A1(n15896), .A2(n19505), .ZN(n15898) );
  OAI211_X1 U18984 ( .C1(n19508), .C2(n15899), .A(n15898), .B(n15897), .ZN(
        n15900) );
  AOI211_X1 U18985 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15902), .A(
        n15901), .B(n15900), .ZN(n15905) );
  OR2_X1 U18986 ( .A1(n15903), .A2(n19515), .ZN(n15904) );
  OAI211_X1 U18987 ( .C1(n15906), .C2(n19502), .A(n15905), .B(n15904), .ZN(
        P2_U3018) );
  INV_X1 U18988 ( .A(n15907), .ZN(n15911) );
  OAI21_X1 U18989 ( .B1(n19508), .B2(n15909), .A(n15908), .ZN(n15910) );
  AOI21_X1 U18990 ( .B1(n15911), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15910), .ZN(n15913) );
  OAI211_X1 U18991 ( .C1(n15914), .C2(n16547), .A(n15913), .B(n15912), .ZN(
        n15915) );
  AOI21_X1 U18992 ( .B1(n15916), .B2(n16550), .A(n15915), .ZN(n15917) );
  OAI21_X1 U18993 ( .B1(n15918), .B2(n19502), .A(n15917), .ZN(P2_U3019) );
  NAND2_X1 U18994 ( .A1(n16452), .A2(n19505), .ZN(n15920) );
  OAI211_X1 U18995 ( .C1(n19508), .C2(n16448), .A(n15920), .B(n15919), .ZN(
        n15927) );
  INV_X1 U18996 ( .A(n15953), .ZN(n15921) );
  NAND3_X1 U18997 ( .A1(n15921), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15937), .ZN(n15939) );
  AOI21_X1 U18998 ( .B1(n15939), .B2(n15938), .A(n15922), .ZN(n15926) );
  INV_X1 U18999 ( .A(n15923), .ZN(n15924) );
  NOR3_X1 U19000 ( .A1(n15953), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15924), .ZN(n15925) );
  NOR3_X1 U19001 ( .A1(n15927), .A2(n15926), .A3(n15925), .ZN(n15930) );
  NAND2_X1 U19002 ( .A1(n15928), .A2(n16568), .ZN(n15929) );
  OAI211_X1 U19003 ( .C1(n15931), .C2(n19515), .A(n15930), .B(n15929), .ZN(
        P2_U3020) );
  NAND3_X1 U19004 ( .A1(n15932), .A2(n16550), .A3(n15721), .ZN(n15944) );
  INV_X1 U19005 ( .A(n15933), .ZN(n15942) );
  NAND2_X1 U19006 ( .A1(n16544), .A2(n15934), .ZN(n15935) );
  OAI211_X1 U19007 ( .C1(n15938), .C2(n15937), .A(n15936), .B(n15935), .ZN(
        n15941) );
  INV_X1 U19008 ( .A(n15939), .ZN(n15940) );
  AOI211_X1 U19009 ( .C1(n19505), .C2(n15942), .A(n15941), .B(n15940), .ZN(
        n15943) );
  OAI211_X1 U19010 ( .C1(n15945), .C2(n19502), .A(n15944), .B(n15943), .ZN(
        P2_U3021) );
  INV_X1 U19011 ( .A(n15946), .ZN(n16469) );
  NOR2_X1 U19012 ( .A1(n15948), .A2(n15947), .ZN(n15951) );
  OAI21_X1 U19013 ( .B1(n19508), .B2(n16467), .A(n15949), .ZN(n15950) );
  AOI211_X1 U19014 ( .C1(n16469), .C2(n19505), .A(n15951), .B(n15950), .ZN(
        n15952) );
  OAI21_X1 U19015 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15953), .A(
        n15952), .ZN(n15954) );
  AOI21_X1 U19016 ( .B1(n15955), .B2(n16568), .A(n15954), .ZN(n15956) );
  OAI21_X1 U19017 ( .B1(n15957), .B2(n19515), .A(n15956), .ZN(P2_U3022) );
  NAND2_X1 U19018 ( .A1(n15958), .A2(n16550), .ZN(n15972) );
  NOR2_X1 U19019 ( .A1(n15989), .A2(n15959), .ZN(n15988) );
  NAND2_X1 U19020 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15988), .ZN(
        n15979) );
  AOI221_X1 U19021 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C1(n15960), .C2(n15977), .A(
        n15979), .ZN(n15961) );
  AOI21_X1 U19022 ( .B1(n19303), .B2(P2_REIP_REG_23__SCAN_IN), .A(n15961), 
        .ZN(n15962) );
  OAI21_X1 U19023 ( .B1(n19508), .B2(n15963), .A(n15962), .ZN(n15964) );
  AOI21_X1 U19024 ( .B1(n15965), .B2(n19505), .A(n15964), .ZN(n15971) );
  OR3_X1 U19025 ( .A1(n15967), .A2(n15966), .A3(n19502), .ZN(n15970) );
  OAI21_X1 U19026 ( .B1(n16093), .B2(n15968), .A(n16172), .ZN(n15985) );
  NAND2_X1 U19027 ( .A1(n15985), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15969) );
  NAND4_X1 U19028 ( .A1(n15972), .A2(n15971), .A3(n15970), .A4(n15969), .ZN(
        P2_U3023) );
  NAND2_X1 U19029 ( .A1(n15974), .A2(n15973), .ZN(n15976) );
  XOR2_X1 U19030 ( .A(n15976), .B(n15975), .Z(n16486) );
  AOI21_X1 U19031 ( .B1(n15977), .B2(n15778), .A(n15752), .ZN(n16488) );
  NAND2_X1 U19032 ( .A1(n16488), .A2(n16550), .ZN(n15987) );
  INV_X1 U19033 ( .A(n15978), .ZN(n15982) );
  NOR2_X1 U19034 ( .A1(n10767), .A2(n19277), .ZN(n15981) );
  NOR2_X1 U19035 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15979), .ZN(
        n15980) );
  AOI211_X1 U19036 ( .C1(n16544), .C2(n15982), .A(n15981), .B(n15980), .ZN(
        n15983) );
  OAI21_X1 U19037 ( .B1(n16485), .B2(n16547), .A(n15983), .ZN(n15984) );
  AOI21_X1 U19038 ( .B1(n15985), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15984), .ZN(n15986) );
  OAI211_X1 U19039 ( .C1(n16486), .C2(n19502), .A(n15987), .B(n15986), .ZN(
        P2_U3024) );
  NAND2_X1 U19040 ( .A1(n15988), .A2(n15781), .ZN(n15994) );
  INV_X1 U19041 ( .A(n16172), .ZN(n16092) );
  AOI21_X1 U19042 ( .B1(n15989), .B2(n19499), .A(n16092), .ZN(n15990) );
  NOR2_X1 U19043 ( .A1(n15990), .A2(n15781), .ZN(n15991) );
  AOI211_X1 U19044 ( .C1(n16544), .C2(n19163), .A(n15992), .B(n15991), .ZN(
        n15993) );
  OAI211_X1 U19045 ( .C1(n19165), .C2(n16547), .A(n15994), .B(n15993), .ZN(
        n15995) );
  AOI21_X1 U19046 ( .B1(n15996), .B2(n16550), .A(n15995), .ZN(n15997) );
  OAI21_X1 U19047 ( .B1(n15998), .B2(n19502), .A(n15997), .ZN(P2_U3025) );
  NOR2_X1 U19048 ( .A1(n15657), .A2(n15999), .ZN(n16000) );
  OR2_X1 U19049 ( .A1(n16001), .A2(n16000), .ZN(n19171) );
  NAND2_X1 U19050 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16164), .ZN(
        n16157) );
  INV_X1 U19051 ( .A(n16157), .ZN(n16090) );
  NAND2_X1 U19052 ( .A1(n16002), .A2(n16090), .ZN(n16071) );
  INV_X1 U19053 ( .A(n16071), .ZN(n16054) );
  NAND4_X1 U19054 ( .A1(n16054), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n10154), .A4(n16010), .ZN(n16004) );
  OAI211_X1 U19055 ( .C1(n19508), .C2(n19171), .A(n16004), .B(n16003), .ZN(
        n16012) );
  NAND2_X1 U19056 ( .A1(n19499), .A2(n16005), .ZN(n16006) );
  AND2_X1 U19057 ( .A1(n16172), .A2(n16006), .ZN(n16077) );
  NAND2_X1 U19058 ( .A1(n19499), .A2(n16008), .ZN(n16007) );
  AND2_X1 U19059 ( .A1(n16077), .A2(n16007), .ZN(n16041) );
  NOR2_X1 U19060 ( .A1(n16008), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16009) );
  NAND2_X1 U19061 ( .A1(n16054), .A2(n16009), .ZN(n16018) );
  AOI21_X1 U19062 ( .B1(n16041), .B2(n16018), .A(n16010), .ZN(n16011) );
  AOI211_X1 U19063 ( .C1(n19505), .C2(n19173), .A(n16012), .B(n16011), .ZN(
        n16015) );
  NAND2_X1 U19064 ( .A1(n16013), .A2(n16550), .ZN(n16014) );
  OAI211_X1 U19065 ( .C1(n16016), .C2(n19502), .A(n16015), .B(n16014), .ZN(
        P2_U3026) );
  NAND2_X1 U19066 ( .A1(n16017), .A2(n16568), .ZN(n16025) );
  INV_X1 U19067 ( .A(n16041), .ZN(n16023) );
  INV_X1 U19068 ( .A(n16018), .ZN(n16019) );
  AOI21_X1 U19069 ( .B1(n19303), .B2(P2_REIP_REG_19__SCAN_IN), .A(n16019), 
        .ZN(n16020) );
  OAI21_X1 U19070 ( .B1(n19508), .B2(n19197), .A(n16020), .ZN(n16022) );
  NOR2_X1 U19071 ( .A1(n19193), .A2(n16547), .ZN(n16021) );
  AOI211_X1 U19072 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16023), .A(
        n16022), .B(n16021), .ZN(n16024) );
  OAI211_X1 U19073 ( .C1(n16026), .C2(n19515), .A(n16025), .B(n16024), .ZN(
        P2_U3027) );
  NAND2_X1 U19074 ( .A1(n16028), .A2(n16027), .ZN(n16029) );
  XNOR2_X1 U19075 ( .A(n16030), .B(n16029), .ZN(n16493) );
  INV_X1 U19076 ( .A(n16493), .ZN(n16044) );
  INV_X1 U19077 ( .A(n15800), .ZN(n16032) );
  OAI21_X1 U19078 ( .B1(n16050), .B2(n16033), .A(n16040), .ZN(n16031) );
  NOR2_X1 U19079 ( .A1(n10756), .A2(n19277), .ZN(n16036) );
  NOR3_X1 U19080 ( .A1(n16033), .A2(n16055), .A3(n16071), .ZN(n16034) );
  AND2_X1 U19081 ( .A1(n16040), .A2(n16034), .ZN(n16035) );
  NOR2_X1 U19082 ( .A1(n16036), .A2(n16035), .ZN(n16037) );
  OAI21_X1 U19083 ( .B1(n19508), .B2(n19211), .A(n16037), .ZN(n16038) );
  AOI21_X1 U19084 ( .B1(n19205), .B2(n19505), .A(n16038), .ZN(n16039) );
  OAI21_X1 U19085 ( .B1(n16041), .B2(n16040), .A(n16039), .ZN(n16042) );
  AOI21_X1 U19086 ( .B1(n16492), .B2(n16550), .A(n16042), .ZN(n16043) );
  OAI21_X1 U19087 ( .B1(n16044), .B2(n19502), .A(n16043), .ZN(P2_U3028) );
  OR2_X1 U19088 ( .A1(n16045), .A2(n16550), .ZN(n16049) );
  NAND2_X1 U19089 ( .A1(n16046), .A2(n16076), .ZN(n16047) );
  NAND2_X1 U19090 ( .A1(n16077), .A2(n16047), .ZN(n16048) );
  AOI21_X1 U19091 ( .B1(n16050), .B2(n16049), .A(n16048), .ZN(n16067) );
  OAI21_X1 U19092 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16093), .A(
        n16067), .ZN(n16058) );
  INV_X1 U19093 ( .A(n19213), .ZN(n16051) );
  NAND2_X1 U19094 ( .A1(n16051), .A2(n19505), .ZN(n16053) );
  OAI211_X1 U19095 ( .C1(n19508), .C2(n19212), .A(n16053), .B(n16052), .ZN(
        n16057) );
  INV_X1 U19096 ( .A(n15816), .ZN(n16087) );
  AOI21_X1 U19097 ( .B1(n16087), .B2(n16550), .A(n16054), .ZN(n16063) );
  NOR3_X1 U19098 ( .A1(n16063), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n16055), .ZN(n16056) );
  AOI211_X1 U19099 ( .C1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n16058), .A(
        n16057), .B(n16056), .ZN(n16059) );
  OAI21_X1 U19100 ( .B1(n16060), .B2(n19502), .A(n16059), .ZN(P2_U3029) );
  INV_X1 U19101 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16066) );
  OAI22_X1 U19102 ( .A1(n19508), .A2(n19341), .B1(n20141), .B2(n19277), .ZN(
        n16061) );
  AOI21_X1 U19103 ( .B1(n16062), .B2(n19505), .A(n16061), .ZN(n16065) );
  OR3_X1 U19104 ( .A1(n16063), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n16076), .ZN(n16064) );
  OAI211_X1 U19105 ( .C1(n16067), .C2(n16066), .A(n16065), .B(n16064), .ZN(
        n16068) );
  INV_X1 U19106 ( .A(n16068), .ZN(n16069) );
  OAI21_X1 U19107 ( .B1(n16070), .B2(n19502), .A(n16069), .ZN(P2_U3030) );
  NOR2_X1 U19108 ( .A1(n19508), .A2(n19349), .ZN(n16073) );
  OAI22_X1 U19109 ( .A1(n19277), .A2(n15841), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16071), .ZN(n16072) );
  AOI211_X1 U19110 ( .C1(n16074), .C2(n19505), .A(n16073), .B(n16072), .ZN(
        n16075) );
  OAI21_X1 U19111 ( .B1(n16077), .B2(n16076), .A(n16075), .ZN(n16078) );
  AOI21_X1 U19112 ( .B1(n16079), .B2(n16550), .A(n16078), .ZN(n16080) );
  OAI21_X1 U19113 ( .B1(n16081), .B2(n19502), .A(n16080), .ZN(P2_U3031) );
  INV_X1 U19114 ( .A(n16082), .ZN(n16083) );
  NOR2_X1 U19115 ( .A1(n16084), .A2(n16083), .ZN(n16085) );
  XNOR2_X1 U19116 ( .A(n16086), .B(n16085), .ZN(n16499) );
  INV_X1 U19117 ( .A(n16499), .ZN(n16105) );
  INV_X1 U19118 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16088) );
  AOI21_X1 U19119 ( .B1(n16089), .B2(n16088), .A(n16087), .ZN(n16498) );
  NAND2_X1 U19120 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16094) );
  NAND2_X1 U19121 ( .A1(n16138), .A2(n16090), .ZN(n16091) );
  NOR2_X1 U19122 ( .A1(n16094), .A2(n16091), .ZN(n16096) );
  INV_X1 U19123 ( .A(n16091), .ZN(n16129) );
  AOI21_X1 U19124 ( .B1(n16171), .B2(n19499), .A(n16092), .ZN(n16155) );
  OAI21_X1 U19125 ( .B1(n16138), .B2(n16093), .A(n16155), .ZN(n16127) );
  AOI21_X1 U19126 ( .B1(n16129), .B2(n16094), .A(n16127), .ZN(n16115) );
  INV_X1 U19127 ( .A(n16115), .ZN(n16095) );
  MUX2_X1 U19128 ( .A(n16096), .B(n16095), .S(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n16103) );
  NOR2_X1 U19129 ( .A1(n16098), .A2(n16097), .ZN(n16100) );
  NOR2_X1 U19130 ( .A1(n16100), .A2(n16099), .ZN(n19231) );
  AOI22_X1 U19131 ( .A1(n16544), .A2(n19231), .B1(n19303), .B2(
        P2_REIP_REG_14__SCAN_IN), .ZN(n16101) );
  OAI21_X1 U19132 ( .B1(n16547), .B2(n19232), .A(n16101), .ZN(n16102) );
  AOI211_X1 U19133 ( .C1(n16498), .C2(n16550), .A(n16103), .B(n16102), .ZN(
        n16104) );
  OAI21_X1 U19134 ( .B1(n16105), .B2(n19502), .A(n16104), .ZN(P2_U3032) );
  AOI21_X1 U19135 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16129), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16114) );
  INV_X1 U19136 ( .A(n16097), .ZN(n16106) );
  OAI21_X1 U19137 ( .B1(n16108), .B2(n16107), .A(n16106), .ZN(n19354) );
  OAI22_X1 U19138 ( .A1(n19508), .A2(n19354), .B1(n16109), .B2(n19277), .ZN(
        n16110) );
  INV_X1 U19139 ( .A(n16110), .ZN(n16113) );
  INV_X1 U19140 ( .A(n16111), .ZN(n19247) );
  NAND2_X1 U19141 ( .A1(n19505), .A2(n19247), .ZN(n16112) );
  OAI211_X1 U19142 ( .C1(n16115), .C2(n16114), .A(n16113), .B(n16112), .ZN(
        n16116) );
  AOI21_X1 U19143 ( .B1(n16117), .B2(n16550), .A(n16116), .ZN(n16118) );
  OAI21_X1 U19144 ( .B1(n19502), .B2(n16119), .A(n16118), .ZN(P2_U3033) );
  AOI21_X1 U19145 ( .B1(n16128), .B2(n16121), .A(n16120), .ZN(n16506) );
  INV_X1 U19146 ( .A(n16506), .ZN(n16134) );
  XNOR2_X1 U19147 ( .A(n16122), .B(n16128), .ZN(n16123) );
  XNOR2_X1 U19148 ( .A(n15763), .B(n16123), .ZN(n16505) );
  XNOR2_X1 U19149 ( .A(n16125), .B(n16124), .ZN(n19357) );
  INV_X1 U19150 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20136) );
  NOR2_X1 U19151 ( .A1(n20136), .A2(n19277), .ZN(n16126) );
  AOI221_X1 U19152 ( .B1(n16129), .B2(n16128), .C1(n16127), .C2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n16126), .ZN(n16131) );
  NAND2_X1 U19153 ( .A1(n19505), .A2(n16504), .ZN(n16130) );
  OAI211_X1 U19154 ( .C1(n19357), .C2(n19508), .A(n16131), .B(n16130), .ZN(
        n16132) );
  AOI21_X1 U19155 ( .B1(n16505), .B2(n16568), .A(n16132), .ZN(n16133) );
  OAI21_X1 U19156 ( .B1(n16134), .B2(n19515), .A(n16133), .ZN(P2_U3034) );
  INV_X1 U19157 ( .A(n16135), .ZN(n16136) );
  AOI22_X1 U19158 ( .A1(n19505), .A2(n16136), .B1(n19303), .B2(
        P2_REIP_REG_11__SCAN_IN), .ZN(n16141) );
  OAI22_X1 U19159 ( .A1(n16138), .A2(n16157), .B1(n16155), .B2(n16137), .ZN(
        n16139) );
  OAI21_X1 U19160 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16139), .ZN(n16140) );
  OAI211_X1 U19161 ( .C1(n19359), .C2(n19508), .A(n16141), .B(n16140), .ZN(
        n16142) );
  AOI21_X1 U19162 ( .B1(n16143), .B2(n16568), .A(n16142), .ZN(n16144) );
  OAI21_X1 U19163 ( .B1(n16145), .B2(n19515), .A(n16144), .ZN(P2_U3035) );
  XNOR2_X1 U19164 ( .A(n15850), .B(n16156), .ZN(n16509) );
  INV_X1 U19165 ( .A(n16509), .ZN(n16163) );
  INV_X1 U19166 ( .A(n16146), .ZN(n16148) );
  OAI21_X1 U19167 ( .B1(n16149), .B2(n16148), .A(n16147), .ZN(n16153) );
  NAND2_X1 U19168 ( .A1(n16151), .A2(n16150), .ZN(n16152) );
  XNOR2_X1 U19169 ( .A(n16153), .B(n16152), .ZN(n16511) );
  NAND2_X1 U19170 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19303), .ZN(n16154) );
  OAI221_X1 U19171 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16157), 
        .C1(n16156), .C2(n16155), .A(n16154), .ZN(n16161) );
  INV_X1 U19172 ( .A(n16510), .ZN(n16159) );
  INV_X1 U19173 ( .A(n16158), .ZN(n19362) );
  OAI22_X1 U19174 ( .A1(n16547), .A2(n16159), .B1(n19508), .B2(n19362), .ZN(
        n16160) );
  AOI211_X1 U19175 ( .C1(n16511), .C2(n16568), .A(n16161), .B(n16160), .ZN(
        n16162) );
  OAI21_X1 U19176 ( .B1(n16163), .B2(n19515), .A(n16162), .ZN(P2_U3036) );
  NAND2_X1 U19177 ( .A1(n16164), .A2(n16171), .ZN(n16170) );
  OAI21_X1 U19178 ( .B1(n16167), .B2(n16166), .A(n16165), .ZN(n19364) );
  OAI22_X1 U19179 ( .A1(n19508), .A2(n19364), .B1(n20132), .B2(n19277), .ZN(
        n16168) );
  AOI21_X1 U19180 ( .B1(n19505), .B2(n19269), .A(n16168), .ZN(n16169) );
  OAI211_X1 U19181 ( .C1(n16172), .C2(n16171), .A(n16170), .B(n16169), .ZN(
        n16173) );
  AOI21_X1 U19182 ( .B1(n16174), .B2(n16568), .A(n16173), .ZN(n16175) );
  OAI21_X1 U19183 ( .B1(n16176), .B2(n19515), .A(n16175), .ZN(P2_U3037) );
  AOI22_X1 U19184 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16180) );
  AOI22_X1 U19185 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9689), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16179) );
  AOI22_X1 U19186 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16178) );
  AOI22_X1 U19187 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16177) );
  NAND4_X1 U19188 ( .A1(n16180), .A2(n16179), .A3(n16178), .A4(n16177), .ZN(
        n16187) );
  AOI22_X1 U19189 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16185) );
  AOI22_X1 U19190 ( .A1(n17423), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16184) );
  AOI22_X1 U19191 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16183) );
  AOI22_X1 U19192 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16182) );
  NAND4_X1 U19193 ( .A1(n16185), .A2(n16184), .A3(n16183), .A4(n16182), .ZN(
        n16186) );
  NOR2_X1 U19194 ( .A1(n16187), .A2(n16186), .ZN(n17584) );
  INV_X1 U19195 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17043) );
  AOI21_X1 U19196 ( .B1(n17470), .B2(n17403), .A(n17043), .ZN(n17391) );
  OAI22_X1 U19197 ( .A1(n17482), .A2(n17391), .B1(P3_EBX_REG_13__SCAN_IN), 
        .B2(n17484), .ZN(n17375) );
  OAI21_X1 U19198 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17391), .A(n17375), .ZN(
        n16188) );
  OAI21_X1 U19199 ( .B1(n17584), .B2(n17470), .A(n16188), .ZN(P3_U2690) );
  NAND2_X1 U19200 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18362) );
  NOR2_X1 U19201 ( .A1(n18360), .A2(n18362), .ZN(n18234) );
  NAND3_X1 U19202 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18233) );
  NAND2_X1 U19203 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18406) );
  NOR2_X1 U19204 ( .A1(n18233), .A2(n18406), .ZN(n18355) );
  NAND2_X1 U19205 ( .A1(n18234), .A2(n18355), .ZN(n18281) );
  NOR2_X1 U19206 ( .A1(n16189), .A2(n18281), .ZN(n18186) );
  NAND2_X1 U19207 ( .A1(n18178), .A2(n18186), .ZN(n18132) );
  AOI21_X1 U19208 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18428) );
  NOR2_X1 U19209 ( .A1(n18428), .A2(n18233), .ZN(n18356) );
  NAND2_X1 U19210 ( .A1(n18356), .A2(n18234), .ZN(n18256) );
  NOR3_X1 U19211 ( .A1(n18242), .A2(n16189), .A3(n18256), .ZN(n18240) );
  NAND2_X1 U19212 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18240), .ZN(
        n18188) );
  NOR2_X1 U19213 ( .A1(n16190), .A2(n18188), .ZN(n16202) );
  INV_X1 U19214 ( .A(n16202), .ZN(n18172) );
  OAI22_X1 U19215 ( .A1(n18937), .A2(n18132), .B1(n18924), .B2(n18172), .ZN(
        n16191) );
  NOR2_X1 U19216 ( .A1(n19091), .A2(n18281), .ZN(n18347) );
  NAND2_X1 U19217 ( .A1(n18237), .A2(n18347), .ZN(n18257) );
  OR2_X1 U19218 ( .A1(n18204), .A2(n18257), .ZN(n18205) );
  NOR2_X1 U19219 ( .A1(n16190), .A2(n18205), .ZN(n18191) );
  OAI221_X1 U19220 ( .B1(n16191), .B2(n18191), .C1(n16191), .C2(n9660), .A(
        n18133), .ZN(n18152) );
  NOR2_X1 U19221 ( .A1(n16203), .A2(n18152), .ZN(n16666) );
  AOI22_X1 U19222 ( .A1(n18906), .A2(n18131), .B1(n18139), .B2(n18323), .ZN(
        n16192) );
  INV_X1 U19223 ( .A(n16192), .ZN(n16201) );
  OAI21_X1 U19224 ( .B1(n16824), .B2(n16193), .A(n19113), .ZN(n16791) );
  NOR2_X1 U19225 ( .A1(n16786), .A2(n16791), .ZN(n16197) );
  AND4_X1 U19226 ( .A1(n16828), .A2(n16194), .A3(n18911), .A4(n18485), .ZN(
        n16196) );
  AOI211_X1 U19227 ( .C1(n16197), .C2(n16200), .A(n16196), .B(n16195), .ZN(
        n16199) );
  AOI221_X4 U19228 ( .B1(n16200), .B2(n16199), .C1(n16198), .C2(n16199), .A(
        n18967), .ZN(n18451) );
  OAI211_X1 U19229 ( .C1(n16666), .C2(n16201), .A(n18451), .B(n16252), .ZN(
        n16258) );
  NOR2_X1 U19230 ( .A1(n9803), .A2(n18433), .ZN(n18446) );
  INV_X1 U19231 ( .A(n18337), .ZN(n16206) );
  NOR3_X1 U19232 ( .A1(n18140), .A2(n18257), .A3(n16680), .ZN(n16205) );
  AOI21_X1 U19233 ( .B1(n16202), .B2(n18133), .A(n18924), .ZN(n18154) );
  AOI21_X1 U19234 ( .B1(n18933), .B2(n16203), .A(n18154), .ZN(n18134) );
  INV_X1 U19235 ( .A(n18186), .ZN(n18238) );
  OAI21_X1 U19236 ( .B1(n16680), .B2(n18238), .A(n18921), .ZN(n16204) );
  OAI211_X1 U19237 ( .C1(n18330), .C2(n16205), .A(n18134), .B(n16204), .ZN(
        n16253) );
  AOI211_X1 U19238 ( .C1(n16206), .C2(n18140), .A(n18433), .B(n16253), .ZN(
        n16689) );
  NAND2_X1 U19239 ( .A1(n18906), .A2(n18451), .ZN(n18457) );
  INV_X1 U19240 ( .A(n18457), .ZN(n18443) );
  NAND2_X1 U19241 ( .A1(n18451), .A2(n18323), .ZN(n18165) );
  INV_X1 U19242 ( .A(n18165), .ZN(n18368) );
  AOI22_X1 U19243 ( .A1(n18443), .A2(n16207), .B1(n18368), .B2(n16646), .ZN(
        n16254) );
  OAI21_X1 U19244 ( .B1(n18385), .B2(n16689), .A(n16254), .ZN(n16208) );
  AOI21_X1 U19245 ( .B1(n18446), .B2(n17755), .A(n16208), .ZN(n16210) );
  NOR3_X2 U19246 ( .A1(n18912), .A2(n18433), .A3(n17605), .ZN(n18367) );
  OAI221_X1 U19247 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16258), 
        .C1(n12306), .C2(n16210), .A(n16209), .ZN(P3_U2833) );
  INV_X1 U19248 ( .A(n16211), .ZN(n16214) );
  INV_X1 U19249 ( .A(n16212), .ZN(n16213) );
  OAI211_X1 U19250 ( .C1(n16215), .C2(n16214), .A(n16213), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n16219) );
  INV_X1 U19251 ( .A(n16216), .ZN(n16218) );
  OAI211_X1 U19252 ( .C1(n20722), .C2(n16219), .A(n16218), .B(n16217), .ZN(
        n16221) );
  NAND2_X1 U19253 ( .A1(n16219), .A2(n20722), .ZN(n16220) );
  NAND2_X1 U19254 ( .A1(n16221), .A2(n16220), .ZN(n16222) );
  AOI222_X1 U19255 ( .A1(n16223), .A2(n20787), .B1(n16223), .B2(n16222), .C1(
        n20787), .C2(n16222), .ZN(n16224) );
  AOI222_X1 U19256 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16225), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16224), .C1(n16225), 
        .C2(n16224), .ZN(n16233) );
  OAI21_X1 U19257 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n16226), .ZN(n16227) );
  NAND4_X1 U19258 ( .A1(n16230), .A2(n16229), .A3(n16228), .A4(n16227), .ZN(
        n16231) );
  AOI211_X1 U19259 ( .C1(n16233), .C2(n20418), .A(n16232), .B(n16231), .ZN(
        n16234) );
  INV_X1 U19260 ( .A(n16234), .ZN(n16242) );
  NAND2_X1 U19261 ( .A1(n16235), .A2(n20852), .ZN(n21052) );
  NOR3_X1 U19262 ( .A1(n16236), .A2(n12149), .A3(n21052), .ZN(n16240) );
  INV_X1 U19263 ( .A(n16237), .ZN(n16238) );
  AOI21_X1 U19264 ( .B1(n20976), .B2(n16238), .A(n16243), .ZN(n16239) );
  OR2_X1 U19265 ( .A1(n16240), .A2(n16239), .ZN(n16426) );
  AOI221_X1 U19266 ( .B1(n20963), .B2(n20962), .C1(n16242), .C2(n20962), .A(
        n16426), .ZN(n16431) );
  AOI21_X1 U19267 ( .B1(n16243), .B2(n16242), .A(n16241), .ZN(n16245) );
  OAI211_X1 U19268 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21050), .A(n16245), 
        .B(n16244), .ZN(n16246) );
  NOR2_X1 U19269 ( .A1(n16431), .A2(n16246), .ZN(n16250) );
  NAND2_X1 U19270 ( .A1(n21054), .A2(n16247), .ZN(n16248) );
  NAND2_X1 U19271 ( .A1(n20963), .A2(n16248), .ZN(n16249) );
  OAI22_X1 U19272 ( .A1(n16250), .A2(n20963), .B1(n16431), .B2(n16249), .ZN(
        P1_U3161) );
  INV_X1 U19273 ( .A(n16251), .ZN(n16259) );
  OR2_X1 U19274 ( .A1(n18445), .A2(n18446), .ZN(n18408) );
  NAND3_X1 U19275 ( .A1(n16252), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n18451), .ZN(n16665) );
  AOI22_X1 U19276 ( .A1(n18451), .A2(n16253), .B1(n18408), .B2(n16665), .ZN(
        n16670) );
  AOI21_X1 U19277 ( .B1(n16670), .B2(n16254), .A(n16628), .ZN(n16255) );
  AOI21_X1 U19278 ( .B1(n18367), .B2(n9726), .A(n16255), .ZN(n16257) );
  OAI211_X1 U19279 ( .C1(n16259), .C2(n16258), .A(n16257), .B(n16256), .ZN(
        P3_U2832) );
  NAND2_X1 U19280 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20973) );
  INV_X1 U19281 ( .A(n20973), .ZN(n16260) );
  INV_X1 U19282 ( .A(HOLD), .ZN(n20110) );
  NOR2_X1 U19283 ( .A1(n16263), .A2(n20110), .ZN(n20971) );
  INV_X1 U19284 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20982) );
  OAI22_X1 U19285 ( .A1(n16260), .A2(n20971), .B1(n20982), .B2(n20110), .ZN(
        n16261) );
  OAI211_X1 U19286 ( .C1(n21050), .C2(n16263), .A(n16262), .B(n16261), .ZN(
        P1_U3195) );
  AND2_X1 U19287 ( .A1(n16264), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U19288 ( .A1(n20114), .A2(n16267), .ZN(n20096) );
  AOI211_X1 U19289 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n16267), .A(
        P2_STATE2_REG_2__SCAN_IN), .B(n20096), .ZN(n16265) );
  NOR3_X1 U19290 ( .A1(n16617), .A2(n16610), .A3(n16265), .ZN(P2_U3178) );
  INV_X1 U19291 ( .A(n16610), .ZN(n16624) );
  NOR2_X1 U19292 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16617), .ZN(n20225) );
  AOI21_X4 U19293 ( .B1(n9681), .B2(n16616), .A(n16266), .ZN(n19956) );
  OAI221_X1 U19294 ( .B1(n10688), .B2(n16624), .C1(n20217), .C2(n16624), .A(
        n19956), .ZN(n20207) );
  NOR2_X1 U19295 ( .A1(n16268), .A2(n20207), .ZN(P2_U3047) );
  NOR3_X1 U19296 ( .A1(n16269), .A2(n17642), .A3(n16828), .ZN(n16270) );
  INV_X1 U19297 ( .A(n17487), .ZN(n16272) );
  INV_X1 U19298 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18471) );
  INV_X1 U19299 ( .A(n18124), .ZN(n16274) );
  NOR2_X1 U19300 ( .A1(n17597), .A2(n17487), .ZN(n17490) );
  NAND2_X1 U19301 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17490), .ZN(n17639) );
  NAND2_X1 U19302 ( .A1(n17622), .A2(n17639), .ZN(n17638) );
  NOR2_X1 U19303 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17490), .ZN(n16273) );
  OAI222_X1 U19304 ( .A1(n17633), .A2(n18471), .B1(n17630), .B2(n16274), .C1(
        n17638), .C2(n16273), .ZN(P3_U2735) );
  AOI21_X1 U19305 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n16275), .A(
        P1_REIP_REG_17__SCAN_IN), .ZN(n16283) );
  INV_X1 U19306 ( .A(n16276), .ZN(n16282) );
  OAI22_X1 U19307 ( .A1(n20308), .A2(n21212), .B1(n20279), .B2(n16277), .ZN(
        n16278) );
  AOI211_X1 U19308 ( .C1(n20339), .C2(n16279), .A(n20310), .B(n16278), .ZN(
        n16281) );
  AOI22_X1 U19309 ( .A1(n16307), .A2(n20317), .B1(n20334), .B2(n16306), .ZN(
        n16280) );
  OAI211_X1 U19310 ( .C1(n16283), .C2(n16282), .A(n16281), .B(n16280), .ZN(
        P1_U2823) );
  INV_X1 U19311 ( .A(n16284), .ZN(n16289) );
  INV_X1 U19312 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16285) );
  OAI21_X1 U19313 ( .B1(n20279), .B2(n16285), .A(n20322), .ZN(n16287) );
  AOI211_X1 U19314 ( .C1(n20335), .C2(P1_EBX_REG_15__SCAN_IN), .A(n16287), .B(
        n16286), .ZN(n16288) );
  OAI21_X1 U19315 ( .B1(n16289), .B2(n21003), .A(n16288), .ZN(n16290) );
  AOI21_X1 U19316 ( .B1(n16316), .B2(n20317), .A(n16290), .ZN(n16292) );
  NAND2_X1 U19317 ( .A1(n16315), .A2(n20339), .ZN(n16291) );
  OAI211_X1 U19318 ( .C1(n16348), .C2(n20325), .A(n16292), .B(n16291), .ZN(
        P1_U2825) );
  AOI21_X1 U19319 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16303), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16298) );
  OAI22_X1 U19320 ( .A1(n20308), .A2(n16311), .B1(n16293), .B2(n20279), .ZN(
        n16294) );
  AOI211_X1 U19321 ( .C1(n16309), .C2(n20334), .A(n20310), .B(n16294), .ZN(
        n16296) );
  AOI22_X1 U19322 ( .A1(n16320), .A2(n20339), .B1(n20317), .B2(n16319), .ZN(
        n16295) );
  OAI211_X1 U19323 ( .C1(n16298), .C2(n16297), .A(n16296), .B(n16295), .ZN(
        P1_U2828) );
  AOI21_X1 U19324 ( .B1(n20340), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20310), .ZN(n16300) );
  NAND2_X1 U19325 ( .A1(n20335), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n16299) );
  OAI211_X1 U19326 ( .C1(n16379), .C2(n20325), .A(n16300), .B(n16299), .ZN(
        n16301) );
  AOI21_X1 U19327 ( .B1(n16302), .B2(P1_REIP_REG_11__SCAN_IN), .A(n16301), 
        .ZN(n16305) );
  INV_X1 U19328 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20998) );
  AOI22_X1 U19329 ( .A1(n16328), .A2(n20317), .B1(n16303), .B2(n20998), .ZN(
        n16304) );
  OAI211_X1 U19330 ( .C1(n16331), .C2(n20330), .A(n16305), .B(n16304), .ZN(
        P1_U2829) );
  AOI22_X1 U19331 ( .A1(n16307), .A2(n20352), .B1(n20351), .B2(n16306), .ZN(
        n16308) );
  OAI21_X1 U19332 ( .B1(n20356), .B2(n21212), .A(n16308), .ZN(P1_U2855) );
  AOI22_X1 U19333 ( .A1(n16319), .A2(n20352), .B1(n20351), .B2(n16309), .ZN(
        n16310) );
  OAI21_X1 U19334 ( .B1(n20356), .B2(n16311), .A(n16310), .ZN(P1_U2860) );
  XNOR2_X1 U19335 ( .A(n15011), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16313) );
  XNOR2_X1 U19336 ( .A(n16314), .B(n16313), .ZN(n16349) );
  AOI22_X1 U19337 ( .A1(n20357), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20407), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16318) );
  AOI22_X1 U19338 ( .A1(n16316), .A2(n16332), .B1(n16315), .B2(n16321), .ZN(
        n16317) );
  OAI211_X1 U19339 ( .C1(n16349), .C2(n20363), .A(n16318), .B(n16317), .ZN(
        P1_U2984) );
  AOI22_X1 U19340 ( .A1(n20357), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20407), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16323) );
  AOI22_X1 U19341 ( .A1(n16321), .A2(n16320), .B1(n16332), .B2(n16319), .ZN(
        n16322) );
  OAI211_X1 U19342 ( .C1(n16324), .C2(n20363), .A(n16323), .B(n16322), .ZN(
        P1_U2987) );
  AOI22_X1 U19343 ( .A1(n20357), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20407), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16330) );
  NOR2_X1 U19344 ( .A1(n15197), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16326) );
  NOR2_X1 U19345 ( .A1(n15149), .A2(n15006), .ZN(n16325) );
  MUX2_X1 U19346 ( .A(n16326), .B(n16325), .S(n15011), .Z(n16327) );
  XNOR2_X1 U19347 ( .A(n16327), .B(n15005), .ZN(n16376) );
  AOI22_X1 U19348 ( .A1(n16345), .A2(n16376), .B1(n16332), .B2(n16328), .ZN(
        n16329) );
  OAI211_X1 U19349 ( .C1(n20368), .C2(n16331), .A(n16330), .B(n16329), .ZN(
        P1_U2988) );
  AOI22_X1 U19350 ( .A1(n20357), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20407), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16335) );
  AOI22_X1 U19351 ( .A1(n16333), .A2(n16345), .B1(n16332), .B2(n20297), .ZN(
        n16334) );
  OAI211_X1 U19352 ( .C1(n20368), .C2(n20307), .A(n16335), .B(n16334), .ZN(
        P1_U2992) );
  AOI22_X1 U19353 ( .A1(n20357), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20407), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16340) );
  XNOR2_X1 U19354 ( .A(n16337), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16338) );
  XNOR2_X1 U19355 ( .A(n16336), .B(n16338), .ZN(n16402) );
  AOI22_X1 U19356 ( .A1(n16402), .A2(n16345), .B1(n16332), .B2(n20353), .ZN(
        n16339) );
  OAI211_X1 U19357 ( .C1(n20368), .C2(n20319), .A(n16340), .B(n16339), .ZN(
        P1_U2993) );
  AOI22_X1 U19358 ( .A1(n20357), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20407), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16347) );
  OAI21_X1 U19359 ( .B1(n16343), .B2(n16342), .A(n16341), .ZN(n16344) );
  INV_X1 U19360 ( .A(n16344), .ZN(n16408) );
  AOI22_X1 U19361 ( .A1(n16408), .A2(n16345), .B1(n16332), .B2(n20327), .ZN(
        n16346) );
  OAI211_X1 U19362 ( .C1(n20368), .C2(n20331), .A(n16347), .B(n16346), .ZN(
        P1_U2994) );
  NOR2_X1 U19363 ( .A1(n20393), .A2(n21003), .ZN(n16351) );
  OAI22_X1 U19364 ( .A1(n16349), .A2(n20408), .B1(n16412), .B2(n16348), .ZN(
        n16350) );
  AOI211_X1 U19365 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16352), .A(
        n16351), .B(n16350), .ZN(n16353) );
  OAI21_X1 U19366 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16354), .A(
        n16353), .ZN(P1_U3016) );
  INV_X1 U19367 ( .A(n16355), .ZN(n16360) );
  AOI22_X1 U19368 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16367), .B1(
        n20407), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16359) );
  AOI22_X1 U19369 ( .A1(n16357), .A2(n20399), .B1(n20406), .B2(n16356), .ZN(
        n16358) );
  OAI211_X1 U19370 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16360), .A(
        n16359), .B(n16358), .ZN(P1_U3017) );
  NAND2_X1 U19371 ( .A1(n16362), .A2(n16361), .ZN(n16365) );
  OAI211_X1 U19372 ( .C1(n16365), .C2(n16364), .A(n16363), .B(n15008), .ZN(
        n16366) );
  AOI22_X1 U19373 ( .A1(n16368), .A2(n20399), .B1(n16367), .B2(n16366), .ZN(
        n16370) );
  NAND2_X1 U19374 ( .A1(n20407), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n16369) );
  OAI211_X1 U19375 ( .C1(n16412), .C2(n16371), .A(n16370), .B(n16369), .ZN(
        P1_U3018) );
  INV_X1 U19376 ( .A(n16372), .ZN(n20388) );
  OAI22_X1 U19377 ( .A1(n20388), .A2(n16374), .B1(n16373), .B2(n15005), .ZN(
        n16375) );
  AOI21_X1 U19378 ( .B1(n16376), .B2(n20399), .A(n16375), .ZN(n16378) );
  NAND2_X1 U19379 ( .A1(n20407), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n16377) );
  OAI211_X1 U19380 ( .C1(n16412), .C2(n16379), .A(n16378), .B(n16377), .ZN(
        P1_U3020) );
  AOI22_X1 U19381 ( .A1(n20407), .A2(P1_REIP_REG_10__SCAN_IN), .B1(n20406), 
        .B2(n16380), .ZN(n16387) );
  AOI22_X1 U19382 ( .A1(n16382), .A2(n20399), .B1(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16381), .ZN(n16386) );
  OAI221_X1 U19383 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n15006), .C2(n16384), .A(
        n16383), .ZN(n16385) );
  NAND3_X1 U19384 ( .A1(n16387), .A2(n16386), .A3(n16385), .ZN(P1_U3021) );
  AOI22_X1 U19385 ( .A1(n20407), .A2(P1_REIP_REG_8__SCAN_IN), .B1(n20406), 
        .B2(n20284), .ZN(n16395) );
  AOI22_X1 U19386 ( .A1(n16389), .A2(n20399), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16388), .ZN(n16394) );
  INV_X1 U19387 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16392) );
  OAI221_X1 U19388 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16392), .C2(n16391), .A(
        n16390), .ZN(n16393) );
  NAND3_X1 U19389 ( .A1(n16395), .A2(n16394), .A3(n16393), .ZN(P1_U3023) );
  AND2_X1 U19390 ( .A1(n16397), .A2(n16396), .ZN(n16405) );
  NAND2_X1 U19391 ( .A1(n16399), .A2(n16398), .ZN(n16400) );
  NAND2_X1 U19392 ( .A1(n16401), .A2(n16400), .ZN(n20312) );
  INV_X1 U19393 ( .A(n20312), .ZN(n20350) );
  AOI22_X1 U19394 ( .A1(n16402), .A2(n20399), .B1(n20406), .B2(n20350), .ZN(
        n16404) );
  NAND2_X1 U19395 ( .A1(n20407), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n16403) );
  OAI211_X1 U19396 ( .C1(n16406), .C2(n16405), .A(n16404), .B(n16403), .ZN(
        P1_U3025) );
  AOI22_X1 U19397 ( .A1(n16408), .A2(n20399), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16407), .ZN(n16416) );
  NAND2_X1 U19398 ( .A1(n20375), .A2(n16409), .ZN(n16410) );
  OAI22_X1 U19399 ( .A1(n16412), .A2(n20324), .B1(n16411), .B2(n16410), .ZN(
        n16413) );
  AOI211_X1 U19400 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n20407), .A(n16414), .B(
        n16413), .ZN(n16415) );
  NAND2_X1 U19401 ( .A1(n16416), .A2(n16415), .ZN(P1_U3026) );
  INV_X1 U19402 ( .A(n16417), .ZN(n16423) );
  NAND3_X1 U19403 ( .A1(n16420), .A2(n16419), .A3(n16418), .ZN(n16421) );
  OAI21_X1 U19404 ( .B1(n16423), .B2(n16422), .A(n16421), .ZN(P1_U3468) );
  NAND4_X1 U19405 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20966), .A4(n21050), .ZN(n16424) );
  NAND2_X1 U19406 ( .A1(n16425), .A2(n16424), .ZN(n20964) );
  OAI21_X1 U19407 ( .B1(n16427), .B2(n20964), .A(n16426), .ZN(n16428) );
  OAI221_X1 U19408 ( .B1(n16429), .B2(n20674), .C1(n16429), .C2(n21050), .A(
        n16428), .ZN(n16430) );
  AOI221_X1 U19409 ( .B1(n16431), .B2(n20962), .C1(n20963), .C2(n20962), .A(
        n16430), .ZN(P1_U3162) );
  NOR2_X1 U19410 ( .A1(n16431), .A2(n20963), .ZN(n16433) );
  OAI22_X1 U19411 ( .A1(n20674), .A2(n16433), .B1(n16432), .B2(n20963), .ZN(
        P1_U3466) );
  AOI21_X1 U19412 ( .B1(n16435), .B2(n16434), .A(n20099), .ZN(n16436) );
  INV_X1 U19413 ( .A(n16436), .ZN(n16444) );
  AOI22_X1 U19414 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19298), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19320), .ZN(n16437) );
  OAI21_X1 U19415 ( .B1(n19260), .B2(n20160), .A(n16437), .ZN(n16438) );
  AOI21_X1 U19416 ( .B1(n16439), .B2(n19317), .A(n16438), .ZN(n16440) );
  OAI21_X1 U19417 ( .B1(n16441), .B2(n19292), .A(n16440), .ZN(n16442) );
  INV_X1 U19418 ( .A(n16442), .ZN(n16443) );
  INV_X1 U19419 ( .A(n16445), .ZN(n16446) );
  OAI21_X1 U19420 ( .B1(n16447), .B2(n19312), .A(n16446), .ZN(P2_U2826) );
  INV_X1 U19421 ( .A(n16448), .ZN(n16462) );
  AOI211_X1 U19422 ( .C1(n16451), .C2(n16449), .A(n16450), .B(n20099), .ZN(
        n16461) );
  INV_X1 U19423 ( .A(n16452), .ZN(n16459) );
  INV_X1 U19424 ( .A(n16453), .ZN(n16457) );
  AOI22_X1 U19425 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19298), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19320), .ZN(n16454) );
  OAI21_X1 U19426 ( .B1(n19260), .B2(n16455), .A(n16454), .ZN(n16456) );
  AOI21_X1 U19427 ( .B1(n16457), .B2(n19317), .A(n16456), .ZN(n16458) );
  OAI21_X1 U19428 ( .B1(n16459), .B2(n19292), .A(n16458), .ZN(n16460) );
  AOI211_X1 U19429 ( .C1(n19319), .C2(n16462), .A(n16461), .B(n16460), .ZN(
        n16463) );
  INV_X1 U19430 ( .A(n16463), .ZN(P2_U2829) );
  AOI22_X1 U19431 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19320), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19318), .ZN(n16477) );
  OAI22_X1 U19432 ( .A1(n16465), .A2(n19300), .B1(n19326), .B2(n16464), .ZN(
        n16466) );
  INV_X1 U19433 ( .A(n16466), .ZN(n16476) );
  INV_X1 U19434 ( .A(n16467), .ZN(n16468) );
  AOI22_X1 U19435 ( .A1(n16469), .A2(n19313), .B1(n19319), .B2(n16468), .ZN(
        n16475) );
  AOI21_X1 U19436 ( .B1(n16472), .B2(n16471), .A(n16470), .ZN(n16473) );
  NAND2_X1 U19437 ( .A1(n19308), .A2(n16473), .ZN(n16474) );
  NAND4_X1 U19438 ( .A1(n16477), .A2(n16476), .A3(n16475), .A4(n16474), .ZN(
        P2_U2831) );
  INV_X1 U19439 ( .A(n19550), .ZN(n16478) );
  AOI22_X1 U19440 ( .A1(n19338), .A2(n16478), .B1(n19399), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16484) );
  AOI22_X1 U19441 ( .A1(n19340), .A2(BUF2_REG_20__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16483) );
  OAI22_X1 U19442 ( .A1(n16480), .A2(n16479), .B1(n19342), .B2(n19171), .ZN(
        n16481) );
  INV_X1 U19443 ( .A(n16481), .ZN(n16482) );
  NAND3_X1 U19444 ( .A1(n16484), .A2(n16483), .A3(n16482), .ZN(P2_U2899) );
  AOI22_X1 U19445 ( .A1(n19484), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19303), .ZN(n16490) );
  OAI22_X1 U19446 ( .A1(n16486), .A2(n16537), .B1(n16526), .B2(n16485), .ZN(
        n16487) );
  AOI21_X1 U19447 ( .B1(n16488), .B2(n16529), .A(n16487), .ZN(n16489) );
  OAI211_X1 U19448 ( .C1(n19496), .C2(n16491), .A(n16490), .B(n16489), .ZN(
        P2_U2992) );
  AOI22_X1 U19449 ( .A1(n19484), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19303), .ZN(n16495) );
  AOI222_X1 U19450 ( .A1(n16493), .A2(n10990), .B1(n16529), .B2(n16492), .C1(
        n19486), .C2(n19205), .ZN(n16494) );
  OAI211_X1 U19451 ( .C1(n19496), .C2(n16496), .A(n16495), .B(n16494), .ZN(
        P2_U2996) );
  AOI22_X1 U19452 ( .A1(n19484), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19303), .ZN(n16503) );
  NOR2_X1 U19453 ( .A1(n19232), .A2(n16526), .ZN(n16497) );
  AOI21_X1 U19454 ( .B1(n16498), .B2(n16529), .A(n16497), .ZN(n16501) );
  NAND2_X1 U19455 ( .A1(n16499), .A2(n10990), .ZN(n16500) );
  AND2_X1 U19456 ( .A1(n16501), .A2(n16500), .ZN(n16502) );
  OAI211_X1 U19457 ( .C1(n19496), .C2(n19225), .A(n16503), .B(n16502), .ZN(
        P2_U3000) );
  AOI22_X1 U19458 ( .A1(n19484), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19303), .ZN(n16508) );
  AOI222_X1 U19459 ( .A1(n16506), .A2(n16529), .B1(n10990), .B2(n16505), .C1(
        n19486), .C2(n16504), .ZN(n16507) );
  OAI211_X1 U19460 ( .C1(n19496), .C2(n19251), .A(n16508), .B(n16507), .ZN(
        P2_U3002) );
  AOI22_X1 U19461 ( .A1(n19484), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19303), .ZN(n16513) );
  AOI222_X1 U19462 ( .A1(n16511), .A2(n10990), .B1(n19486), .B2(n16510), .C1(
        n16529), .C2(n16509), .ZN(n16512) );
  OAI211_X1 U19463 ( .C1(n19496), .C2(n16514), .A(n16513), .B(n16512), .ZN(
        P2_U3004) );
  AOI22_X1 U19464 ( .A1(n19484), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19303), .ZN(n16524) );
  XOR2_X1 U19465 ( .A(n16515), .B(n16516), .Z(n16551) );
  NOR2_X1 U19466 ( .A1(n14233), .A2(n16517), .ZN(n16521) );
  NAND2_X1 U19467 ( .A1(n16519), .A2(n16518), .ZN(n16520) );
  XNOR2_X1 U19468 ( .A(n16521), .B(n16520), .ZN(n16542) );
  INV_X1 U19469 ( .A(n16548), .ZN(n16522) );
  AOI222_X1 U19470 ( .A1(n16551), .A2(n16529), .B1(n10990), .B2(n16542), .C1(
        n19486), .C2(n16522), .ZN(n16523) );
  OAI211_X1 U19471 ( .C1(n19496), .C2(n16525), .A(n16524), .B(n16523), .ZN(
        P2_U3006) );
  AOI22_X1 U19472 ( .A1(n19484), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19303), .ZN(n16532) );
  OAI22_X1 U19473 ( .A1(n16527), .A2(n16537), .B1(n16526), .B2(n19293), .ZN(
        n16528) );
  AOI21_X1 U19474 ( .B1(n16530), .B2(n16529), .A(n16528), .ZN(n16531) );
  OAI211_X1 U19475 ( .C1(n19496), .C2(n19291), .A(n16532), .B(n16531), .ZN(
        P2_U3008) );
  AOI22_X1 U19476 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19303), .B1(n16533), 
        .B2(n19306), .ZN(n16540) );
  INV_X1 U19477 ( .A(n16534), .ZN(n19307) );
  OAI22_X1 U19478 ( .A1(n16537), .A2(n16536), .B1(n16535), .B2(n19490), .ZN(
        n16538) );
  AOI21_X1 U19479 ( .B1(n19486), .B2(n19307), .A(n16538), .ZN(n16539) );
  OAI211_X1 U19480 ( .C1(n16541), .C2(n10719), .A(n16540), .B(n16539), .ZN(
        P2_U3009) );
  INV_X1 U19481 ( .A(n16560), .ZN(n16558) );
  NAND2_X1 U19482 ( .A1(n16542), .A2(n16568), .ZN(n16546) );
  INV_X1 U19483 ( .A(n19368), .ZN(n16543) );
  AOI22_X1 U19484 ( .A1(n16544), .A2(n16543), .B1(n19303), .B2(
        P2_REIP_REG_8__SCAN_IN), .ZN(n16545) );
  OAI211_X1 U19485 ( .C1(n16548), .C2(n16547), .A(n16546), .B(n16545), .ZN(
        n16549) );
  AOI21_X1 U19486 ( .B1(n16551), .B2(n16550), .A(n16549), .ZN(n16556) );
  NOR2_X1 U19487 ( .A1(n16553), .A2(n16552), .ZN(n16561) );
  OAI211_X1 U19488 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16561), .B(n16554), .ZN(n16555) );
  OAI211_X1 U19489 ( .C1(n16558), .C2(n16557), .A(n16556), .B(n16555), .ZN(
        P2_U3038) );
  AOI22_X1 U19490 ( .A1(n16560), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19505), .B2(n16559), .ZN(n16571) );
  INV_X1 U19491 ( .A(n16561), .ZN(n16562) );
  NOR2_X1 U19492 ( .A1(n16562), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16567) );
  OR2_X1 U19493 ( .A1(n16564), .A2(n16563), .ZN(n16565) );
  NAND2_X1 U19494 ( .A1(n16565), .A2(n13599), .ZN(n19369) );
  OAI22_X1 U19495 ( .A1(n19508), .A2(n19369), .B1(n20129), .B2(n19277), .ZN(
        n16566) );
  AOI211_X1 U19496 ( .C1(n16569), .C2(n16568), .A(n16567), .B(n16566), .ZN(
        n16570) );
  OAI211_X1 U19497 ( .C1(n19515), .C2(n16572), .A(n16571), .B(n16570), .ZN(
        P2_U3039) );
  NAND2_X1 U19498 ( .A1(n16589), .A2(n10261), .ZN(n16573) );
  OAI21_X1 U19499 ( .B1(n16574), .B2(n16589), .A(n16573), .ZN(n16588) );
  NAND2_X1 U19500 ( .A1(n16589), .A2(n16575), .ZN(n16576) );
  OAI21_X1 U19501 ( .B1(n16577), .B2(n16589), .A(n16576), .ZN(n16587) );
  OR2_X1 U19502 ( .A1(n16578), .A2(n20208), .ZN(n16579) );
  OAI21_X1 U19503 ( .B1(n16580), .B2(n16579), .A(n20199), .ZN(n16582) );
  NAND2_X1 U19504 ( .A1(n16580), .A2(n16579), .ZN(n16581) );
  AOI21_X1 U19505 ( .B1(n16582), .B2(n16581), .A(n16589), .ZN(n16585) );
  AOI22_X1 U19506 ( .A1(n16587), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n16588), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16584) );
  NOR2_X1 U19507 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19626) );
  INV_X1 U19508 ( .A(n19626), .ZN(n19625) );
  OAI22_X1 U19509 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16588), .B1(
        n19625), .B2(n16587), .ZN(n16583) );
  AOI21_X1 U19510 ( .B1(n16585), .B2(n16584), .A(n16583), .ZN(n16586) );
  OAI22_X1 U19511 ( .A1(n16588), .A2(n16587), .B1(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n16586), .ZN(n16607) );
  NAND2_X1 U19512 ( .A1(n16589), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n16605) );
  INV_X1 U19513 ( .A(n16590), .ZN(n16592) );
  NAND2_X1 U19514 ( .A1(n16592), .A2(n16591), .ZN(n16595) );
  NAND2_X1 U19515 ( .A1(n16597), .A2(n16593), .ZN(n16594) );
  OAI211_X1 U19516 ( .C1(n16597), .C2(n16596), .A(n16595), .B(n16594), .ZN(
        n20211) );
  NOR2_X1 U19517 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n16601) );
  NAND2_X1 U19518 ( .A1(n16598), .A2(n10297), .ZN(n16599) );
  OAI211_X1 U19519 ( .C1(n16602), .C2(n16601), .A(n16600), .B(n16599), .ZN(
        n16603) );
  NOR2_X1 U19520 ( .A1(n20211), .A2(n16603), .ZN(n16604) );
  NAND2_X1 U19521 ( .A1(n16605), .A2(n16604), .ZN(n16606) );
  OR2_X1 U19522 ( .A1(n16607), .A2(n16606), .ZN(n16611) );
  INV_X1 U19523 ( .A(n16611), .ZN(n16623) );
  NOR3_X1 U19524 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n16267), .A3(n20226), 
        .ZN(n16609) );
  AOI211_X1 U19525 ( .C1(n20217), .C2(n16610), .A(n16609), .B(n16608), .ZN(
        n16621) );
  OAI21_X1 U19526 ( .B1(n16611), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16612) );
  OAI21_X1 U19527 ( .B1(n16613), .B2(n12773), .A(n16612), .ZN(n16614) );
  AOI21_X1 U19528 ( .B1(n16617), .B2(n16616), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16619) );
  NAND2_X1 U19529 ( .A1(n20101), .A2(n20114), .ZN(n16618) );
  AOI22_X1 U19530 ( .A1(n20101), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16619), 
        .B2(n16618), .ZN(n16620) );
  OAI211_X1 U19531 ( .C1(n16623), .C2(n16622), .A(n16621), .B(n16620), .ZN(
        P2_U3176) );
  INV_X1 U19532 ( .A(n20101), .ZN(n16625) );
  OAI221_X1 U19533 ( .B1(n20041), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n20041), 
        .C2(n16625), .A(n16624), .ZN(P2_U3593) );
  INV_X1 U19534 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19074) );
  NAND2_X1 U19535 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19074), .ZN(
        n16669) );
  OAI211_X1 U19536 ( .C1(n18038), .C2(n16627), .A(n16669), .B(n10147), .ZN(
        n16632) );
  OAI21_X1 U19537 ( .B1(n17933), .B2(n16628), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16630) );
  NOR2_X1 U19538 ( .A1(n17933), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16633) );
  INV_X1 U19539 ( .A(n16633), .ZN(n16629) );
  AND2_X1 U19540 ( .A1(n16630), .A2(n16629), .ZN(n16631) );
  NAND2_X1 U19541 ( .A1(n16632), .A2(n16631), .ZN(n16639) );
  NAND2_X1 U19542 ( .A1(n16626), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16637) );
  NOR2_X1 U19543 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19074), .ZN(
        n16673) );
  AOI21_X1 U19544 ( .B1(n16673), .B2(n16634), .A(n16633), .ZN(n16635) );
  NAND2_X1 U19545 ( .A1(n16637), .A2(n16636), .ZN(n16638) );
  INV_X1 U19546 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16830) );
  INV_X1 U19547 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19054) );
  NOR2_X1 U19548 ( .A1(n19054), .A2(n18384), .ZN(n16672) );
  NOR2_X1 U19549 ( .A1(n16844), .A2(n16641), .ZN(n16644) );
  INV_X1 U19550 ( .A(n16642), .ZN(n16643) );
  MUX2_X1 U19551 ( .A(n16644), .B(n16643), .S(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .Z(n16645) );
  AOI211_X1 U19552 ( .C1(n17979), .C2(n9942), .A(n16672), .B(n16645), .ZN(
        n16650) );
  INV_X1 U19553 ( .A(n16646), .ZN(n16654) );
  NAND2_X1 U19554 ( .A1(n16654), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16647) );
  XOR2_X1 U19555 ( .A(n16647), .B(n19074), .Z(n16675) );
  NAND2_X1 U19556 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16656), .ZN(
        n16648) );
  XOR2_X1 U19557 ( .A(n19074), .B(n16648), .Z(n16674) );
  AOI22_X1 U19558 ( .A1(n9802), .A2(n16675), .B1(n18115), .B2(n16674), .ZN(
        n16649) );
  OAI211_X1 U19559 ( .C1(n18024), .C2(n16678), .A(n16650), .B(n16649), .ZN(
        P3_U2799) );
  OAI21_X1 U19560 ( .B1(n18507), .B2(n16651), .A(n16862), .ZN(n16652) );
  AOI22_X1 U19561 ( .A1(n18385), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n16653), 
        .B2(n16652), .ZN(n16664) );
  AOI211_X1 U19562 ( .C1(n16655), .C2(n12306), .A(n16654), .B(n17971), .ZN(
        n16658) );
  AOI211_X1 U19563 ( .C1(n12306), .C2(n16691), .A(n16656), .B(n18130), .ZN(
        n16657) );
  AOI211_X1 U19564 ( .C1(n16659), .C2(n18039), .A(n16658), .B(n16657), .ZN(
        n16663) );
  AOI21_X1 U19565 ( .B1(n16862), .B2(n16810), .A(n16660), .ZN(n16856) );
  OAI21_X1 U19566 ( .B1(n16661), .B2(n17979), .A(n16856), .ZN(n16662) );
  NAND3_X1 U19567 ( .A1(n16664), .A2(n16663), .A3(n16662), .ZN(P3_U2801) );
  INV_X1 U19568 ( .A(n16665), .ZN(n16667) );
  NAND2_X1 U19569 ( .A1(n16667), .A2(n16666), .ZN(n16668) );
  OAI22_X1 U19570 ( .A1(n16670), .A2(n19074), .B1(n16669), .B2(n16668), .ZN(
        n16671) );
  AOI211_X1 U19571 ( .C1(n16673), .C2(n18446), .A(n16672), .B(n16671), .ZN(
        n16677) );
  AOI22_X1 U19572 ( .A1(n16675), .A2(n18368), .B1(n16674), .B2(n18443), .ZN(
        n16676) );
  OAI211_X1 U19573 ( .C1(n16678), .C2(n18352), .A(n16677), .B(n16676), .ZN(
        P3_U2831) );
  NOR2_X1 U19574 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18140), .ZN(
        n17765) );
  OAI22_X1 U19575 ( .A1(n18324), .A2(n18303), .B1(n18322), .B2(n18301), .ZN(
        n18235) );
  AOI21_X1 U19576 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n9660), .A(
        n18921), .ZN(n18425) );
  OAI22_X1 U19577 ( .A1(n18924), .A2(n18256), .B1(n18281), .B2(n18425), .ZN(
        n16679) );
  OAI21_X1 U19578 ( .B1(n18235), .B2(n16679), .A(n18237), .ZN(n18145) );
  NOR2_X1 U19579 ( .A1(n16680), .A2(n18145), .ZN(n18141) );
  INV_X1 U19580 ( .A(n17773), .ZN(n16682) );
  INV_X1 U19581 ( .A(n18912), .ZN(n18372) );
  OAI21_X1 U19582 ( .B1(n18038), .B2(n17755), .A(n16683), .ZN(n17768) );
  NAND2_X1 U19583 ( .A1(n17768), .A2(n17767), .ZN(n17766) );
  NAND3_X1 U19584 ( .A1(n18372), .A2(n16681), .A3(n17766), .ZN(n16685) );
  AOI21_X1 U19585 ( .B1(n16683), .B2(n16682), .A(n16685), .ZN(n16684) );
  AOI21_X1 U19586 ( .B1(n17765), .B2(n18141), .A(n16684), .ZN(n16697) );
  INV_X1 U19587 ( .A(n16685), .ZN(n16687) );
  NAND2_X1 U19588 ( .A1(n16687), .A2(n16686), .ZN(n16694) );
  OR2_X1 U19589 ( .A1(n16688), .A2(n18301), .ZN(n16693) );
  INV_X1 U19590 ( .A(n16689), .ZN(n16690) );
  NAND2_X1 U19591 ( .A1(n16694), .A2(n10192), .ZN(n16695) );
  NAND3_X1 U19592 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18384), .A3(
        n16695), .ZN(n16696) );
  NAND2_X1 U19593 ( .A1(n18385), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17760) );
  OAI211_X1 U19594 ( .C1(n16697), .C2(n18433), .A(n16696), .B(n17760), .ZN(
        P3_U2834) );
  INV_X1 U19595 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n21206) );
  NOR4_X1 U19596 ( .A1(P3_BE_N_REG_0__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .A4(n21206), .ZN(n16699) );
  NOR4_X1 U19597 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16698) );
  NAND3_X1 U19598 ( .A1(n16699), .A2(n16698), .A3(U215), .ZN(U213) );
  INV_X1 U19599 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19415) );
  NOR2_X1 U19600 ( .A1(n16743), .A2(n16700), .ZN(n16744) );
  INV_X1 U19601 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16781) );
  OAI222_X1 U19602 ( .A1(U212), .A2(n19415), .B1(n16750), .B2(n16701), .C1(
        U214), .C2(n16781), .ZN(U216) );
  AOI22_X1 U19603 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n16743), .ZN(n16702) );
  OAI21_X1 U19604 ( .B1(n14900), .B2(n16750), .A(n16702), .ZN(U217) );
  AOI22_X1 U19605 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16743), .ZN(n16703) );
  OAI21_X1 U19606 ( .B1(n14331), .B2(n16750), .A(n16703), .ZN(U218) );
  INV_X1 U19607 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n21094) );
  AOI22_X1 U19608 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16743), .ZN(n16704) );
  OAI21_X1 U19609 ( .B1(n21094), .B2(n16750), .A(n16704), .ZN(U219) );
  INV_X1 U19610 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16706) );
  AOI22_X1 U19611 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16743), .ZN(n16705) );
  OAI21_X1 U19612 ( .B1(n16706), .B2(n16750), .A(n16705), .ZN(U220) );
  INV_X1 U19613 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16708) );
  AOI22_X1 U19614 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16743), .ZN(n16707) );
  OAI21_X1 U19615 ( .B1(n16708), .B2(n16750), .A(n16707), .ZN(U221) );
  INV_X1 U19616 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16710) );
  AOI22_X1 U19617 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16743), .ZN(n16709) );
  OAI21_X1 U19618 ( .B1(n16710), .B2(n16750), .A(n16709), .ZN(U222) );
  INV_X1 U19619 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16712) );
  AOI22_X1 U19620 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16743), .ZN(n16711) );
  OAI21_X1 U19621 ( .B1(n16712), .B2(n16750), .A(n16711), .ZN(U223) );
  INV_X1 U19622 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16714) );
  AOI22_X1 U19623 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16743), .ZN(n16713) );
  OAI21_X1 U19624 ( .B1(n16714), .B2(n16750), .A(n16713), .ZN(U224) );
  INV_X1 U19625 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n19559) );
  AOI22_X1 U19626 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16743), .ZN(n16715) );
  OAI21_X1 U19627 ( .B1(n19559), .B2(n16750), .A(n16715), .ZN(U225) );
  AOI22_X1 U19628 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16743), .ZN(n16716) );
  OAI21_X1 U19629 ( .B1(n16717), .B2(n16750), .A(n16716), .ZN(U226) );
  INV_X1 U19630 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16719) );
  AOI22_X1 U19631 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16743), .ZN(n16718) );
  OAI21_X1 U19632 ( .B1(n16719), .B2(n16750), .A(n16718), .ZN(U227) );
  INV_X1 U19633 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n19544) );
  AOI22_X1 U19634 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16743), .ZN(n16720) );
  OAI21_X1 U19635 ( .B1(n19544), .B2(n16750), .A(n16720), .ZN(U228) );
  INV_X1 U19636 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16722) );
  AOI22_X1 U19637 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16743), .ZN(n16721) );
  OAI21_X1 U19638 ( .B1(n16722), .B2(n16750), .A(n16721), .ZN(U229) );
  AOI22_X1 U19639 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16743), .ZN(n16723) );
  OAI21_X1 U19640 ( .B1(n16724), .B2(n16750), .A(n16723), .ZN(U230) );
  INV_X1 U19641 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16727) );
  AOI22_X1 U19642 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16725), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16743), .ZN(n16726) );
  OAI21_X1 U19643 ( .B1(n16727), .B2(n16750), .A(n16726), .ZN(U231) );
  AOI22_X1 U19644 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16743), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16725), .ZN(n16728) );
  OAI21_X1 U19645 ( .B1(n13099), .B2(n16750), .A(n16728), .ZN(U232) );
  AOI22_X1 U19646 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16743), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16725), .ZN(n16729) );
  OAI21_X1 U19647 ( .B1(n12860), .B2(n16750), .A(n16729), .ZN(U233) );
  AOI22_X1 U19648 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16743), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16725), .ZN(n16730) );
  OAI21_X1 U19649 ( .B1(n16731), .B2(n16750), .A(n16730), .ZN(U234) );
  AOI22_X1 U19650 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16743), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16725), .ZN(n16732) );
  OAI21_X1 U19651 ( .B1(n16733), .B2(n16750), .A(n16732), .ZN(U235) );
  INV_X1 U19652 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n21219) );
  AOI22_X1 U19653 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16744), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16743), .ZN(n16734) );
  OAI21_X1 U19654 ( .B1(n21219), .B2(U212), .A(n16734), .ZN(U236) );
  AOI222_X1 U19655 ( .A1(n16725), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n16744), 
        .B2(BUF1_REG_10__SCAN_IN), .C1(n16743), .C2(P1_DATAO_REG_10__SCAN_IN), 
        .ZN(n16735) );
  INV_X1 U19656 ( .A(n16735), .ZN(U237) );
  INV_X1 U19657 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16761) );
  AOI22_X1 U19658 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16744), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16743), .ZN(n16736) );
  OAI21_X1 U19659 ( .B1(n16761), .B2(U212), .A(n16736), .ZN(U238) );
  AOI22_X1 U19660 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16743), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16725), .ZN(n16737) );
  OAI21_X1 U19661 ( .B1(n16738), .B2(n16750), .A(n16737), .ZN(U239) );
  INV_X1 U19662 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16759) );
  AOI22_X1 U19663 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16744), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16743), .ZN(n16739) );
  OAI21_X1 U19664 ( .B1(n16759), .B2(U212), .A(n16739), .ZN(U240) );
  INV_X1 U19665 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16758) );
  AOI22_X1 U19666 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16744), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16743), .ZN(n16740) );
  OAI21_X1 U19667 ( .B1(n16758), .B2(U212), .A(n16740), .ZN(U241) );
  INV_X1 U19668 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16757) );
  AOI22_X1 U19669 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16744), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16743), .ZN(n16741) );
  OAI21_X1 U19670 ( .B1(n16757), .B2(U212), .A(n16741), .ZN(U242) );
  INV_X1 U19671 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n21194) );
  AOI22_X1 U19672 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16743), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16725), .ZN(n16742) );
  OAI21_X1 U19673 ( .B1(n21194), .B2(n16750), .A(n16742), .ZN(U243) );
  INV_X1 U19674 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16755) );
  AOI22_X1 U19675 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16744), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16743), .ZN(n16745) );
  OAI21_X1 U19676 ( .B1(n16755), .B2(U212), .A(n16745), .ZN(U244) );
  INV_X1 U19677 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n21098) );
  AOI22_X1 U19678 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16743), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16725), .ZN(n16746) );
  OAI21_X1 U19679 ( .B1(n21098), .B2(n16750), .A(n16746), .ZN(U245) );
  INV_X1 U19680 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16748) );
  AOI22_X1 U19681 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16743), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16725), .ZN(n16747) );
  OAI21_X1 U19682 ( .B1(n16748), .B2(n16750), .A(n16747), .ZN(U246) );
  INV_X1 U19683 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16751) );
  AOI22_X1 U19684 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16743), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16725), .ZN(n16749) );
  OAI21_X1 U19685 ( .B1(n16751), .B2(n16750), .A(n16749), .ZN(U247) );
  OAI22_X1 U19686 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n21255), .ZN(n16752) );
  INV_X1 U19687 ( .A(n16752), .ZN(U251) );
  OAI22_X1 U19688 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n21255), .ZN(n16753) );
  INV_X1 U19689 ( .A(n16753), .ZN(U252) );
  OAI22_X1 U19690 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n21255), .ZN(n16754) );
  INV_X1 U19691 ( .A(n16754), .ZN(U253) );
  INV_X1 U19692 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18489) );
  AOI22_X1 U19693 ( .A1(n21255), .A2(n16755), .B1(n18489), .B2(U215), .ZN(U254) );
  OAI22_X1 U19694 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n21255), .ZN(n16756) );
  INV_X1 U19695 ( .A(n16756), .ZN(U255) );
  INV_X1 U19696 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18501) );
  AOI22_X1 U19697 ( .A1(n21255), .A2(n16757), .B1(n18501), .B2(U215), .ZN(U256) );
  INV_X1 U19698 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18509) );
  AOI22_X1 U19699 ( .A1(n21255), .A2(n16758), .B1(n18509), .B2(U215), .ZN(U257) );
  INV_X1 U19700 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18514) );
  AOI22_X1 U19701 ( .A1(n21255), .A2(n16759), .B1(n18514), .B2(U215), .ZN(U258) );
  OAI22_X1 U19702 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16778), .ZN(n16760) );
  INV_X1 U19703 ( .A(n16760), .ZN(U259) );
  INV_X1 U19704 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17736) );
  AOI22_X1 U19705 ( .A1(n21255), .A2(n16761), .B1(n17736), .B2(U215), .ZN(U260) );
  INV_X1 U19706 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n19458) );
  INV_X1 U19707 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17738) );
  AOI22_X1 U19708 ( .A1(n21255), .A2(n19458), .B1(n17738), .B2(U215), .ZN(U261) );
  INV_X1 U19709 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17740) );
  AOI22_X1 U19710 ( .A1(n21255), .A2(n21219), .B1(n17740), .B2(U215), .ZN(U262) );
  OAI22_X1 U19711 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16778), .ZN(n16762) );
  INV_X1 U19712 ( .A(n16762), .ZN(U263) );
  OAI22_X1 U19713 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16778), .ZN(n16763) );
  INV_X1 U19714 ( .A(n16763), .ZN(U264) );
  OAI22_X1 U19715 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16778), .ZN(n16764) );
  INV_X1 U19716 ( .A(n16764), .ZN(U265) );
  OAI22_X1 U19717 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n21255), .ZN(n16765) );
  INV_X1 U19718 ( .A(n16765), .ZN(U266) );
  OAI22_X1 U19719 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n21255), .ZN(n16766) );
  INV_X1 U19720 ( .A(n16766), .ZN(U267) );
  OAI22_X1 U19721 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n21255), .ZN(n16767) );
  INV_X1 U19722 ( .A(n16767), .ZN(U268) );
  OAI22_X1 U19723 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n21255), .ZN(n16768) );
  INV_X1 U19724 ( .A(n16768), .ZN(U269) );
  INV_X1 U19725 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n21099) );
  INV_X1 U19726 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n19543) );
  AOI22_X1 U19727 ( .A1(n21255), .A2(n21099), .B1(n19543), .B2(U215), .ZN(U270) );
  OAI22_X1 U19728 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n21255), .ZN(n16769) );
  INV_X1 U19729 ( .A(n16769), .ZN(U271) );
  OAI22_X1 U19730 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n21255), .ZN(n16770) );
  INV_X1 U19731 ( .A(n16770), .ZN(U272) );
  INV_X1 U19732 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n21211) );
  INV_X1 U19733 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19557) );
  AOI22_X1 U19734 ( .A1(n21255), .A2(n21211), .B1(n19557), .B2(U215), .ZN(U273) );
  OAI22_X1 U19735 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n21255), .ZN(n16771) );
  INV_X1 U19736 ( .A(n16771), .ZN(U274) );
  OAI22_X1 U19737 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n21255), .ZN(n16772) );
  INV_X1 U19738 ( .A(n16772), .ZN(U275) );
  OAI22_X1 U19739 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16778), .ZN(n16773) );
  INV_X1 U19740 ( .A(n16773), .ZN(U276) );
  OAI22_X1 U19741 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16778), .ZN(n16774) );
  INV_X1 U19742 ( .A(n16774), .ZN(U277) );
  OAI22_X1 U19743 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16778), .ZN(n16775) );
  INV_X1 U19744 ( .A(n16775), .ZN(U278) );
  OAI22_X1 U19745 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16778), .ZN(n16776) );
  INV_X1 U19746 ( .A(n16776), .ZN(U279) );
  OAI22_X1 U19747 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16778), .ZN(n16777) );
  INV_X1 U19748 ( .A(n16777), .ZN(U280) );
  OAI22_X1 U19749 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16778), .ZN(n16779) );
  INV_X1 U19750 ( .A(n16779), .ZN(U281) );
  INV_X1 U19751 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16780) );
  AOI222_X1 U19752 ( .A1(n19415), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16781), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16780), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16782) );
  INV_X2 U19753 ( .A(n16784), .ZN(n16783) );
  INV_X1 U19754 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19015) );
  INV_X1 U19755 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20134) );
  AOI22_X1 U19756 ( .A1(n16783), .A2(n19015), .B1(n20134), .B2(n16784), .ZN(
        U347) );
  INV_X1 U19757 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19014) );
  INV_X1 U19758 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20133) );
  AOI22_X1 U19759 ( .A1(n16783), .A2(n19014), .B1(n20133), .B2(n16784), .ZN(
        U348) );
  INV_X1 U19760 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19011) );
  INV_X1 U19761 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20131) );
  AOI22_X1 U19762 ( .A1(n16783), .A2(n19011), .B1(n20131), .B2(n16784), .ZN(
        U349) );
  INV_X1 U19763 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19010) );
  INV_X1 U19764 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20130) );
  AOI22_X1 U19765 ( .A1(n16783), .A2(n19010), .B1(n20130), .B2(n16784), .ZN(
        U350) );
  INV_X1 U19766 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19008) );
  INV_X1 U19767 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20128) );
  AOI22_X1 U19768 ( .A1(n16783), .A2(n19008), .B1(n20128), .B2(n16784), .ZN(
        U351) );
  INV_X1 U19769 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19006) );
  INV_X1 U19770 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20126) );
  AOI22_X1 U19771 ( .A1(n16783), .A2(n19006), .B1(n20126), .B2(n16784), .ZN(
        U352) );
  INV_X1 U19772 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19004) );
  INV_X1 U19773 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20125) );
  AOI22_X1 U19774 ( .A1(n16783), .A2(n19004), .B1(n20125), .B2(n16784), .ZN(
        U353) );
  INV_X1 U19775 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19001) );
  AOI22_X1 U19776 ( .A1(n16783), .A2(n19001), .B1(n20124), .B2(n16784), .ZN(
        U354) );
  INV_X1 U19777 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19056) );
  INV_X1 U19778 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20164) );
  AOI22_X1 U19779 ( .A1(n16783), .A2(n19056), .B1(n20164), .B2(n16784), .ZN(
        U355) );
  INV_X1 U19780 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19053) );
  INV_X1 U19781 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20161) );
  AOI22_X1 U19782 ( .A1(n16783), .A2(n19053), .B1(n20161), .B2(n16784), .ZN(
        U356) );
  INV_X1 U19783 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19051) );
  INV_X1 U19784 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20159) );
  AOI22_X1 U19785 ( .A1(n16783), .A2(n19051), .B1(n20159), .B2(n16784), .ZN(
        U357) );
  INV_X1 U19786 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19050) );
  INV_X1 U19787 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20156) );
  AOI22_X1 U19788 ( .A1(n16783), .A2(n19050), .B1(n20156), .B2(n16784), .ZN(
        U358) );
  INV_X1 U19789 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19048) );
  INV_X1 U19790 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20155) );
  AOI22_X1 U19791 ( .A1(n16783), .A2(n19048), .B1(n20155), .B2(n16784), .ZN(
        U359) );
  INV_X1 U19792 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19046) );
  INV_X1 U19793 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n21237) );
  AOI22_X1 U19794 ( .A1(n16783), .A2(n19046), .B1(n21237), .B2(n16784), .ZN(
        U360) );
  INV_X1 U19795 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19043) );
  INV_X1 U19796 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20153) );
  AOI22_X1 U19797 ( .A1(n16783), .A2(n19043), .B1(n20153), .B2(n16784), .ZN(
        U361) );
  INV_X1 U19798 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19041) );
  INV_X1 U19799 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20151) );
  AOI22_X1 U19800 ( .A1(n16783), .A2(n19041), .B1(n20151), .B2(n16784), .ZN(
        U362) );
  INV_X1 U19801 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19039) );
  INV_X1 U19802 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20150) );
  AOI22_X1 U19803 ( .A1(n16783), .A2(n19039), .B1(n20150), .B2(n16784), .ZN(
        U363) );
  INV_X1 U19804 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19037) );
  INV_X1 U19805 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20149) );
  AOI22_X1 U19806 ( .A1(n16783), .A2(n19037), .B1(n20149), .B2(n16784), .ZN(
        U364) );
  INV_X1 U19807 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18999) );
  INV_X1 U19808 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20123) );
  AOI22_X1 U19809 ( .A1(n16783), .A2(n18999), .B1(n20123), .B2(n16784), .ZN(
        U365) );
  INV_X1 U19810 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19035) );
  INV_X1 U19811 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20147) );
  AOI22_X1 U19812 ( .A1(n16783), .A2(n19035), .B1(n20147), .B2(n16784), .ZN(
        U366) );
  INV_X1 U19813 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19033) );
  INV_X1 U19814 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20146) );
  AOI22_X1 U19815 ( .A1(n16783), .A2(n19033), .B1(n20146), .B2(n16784), .ZN(
        U367) );
  INV_X1 U19816 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19031) );
  INV_X1 U19817 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20145) );
  AOI22_X1 U19818 ( .A1(n16783), .A2(n19031), .B1(n20145), .B2(n16784), .ZN(
        U368) );
  INV_X1 U19819 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19029) );
  INV_X1 U19820 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20144) );
  AOI22_X1 U19821 ( .A1(n16783), .A2(n19029), .B1(n20144), .B2(n16784), .ZN(
        U369) );
  INV_X1 U19822 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19027) );
  INV_X1 U19823 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20142) );
  AOI22_X1 U19824 ( .A1(n16783), .A2(n19027), .B1(n20142), .B2(n16784), .ZN(
        U370) );
  INV_X1 U19825 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19025) );
  INV_X1 U19826 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20140) );
  AOI22_X1 U19827 ( .A1(n16783), .A2(n19025), .B1(n20140), .B2(n16784), .ZN(
        U371) );
  INV_X1 U19828 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19022) );
  INV_X1 U19829 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20139) );
  AOI22_X1 U19830 ( .A1(n16783), .A2(n19022), .B1(n20139), .B2(n16784), .ZN(
        U372) );
  INV_X1 U19831 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19021) );
  INV_X1 U19832 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20138) );
  AOI22_X1 U19833 ( .A1(n16783), .A2(n19021), .B1(n20138), .B2(n16784), .ZN(
        U373) );
  INV_X1 U19834 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19019) );
  INV_X1 U19835 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20137) );
  AOI22_X1 U19836 ( .A1(n16783), .A2(n19019), .B1(n20137), .B2(n16784), .ZN(
        U374) );
  INV_X1 U19837 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19017) );
  INV_X1 U19838 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20135) );
  AOI22_X1 U19839 ( .A1(n16783), .A2(n19017), .B1(n20135), .B2(n16784), .ZN(
        U375) );
  INV_X1 U19840 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18997) );
  INV_X1 U19841 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20122) );
  AOI22_X1 U19842 ( .A1(n16783), .A2(n18997), .B1(n20122), .B2(n16784), .ZN(
        U376) );
  INV_X1 U19843 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18994) );
  NOR2_X1 U19844 ( .A1(n18982), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18985) );
  OAI22_X1 U19845 ( .A1(n18994), .A2(n18985), .B1(n18982), .B2(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18978) );
  INV_X1 U19846 ( .A(n18978), .ZN(n19065) );
  AOI21_X1 U19847 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19065), .ZN(n16785) );
  INV_X1 U19848 ( .A(n16785), .ZN(P3_U2633) );
  NOR2_X1 U19849 ( .A1(n17706), .A2(n16792), .ZN(n16787) );
  OAI21_X1 U19850 ( .B1(n16787), .B2(n17641), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16788) );
  OAI21_X1 U19851 ( .B1(n16789), .B2(n18970), .A(n16788), .ZN(P3_U2634) );
  INV_X1 U19852 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18996) );
  AOI21_X1 U19853 ( .B1(n18994), .B2(n18996), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16790) );
  AOI22_X1 U19854 ( .A1(n19121), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16790), 
        .B2(n19120), .ZN(P3_U2635) );
  OAI21_X1 U19855 ( .B1(n18980), .B2(BS16), .A(n19065), .ZN(n19063) );
  OAI21_X1 U19856 ( .B1(n19065), .B2(n19111), .A(n19063), .ZN(P3_U2636) );
  OAI211_X1 U19857 ( .C1(n17706), .C2(n16792), .A(n16791), .B(n18910), .ZN(
        n16793) );
  INV_X1 U19858 ( .A(n16793), .ZN(n18913) );
  NOR2_X1 U19859 ( .A1(n18913), .A2(n18967), .ZN(n19104) );
  OAI21_X1 U19860 ( .B1(n19104), .B2(n18460), .A(n16794), .ZN(P3_U2637) );
  NOR4_X1 U19861 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16798) );
  NOR4_X1 U19862 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16797) );
  NOR4_X1 U19863 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16796) );
  NOR4_X1 U19864 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16795) );
  NAND4_X1 U19865 ( .A1(n16798), .A2(n16797), .A3(n16796), .A4(n16795), .ZN(
        n16804) );
  NOR4_X1 U19866 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16802) );
  AOI211_X1 U19867 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_16__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16801) );
  NOR4_X1 U19868 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16800) );
  NOR4_X1 U19869 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16799) );
  NAND4_X1 U19870 ( .A1(n16802), .A2(n16801), .A3(n16800), .A4(n16799), .ZN(
        n16803) );
  NOR2_X1 U19871 ( .A1(n16804), .A2(n16803), .ZN(n19102) );
  INV_X1 U19872 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16806) );
  NOR3_X1 U19873 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16807) );
  OAI21_X1 U19874 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16807), .A(n19102), .ZN(
        n16805) );
  OAI21_X1 U19875 ( .B1(n19102), .B2(n16806), .A(n16805), .ZN(P3_U2638) );
  INV_X1 U19876 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19095) );
  INV_X1 U19877 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19064) );
  AOI21_X1 U19878 ( .B1(n19095), .B2(n19064), .A(n16807), .ZN(n16809) );
  INV_X1 U19879 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16808) );
  INV_X1 U19880 ( .A(n19102), .ZN(n19097) );
  AOI22_X1 U19881 ( .A1(n19102), .A2(n16809), .B1(n16808), .B2(n19097), .ZN(
        P3_U2639) );
  INV_X1 U19882 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16812) );
  NAND2_X1 U19883 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n9777), .ZN(
        n16813) );
  INV_X1 U19884 ( .A(n16810), .ZN(n16811) );
  AOI21_X1 U19885 ( .B1(n16812), .B2(n16813), .A(n16811), .ZN(n17759) );
  OAI21_X1 U19886 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n9777), .A(
        n16813), .ZN(n17780) );
  INV_X1 U19887 ( .A(n17780), .ZN(n16876) );
  AOI21_X1 U19888 ( .B1(n21234), .B2(n17758), .A(n9777), .ZN(n17785) );
  INV_X1 U19889 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17811) );
  INV_X1 U19890 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17844) );
  INV_X1 U19891 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17906) );
  NAND2_X1 U19892 ( .A1(n17903), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16996) );
  NAND2_X1 U19893 ( .A1(n12457), .A2(n17877), .ZN(n17838) );
  NAND2_X1 U19894 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16819), .ZN(
        n16817) );
  NAND2_X1 U19895 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17823), .ZN(
        n16815) );
  NOR2_X1 U19896 ( .A1(n17811), .A2(n16815), .ZN(n16814) );
  OAI21_X1 U19897 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16814), .A(
        n17758), .ZN(n17798) );
  INV_X1 U19898 ( .A(n17798), .ZN(n16896) );
  AOI21_X1 U19899 ( .B1(n17811), .B2(n16815), .A(n16814), .ZN(n17807) );
  INV_X1 U19900 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16916) );
  INV_X1 U19901 ( .A(n17823), .ZN(n16816) );
  INV_X1 U19902 ( .A(n16815), .ZN(n17793) );
  AOI21_X1 U19903 ( .B1(n16916), .B2(n16816), .A(n17793), .ZN(n17827) );
  AOI21_X1 U19904 ( .B1(n17844), .B2(n16817), .A(n17823), .ZN(n17847) );
  OAI21_X1 U19905 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n16819), .A(
        n16817), .ZN(n16818) );
  INV_X1 U19906 ( .A(n16818), .ZN(n17859) );
  AOI21_X1 U19907 ( .B1(n17863), .B2(n17838), .A(n16819), .ZN(n17867) );
  NAND2_X1 U19908 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17877), .ZN(
        n16967) );
  INV_X1 U19909 ( .A(n16967), .ZN(n16956) );
  INV_X1 U19910 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18121) );
  NOR2_X1 U19911 ( .A1(n17919), .A2(n18121), .ZN(n17920) );
  NAND2_X1 U19912 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17920), .ZN(
        n17002) );
  INV_X1 U19913 ( .A(n17002), .ZN(n16997) );
  INV_X1 U19914 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17180) );
  AOI21_X1 U19915 ( .B1(n16997), .B2(n17180), .A(n16820), .ZN(n17005) );
  INV_X1 U19916 ( .A(n17005), .ZN(n16998) );
  OAI21_X1 U19917 ( .B1(n17144), .B2(n16956), .A(n16998), .ZN(n16957) );
  INV_X1 U19918 ( .A(n16957), .ZN(n16959) );
  NOR2_X1 U19919 ( .A1(n16936), .A2(n17144), .ZN(n16929) );
  NOR2_X1 U19920 ( .A1(n17847), .A2(n16929), .ZN(n16928) );
  NOR2_X1 U19921 ( .A1(n16928), .A2(n17144), .ZN(n16915) );
  NOR2_X1 U19922 ( .A1(n16896), .A2(n16895), .ZN(n16894) );
  NOR2_X1 U19923 ( .A1(n16894), .A2(n17144), .ZN(n16887) );
  NOR2_X1 U19924 ( .A1(n17785), .A2(n16887), .ZN(n16886) );
  NOR2_X1 U19925 ( .A1(n16886), .A2(n17144), .ZN(n16875) );
  NOR2_X1 U19926 ( .A1(n16876), .A2(n16875), .ZN(n16874) );
  NOR2_X1 U19927 ( .A1(n16874), .A2(n17144), .ZN(n16866) );
  NAND2_X1 U19928 ( .A1(n16841), .A2(n16842), .ZN(n16839) );
  NAND3_X1 U19929 ( .A1(n21075), .A2(n19123), .A3(n19111), .ZN(n18976) );
  NOR2_X1 U19930 ( .A1(n19075), .A2(n18976), .ZN(n17164) );
  INV_X1 U19931 ( .A(n17164), .ZN(n18974) );
  NOR2_X1 U19932 ( .A1(n17144), .A2(n18974), .ZN(n17039) );
  INV_X1 U19933 ( .A(n17039), .ZN(n17179) );
  NAND2_X1 U19934 ( .A1(n19122), .A2(n17642), .ZN(n16826) );
  NAND2_X1 U19935 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16828), .ZN(n16823) );
  AOI211_X4 U19936 ( .C1(n19111), .C2(n19113), .A(n16826), .B(n16823), .ZN(
        n17191) );
  NOR2_X1 U19937 ( .A1(n17169), .A2(P3_EBX_REG_3__SCAN_IN), .ZN(n17149) );
  INV_X1 U19938 ( .A(n17149), .ZN(n17133) );
  INV_X1 U19939 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17119) );
  NAND2_X1 U19940 ( .A1(n17132), .A2(n17119), .ZN(n17118) );
  INV_X1 U19941 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17335) );
  NAND2_X1 U19942 ( .A1(n17109), .A2(n17335), .ZN(n17096) );
  NAND2_X1 U19943 ( .A1(n17083), .A2(n17078), .ZN(n17077) );
  INV_X1 U19944 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17056) );
  NAND2_X1 U19945 ( .A1(n17059), .A2(n17056), .ZN(n17055) );
  INV_X1 U19946 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17032) );
  NAND2_X1 U19947 ( .A1(n17037), .A2(n17032), .ZN(n17029) );
  INV_X1 U19948 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17360) );
  NAND2_X1 U19949 ( .A1(n17016), .A2(n17360), .ZN(n17003) );
  INV_X1 U19950 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16986) );
  NAND2_X1 U19951 ( .A1(n16990), .A2(n16986), .ZN(n16985) );
  INV_X1 U19952 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16963) );
  NAND2_X1 U19953 ( .A1(n16969), .A2(n16963), .ZN(n16962) );
  INV_X1 U19954 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17277) );
  NAND2_X1 U19955 ( .A1(n16948), .A2(n17277), .ZN(n16940) );
  INV_X1 U19956 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16922) );
  NAND2_X1 U19957 ( .A1(n16927), .A2(n16922), .ZN(n16921) );
  NOR2_X1 U19958 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16921), .ZN(n16908) );
  NAND2_X1 U19959 ( .A1(n16908), .A2(n16902), .ZN(n16901) );
  NOR2_X1 U19960 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16901), .ZN(n16885) );
  INV_X1 U19961 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17233) );
  NAND2_X1 U19962 ( .A1(n16885), .A2(n17233), .ZN(n16881) );
  NOR2_X1 U19963 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16881), .ZN(n16864) );
  INV_X1 U19964 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17226) );
  NAND2_X1 U19965 ( .A1(n16864), .A2(n17226), .ZN(n16840) );
  NOR2_X1 U19966 ( .A1(n17181), .A2(n16840), .ZN(n16848) );
  INV_X1 U19967 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16833) );
  INV_X1 U19968 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19057) );
  INV_X1 U19969 ( .A(n16824), .ZN(n19110) );
  AOI211_X1 U19970 ( .C1(n19112), .C2(n19110), .A(n18988), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16827) );
  INV_X1 U19971 ( .A(n16827), .ZN(n18959) );
  INV_X1 U19972 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19045) );
  INV_X1 U19973 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19040) );
  INV_X1 U19974 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19038) );
  INV_X1 U19975 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19036) );
  INV_X1 U19976 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19023) );
  INV_X1 U19977 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19018) );
  INV_X1 U19978 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19012) );
  INV_X1 U19979 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19009) );
  INV_X1 U19980 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19005) );
  NAND2_X1 U19981 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17167) );
  NOR2_X1 U19982 ( .A1(n19000), .A2(n17167), .ZN(n17134) );
  NAND2_X1 U19983 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17134), .ZN(n17122) );
  NOR2_X1 U19984 ( .A1(n19005), .A2(n17122), .ZN(n17117) );
  NAND2_X1 U19985 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17117), .ZN(n17085) );
  NOR3_X1 U19986 ( .A1(n19012), .A2(n19009), .A3(n17085), .ZN(n17061) );
  NAND4_X1 U19987 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n17061), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n17041) );
  NOR2_X1 U19988 ( .A1(n19018), .A2(n17041), .ZN(n17026) );
  NAND2_X1 U19989 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17026), .ZN(n17013) );
  NOR2_X1 U19990 ( .A1(n19023), .A2(n17013), .ZN(n16954) );
  INV_X1 U19991 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19032) );
  INV_X1 U19992 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19030) );
  NAND3_X1 U19993 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16955) );
  NOR3_X1 U19994 ( .A1(n19032), .A2(n19030), .A3(n16955), .ZN(n16945) );
  NAND3_X1 U19995 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16954), .A3(n16945), 
        .ZN(n16925) );
  NOR4_X1 U19996 ( .A1(n19040), .A2(n19038), .A3(n19036), .A4(n16925), .ZN(
        n16907) );
  NAND2_X1 U19997 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16907), .ZN(n16898) );
  NOR2_X1 U19998 ( .A1(n19045), .A2(n16898), .ZN(n16884) );
  NAND2_X1 U19999 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16884), .ZN(n16835) );
  NOR2_X1 U20000 ( .A1(n17182), .A2(n16835), .ZN(n16880) );
  NAND4_X1 U20001 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16880), .ZN(n16834) );
  NOR3_X1 U20002 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19057), .A3(n16834), 
        .ZN(n16832) );
  NOR2_X1 U20003 ( .A1(n19068), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18971) );
  INV_X1 U20004 ( .A(n18971), .ZN(n18964) );
  NOR2_X1 U20005 ( .A1(n18385), .A2(n17164), .ZN(n16825) );
  INV_X1 U20006 ( .A(n19122), .ZN(n19126) );
  NOR2_X2 U20007 ( .A1(n19068), .A2(n17177), .ZN(n17146) );
  INV_X1 U20008 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16829) );
  AOI211_X4 U20009 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16828), .A(n16827), .B(
        n16826), .ZN(n17192) );
  OAI22_X1 U20010 ( .A1(n16830), .A2(n17178), .B1(n16829), .B2(n17157), .ZN(
        n16831) );
  AOI211_X1 U20011 ( .C1(n16848), .C2(n16833), .A(n16832), .B(n16831), .ZN(
        n16838) );
  NOR2_X1 U20012 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16834), .ZN(n16846) );
  NAND3_X1 U20013 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16836) );
  OR2_X1 U20014 ( .A1(n16835), .A2(n17177), .ZN(n16863) );
  NOR2_X1 U20015 ( .A1(n17168), .A2(n17177), .ZN(n16979) );
  INV_X1 U20016 ( .A(n16979), .ZN(n17189) );
  OAI21_X1 U20017 ( .B1(n16836), .B2(n16863), .A(n17189), .ZN(n16843) );
  INV_X1 U20018 ( .A(n16843), .ZN(n16859) );
  OAI21_X1 U20019 ( .B1(n16846), .B2(n16859), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16837) );
  OAI211_X1 U20020 ( .C1(n16839), .C2(n17179), .A(n16838), .B(n16837), .ZN(
        P3_U2640) );
  NAND2_X1 U20021 ( .A1(n17191), .A2(n16840), .ZN(n16852) );
  XOR2_X1 U20022 ( .A(n16842), .B(n16841), .Z(n16847) );
  OAI22_X1 U20023 ( .A1(n16844), .A2(n17178), .B1(n19057), .B2(n16843), .ZN(
        n16845) );
  AOI211_X1 U20024 ( .C1(n16847), .C2(n17164), .A(n16846), .B(n16845), .ZN(
        n16850) );
  OAI21_X1 U20025 ( .B1(n17192), .B2(n16848), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16849) );
  OAI211_X1 U20026 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16852), .A(n16850), .B(
        n16849), .ZN(P3_U2641) );
  NAND2_X1 U20027 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16870) );
  NOR2_X1 U20028 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16870), .ZN(n16851) );
  AOI22_X1 U20029 ( .A1(n17192), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n16880), 
        .B2(n16851), .ZN(n16861) );
  INV_X1 U20030 ( .A(n16864), .ZN(n16853) );
  AOI21_X1 U20031 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16853), .A(n16852), .ZN(
        n16858) );
  AOI211_X1 U20032 ( .C1(n16856), .C2(n16855), .A(n16854), .B(n18974), .ZN(
        n16857) );
  AOI211_X1 U20033 ( .C1(n16859), .C2(P3_REIP_REG_29__SCAN_IN), .A(n16858), 
        .B(n16857), .ZN(n16860) );
  OAI211_X1 U20034 ( .C1(n16862), .C2(n17178), .A(n16861), .B(n16860), .ZN(
        P3_U2642) );
  AOI22_X1 U20035 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17146), .B1(
        n17192), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16873) );
  NAND2_X1 U20036 ( .A1(n17189), .A2(n16863), .ZN(n16892) );
  INV_X1 U20037 ( .A(n16892), .ZN(n16869) );
  AOI211_X1 U20038 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16881), .A(n16864), .B(
        n17181), .ZN(n16868) );
  AOI211_X1 U20039 ( .C1(n17759), .C2(n16866), .A(n16865), .B(n18974), .ZN(
        n16867) );
  AOI211_X1 U20040 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16869), .A(n16868), 
        .B(n16867), .ZN(n16872) );
  OAI211_X1 U20041 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16880), .B(n16870), .ZN(n16871) );
  NAND3_X1 U20042 ( .A1(n16873), .A2(n16872), .A3(n16871), .ZN(P3_U2643) );
  INV_X1 U20043 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19049) );
  AOI211_X1 U20044 ( .C1(n16876), .C2(n16875), .A(n16874), .B(n18974), .ZN(
        n16879) );
  INV_X1 U20045 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16877) );
  OAI22_X1 U20046 ( .A1(n16877), .A2(n17178), .B1(n17157), .B2(n17233), .ZN(
        n16878) );
  AOI211_X1 U20047 ( .C1(n16880), .C2(n19049), .A(n16879), .B(n16878), .ZN(
        n16883) );
  OAI211_X1 U20048 ( .C1(n16885), .C2(n17233), .A(n17191), .B(n16881), .ZN(
        n16882) );
  OAI211_X1 U20049 ( .C1(n16892), .C2(n19049), .A(n16883), .B(n16882), .ZN(
        P3_U2644) );
  AOI21_X1 U20050 ( .B1(n17168), .B2(n16884), .A(P3_REIP_REG_26__SCAN_IN), 
        .ZN(n16893) );
  AOI22_X1 U20051 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17146), .B1(
        n17192), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16891) );
  AOI211_X1 U20052 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16901), .A(n16885), .B(
        n17181), .ZN(n16889) );
  AOI211_X1 U20053 ( .C1(n17785), .C2(n16887), .A(n16886), .B(n18974), .ZN(
        n16888) );
  NOR2_X1 U20054 ( .A1(n16889), .A2(n16888), .ZN(n16890) );
  OAI211_X1 U20055 ( .C1(n16893), .C2(n16892), .A(n16891), .B(n16890), .ZN(
        P3_U2645) );
  INV_X1 U20056 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19042) );
  OAI21_X1 U20057 ( .B1(n16907), .B2(n17182), .A(n17190), .ZN(n16920) );
  AOI21_X1 U20058 ( .B1(n17168), .B2(n19042), .A(n16920), .ZN(n16905) );
  AOI211_X1 U20059 ( .C1(n16896), .C2(n16895), .A(n16894), .B(n18974), .ZN(
        n16900) );
  NAND2_X1 U20060 ( .A1(n17168), .A2(n19045), .ZN(n16897) );
  OAI22_X1 U20061 ( .A1(n17157), .A2(n16902), .B1(n16898), .B2(n16897), .ZN(
        n16899) );
  AOI211_X1 U20062 ( .C1(n17146), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16900), .B(n16899), .ZN(n16904) );
  OAI211_X1 U20063 ( .C1(n16908), .C2(n16902), .A(n17191), .B(n16901), .ZN(
        n16903) );
  OAI211_X1 U20064 ( .C1(n16905), .C2(n19045), .A(n16904), .B(n16903), .ZN(
        P3_U2646) );
  NOR2_X1 U20065 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17182), .ZN(n16906) );
  AOI22_X1 U20066 ( .A1(n17192), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16907), 
        .B2(n16906), .ZN(n16913) );
  AOI211_X1 U20067 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16921), .A(n16908), .B(
        n17181), .ZN(n16911) );
  AOI211_X1 U20068 ( .C1(n17807), .C2(n9768), .A(n16909), .B(n18974), .ZN(
        n16910) );
  AOI211_X1 U20069 ( .C1(n16920), .C2(P3_REIP_REG_24__SCAN_IN), .A(n16911), 
        .B(n16910), .ZN(n16912) );
  OAI211_X1 U20070 ( .C1(n17811), .C2(n17178), .A(n16913), .B(n16912), .ZN(
        P3_U2647) );
  NOR2_X1 U20071 ( .A1(n17182), .A2(n16925), .ZN(n16926) );
  NAND2_X1 U20072 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16926), .ZN(n16935) );
  OAI21_X1 U20073 ( .B1(n19038), .B2(n16935), .A(n19040), .ZN(n16919) );
  AOI211_X1 U20074 ( .C1(n17827), .C2(n16915), .A(n16914), .B(n18974), .ZN(
        n16918) );
  OAI22_X1 U20075 ( .A1(n16916), .A2(n17178), .B1(n17157), .B2(n16922), .ZN(
        n16917) );
  AOI211_X1 U20076 ( .C1(n16920), .C2(n16919), .A(n16918), .B(n16917), .ZN(
        n16924) );
  OAI211_X1 U20077 ( .C1(n16927), .C2(n16922), .A(n17191), .B(n16921), .ZN(
        n16923) );
  NAND2_X1 U20078 ( .A1(n16924), .A2(n16923), .ZN(P3_U2648) );
  AOI22_X1 U20079 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17146), .B1(
        n17192), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16934) );
  AOI21_X1 U20080 ( .B1(n17168), .B2(n16925), .A(n17177), .ZN(n16953) );
  NAND2_X1 U20081 ( .A1(n16926), .A2(n19036), .ZN(n16942) );
  AOI21_X1 U20082 ( .B1(n16953), .B2(n16942), .A(n19038), .ZN(n16932) );
  AOI211_X1 U20083 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16940), .A(n16927), .B(
        n17181), .ZN(n16931) );
  AOI211_X1 U20084 ( .C1(n17847), .C2(n16929), .A(n16928), .B(n18974), .ZN(
        n16930) );
  NOR3_X1 U20085 ( .A1(n16932), .A2(n16931), .A3(n16930), .ZN(n16933) );
  OAI211_X1 U20086 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16935), .A(n16934), 
        .B(n16933), .ZN(P3_U2649) );
  INV_X1 U20087 ( .A(n16953), .ZN(n16939) );
  AOI211_X1 U20088 ( .C1(n17859), .C2(n9782), .A(n16936), .B(n18974), .ZN(
        n16938) );
  INV_X1 U20089 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17856) );
  OAI22_X1 U20090 ( .A1(n17856), .A2(n17178), .B1(n17157), .B2(n17277), .ZN(
        n16937) );
  AOI211_X1 U20091 ( .C1(n16939), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16938), 
        .B(n16937), .ZN(n16943) );
  OAI211_X1 U20092 ( .C1(n16948), .C2(n17277), .A(n17191), .B(n16940), .ZN(
        n16941) );
  NAND3_X1 U20093 ( .A1(n16943), .A2(n16942), .A3(n16941), .ZN(P3_U2650) );
  INV_X1 U20094 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19034) );
  NAND2_X1 U20095 ( .A1(n17168), .A2(n16954), .ZN(n17007) );
  NOR2_X1 U20096 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17007), .ZN(n16944) );
  AOI22_X1 U20097 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17146), .B1(
        n16945), .B2(n16944), .ZN(n16952) );
  AOI211_X1 U20098 ( .C1(n17867), .C2(n16947), .A(n16946), .B(n18974), .ZN(
        n16950) );
  AOI211_X1 U20099 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16962), .A(n16948), .B(
        n17181), .ZN(n16949) );
  AOI211_X1 U20100 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17192), .A(n16950), .B(
        n16949), .ZN(n16951) );
  OAI211_X1 U20101 ( .C1(n19034), .C2(n16953), .A(n16952), .B(n16951), .ZN(
        P3_U2651) );
  AOI22_X1 U20102 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17146), .B1(
        n17192), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16966) );
  NAND2_X1 U20103 ( .A1(n16954), .A2(n17190), .ZN(n17012) );
  NOR2_X1 U20104 ( .A1(n16955), .A2(n17012), .ZN(n16978) );
  AOI21_X1 U20105 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16978), .A(n16979), 
        .ZN(n16971) );
  NAND2_X1 U20106 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16991) );
  NOR2_X1 U20107 ( .A1(n16991), .A2(n17007), .ZN(n16983) );
  NAND2_X1 U20108 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16983), .ZN(n16970) );
  NOR2_X1 U20109 ( .A1(n19030), .A2(n16970), .ZN(n16961) );
  OAI21_X1 U20110 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16956), .A(
        n17838), .ZN(n16958) );
  INV_X1 U20111 ( .A(n16958), .ZN(n17878) );
  AOI221_X1 U20112 ( .B1(n16959), .B2(n16958), .C1(n16957), .C2(n17878), .A(
        n18974), .ZN(n16960) );
  AOI221_X1 U20113 ( .B1(n16971), .B2(P3_REIP_REG_19__SCAN_IN), .C1(n16961), 
        .C2(n19032), .A(n16960), .ZN(n16965) );
  OAI211_X1 U20114 ( .C1(n16969), .C2(n16963), .A(n17191), .B(n16962), .ZN(
        n16964) );
  NAND4_X1 U20115 ( .A1(n16966), .A2(n16965), .A3(n18384), .A4(n16964), .ZN(
        P3_U2652) );
  OAI21_X1 U20116 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17877), .A(
        n16967), .ZN(n17888) );
  NOR2_X1 U20117 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18121), .ZN(
        n17166) );
  AOI21_X1 U20118 ( .B1(n17876), .B2(n17166), .A(n17144), .ZN(n16968) );
  XOR2_X1 U20119 ( .A(n17888), .B(n16968), .Z(n16977) );
  AOI211_X1 U20120 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16985), .A(n16969), .B(
        n17181), .ZN(n16975) );
  INV_X1 U20121 ( .A(n16970), .ZN(n16972) );
  OAI21_X1 U20122 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16972), .A(n16971), 
        .ZN(n16973) );
  OAI211_X1 U20123 ( .C1(n17157), .C2(n17305), .A(n18384), .B(n16973), .ZN(
        n16974) );
  AOI211_X1 U20124 ( .C1(n17146), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16975), .B(n16974), .ZN(n16976) );
  OAI21_X1 U20125 ( .B1(n18974), .B2(n16977), .A(n16976), .ZN(P3_U2653) );
  AOI22_X1 U20126 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17146), .B1(
        n17192), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16989) );
  NOR2_X1 U20127 ( .A1(n16979), .A2(n16978), .ZN(n16984) );
  INV_X1 U20128 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19028) );
  AOI21_X1 U20129 ( .B1(n17906), .B2(n16996), .A(n17877), .ZN(n17908) );
  AOI21_X1 U20130 ( .B1(n17903), .B2(n17166), .A(n17144), .ZN(n16981) );
  OAI21_X1 U20131 ( .B1(n17908), .B2(n16981), .A(n17164), .ZN(n16980) );
  AOI21_X1 U20132 ( .B1(n17908), .B2(n16981), .A(n16980), .ZN(n16982) );
  AOI221_X1 U20133 ( .B1(n16984), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16983), 
        .C2(n19028), .A(n16982), .ZN(n16988) );
  OAI211_X1 U20134 ( .C1(n16990), .C2(n16986), .A(n17191), .B(n16985), .ZN(
        n16987) );
  NAND4_X1 U20135 ( .A1(n16989), .A2(n16988), .A3(n18384), .A4(n16987), .ZN(
        P3_U2654) );
  NAND2_X1 U20136 ( .A1(n17189), .A2(n17012), .ZN(n17024) );
  INV_X1 U20137 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19026) );
  AOI211_X1 U20138 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17003), .A(n16990), .B(
        n17181), .ZN(n16995) );
  INV_X1 U20139 ( .A(n17007), .ZN(n16992) );
  OAI211_X1 U20140 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16992), .B(n16991), .ZN(n16993) );
  OAI211_X1 U20141 ( .C1(n17917), .C2(n17178), .A(n18384), .B(n16993), .ZN(
        n16994) );
  AOI211_X1 U20142 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17192), .A(n16995), .B(
        n16994), .ZN(n17001) );
  OAI21_X1 U20143 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16997), .A(
        n16996), .ZN(n17922) );
  INV_X1 U20144 ( .A(n17922), .ZN(n16999) );
  OAI221_X1 U20145 ( .B1(n17005), .B2(n16999), .C1(n16998), .C2(n17922), .A(
        n17164), .ZN(n17000) );
  OAI211_X1 U20146 ( .C1(n17024), .C2(n19026), .A(n17001), .B(n17000), .ZN(
        P3_U2655) );
  OAI21_X1 U20147 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17920), .A(
        n17002), .ZN(n17928) );
  AOI21_X1 U20148 ( .B1(n9942), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18974), .ZN(n17184) );
  OAI21_X1 U20149 ( .B1(n17144), .B2(n17918), .A(n17184), .ZN(n17011) );
  OAI211_X1 U20150 ( .C1(n17016), .C2(n17360), .A(n17191), .B(n17003), .ZN(
        n17004) );
  OAI211_X1 U20151 ( .C1(n17157), .C2(n17360), .A(n18384), .B(n17004), .ZN(
        n17009) );
  INV_X1 U20152 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19024) );
  NAND3_X1 U20153 ( .A1(n17005), .A2(n17164), .A3(n17928), .ZN(n17006) );
  OAI221_X1 U20154 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n17007), .C1(n19024), 
        .C2(n17024), .A(n17006), .ZN(n17008) );
  AOI211_X1 U20155 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17146), .A(
        n17009), .B(n17008), .ZN(n17010) );
  OAI21_X1 U20156 ( .B1(n17928), .B2(n17011), .A(n17010), .ZN(P3_U2656) );
  INV_X1 U20157 ( .A(n17012), .ZN(n17014) );
  NOR3_X1 U20158 ( .A1(n17014), .A2(n17013), .A3(n17182), .ZN(n17015) );
  AOI211_X1 U20159 ( .C1(n17192), .C2(P3_EBX_REG_14__SCAN_IN), .A(n18385), .B(
        n17015), .ZN(n17023) );
  INV_X1 U20160 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17964) );
  INV_X1 U20161 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17963) );
  INV_X1 U20162 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18014) );
  INV_X1 U20163 ( .A(n18029), .ZN(n18046) );
  NOR3_X1 U20164 ( .A1(n18046), .A2(n18048), .A3(n18121), .ZN(n17094) );
  NAND2_X1 U20165 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17094), .ZN(
        n17086) );
  NOR2_X1 U20166 ( .A1(n18014), .A2(n17086), .ZN(n17072) );
  NAND2_X1 U20167 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17072), .ZN(
        n17062) );
  NOR2_X1 U20168 ( .A1(n17995), .A2(n17062), .ZN(n17049) );
  INV_X1 U20169 ( .A(n17049), .ZN(n17961) );
  NOR3_X1 U20170 ( .A1(n17964), .A2(n17963), .A3(n17961), .ZN(n17017) );
  INV_X1 U20171 ( .A(n17017), .ZN(n17025) );
  AOI21_X1 U20172 ( .B1(n17947), .B2(n17025), .A(n17920), .ZN(n17949) );
  INV_X1 U20173 ( .A(n17949), .ZN(n17021) );
  AOI21_X1 U20174 ( .B1(n17017), .B2(n17180), .A(n17179), .ZN(n17035) );
  AOI211_X1 U20175 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17029), .A(n17016), .B(
        n17181), .ZN(n17020) );
  OAI221_X1 U20176 ( .B1(n17144), .B2(n17017), .C1(n17144), .C2(n17180), .A(
        n17164), .ZN(n17018) );
  OAI22_X1 U20177 ( .A1(n17018), .A2(n17021), .B1(n17947), .B2(n17178), .ZN(
        n17019) );
  AOI211_X1 U20178 ( .C1(n17021), .C2(n17035), .A(n17020), .B(n17019), .ZN(
        n17022) );
  OAI211_X1 U20179 ( .C1(n19023), .C2(n17024), .A(n17023), .B(n17022), .ZN(
        P3_U2657) );
  INV_X1 U20180 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19020) );
  AOI21_X1 U20181 ( .B1(n17168), .B2(n17041), .A(n17177), .ZN(n17052) );
  NAND2_X1 U20182 ( .A1(n17168), .A2(n19018), .ZN(n17040) );
  NOR2_X1 U20183 ( .A1(n17964), .A2(n17961), .ZN(n17038) );
  OAI21_X1 U20184 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17038), .A(
        n17025), .ZN(n17966) );
  NAND3_X1 U20185 ( .A1(n17168), .A2(n17026), .A3(n19020), .ZN(n17027) );
  OAI211_X1 U20186 ( .C1(n17963), .C2(n17178), .A(n18384), .B(n17027), .ZN(
        n17034) );
  INV_X1 U20187 ( .A(n17966), .ZN(n17028) );
  OAI211_X1 U20188 ( .C1(n17144), .C2(n17963), .A(n17028), .B(n17184), .ZN(
        n17031) );
  OAI211_X1 U20189 ( .C1(n17037), .C2(n17032), .A(n17191), .B(n17029), .ZN(
        n17030) );
  OAI211_X1 U20190 ( .C1(n17032), .C2(n17157), .A(n17031), .B(n17030), .ZN(
        n17033) );
  AOI211_X1 U20191 ( .C1(n17966), .C2(n17035), .A(n17034), .B(n17033), .ZN(
        n17036) );
  OAI221_X1 U20192 ( .B1(n19020), .B2(n17052), .C1(n19020), .C2(n17040), .A(
        n17036), .ZN(P3_U2658) );
  AOI211_X1 U20193 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17055), .A(n17037), .B(
        n17181), .ZN(n17046) );
  AOI21_X1 U20194 ( .B1(n17964), .B2(n17961), .A(n17038), .ZN(n17978) );
  OAI21_X1 U20195 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17964), .A(
        n17039), .ZN(n17042) );
  OAI22_X1 U20196 ( .A1(n17978), .A2(n17042), .B1(n17041), .B2(n17040), .ZN(
        n17045) );
  OAI22_X1 U20197 ( .A1(n17964), .A2(n17178), .B1(n17157), .B2(n17043), .ZN(
        n17044) );
  NOR4_X1 U20198 ( .A1(n18385), .A2(n17046), .A3(n17045), .A4(n17044), .ZN(
        n17048) );
  OAI211_X1 U20199 ( .C1(n17049), .C2(n17144), .A(n17978), .B(n17184), .ZN(
        n17047) );
  OAI211_X1 U20200 ( .C1(n17052), .C2(n19018), .A(n17048), .B(n17047), .ZN(
        P3_U2659) );
  INV_X1 U20201 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n21188) );
  INV_X1 U20202 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19013) );
  NOR2_X1 U20203 ( .A1(n21188), .A2(n19013), .ZN(n17066) );
  NOR4_X1 U20204 ( .A1(n17182), .A2(n19012), .A3(n19009), .A4(n17085), .ZN(
        n17071) );
  AOI21_X1 U20205 ( .B1(n17066), .B2(n17071), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17053) );
  AOI21_X1 U20206 ( .B1(n17995), .B2(n17062), .A(n17049), .ZN(n17993) );
  OAI21_X1 U20207 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17062), .A(
        n9942), .ZN(n17050) );
  XOR2_X1 U20208 ( .A(n17993), .B(n17050), .Z(n17051) );
  OAI22_X1 U20209 ( .A1(n17053), .A2(n17052), .B1(n18974), .B2(n17051), .ZN(
        n17054) );
  AOI211_X1 U20210 ( .C1(n17192), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18385), .B(
        n17054), .ZN(n17058) );
  OAI211_X1 U20211 ( .C1(n17059), .C2(n17056), .A(n17191), .B(n17055), .ZN(
        n17057) );
  OAI211_X1 U20212 ( .C1(n17178), .C2(n17995), .A(n17058), .B(n17057), .ZN(
        P3_U2660) );
  INV_X1 U20213 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18009) );
  AOI211_X1 U20214 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17077), .A(n17059), .B(
        n17181), .ZN(n17060) );
  AOI211_X1 U20215 ( .C1(n17192), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18385), .B(
        n17060), .ZN(n17070) );
  OAI21_X1 U20216 ( .B1(n17061), .B2(n17182), .A(n17190), .ZN(n17084) );
  OAI21_X1 U20217 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17072), .A(
        n17062), .ZN(n18002) );
  AOI21_X1 U20218 ( .B1(n17180), .B2(n17072), .A(n17144), .ZN(n17063) );
  INV_X1 U20219 ( .A(n17063), .ZN(n17075) );
  OAI21_X1 U20220 ( .B1(n18002), .B2(n17075), .A(n17164), .ZN(n17064) );
  AOI21_X1 U20221 ( .B1(n18002), .B2(n17075), .A(n17064), .ZN(n17068) );
  INV_X1 U20222 ( .A(n17071), .ZN(n17065) );
  AOI211_X1 U20223 ( .C1(n21188), .C2(n19013), .A(n17066), .B(n17065), .ZN(
        n17067) );
  AOI211_X1 U20224 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n17084), .A(n17068), 
        .B(n17067), .ZN(n17069) );
  OAI211_X1 U20225 ( .C1(n18009), .C2(n17178), .A(n17070), .B(n17069), .ZN(
        P3_U2661) );
  AOI22_X1 U20226 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17146), .B1(
        n17192), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20227 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17084), .B1(n17071), 
        .B2(n19013), .ZN(n17081) );
  AOI21_X1 U20228 ( .B1(n18014), .B2(n17086), .A(n17072), .ZN(n18018) );
  INV_X1 U20229 ( .A(n18018), .ZN(n17074) );
  NAND2_X1 U20230 ( .A1(n18029), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17104) );
  NOR2_X1 U20231 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17104), .ZN(
        n17107) );
  NAND3_X1 U20232 ( .A1(n18027), .A2(n17107), .A3(n18014), .ZN(n17073) );
  OAI221_X1 U20233 ( .B1(n18018), .B2(n17075), .C1(n17074), .C2(n9942), .A(
        n17073), .ZN(n17076) );
  AOI21_X1 U20234 ( .B1(n17164), .B2(n17076), .A(n18385), .ZN(n17080) );
  OAI211_X1 U20235 ( .C1(n17083), .C2(n17078), .A(n17191), .B(n17077), .ZN(
        n17079) );
  NAND4_X1 U20236 ( .A1(n17082), .A2(n17081), .A3(n17080), .A4(n17079), .ZN(
        P3_U2662) );
  AOI211_X1 U20237 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17096), .A(n17083), .B(
        n17181), .ZN(n17092) );
  INV_X1 U20238 ( .A(n17084), .ZN(n17090) );
  NOR2_X1 U20239 ( .A1(n17182), .A2(n17085), .ZN(n17100) );
  AOI21_X1 U20240 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n17100), .A(
        P3_REIP_REG_8__SCAN_IN), .ZN(n17089) );
  AOI21_X1 U20241 ( .B1(n17094), .B2(n17180), .A(n17144), .ZN(n17087) );
  OAI21_X1 U20242 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17094), .A(
        n17086), .ZN(n18033) );
  XOR2_X1 U20243 ( .A(n17087), .B(n18033), .Z(n17088) );
  OAI22_X1 U20244 ( .A1(n17090), .A2(n17089), .B1(n18974), .B2(n17088), .ZN(
        n17091) );
  AOI211_X1 U20245 ( .C1(n17146), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17092), .B(n17091), .ZN(n17093) );
  OAI211_X1 U20246 ( .C1(n17157), .C2(n17451), .A(n17093), .B(n18384), .ZN(
        P3_U2663) );
  AOI21_X1 U20247 ( .B1(n18048), .B2(n17104), .A(n17094), .ZN(n18052) );
  NOR2_X1 U20248 ( .A1(n17107), .A2(n17144), .ZN(n17095) );
  XNOR2_X1 U20249 ( .A(n18052), .B(n17095), .ZN(n17103) );
  AOI22_X1 U20250 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17146), .B1(
        n17192), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n17102) );
  OAI221_X1 U20251 ( .B1(n17182), .B2(P3_REIP_REG_6__SCAN_IN), .C1(n17182), 
        .C2(n17117), .A(n17190), .ZN(n17099) );
  OAI211_X1 U20252 ( .C1(n17109), .C2(n17335), .A(n17191), .B(n17096), .ZN(
        n17097) );
  NAND2_X1 U20253 ( .A1(n18384), .A2(n17097), .ZN(n17098) );
  AOI221_X1 U20254 ( .B1(n17100), .B2(n19009), .C1(n17099), .C2(
        P3_REIP_REG_7__SCAN_IN), .A(n17098), .ZN(n17101) );
  OAI211_X1 U20255 ( .C1(n18974), .C2(n17103), .A(n17102), .B(n17101), .ZN(
        P3_U2664) );
  NOR2_X1 U20256 ( .A1(n18061), .A2(n18121), .ZN(n17115) );
  OAI21_X1 U20257 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17115), .A(
        n17104), .ZN(n18063) );
  OAI21_X1 U20258 ( .B1(n17144), .B2(n18062), .A(n17184), .ZN(n17114) );
  INV_X1 U20259 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17457) );
  INV_X1 U20260 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19007) );
  NAND3_X1 U20261 ( .A1(n17168), .A2(n17117), .A3(n19007), .ZN(n17105) );
  OAI211_X1 U20262 ( .C1(n17157), .C2(n17457), .A(n18384), .B(n17105), .ZN(
        n17106) );
  AOI21_X1 U20263 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17146), .A(
        n17106), .ZN(n17113) );
  OAI21_X1 U20264 ( .B1(n17117), .B2(n17182), .A(n17190), .ZN(n17124) );
  INV_X1 U20265 ( .A(n18063), .ZN(n17108) );
  NOR3_X1 U20266 ( .A1(n17108), .A2(n17107), .A3(n17179), .ZN(n17111) );
  AOI211_X1 U20267 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17118), .A(n17109), .B(
        n17181), .ZN(n17110) );
  AOI211_X1 U20268 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n17124), .A(n17111), .B(
        n17110), .ZN(n17112) );
  OAI211_X1 U20269 ( .C1(n18063), .C2(n17114), .A(n17113), .B(n17112), .ZN(
        P3_U2665) );
  AOI21_X1 U20270 ( .B1(n18073), .B2(n17166), .A(n17144), .ZN(n17130) );
  NOR3_X1 U20271 ( .A1(n18085), .A2(n18093), .A3(n18121), .ZN(n17128) );
  INV_X1 U20272 ( .A(n17115), .ZN(n17116) );
  OAI21_X1 U20273 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17128), .A(
        n17116), .ZN(n18076) );
  XOR2_X1 U20274 ( .A(n17130), .B(n18076), .Z(n17127) );
  AOI22_X1 U20275 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17146), .B1(
        n17192), .B2(P3_EBX_REG_5__SCAN_IN), .ZN(n17126) );
  OR2_X1 U20276 ( .A1(n17182), .A2(n17117), .ZN(n17121) );
  OAI211_X1 U20277 ( .C1(n17132), .C2(n17119), .A(n17191), .B(n17118), .ZN(
        n17120) );
  OAI211_X1 U20278 ( .C1(n17122), .C2(n17121), .A(n18384), .B(n17120), .ZN(
        n17123) );
  AOI21_X1 U20279 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n17124), .A(n17123), .ZN(
        n17125) );
  OAI211_X1 U20280 ( .C1(n18974), .C2(n17127), .A(n17126), .B(n17125), .ZN(
        P3_U2666) );
  NOR2_X1 U20281 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18085), .ZN(
        n17131) );
  OR2_X1 U20282 ( .A1(n18085), .A2(n18121), .ZN(n17145) );
  AOI21_X1 U20283 ( .B1(n18093), .B2(n17145), .A(n17128), .ZN(n18090) );
  INV_X1 U20284 ( .A(n18090), .ZN(n17129) );
  AOI22_X1 U20285 ( .A1(n17166), .A2(n17131), .B1(n17130), .B2(n17129), .ZN(
        n17143) );
  NOR2_X1 U20286 ( .A1(n9942), .A2(n18974), .ZN(n17162) );
  AOI211_X1 U20287 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17133), .A(n17132), .B(
        n17181), .ZN(n17141) );
  NAND2_X1 U20288 ( .A1(n17168), .A2(n17134), .ZN(n17139) );
  INV_X1 U20289 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19003) );
  OAI21_X1 U20290 ( .B1(n17182), .B2(n17134), .A(n17190), .ZN(n17135) );
  INV_X1 U20291 ( .A(n17135), .ZN(n17150) );
  NAND2_X1 U20292 ( .A1(n18475), .A2(n19122), .ZN(n17188) );
  INV_X1 U20293 ( .A(n17188), .ZN(n19129) );
  OAI22_X1 U20294 ( .A1(n18093), .A2(n17178), .B1(n17157), .B2(n17136), .ZN(
        n17137) );
  AOI221_X1 U20295 ( .B1(n17319), .B2(n19129), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n19129), .A(n17137), .ZN(
        n17138) );
  OAI221_X1 U20296 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n17139), .C1(n19003), 
        .C2(n17150), .A(n17138), .ZN(n17140) );
  AOI211_X1 U20297 ( .C1(n17162), .C2(n18090), .A(n17141), .B(n17140), .ZN(
        n17142) );
  OAI211_X1 U20298 ( .C1(n17143), .C2(n18974), .A(n17142), .B(n18384), .ZN(
        P3_U2667) );
  INV_X1 U20299 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17158) );
  NOR2_X1 U20300 ( .A1(n17158), .A2(n18121), .ZN(n17156) );
  AOI21_X1 U20301 ( .B1(n17156), .B2(n17180), .A(n17144), .ZN(n17163) );
  OAI21_X1 U20302 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17156), .A(
        n17145), .ZN(n18100) );
  XOR2_X1 U20303 ( .A(n17163), .B(n18100), .Z(n17155) );
  AOI22_X1 U20304 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n17146), .B1(
        n17192), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n17154) );
  NAND2_X1 U20305 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18922) );
  NOR2_X1 U20306 ( .A1(n17147), .A2(n18922), .ZN(n17159) );
  OAI21_X1 U20307 ( .B1(n17159), .B2(n19072), .A(n17148), .ZN(n19069) );
  AOI211_X1 U20308 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n17169), .A(n17149), .B(
        n17181), .ZN(n17152) );
  AOI221_X1 U20309 ( .B1(n17182), .B2(n19000), .C1(n17167), .C2(n19000), .A(
        n17150), .ZN(n17151) );
  AOI211_X1 U20310 ( .C1(n19129), .C2(n19069), .A(n17152), .B(n17151), .ZN(
        n17153) );
  OAI211_X1 U20311 ( .C1(n18974), .C2(n17155), .A(n17154), .B(n17153), .ZN(
        P3_U2668) );
  AOI21_X1 U20312 ( .B1(n17158), .B2(n18121), .A(n17156), .ZN(n18109) );
  INV_X1 U20313 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17473) );
  OAI22_X1 U20314 ( .A1(n17158), .A2(n17178), .B1(n17157), .B2(n17473), .ZN(
        n17161) );
  INV_X1 U20315 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18998) );
  AND2_X1 U20316 ( .A1(n12320), .A2(n17176), .ZN(n18923) );
  OR2_X1 U20317 ( .A1(n18923), .A2(n17159), .ZN(n19076) );
  OAI22_X1 U20318 ( .A1(n18998), .A2(n17190), .B1(n19076), .B2(n17188), .ZN(
        n17160) );
  AOI211_X1 U20319 ( .C1(n18109), .C2(n17162), .A(n17161), .B(n17160), .ZN(
        n17174) );
  INV_X1 U20320 ( .A(n18109), .ZN(n17165) );
  OAI211_X1 U20321 ( .C1(n17166), .C2(n17165), .A(n17164), .B(n17163), .ZN(
        n17173) );
  OAI211_X1 U20322 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17168), .B(n17167), .ZN(n17172) );
  NOR2_X1 U20323 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17170) );
  OAI211_X1 U20324 ( .C1(n17170), .C2(n17473), .A(n17191), .B(n17169), .ZN(
        n17171) );
  NAND4_X1 U20325 ( .A1(n17174), .A2(n17173), .A3(n17172), .A4(n17171), .ZN(
        P3_U2669) );
  NAND2_X1 U20326 ( .A1(n17176), .A2(n17175), .ZN(n19083) );
  AOI22_X1 U20327 ( .A1(n17192), .A2(P3_EBX_REG_1__SCAN_IN), .B1(
        P3_REIP_REG_1__SCAN_IN), .B2(n17177), .ZN(n17187) );
  OAI21_X1 U20328 ( .B1(n17180), .B2(n17179), .A(n17178), .ZN(n17185) );
  NAND2_X1 U20329 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17474) );
  OAI21_X1 U20330 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17474), .ZN(n17480) );
  OAI22_X1 U20331 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17182), .B1(n17181), 
        .B2(n17480), .ZN(n17183) );
  AOI221_X1 U20332 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17185), .C1(
        n18121), .C2(n17184), .A(n17183), .ZN(n17186) );
  OAI211_X1 U20333 ( .C1(n19083), .C2(n17188), .A(n17187), .B(n17186), .ZN(
        P3_U2670) );
  AOI22_X1 U20334 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17189), .B1(n19129), 
        .B2(n17147), .ZN(n17195) );
  NAND3_X1 U20335 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19078), .A3(
        n17190), .ZN(n17194) );
  OAI21_X1 U20336 ( .B1(n17192), .B2(n17191), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n17193) );
  NAND3_X1 U20337 ( .A1(n17195), .A2(n17194), .A3(n17193), .ZN(P3_U2671) );
  AOI22_X1 U20338 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n16181), .ZN(n17200) );
  AOI22_X1 U20339 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17392), .ZN(n17199) );
  AOI22_X1 U20340 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17423), .ZN(n17198) );
  AOI22_X1 U20341 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17197) );
  NAND4_X1 U20342 ( .A1(n17200), .A2(n17199), .A3(n17198), .A4(n17197), .ZN(
        n17206) );
  AOI22_X1 U20343 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n14205), .B1(
        n9687), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17204) );
  AOI22_X1 U20344 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n9689), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17441), .ZN(n17203) );
  AOI22_X1 U20345 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17348), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U20346 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17406), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n9673), .ZN(n17201) );
  NAND4_X1 U20347 ( .A1(n17204), .A2(n17203), .A3(n17202), .A4(n17201), .ZN(
        n17205) );
  NOR2_X1 U20348 ( .A1(n17206), .A2(n17205), .ZN(n17219) );
  AOI22_X1 U20349 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20350 ( .A1(n12239), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20351 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17207) );
  OAI21_X1 U20352 ( .B1(n17208), .B2(n18513), .A(n17207), .ZN(n17215) );
  AOI22_X1 U20353 ( .A1(n17423), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17213) );
  AOI22_X1 U20354 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9689), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20355 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12249), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20356 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17210) );
  NAND4_X1 U20357 ( .A1(n17213), .A2(n17212), .A3(n17211), .A4(n17210), .ZN(
        n17214) );
  AOI211_X1 U20358 ( .C1(n17422), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n17215), .B(n17214), .ZN(n17216) );
  NAND3_X1 U20359 ( .A1(n17218), .A2(n17217), .A3(n17216), .ZN(n17224) );
  NAND2_X1 U20360 ( .A1(n17225), .A2(n17224), .ZN(n17223) );
  XNOR2_X1 U20361 ( .A(n17219), .B(n17223), .ZN(n17496) );
  NOR2_X1 U20362 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n17220), .ZN(n17222) );
  OAI22_X1 U20363 ( .A1(n17496), .A2(n17470), .B1(n17222), .B2(n17221), .ZN(
        P3_U2673) );
  OAI21_X1 U20364 ( .B1(n17225), .B2(n17224), .A(n17223), .ZN(n17504) );
  NAND4_X1 U20365 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17243), .A3(n17227), 
        .A4(n17226), .ZN(n17230) );
  NAND2_X1 U20366 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17228), .ZN(n17229) );
  OAI211_X1 U20367 ( .C1(n17470), .C2(n17504), .A(n17230), .B(n17229), .ZN(
        P3_U2674) );
  OAI211_X1 U20368 ( .C1(n17511), .C2(n17510), .A(n17482), .B(n17509), .ZN(
        n17231) );
  OAI221_X1 U20369 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17234), .C1(n17233), 
        .C2(n17232), .A(n17231), .ZN(P3_U2676) );
  AOI21_X1 U20370 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17470), .A(n17243), .ZN(
        n17236) );
  XNOR2_X1 U20371 ( .A(n17235), .B(n17239), .ZN(n17520) );
  OAI22_X1 U20372 ( .A1(n17237), .A2(n17236), .B1(n17470), .B2(n17520), .ZN(
        P3_U2677) );
  INV_X1 U20373 ( .A(n17238), .ZN(n17246) );
  AOI21_X1 U20374 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17470), .A(n17246), .ZN(
        n17242) );
  OAI21_X1 U20375 ( .B1(n17241), .B2(n17240), .A(n17239), .ZN(n17525) );
  OAI22_X1 U20376 ( .A1(n17243), .A2(n17242), .B1(n17470), .B2(n17525), .ZN(
        P3_U2678) );
  AOI21_X1 U20377 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17470), .A(n17251), .ZN(
        n17245) );
  XNOR2_X1 U20378 ( .A(n17244), .B(n17247), .ZN(n17531) );
  OAI22_X1 U20379 ( .A1(n17246), .A2(n17245), .B1(n17470), .B2(n17531), .ZN(
        P3_U2679) );
  INV_X1 U20380 ( .A(n17262), .ZN(n17278) );
  AOI21_X1 U20381 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17470), .A(n17265), .ZN(
        n17250) );
  OAI21_X1 U20382 ( .B1(n17249), .B2(n17248), .A(n17247), .ZN(n17537) );
  OAI22_X1 U20383 ( .A1(n17251), .A2(n17250), .B1(n17470), .B2(n17537), .ZN(
        P3_U2680) );
  AOI22_X1 U20384 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12249), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17255) );
  AOI22_X1 U20385 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U20386 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17253) );
  AOI22_X1 U20387 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17252) );
  NAND4_X1 U20388 ( .A1(n17255), .A2(n17254), .A3(n17253), .A4(n17252), .ZN(
        n17261) );
  AOI22_X1 U20389 ( .A1(n12239), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U20390 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9687), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17258) );
  AOI22_X1 U20391 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17257) );
  AOI22_X1 U20392 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17256) );
  NAND4_X1 U20393 ( .A1(n17259), .A2(n17258), .A3(n17257), .A4(n17256), .ZN(
        n17260) );
  NOR2_X1 U20394 ( .A1(n17261), .A2(n17260), .ZN(n17539) );
  NOR2_X1 U20395 ( .A1(n17277), .A2(n17262), .ZN(n17263) );
  AOI21_X1 U20396 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17470), .A(n17263), .ZN(
        n17264) );
  OAI22_X1 U20397 ( .A1(n17539), .A2(n17470), .B1(n17265), .B2(n17264), .ZN(
        P3_U2681) );
  AOI22_X1 U20398 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U20399 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17268) );
  AOI22_X1 U20400 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17267) );
  AOI22_X1 U20401 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17266) );
  NAND4_X1 U20402 ( .A1(n17269), .A2(n17268), .A3(n17267), .A4(n17266), .ZN(
        n17275) );
  AOI22_X1 U20403 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9689), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17273) );
  AOI22_X1 U20404 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17272) );
  AOI22_X1 U20405 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9687), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20406 ( .A1(n12239), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17270) );
  NAND4_X1 U20407 ( .A1(n17273), .A2(n17272), .A3(n17271), .A4(n17270), .ZN(
        n17274) );
  NOR2_X1 U20408 ( .A1(n17275), .A2(n17274), .ZN(n17547) );
  NOR2_X1 U20409 ( .A1(n17482), .A2(n17276), .ZN(n17290) );
  AOI22_X1 U20410 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17290), .B1(n17278), 
        .B2(n17277), .ZN(n17279) );
  OAI21_X1 U20411 ( .B1(n17547), .B2(n17470), .A(n17279), .ZN(P3_U2682) );
  AOI22_X1 U20412 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20413 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U20414 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U20415 ( .A1(n17406), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17280) );
  NAND4_X1 U20416 ( .A1(n17283), .A2(n17282), .A3(n17281), .A4(n17280), .ZN(
        n17289) );
  AOI22_X1 U20417 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20418 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20419 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9689), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17285) );
  AOI22_X1 U20420 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17284) );
  NAND4_X1 U20421 ( .A1(n17287), .A2(n17286), .A3(n17285), .A4(n17284), .ZN(
        n17288) );
  NOR2_X1 U20422 ( .A1(n17289), .A2(n17288), .ZN(n17551) );
  OAI21_X1 U20423 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17291), .A(n17290), .ZN(
        n17292) );
  OAI21_X1 U20424 ( .B1(n17551), .B2(n17470), .A(n17292), .ZN(P3_U2683) );
  AOI22_X1 U20425 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9689), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U20426 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U20427 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17294) );
  AOI22_X1 U20428 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17293) );
  NAND4_X1 U20429 ( .A1(n17296), .A2(n17295), .A3(n17294), .A4(n17293), .ZN(
        n17302) );
  AOI22_X1 U20430 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U20431 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17299) );
  AOI22_X1 U20432 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17298) );
  AOI22_X1 U20433 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17297) );
  NAND4_X1 U20434 ( .A1(n17300), .A2(n17299), .A3(n17298), .A4(n17297), .ZN(
        n17301) );
  NOR2_X1 U20435 ( .A1(n17302), .A2(n17301), .ZN(n17556) );
  OAI21_X1 U20436 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17318), .A(n17303), .ZN(
        n17304) );
  AOI22_X1 U20437 ( .A1(n17482), .A2(n17556), .B1(n17304), .B2(n17470), .ZN(
        P3_U2684) );
  AOI21_X1 U20438 ( .B1(n17305), .B2(n17330), .A(n17482), .ZN(n17306) );
  INV_X1 U20439 ( .A(n17306), .ZN(n17317) );
  AOI22_X1 U20440 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17310) );
  AOI22_X1 U20441 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20442 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U20443 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17307) );
  NAND4_X1 U20444 ( .A1(n17310), .A2(n17309), .A3(n17308), .A4(n17307), .ZN(
        n17316) );
  AOI22_X1 U20445 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17314) );
  AOI22_X1 U20446 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17313) );
  AOI22_X1 U20447 ( .A1(n17353), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17312) );
  AOI22_X1 U20448 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17311) );
  NAND4_X1 U20449 ( .A1(n17314), .A2(n17313), .A3(n17312), .A4(n17311), .ZN(
        n17315) );
  NOR2_X1 U20450 ( .A1(n17316), .A2(n17315), .ZN(n17561) );
  OAI22_X1 U20451 ( .A1(n17318), .A2(n17317), .B1(n17561), .B2(n17470), .ZN(
        P3_U2685) );
  AOI22_X1 U20452 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17323) );
  AOI22_X1 U20453 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17322) );
  AOI22_X1 U20454 ( .A1(n17406), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17321) );
  AOI22_X1 U20455 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17320) );
  NAND4_X1 U20456 ( .A1(n17323), .A2(n17322), .A3(n17321), .A4(n17320), .ZN(
        n17329) );
  AOI22_X1 U20457 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17327) );
  AOI22_X1 U20458 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17326) );
  AOI22_X1 U20459 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U20460 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17324) );
  NAND4_X1 U20461 ( .A1(n17327), .A2(n17326), .A3(n17325), .A4(n17324), .ZN(
        n17328) );
  NOR2_X1 U20462 ( .A1(n17329), .A2(n17328), .ZN(n17565) );
  OAI21_X1 U20463 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17331), .A(n17330), .ZN(
        n17332) );
  AOI22_X1 U20464 ( .A1(n17482), .A2(n17565), .B1(n17332), .B2(n17470), .ZN(
        P3_U2686) );
  INV_X1 U20465 ( .A(n17333), .ZN(n17336) );
  NAND3_X1 U20466 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17465), .A3(n17464), .ZN(
        n17461) );
  NOR2_X1 U20467 ( .A1(n17457), .A2(n17461), .ZN(n17460) );
  NAND4_X1 U20468 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(n17460), .ZN(n17334) );
  NOR3_X1 U20469 ( .A1(n17419), .A2(n17335), .A3(n17334), .ZN(n17389) );
  NAND2_X1 U20470 ( .A1(n17336), .A2(n17389), .ZN(n17362) );
  AOI22_X1 U20471 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17340) );
  AOI22_X1 U20472 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17339) );
  AOI22_X1 U20473 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12249), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U20474 ( .A1(n17406), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17337) );
  NAND4_X1 U20475 ( .A1(n17340), .A2(n17339), .A3(n17338), .A4(n17337), .ZN(
        n17346) );
  AOI22_X1 U20476 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17344) );
  AOI22_X1 U20477 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17343) );
  AOI22_X1 U20478 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17342) );
  AOI22_X1 U20479 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17341) );
  NAND4_X1 U20480 ( .A1(n17344), .A2(n17343), .A3(n17342), .A4(n17341), .ZN(
        n17345) );
  NOR2_X1 U20481 ( .A1(n17346), .A2(n17345), .ZN(n17572) );
  NAND3_X1 U20482 ( .A1(n17362), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17470), 
        .ZN(n17347) );
  OAI221_X1 U20483 ( .B1(n17362), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n17470), 
        .C2(n17572), .A(n17347), .ZN(P3_U2687) );
  AOI22_X1 U20484 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9687), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U20485 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17348), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17351) );
  AOI22_X1 U20486 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17423), .ZN(n17350) );
  AOI22_X1 U20487 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n14166), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17406), .ZN(n17349) );
  NAND4_X1 U20488 ( .A1(n17352), .A2(n17351), .A3(n17350), .A4(n17349), .ZN(
        n17359) );
  AOI22_X1 U20489 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17353), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U20490 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9689), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17356) );
  AOI22_X1 U20491 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17441), .ZN(n17355) );
  AOI22_X1 U20492 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n9673), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n16181), .ZN(n17354) );
  NAND4_X1 U20493 ( .A1(n17357), .A2(n17356), .A3(n17355), .A4(n17354), .ZN(
        n17358) );
  NOR2_X1 U20494 ( .A1(n17359), .A2(n17358), .ZN(n17576) );
  NAND3_X1 U20495 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .ZN(n17361) );
  OAI21_X1 U20496 ( .B1(n17403), .B2(n17361), .A(n17360), .ZN(n17363) );
  NAND3_X1 U20497 ( .A1(n17363), .A2(n17362), .A3(n17470), .ZN(n17364) );
  OAI21_X1 U20498 ( .B1(n17576), .B2(n17470), .A(n17364), .ZN(P3_U2688) );
  NAND3_X1 U20499 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n17389), .ZN(n17377) );
  AOI22_X1 U20500 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17374) );
  AOI22_X1 U20501 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17373) );
  AOI22_X1 U20502 ( .A1(n17392), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17365) );
  OAI21_X1 U20503 ( .B1(n12237), .B2(n18513), .A(n17365), .ZN(n17371) );
  AOI22_X1 U20504 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U20505 ( .A1(n12239), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17368) );
  AOI22_X1 U20506 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17367) );
  AOI22_X1 U20507 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9689), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17366) );
  NAND4_X1 U20508 ( .A1(n17369), .A2(n17368), .A3(n17367), .A4(n17366), .ZN(
        n17370) );
  AOI211_X1 U20509 ( .C1(n9673), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n17371), .B(n17370), .ZN(n17372) );
  NAND3_X1 U20510 ( .A1(n17374), .A2(n17373), .A3(n17372), .ZN(n17578) );
  AOI22_X1 U20511 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17375), .B1(n17482), 
        .B2(n17578), .ZN(n17376) );
  OAI21_X1 U20512 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17377), .A(n17376), .ZN(
        P3_U2689) );
  AOI22_X1 U20513 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U20514 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9673), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17380) );
  AOI22_X1 U20515 ( .A1(n17392), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17379) );
  AOI22_X1 U20516 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17378) );
  NAND4_X1 U20517 ( .A1(n17381), .A2(n17380), .A3(n17379), .A4(n17378), .ZN(
        n17388) );
  AOI22_X1 U20518 ( .A1(n17441), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17386) );
  AOI22_X1 U20519 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9689), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17385) );
  AOI22_X1 U20520 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17384) );
  AOI22_X1 U20521 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17383) );
  NAND4_X1 U20522 ( .A1(n17386), .A2(n17385), .A3(n17384), .A4(n17383), .ZN(
        n17387) );
  NOR2_X1 U20523 ( .A1(n17388), .A2(n17387), .ZN(n17588) );
  NOR2_X1 U20524 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17389), .ZN(n17390) );
  OAI22_X1 U20525 ( .A1(n17588), .A2(n17470), .B1(n17391), .B2(n17390), .ZN(
        P3_U2691) );
  AOI22_X1 U20526 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U20527 ( .A1(n17392), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U20528 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17394) );
  AOI22_X1 U20529 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17393) );
  NAND4_X1 U20530 ( .A1(n17396), .A2(n17395), .A3(n17394), .A4(n17393), .ZN(
        n17402) );
  AOI22_X1 U20531 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17400) );
  AOI22_X1 U20532 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U20533 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12249), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17398) );
  AOI22_X1 U20534 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17397) );
  NAND4_X1 U20535 ( .A1(n17400), .A2(n17399), .A3(n17398), .A4(n17397), .ZN(
        n17401) );
  NOR2_X1 U20536 ( .A1(n17402), .A2(n17401), .ZN(n17591) );
  OAI211_X1 U20537 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n17404), .A(n17403), .B(
        n17470), .ZN(n17405) );
  OAI21_X1 U20538 ( .B1(n17591), .B2(n17470), .A(n17405), .ZN(P3_U2692) );
  AOI22_X1 U20539 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U20540 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17409) );
  AOI22_X1 U20541 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U20542 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17406), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17407) );
  NAND4_X1 U20543 ( .A1(n17410), .A2(n17409), .A3(n17408), .A4(n17407), .ZN(
        n17417) );
  AOI22_X1 U20544 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17415) );
  AOI22_X1 U20545 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17414) );
  AOI22_X1 U20546 ( .A1(n12239), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17319), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U20547 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17412) );
  NAND4_X1 U20548 ( .A1(n17415), .A2(n17414), .A3(n17413), .A4(n17412), .ZN(
        n17416) );
  NOR2_X1 U20549 ( .A1(n17417), .A2(n17416), .ZN(n17594) );
  OAI33_X1 U20550 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17597), .A3(n17435), 
        .B1(n17419), .B2(n17482), .B3(n17418), .ZN(n17420) );
  INV_X1 U20551 ( .A(n17420), .ZN(n17421) );
  OAI21_X1 U20552 ( .B1(n17594), .B2(n17470), .A(n17421), .ZN(P3_U2693) );
  AOI22_X1 U20553 ( .A1(n9683), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9689), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17427) );
  AOI22_X1 U20554 ( .A1(n17422), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14205), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17426) );
  AOI22_X1 U20555 ( .A1(n17411), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17423), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17425) );
  AOI22_X1 U20556 ( .A1(n17406), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17424) );
  NAND4_X1 U20557 ( .A1(n17427), .A2(n17426), .A3(n17425), .A4(n17424), .ZN(
        n17434) );
  AOI22_X1 U20558 ( .A1(n9687), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(n9673), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U20559 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17431) );
  AOI22_X1 U20560 ( .A1(n17319), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U20561 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17429) );
  NAND4_X1 U20562 ( .A1(n17432), .A2(n17431), .A3(n17430), .A4(n17429), .ZN(
        n17433) );
  NOR2_X1 U20563 ( .A1(n17434), .A2(n17433), .ZN(n17598) );
  INV_X1 U20564 ( .A(n17452), .ZN(n17456) );
  AOI21_X1 U20565 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17456), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n17437) );
  NAND2_X1 U20566 ( .A1(n17470), .A2(n17435), .ZN(n17436) );
  OAI22_X1 U20567 ( .A1(n17598), .A2(n17470), .B1(n17437), .B2(n17436), .ZN(
        P3_U2694) );
  AOI22_X1 U20568 ( .A1(n9688), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17411), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17450) );
  AOI22_X1 U20569 ( .A1(n17353), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17449) );
  AOI22_X1 U20570 ( .A1(n9673), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16181), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17439) );
  OAI21_X1 U20571 ( .B1(n12237), .B2(n18478), .A(n17439), .ZN(n17447) );
  AOI22_X1 U20572 ( .A1(n9658), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9683), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17445) );
  AOI22_X1 U20573 ( .A1(n14205), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9689), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20574 ( .A1(n17428), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17441), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U20575 ( .A1(n17348), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17442) );
  NAND4_X1 U20576 ( .A1(n17445), .A2(n17444), .A3(n17443), .A4(n17442), .ZN(
        n17446) );
  AOI211_X1 U20577 ( .C1(n17319), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n17447), .B(n17446), .ZN(n17448) );
  NAND3_X1 U20578 ( .A1(n17450), .A2(n17449), .A3(n17448), .ZN(n17601) );
  INV_X1 U20579 ( .A(n17601), .ZN(n17454) );
  AOI22_X1 U20580 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17452), .B1(n17456), .B2(
        n17451), .ZN(n17453) );
  AOI22_X1 U20581 ( .A1(n17482), .A2(n17454), .B1(n17453), .B2(n17470), .ZN(
        P3_U2695) );
  OAI21_X1 U20582 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17460), .A(n17470), .ZN(
        n17455) );
  INV_X1 U20583 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18522) );
  OAI22_X1 U20584 ( .A1(n17456), .A2(n17455), .B1(n18522), .B2(n17470), .ZN(
        P3_U2696) );
  OAI21_X1 U20585 ( .B1(n17457), .B2(n17482), .A(n17461), .ZN(n17458) );
  INV_X1 U20586 ( .A(n17458), .ZN(n17459) );
  OAI22_X1 U20587 ( .A1(n17460), .A2(n17459), .B1(n18513), .B2(n17470), .ZN(
        P3_U2697) );
  INV_X1 U20588 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18506) );
  OAI21_X1 U20589 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17462), .A(n17461), .ZN(
        n17463) );
  AOI22_X1 U20590 ( .A1(n17482), .A2(n18506), .B1(n17463), .B2(n17470), .ZN(
        P3_U2698) );
  AND2_X1 U20591 ( .A1(n17465), .A2(n17464), .ZN(n17468) );
  NOR3_X1 U20592 ( .A1(n17466), .A2(n17469), .A3(n17484), .ZN(n17472) );
  AOI21_X1 U20593 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17470), .A(n17472), .ZN(
        n17467) );
  OAI22_X1 U20594 ( .A1(n17468), .A2(n17467), .B1(n18500), .B2(n17470), .ZN(
        P3_U2699) );
  NOR2_X1 U20595 ( .A1(n17469), .A2(n17484), .ZN(n17476) );
  AOI21_X1 U20596 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17470), .A(n17476), .ZN(
        n17471) );
  INV_X1 U20597 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18494) );
  OAI22_X1 U20598 ( .A1(n17472), .A2(n17471), .B1(n18494), .B2(n17470), .ZN(
        P3_U2700) );
  OAI221_X1 U20599 ( .B1(n17474), .B2(n17481), .C1(n18518), .C2(n17481), .A(
        n17473), .ZN(n17475) );
  INV_X1 U20600 ( .A(n17475), .ZN(n17477) );
  AOI211_X1 U20601 ( .C1(n17482), .C2(n18488), .A(n17477), .B(n17476), .ZN(
        P3_U2701) );
  INV_X1 U20602 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17479) );
  OAI222_X1 U20603 ( .A1(n17480), .A2(n17484), .B1(n17479), .B2(n17478), .C1(
        n18482), .C2(n17470), .ZN(P3_U2702) );
  AOI22_X1 U20604 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17482), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17481), .ZN(n17483) );
  OAI21_X1 U20605 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17484), .A(n17483), .ZN(
        P3_U2703) );
  INV_X1 U20606 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18516) );
  NOR2_X2 U20607 ( .A1(n17622), .A2(n18510), .ZN(n17566) );
  INV_X1 U20608 ( .A(n17566), .ZN(n17538) );
  INV_X1 U20609 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17649) );
  INV_X1 U20610 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17653) );
  INV_X1 U20611 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17655) );
  INV_X1 U20612 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17657) );
  INV_X1 U20613 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17671) );
  NAND4_X1 U20614 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n17488)
         );
  NAND4_X1 U20615 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17486) );
  NAND4_X1 U20616 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_1__SCAN_IN), .A4(P3_EAX_REG_0__SCAN_IN), .ZN(n17485) );
  INV_X1 U20617 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17663) );
  INV_X1 U20618 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17665) );
  INV_X1 U20619 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17667) );
  INV_X1 U20620 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17709) );
  NOR4_X1 U20621 ( .A1(n17663), .A2(n17665), .A3(n17667), .A4(n17709), .ZN(
        n17489) );
  NAND4_X1 U20622 ( .A1(n17568), .A2(P3_EAX_REG_22__SCAN_IN), .A3(
        P3_EAX_REG_21__SCAN_IN), .A4(n17489), .ZN(n17533) );
  NAND2_X1 U20623 ( .A1(n18518), .A2(n17532), .ZN(n17526) );
  NAND2_X1 U20624 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17501), .ZN(n17500) );
  NOR2_X1 U20625 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17500), .ZN(n17493) );
  INV_X1 U20626 ( .A(n17490), .ZN(n17491) );
  NAND2_X1 U20627 ( .A1(n17622), .A2(n17500), .ZN(n17499) );
  OAI21_X1 U20628 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17491), .A(n17499), .ZN(
        n17492) );
  AOI22_X1 U20629 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17493), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17492), .ZN(n17494) );
  OAI21_X1 U20630 ( .B1(n18516), .B2(n17538), .A(n17494), .ZN(P3_U2704) );
  INV_X1 U20631 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17723) );
  NOR2_X2 U20632 ( .A1(n17495), .A2(n17622), .ZN(n17567) );
  INV_X1 U20633 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18508) );
  OAI22_X1 U20634 ( .A1(n17496), .A2(n17614), .B1(n18508), .B2(n17538), .ZN(
        n17497) );
  AOI21_X1 U20635 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17567), .A(n17497), .ZN(
        n17498) );
  OAI221_X1 U20636 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17500), .C1(n17723), 
        .C2(n17499), .A(n17498), .ZN(P3_U2705) );
  AOI22_X1 U20637 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17566), .ZN(n17503) );
  OAI211_X1 U20638 ( .C1(n17501), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17622), .B(
        n17500), .ZN(n17502) );
  OAI211_X1 U20639 ( .C1(n17504), .C2(n17630), .A(n17503), .B(n17502), .ZN(
        P3_U2706) );
  INV_X1 U20640 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18496) );
  AOI22_X1 U20641 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17567), .B1(n17635), .B2(
        n17505), .ZN(n17508) );
  OAI211_X1 U20642 ( .C1(n17512), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17622), .B(
        n17506), .ZN(n17507) );
  OAI211_X1 U20643 ( .C1(n17538), .C2(n18496), .A(n17508), .B(n17507), .ZN(
        P3_U2707) );
  OAI21_X1 U20644 ( .B1(n17511), .B2(n17510), .A(n17509), .ZN(n17516) );
  AOI22_X1 U20645 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17566), .ZN(n17515) );
  AOI211_X1 U20646 ( .C1(n17649), .C2(n17517), .A(n17512), .B(n17580), .ZN(
        n17513) );
  INV_X1 U20647 ( .A(n17513), .ZN(n17514) );
  OAI211_X1 U20648 ( .C1(n17516), .C2(n17614), .A(n17515), .B(n17514), .ZN(
        P3_U2708) );
  AOI22_X1 U20649 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17566), .ZN(n17519) );
  OAI211_X1 U20650 ( .C1(n17521), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17622), .B(
        n17517), .ZN(n17518) );
  OAI211_X1 U20651 ( .C1(n17520), .C2(n17630), .A(n17519), .B(n17518), .ZN(
        P3_U2709) );
  AOI22_X1 U20652 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17566), .ZN(n17524) );
  AOI211_X1 U20653 ( .C1(n17653), .C2(n17527), .A(n17521), .B(n17580), .ZN(
        n17522) );
  INV_X1 U20654 ( .A(n17522), .ZN(n17523) );
  OAI211_X1 U20655 ( .C1(n17525), .C2(n17630), .A(n17524), .B(n17523), .ZN(
        P3_U2710) );
  AOI22_X1 U20656 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17566), .ZN(n17530) );
  OAI21_X1 U20657 ( .B1(n17655), .B2(n17580), .A(n17526), .ZN(n17528) );
  NAND2_X1 U20658 ( .A1(n17528), .A2(n17527), .ZN(n17529) );
  OAI211_X1 U20659 ( .C1(n17531), .C2(n17614), .A(n17530), .B(n17529), .ZN(
        P3_U2711) );
  AOI211_X1 U20660 ( .C1(n17657), .C2(n17533), .A(n17580), .B(n17532), .ZN(
        n17534) );
  AOI21_X1 U20661 ( .B1(n17566), .B2(BUF2_REG_23__SCAN_IN), .A(n17534), .ZN(
        n17536) );
  NAND2_X1 U20662 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17567), .ZN(n17535) );
  OAI211_X1 U20663 ( .C1(n17537), .C2(n17614), .A(n17536), .B(n17535), .ZN(
        P3_U2712) );
  NAND3_X1 U20664 ( .A1(n18518), .A2(n17568), .A3(P3_EAX_REG_17__SCAN_IN), 
        .ZN(n17562) );
  NAND2_X1 U20665 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17558), .ZN(n17557) );
  NAND2_X1 U20666 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17552), .ZN(n17548) );
  NAND2_X1 U20667 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17544), .ZN(n17543) );
  NAND2_X1 U20668 ( .A1(n17543), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17542) );
  OAI22_X1 U20669 ( .A1(n17539), .A2(n17614), .B1(n19557), .B2(n17538), .ZN(
        n17540) );
  AOI21_X1 U20670 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17567), .A(n17540), .ZN(
        n17541) );
  OAI221_X1 U20671 ( .B1(n17543), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17542), 
        .C2(n17580), .A(n17541), .ZN(P3_U2713) );
  AOI22_X1 U20672 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17566), .ZN(n17546) );
  OAI211_X1 U20673 ( .C1(n17544), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17622), .B(
        n17543), .ZN(n17545) );
  OAI211_X1 U20674 ( .C1(n17547), .C2(n17614), .A(n17546), .B(n17545), .ZN(
        P3_U2714) );
  AOI22_X1 U20675 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17566), .ZN(n17550) );
  OAI211_X1 U20676 ( .C1(n17552), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17622), .B(
        n17548), .ZN(n17549) );
  OAI211_X1 U20677 ( .C1(n17551), .C2(n17614), .A(n17550), .B(n17549), .ZN(
        P3_U2715) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17566), .ZN(n17555) );
  AOI211_X1 U20679 ( .C1(n17665), .C2(n17557), .A(n17552), .B(n17580), .ZN(
        n17553) );
  INV_X1 U20680 ( .A(n17553), .ZN(n17554) );
  OAI211_X1 U20681 ( .C1(n17556), .C2(n17614), .A(n17555), .B(n17554), .ZN(
        P3_U2716) );
  AOI22_X1 U20682 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17566), .ZN(n17560) );
  OAI211_X1 U20683 ( .C1(n17558), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17622), .B(
        n17557), .ZN(n17559) );
  OAI211_X1 U20684 ( .C1(n17561), .C2(n17614), .A(n17560), .B(n17559), .ZN(
        P3_U2717) );
  AOI22_X1 U20685 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17566), .ZN(n17564) );
  OAI211_X1 U20686 ( .C1(n17568), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17622), .B(
        n17562), .ZN(n17563) );
  OAI211_X1 U20687 ( .C1(n17565), .C2(n17614), .A(n17564), .B(n17563), .ZN(
        P3_U2718) );
  AOI22_X1 U20688 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17566), .ZN(n17571) );
  AOI211_X1 U20689 ( .C1(n17671), .C2(n17573), .A(n17580), .B(n17568), .ZN(
        n17569) );
  INV_X1 U20690 ( .A(n17569), .ZN(n17570) );
  OAI211_X1 U20691 ( .C1(n17572), .C2(n17614), .A(n17571), .B(n17570), .ZN(
        P3_U2719) );
  NAND2_X1 U20692 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17636), .ZN(n17575) );
  OAI211_X1 U20693 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17579), .A(n17627), .B(
        n17573), .ZN(n17574) );
  OAI211_X1 U20694 ( .C1(n17576), .C2(n17614), .A(n17575), .B(n17574), .ZN(
        P3_U2720) );
  INV_X1 U20695 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17678) );
  INV_X1 U20696 ( .A(n17577), .ZN(n17602) );
  INV_X1 U20697 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n21224) );
  INV_X1 U20698 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17685) );
  NOR4_X1 U20699 ( .A1(n17597), .A2(n17602), .A3(n21224), .A4(n17685), .ZN(
        n17600) );
  AND2_X1 U20700 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17600), .ZN(n17596) );
  NAND2_X1 U20701 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17596), .ZN(n17587) );
  NOR2_X1 U20702 ( .A1(n17678), .A2(n17587), .ZN(n17590) );
  NAND2_X1 U20703 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17590), .ZN(n17583) );
  AOI22_X1 U20704 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17636), .B1(n17635), .B2(
        n17578), .ZN(n17582) );
  INV_X1 U20705 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17749) );
  OR3_X1 U20706 ( .A1(n17749), .A2(n17580), .A3(n17579), .ZN(n17581) );
  OAI211_X1 U20707 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17583), .A(n17582), .B(
        n17581), .ZN(P3_U2721) );
  INV_X1 U20708 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17746) );
  INV_X1 U20709 ( .A(n17583), .ZN(n17586) );
  AOI21_X1 U20710 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17627), .A(n17590), .ZN(
        n17585) );
  OAI222_X1 U20711 ( .A1(n17633), .A2(n17746), .B1(n17586), .B2(n17585), .C1(
        n17630), .C2(n17584), .ZN(P3_U2722) );
  INV_X1 U20712 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17742) );
  INV_X1 U20713 ( .A(n17587), .ZN(n17593) );
  AOI21_X1 U20714 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17627), .A(n17593), .ZN(
        n17589) );
  OAI222_X1 U20715 ( .A1(n17633), .A2(n17742), .B1(n17590), .B2(n17589), .C1(
        n17630), .C2(n17588), .ZN(P3_U2723) );
  AOI21_X1 U20716 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17627), .A(n17596), .ZN(
        n17592) );
  OAI222_X1 U20717 ( .A1(n17633), .A2(n17740), .B1(n17593), .B2(n17592), .C1(
        n17630), .C2(n17591), .ZN(P3_U2724) );
  AOI21_X1 U20718 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(n17627), .A(n17600), .ZN(
        n17595) );
  OAI222_X1 U20719 ( .A1(n17633), .A2(n17738), .B1(n17596), .B2(n17595), .C1(
        n17630), .C2(n17594), .ZN(P3_U2725) );
  NOR2_X1 U20720 ( .A1(n17597), .A2(n17602), .ZN(n17607) );
  AOI22_X1 U20721 ( .A1(n17607), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17622), .ZN(n17599) );
  OAI222_X1 U20722 ( .A1(n17633), .A2(n17736), .B1(n17600), .B2(n17599), .C1(
        n17630), .C2(n17598), .ZN(P3_U2726) );
  INV_X1 U20723 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17734) );
  AOI22_X1 U20724 ( .A1(n17635), .A2(n17601), .B1(n17607), .B2(n17685), .ZN(
        n17604) );
  NAND3_X1 U20725 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17627), .A3(n17602), .ZN(
        n17603) );
  OAI211_X1 U20726 ( .C1(n17633), .C2(n17734), .A(n17604), .B(n17603), .ZN(
        P3_U2727) );
  INV_X1 U20727 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17690) );
  INV_X1 U20728 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17694) );
  INV_X1 U20729 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17726) );
  NOR2_X1 U20730 ( .A1(n17726), .A2(n17639), .ZN(n17626) );
  NAND3_X1 U20731 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(n17626), .ZN(n17617) );
  NOR2_X1 U20732 ( .A1(n17694), .A2(n17617), .ZN(n17621) );
  NAND2_X1 U20733 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17621), .ZN(n17608) );
  NOR2_X1 U20734 ( .A1(n17690), .A2(n17608), .ZN(n17612) );
  AOI21_X1 U20735 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17627), .A(n17612), .ZN(
        n17606) );
  OAI222_X1 U20736 ( .A1(n18514), .A2(n17633), .B1(n17607), .B2(n17606), .C1(
        n17630), .C2(n17605), .ZN(P3_U2728) );
  INV_X1 U20737 ( .A(n17608), .ZN(n17616) );
  AOI21_X1 U20738 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17627), .A(n17616), .ZN(
        n17611) );
  INV_X1 U20739 ( .A(n17609), .ZN(n17610) );
  OAI222_X1 U20740 ( .A1(n18509), .A2(n17633), .B1(n17612), .B2(n17611), .C1(
        n17630), .C2(n17610), .ZN(P3_U2729) );
  AOI21_X1 U20741 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17627), .A(n17621), .ZN(
        n17615) );
  OAI222_X1 U20742 ( .A1(n18501), .A2(n17633), .B1(n17616), .B2(n17615), .C1(
        n17614), .C2(n17613), .ZN(P3_U2730) );
  INV_X1 U20743 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18495) );
  INV_X1 U20744 ( .A(n17617), .ZN(n17625) );
  AOI21_X1 U20745 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17627), .A(n17625), .ZN(
        n17620) );
  INV_X1 U20746 ( .A(n17618), .ZN(n17619) );
  OAI222_X1 U20747 ( .A1(n18495), .A2(n17633), .B1(n17621), .B2(n17620), .C1(
        n17630), .C2(n17619), .ZN(P3_U2731) );
  AOI22_X1 U20748 ( .A1(n17626), .A2(P3_EAX_REG_2__SCAN_IN), .B1(
        P3_EAX_REG_3__SCAN_IN), .B2(n17622), .ZN(n17624) );
  OAI222_X1 U20749 ( .A1(n18489), .A2(n17633), .B1(n17625), .B2(n17624), .C1(
        n17630), .C2(n17623), .ZN(P3_U2732) );
  INV_X1 U20750 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18483) );
  AND2_X1 U20751 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17626), .ZN(n17632) );
  AOI21_X1 U20752 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17627), .A(n17626), .ZN(
        n17631) );
  INV_X1 U20753 ( .A(n17628), .ZN(n17629) );
  OAI222_X1 U20754 ( .A1(n18483), .A2(n17633), .B1(n17632), .B2(n17631), .C1(
        n17630), .C2(n17629), .ZN(P3_U2733) );
  AOI22_X1 U20755 ( .A1(n17636), .A2(BUF2_REG_1__SCAN_IN), .B1(n17635), .B2(
        n17634), .ZN(n17637) );
  OAI221_X1 U20756 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17639), .C1(n17726), 
        .C2(n17638), .A(n17637), .ZN(P3_U2734) );
  NOR2_X1 U20757 ( .A1(n19075), .A2(n18126), .ZN(n19109) );
  AND2_X1 U20758 ( .A1(n17688), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20759 ( .A1(n17672), .A2(n17642), .ZN(n17670) );
  AOI22_X1 U20760 ( .A1(n19109), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17643) );
  OAI21_X1 U20761 ( .B1(n17723), .B2(n17670), .A(n17643), .ZN(P3_U2737) );
  INV_X1 U20762 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17645) );
  AOI22_X1 U20763 ( .A1(n19109), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17644) );
  OAI21_X1 U20764 ( .B1(n17645), .B2(n17670), .A(n17644), .ZN(P3_U2738) );
  INV_X1 U20765 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17647) );
  AOI22_X1 U20766 ( .A1(n19109), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17646) );
  OAI21_X1 U20767 ( .B1(n17647), .B2(n17670), .A(n17646), .ZN(P3_U2739) );
  AOI22_X1 U20768 ( .A1(n19109), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17688), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17648) );
  OAI21_X1 U20769 ( .B1(n17649), .B2(n17670), .A(n17648), .ZN(P3_U2740) );
  INV_X1 U20770 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17651) );
  AOI22_X1 U20771 ( .A1(n19109), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17688), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17650) );
  OAI21_X1 U20772 ( .B1(n17651), .B2(n17670), .A(n17650), .ZN(P3_U2741) );
  AOI22_X1 U20773 ( .A1(n19109), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17688), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17652) );
  OAI21_X1 U20774 ( .B1(n17653), .B2(n17670), .A(n17652), .ZN(P3_U2742) );
  AOI22_X1 U20775 ( .A1(n19109), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17688), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17654) );
  OAI21_X1 U20776 ( .B1(n17655), .B2(n17670), .A(n17654), .ZN(P3_U2743) );
  CLKBUF_X1 U20777 ( .A(n19109), .Z(n17701) );
  AOI22_X1 U20778 ( .A1(n17701), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17656) );
  OAI21_X1 U20779 ( .B1(n17657), .B2(n17670), .A(n17656), .ZN(P3_U2744) );
  INV_X1 U20780 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17659) );
  AOI22_X1 U20781 ( .A1(n17701), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17658) );
  OAI21_X1 U20782 ( .B1(n17659), .B2(n17670), .A(n17658), .ZN(P3_U2745) );
  INV_X1 U20783 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17661) );
  AOI22_X1 U20784 ( .A1(n17701), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17660) );
  OAI21_X1 U20785 ( .B1(n17661), .B2(n17670), .A(n17660), .ZN(P3_U2746) );
  AOI22_X1 U20786 ( .A1(n17701), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17662) );
  OAI21_X1 U20787 ( .B1(n17663), .B2(n17670), .A(n17662), .ZN(P3_U2747) );
  AOI22_X1 U20788 ( .A1(n17701), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17664) );
  OAI21_X1 U20789 ( .B1(n17665), .B2(n17670), .A(n17664), .ZN(P3_U2748) );
  AOI22_X1 U20790 ( .A1(n17701), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17666) );
  OAI21_X1 U20791 ( .B1(n17667), .B2(n17670), .A(n17666), .ZN(P3_U2749) );
  AOI22_X1 U20792 ( .A1(n17701), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17668) );
  OAI21_X1 U20793 ( .B1(n17709), .B2(n17670), .A(n17668), .ZN(P3_U2750) );
  AOI22_X1 U20794 ( .A1(n17701), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17669) );
  OAI21_X1 U20795 ( .B1(n17671), .B2(n17670), .A(n17669), .ZN(P3_U2751) );
  INV_X1 U20796 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17754) );
  AOI22_X1 U20797 ( .A1(n17701), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17673) );
  OAI21_X1 U20798 ( .B1(n17754), .B2(n17703), .A(n17673), .ZN(P3_U2752) );
  AOI22_X1 U20799 ( .A1(n17701), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17674) );
  OAI21_X1 U20800 ( .B1(n17749), .B2(n17703), .A(n17674), .ZN(P3_U2753) );
  INV_X1 U20801 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17676) );
  AOI22_X1 U20802 ( .A1(n17701), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17675) );
  OAI21_X1 U20803 ( .B1(n17676), .B2(n17703), .A(n17675), .ZN(P3_U2754) );
  AOI22_X1 U20804 ( .A1(n17701), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17677) );
  OAI21_X1 U20805 ( .B1(n17678), .B2(n17703), .A(n17677), .ZN(P3_U2755) );
  INV_X1 U20806 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17680) );
  AOI22_X1 U20807 ( .A1(n17701), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17688), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17679) );
  OAI21_X1 U20808 ( .B1(n17680), .B2(n17703), .A(n17679), .ZN(P3_U2756) );
  INV_X1 U20809 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17682) );
  AOI22_X1 U20810 ( .A1(n17701), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17688), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17681) );
  OAI21_X1 U20811 ( .B1(n17682), .B2(n17703), .A(n17681), .ZN(P3_U2757) );
  AOI22_X1 U20812 ( .A1(n17701), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17688), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17683) );
  OAI21_X1 U20813 ( .B1(n21224), .B2(n17703), .A(n17683), .ZN(P3_U2758) );
  AOI22_X1 U20814 ( .A1(n17701), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17688), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17684) );
  OAI21_X1 U20815 ( .B1(n17685), .B2(n17703), .A(n17684), .ZN(P3_U2759) );
  INV_X1 U20816 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17687) );
  AOI22_X1 U20817 ( .A1(n17701), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17688), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17686) );
  OAI21_X1 U20818 ( .B1(n17687), .B2(n17703), .A(n17686), .ZN(P3_U2760) );
  AOI22_X1 U20819 ( .A1(n17701), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17688), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17689) );
  OAI21_X1 U20820 ( .B1(n17690), .B2(n17703), .A(n17689), .ZN(P3_U2761) );
  INV_X1 U20821 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17692) );
  AOI22_X1 U20822 ( .A1(n17701), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17691) );
  OAI21_X1 U20823 ( .B1(n17692), .B2(n17703), .A(n17691), .ZN(P3_U2762) );
  AOI22_X1 U20824 ( .A1(n17701), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17693) );
  OAI21_X1 U20825 ( .B1(n17694), .B2(n17703), .A(n17693), .ZN(P3_U2763) );
  INV_X1 U20826 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17696) );
  AOI22_X1 U20827 ( .A1(n17701), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17695) );
  OAI21_X1 U20828 ( .B1(n17696), .B2(n17703), .A(n17695), .ZN(P3_U2764) );
  INV_X1 U20829 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17698) );
  AOI22_X1 U20830 ( .A1(n17701), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17697) );
  OAI21_X1 U20831 ( .B1(n17698), .B2(n17703), .A(n17697), .ZN(P3_U2765) );
  AOI22_X1 U20832 ( .A1(n17701), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17699) );
  OAI21_X1 U20833 ( .B1(n17726), .B2(n17703), .A(n17699), .ZN(P3_U2766) );
  INV_X1 U20834 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17704) );
  AOI22_X1 U20835 ( .A1(n17701), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17700), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17702) );
  OAI21_X1 U20836 ( .B1(n17704), .B2(n17703), .A(n17702), .ZN(P3_U2767) );
  OAI211_X1 U20837 ( .C1(n19113), .C2(n19112), .A(n17706), .B(n17705), .ZN(
        n17747) );
  NAND3_X1 U20838 ( .A1(n19112), .A2(n17706), .A3(n17705), .ZN(n17753) );
  INV_X2 U20839 ( .A(n17753), .ZN(n17743) );
  AOI22_X1 U20840 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17750), .ZN(n17707) );
  OAI21_X1 U20841 ( .B1(n18471), .B2(n17745), .A(n17707), .ZN(P3_U2768) );
  AOI22_X1 U20842 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17751), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17750), .ZN(n17708) );
  OAI21_X1 U20843 ( .B1(n17709), .B2(n17753), .A(n17708), .ZN(P3_U2769) );
  AOI22_X1 U20844 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17750), .ZN(n17710) );
  OAI21_X1 U20845 ( .B1(n18483), .B2(n17745), .A(n17710), .ZN(P3_U2770) );
  AOI22_X1 U20846 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17750), .ZN(n17711) );
  OAI21_X1 U20847 ( .B1(n18489), .B2(n17745), .A(n17711), .ZN(P3_U2771) );
  AOI22_X1 U20848 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17750), .ZN(n17712) );
  OAI21_X1 U20849 ( .B1(n18495), .B2(n17745), .A(n17712), .ZN(P3_U2772) );
  AOI22_X1 U20850 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17750), .ZN(n17713) );
  OAI21_X1 U20851 ( .B1(n18501), .B2(n17745), .A(n17713), .ZN(P3_U2773) );
  AOI22_X1 U20852 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17750), .ZN(n17714) );
  OAI21_X1 U20853 ( .B1(n18509), .B2(n17745), .A(n17714), .ZN(P3_U2774) );
  AOI22_X1 U20854 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17750), .ZN(n17715) );
  OAI21_X1 U20855 ( .B1(n18514), .B2(n17745), .A(n17715), .ZN(P3_U2775) );
  AOI22_X1 U20856 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17750), .ZN(n17716) );
  OAI21_X1 U20857 ( .B1(n17734), .B2(n17745), .A(n17716), .ZN(P3_U2776) );
  AOI22_X1 U20858 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17750), .ZN(n17717) );
  OAI21_X1 U20859 ( .B1(n17736), .B2(n17745), .A(n17717), .ZN(P3_U2777) );
  AOI22_X1 U20860 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17750), .ZN(n17718) );
  OAI21_X1 U20861 ( .B1(n17738), .B2(n17745), .A(n17718), .ZN(P3_U2778) );
  AOI22_X1 U20862 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17750), .ZN(n17719) );
  OAI21_X1 U20863 ( .B1(n17740), .B2(n17745), .A(n17719), .ZN(P3_U2779) );
  AOI22_X1 U20864 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17750), .ZN(n17720) );
  OAI21_X1 U20865 ( .B1(n17742), .B2(n17745), .A(n17720), .ZN(P3_U2780) );
  AOI22_X1 U20866 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17743), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17750), .ZN(n17721) );
  OAI21_X1 U20867 ( .B1(n17746), .B2(n17745), .A(n17721), .ZN(P3_U2781) );
  AOI22_X1 U20868 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17751), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17750), .ZN(n17722) );
  OAI21_X1 U20869 ( .B1(n17723), .B2(n17753), .A(n17722), .ZN(P3_U2782) );
  AOI22_X1 U20870 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17750), .ZN(n17724) );
  OAI21_X1 U20871 ( .B1(n18471), .B2(n17745), .A(n17724), .ZN(P3_U2783) );
  AOI22_X1 U20872 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17751), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17750), .ZN(n17725) );
  OAI21_X1 U20873 ( .B1(n17726), .B2(n17753), .A(n17725), .ZN(P3_U2784) );
  AOI22_X1 U20874 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17750), .ZN(n17727) );
  OAI21_X1 U20875 ( .B1(n18483), .B2(n17745), .A(n17727), .ZN(P3_U2785) );
  AOI22_X1 U20876 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17747), .ZN(n17728) );
  OAI21_X1 U20877 ( .B1(n18489), .B2(n17745), .A(n17728), .ZN(P3_U2786) );
  AOI22_X1 U20878 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17747), .ZN(n17729) );
  OAI21_X1 U20879 ( .B1(n18495), .B2(n17745), .A(n17729), .ZN(P3_U2787) );
  AOI22_X1 U20880 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17747), .ZN(n17730) );
  OAI21_X1 U20881 ( .B1(n18501), .B2(n17745), .A(n17730), .ZN(P3_U2788) );
  AOI22_X1 U20882 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17747), .ZN(n17731) );
  OAI21_X1 U20883 ( .B1(n18509), .B2(n17745), .A(n17731), .ZN(P3_U2789) );
  AOI22_X1 U20884 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17747), .ZN(n17732) );
  OAI21_X1 U20885 ( .B1(n18514), .B2(n17745), .A(n17732), .ZN(P3_U2790) );
  AOI22_X1 U20886 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17747), .ZN(n17733) );
  OAI21_X1 U20887 ( .B1(n17734), .B2(n17745), .A(n17733), .ZN(P3_U2791) );
  AOI22_X1 U20888 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17747), .ZN(n17735) );
  OAI21_X1 U20889 ( .B1(n17736), .B2(n17745), .A(n17735), .ZN(P3_U2792) );
  AOI22_X1 U20890 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17747), .ZN(n17737) );
  OAI21_X1 U20891 ( .B1(n17738), .B2(n17745), .A(n17737), .ZN(P3_U2793) );
  AOI22_X1 U20892 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17747), .ZN(n17739) );
  OAI21_X1 U20893 ( .B1(n17740), .B2(n17745), .A(n17739), .ZN(P3_U2794) );
  AOI22_X1 U20894 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17750), .ZN(n17741) );
  OAI21_X1 U20895 ( .B1(n17742), .B2(n17745), .A(n17741), .ZN(P3_U2795) );
  AOI22_X1 U20896 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17743), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17750), .ZN(n17744) );
  OAI21_X1 U20897 ( .B1(n17746), .B2(n17745), .A(n17744), .ZN(P3_U2796) );
  AOI22_X1 U20898 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17751), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17747), .ZN(n17748) );
  OAI21_X1 U20899 ( .B1(n17749), .B2(n17753), .A(n17748), .ZN(P3_U2797) );
  AOI22_X1 U20900 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17751), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17750), .ZN(n17752) );
  OAI21_X1 U20901 ( .B1(n17754), .B2(n17753), .A(n17752), .ZN(P3_U2798) );
  NOR2_X1 U20902 ( .A1(n9802), .A2(n18115), .ZN(n17869) );
  OAI22_X1 U20903 ( .A1(n18139), .A2(n17971), .B1(n18131), .B2(n18130), .ZN(
        n17789) );
  NOR2_X1 U20904 ( .A1(n18140), .A2(n17789), .ZN(n17756) );
  NOR3_X1 U20905 ( .A1(n17869), .A2(n17756), .A3(n17755), .ZN(n17764) );
  OAI211_X1 U20906 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17772), .B(n17976), .ZN(n17762) );
  INV_X1 U20907 ( .A(n18080), .ZN(n18030) );
  OAI21_X1 U20908 ( .B1(n17772), .B2(n18030), .A(n18125), .ZN(n17757) );
  AOI21_X1 U20909 ( .B1(n17839), .B2(n17758), .A(n17757), .ZN(n17782) );
  OAI21_X1 U20910 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17781), .A(
        n17782), .ZN(n17771) );
  AOI22_X1 U20911 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17771), .B1(
        n17979), .B2(n17759), .ZN(n17761) );
  OAI211_X1 U20912 ( .C1(n10174), .C2(n17762), .A(n17761), .B(n17760), .ZN(
        n17763) );
  AOI211_X1 U20913 ( .C1(n17765), .C2(n17777), .A(n17764), .B(n17763), .ZN(
        n17770) );
  OAI211_X1 U20914 ( .C1(n17768), .C2(n17767), .A(n18039), .B(n17766), .ZN(
        n17769) );
  NAND2_X1 U20915 ( .A1(n17770), .A2(n17769), .ZN(P3_U2802) );
  AOI22_X1 U20916 ( .A1(n18385), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17771), .ZN(n17779) );
  NAND2_X1 U20917 ( .A1(n17772), .A2(n17976), .ZN(n17775) );
  NOR2_X1 U20918 ( .A1(n17773), .A2(n9705), .ZN(n17774) );
  OAI22_X1 U20919 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17775), .B1(
        n18144), .B2(n18024), .ZN(n17776) );
  AOI221_X1 U20920 ( .B1(n17777), .B2(n18140), .C1(n17789), .C2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n17776), .ZN(n17778) );
  OAI211_X1 U20921 ( .C1(n17965), .C2(n17780), .A(n17779), .B(n17778), .ZN(
        P3_U2803) );
  NAND4_X1 U20922 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18178), .A3(
        n18133), .A4(n17787), .ZN(n18151) );
  NAND2_X1 U20923 ( .A1(n17965), .A2(n17781), .ZN(n17902) );
  INV_X1 U20924 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19047) );
  NOR2_X1 U20925 ( .A1(n18384), .A2(n19047), .ZN(n18146) );
  AOI221_X1 U20926 ( .B1(n18507), .B2(n21234), .C1(n17783), .C2(n21234), .A(
        n17782), .ZN(n17784) );
  AOI211_X1 U20927 ( .C1(n17785), .C2(n17902), .A(n18146), .B(n17784), .ZN(
        n17791) );
  OAI21_X1 U20928 ( .B1(n17788), .B2(n17787), .A(n17786), .ZN(n18147) );
  AOI22_X1 U20929 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17789), .B1(
        n18039), .B2(n18147), .ZN(n17790) );
  OAI211_X1 U20930 ( .C1(n17927), .C2(n18151), .A(n17791), .B(n17790), .ZN(
        P3_U2804) );
  XOR2_X1 U20931 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17792), .Z(
        n18158) );
  AOI21_X1 U20932 ( .B1(n18854), .B2(n17794), .A(n18079), .ZN(n17822) );
  OAI21_X1 U20933 ( .B1(n17793), .B2(n18126), .A(n17822), .ZN(n17810) );
  NOR2_X1 U20934 ( .A1(n17880), .A2(n17794), .ZN(n17812) );
  OAI211_X1 U20935 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17812), .B(n17795), .ZN(n17797) );
  NOR2_X1 U20936 ( .A1(n18384), .A2(n19045), .ZN(n18160) );
  INV_X1 U20937 ( .A(n18160), .ZN(n17796) );
  OAI211_X1 U20938 ( .C1(n17965), .C2(n17798), .A(n17797), .B(n17796), .ZN(
        n17804) );
  XOR2_X1 U20939 ( .A(n17799), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18164) );
  OAI21_X1 U20940 ( .B1(n18038), .B2(n17801), .A(n17800), .ZN(n17802) );
  XOR2_X1 U20941 ( .A(n17802), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18157) );
  OAI22_X1 U20942 ( .A1(n17971), .A2(n18164), .B1(n18024), .B2(n18157), .ZN(
        n17803) );
  AOI211_X1 U20943 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17810), .A(
        n17804), .B(n17803), .ZN(n17805) );
  OAI21_X1 U20944 ( .B1(n18130), .B2(n18158), .A(n17805), .ZN(P3_U2805) );
  OR2_X1 U20945 ( .A1(n17806), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18177) );
  AOI22_X1 U20946 ( .A1(n18385), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17979), 
        .B2(n17807), .ZN(n17808) );
  INV_X1 U20947 ( .A(n17808), .ZN(n17809) );
  AOI221_X1 U20948 ( .B1(n17812), .B2(n17811), .C1(n17810), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17809), .ZN(n17817) );
  OAI22_X1 U20949 ( .A1(n17828), .A2(n17971), .B1(n18170), .B2(n18130), .ZN(
        n17832) );
  OAI21_X1 U20950 ( .B1(n17815), .B2(n17814), .A(n17813), .ZN(n18166) );
  AOI22_X1 U20951 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17832), .B1(
        n18039), .B2(n18166), .ZN(n17816) );
  OAI211_X1 U20952 ( .C1(n17927), .C2(n18177), .A(n17817), .B(n17816), .ZN(
        P3_U2806) );
  OAI22_X1 U20953 ( .A1(n17818), .A2(n17835), .B1(n18038), .B2(n18195), .ZN(
        n17820) );
  NOR2_X1 U20954 ( .A1(n17820), .A2(n17819), .ZN(n17821) );
  XOR2_X1 U20955 ( .A(n17821), .B(n18171), .Z(n18183) );
  NOR2_X1 U20956 ( .A1(n18384), .A2(n19040), .ZN(n18179) );
  NAND2_X1 U20957 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17842) );
  NAND2_X1 U20958 ( .A1(n9787), .A2(n17976), .ZN(n17857) );
  NOR2_X1 U20959 ( .A1(n17842), .A2(n17857), .ZN(n17825) );
  OAI21_X1 U20960 ( .B1(n18126), .B2(n17823), .A(n17822), .ZN(n17824) );
  MUX2_X1 U20961 ( .A(n17825), .B(n17824), .S(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .Z(n17826) );
  AOI211_X1 U20962 ( .C1(n17827), .C2(n17979), .A(n18179), .B(n17826), .ZN(
        n17834) );
  INV_X1 U20963 ( .A(n17828), .ZN(n18167) );
  NAND2_X1 U20964 ( .A1(n9802), .A2(n18167), .ZN(n17830) );
  NAND4_X1 U20965 ( .A1(n18115), .A2(n18237), .A3(n18171), .A4(n17939), .ZN(
        n17829) );
  OAI21_X1 U20966 ( .B1(n17830), .B2(n18265), .A(n17829), .ZN(n17831) );
  AOI22_X1 U20967 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17832), .B1(
        n18178), .B2(n17831), .ZN(n17833) );
  OAI211_X1 U20968 ( .C1(n18024), .C2(n18183), .A(n17834), .B(n17833), .ZN(
        P3_U2807) );
  INV_X1 U20969 ( .A(n17835), .ZN(n17836) );
  AOI221_X1 U20970 ( .B1(n17914), .B2(n17836), .C1(n18190), .C2(n17836), .A(
        n17819), .ZN(n17837) );
  XOR2_X1 U20971 ( .A(n18195), .B(n17837), .Z(n18202) );
  NAND2_X1 U20972 ( .A1(n18385), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18201) );
  INV_X1 U20973 ( .A(n18201), .ZN(n17846) );
  AOI21_X1 U20974 ( .B1(n17839), .B2(n17838), .A(n18079), .ZN(n17840) );
  OAI21_X1 U20975 ( .B1(n9787), .B2(n18030), .A(n17840), .ZN(n17866) );
  AOI21_X1 U20976 ( .B1(n17841), .B2(n17863), .A(n17866), .ZN(n17855) );
  OAI21_X1 U20977 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17842), .ZN(n17843) );
  OAI22_X1 U20978 ( .A1(n17855), .A2(n17844), .B1(n17857), .B2(n17843), .ZN(
        n17845) );
  AOI211_X1 U20979 ( .C1(n17847), .C2(n17979), .A(n17846), .B(n17845), .ZN(
        n17850) );
  INV_X1 U20980 ( .A(n18190), .ZN(n18199) );
  AOI22_X1 U20981 ( .A1(n9802), .A2(n18265), .B1(n18115), .B2(n18272), .ZN(
        n17926) );
  OAI21_X1 U20982 ( .B1(n18199), .B2(n17869), .A(n17926), .ZN(n17860) );
  OAI21_X1 U20983 ( .B1(n18190), .B2(n17927), .A(n18195), .ZN(n17848) );
  OAI21_X1 U20984 ( .B1(n18195), .B2(n17860), .A(n17848), .ZN(n17849) );
  OAI211_X1 U20985 ( .C1(n18024), .C2(n18202), .A(n17850), .B(n17849), .ZN(
        P3_U2808) );
  NAND3_X1 U20986 ( .A1(n18038), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17851), .ZN(n17874) );
  INV_X1 U20987 ( .A(n17852), .ZN(n17896) );
  OAI22_X1 U20988 ( .A1(n18207), .A2(n17874), .B1(n17896), .B2(n17853), .ZN(
        n17854) );
  XOR2_X1 U20989 ( .A(n18208), .B(n17854), .Z(n18215) );
  NAND2_X1 U20990 ( .A1(n18385), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18213) );
  OAI221_X1 U20991 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17857), .C1(
        n17856), .C2(n17855), .A(n18213), .ZN(n17858) );
  AOI21_X1 U20992 ( .B1(n17979), .B2(n17859), .A(n17858), .ZN(n17862) );
  NOR2_X1 U20993 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18207), .ZN(
        n18212) );
  NOR2_X1 U20994 ( .A1(n18204), .A2(n17927), .ZN(n17886) );
  AOI22_X1 U20995 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17860), .B1(
        n18212), .B2(n17886), .ZN(n17861) );
  OAI211_X1 U20996 ( .C1(n18215), .C2(n18024), .A(n17862), .B(n17861), .ZN(
        P3_U2809) );
  OAI21_X1 U20997 ( .B1(n18507), .B2(n17864), .A(n17863), .ZN(n17865) );
  AOI22_X1 U20998 ( .A1(n17867), .A2(n17902), .B1(n17866), .B2(n17865), .ZN(
        n17873) );
  NAND2_X1 U20999 ( .A1(n17868), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18217) );
  INV_X1 U21000 ( .A(n18217), .ZN(n18185) );
  OAI21_X1 U21001 ( .B1(n17869), .B2(n18185), .A(n17926), .ZN(n17885) );
  INV_X1 U21002 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18228) );
  AOI221_X1 U21003 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17874), 
        .C1(n18228), .C2(n17894), .A(n17819), .ZN(n17870) );
  XOR2_X1 U21004 ( .A(n17870), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n18222) );
  AOI22_X1 U21005 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17885), .B1(
        n18039), .B2(n18222), .ZN(n17872) );
  NAND3_X1 U21006 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17886), .A3(
        n18225), .ZN(n17871) );
  NAND2_X1 U21007 ( .A1(n18385), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18223) );
  NAND4_X1 U21008 ( .A1(n17873), .A2(n17872), .A3(n17871), .A4(n18223), .ZN(
        P3_U2810) );
  OAI21_X1 U21009 ( .B1(n17894), .B2(n17896), .A(n17874), .ZN(n17875) );
  XOR2_X1 U21010 ( .A(n17875), .B(n18228), .Z(n18232) );
  INV_X1 U21011 ( .A(n18122), .ZN(n18060) );
  OAI21_X1 U21012 ( .B1(n18079), .B2(n17879), .A(n18060), .ZN(n17904) );
  OAI21_X1 U21013 ( .B1(n17877), .B2(n18126), .A(n17904), .ZN(n17890) );
  AOI22_X1 U21014 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17890), .B1(
        n17979), .B2(n17878), .ZN(n17883) );
  NOR2_X1 U21015 ( .A1(n17880), .A2(n17879), .ZN(n17892) );
  OAI211_X1 U21016 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17892), .B(n17881), .ZN(n17882) );
  OAI211_X1 U21017 ( .C1(n19032), .C2(n18384), .A(n17883), .B(n17882), .ZN(
        n17884) );
  AOI221_X1 U21018 ( .B1(n17886), .B2(n18228), .C1(n17885), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17884), .ZN(n17887) );
  OAI21_X1 U21019 ( .B1(n18232), .B2(n18024), .A(n17887), .ZN(P3_U2811) );
  NAND2_X1 U21020 ( .A1(n17893), .A2(n17895), .ZN(n18247) );
  INV_X1 U21021 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17891) );
  OAI22_X1 U21022 ( .A1(n18384), .A2(n19030), .B1(n17965), .B2(n17888), .ZN(
        n17889) );
  AOI221_X1 U21023 ( .B1(n17892), .B2(n17891), .C1(n17890), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17889), .ZN(n17899) );
  OAI21_X1 U21024 ( .B1(n17893), .B2(n17927), .A(n17926), .ZN(n17910) );
  OAI21_X1 U21025 ( .B1(n17933), .B2(n17895), .A(n17894), .ZN(n17897) );
  XOR2_X1 U21026 ( .A(n17897), .B(n17896), .Z(n18243) );
  AOI22_X1 U21027 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17910), .B1(
        n18039), .B2(n18243), .ZN(n17898) );
  OAI211_X1 U21028 ( .C1(n17927), .C2(n18247), .A(n17899), .B(n17898), .ZN(
        P3_U2812) );
  AOI21_X1 U21029 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17901), .A(
        n17900), .ZN(n18255) );
  INV_X1 U21030 ( .A(n17902), .ZN(n18101) );
  NOR2_X1 U21031 ( .A1(n18384), .A2(n19028), .ZN(n18252) );
  INV_X1 U21032 ( .A(n17903), .ZN(n17905) );
  AOI221_X1 U21033 ( .B1(n18507), .B2(n17906), .C1(n17905), .C2(n17906), .A(
        n17904), .ZN(n17907) );
  AOI211_X1 U21034 ( .C1(n17908), .C2(n17902), .A(n18252), .B(n17907), .ZN(
        n17912) );
  INV_X1 U21035 ( .A(n17927), .ZN(n17909) );
  NOR2_X1 U21036 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21233), .ZN(
        n18249) );
  AOI22_X1 U21037 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17910), .B1(
        n17909), .B2(n18249), .ZN(n17911) );
  OAI211_X1 U21038 ( .C1(n18255), .C2(n18024), .A(n17912), .B(n17911), .ZN(
        P3_U2813) );
  AND2_X1 U21039 ( .A1(n18038), .A2(n17913), .ZN(n18010) );
  AOI22_X1 U21040 ( .A1(n18010), .A2(n18237), .B1(n17914), .B2(n17933), .ZN(
        n17915) );
  XOR2_X1 U21041 ( .A(n21233), .B(n17915), .Z(n18261) );
  NAND2_X1 U21042 ( .A1(n17916), .A2(n17976), .ZN(n17929) );
  AOI221_X1 U21043 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C1(n17918), .C2(n17917), .A(
        n17929), .ZN(n17924) );
  AOI21_X1 U21044 ( .B1(n18080), .B2(n17919), .A(n18079), .ZN(n17945) );
  OAI21_X1 U21045 ( .B1(n17920), .B2(n18126), .A(n17945), .ZN(n17932) );
  AOI22_X1 U21046 ( .A1(n18385), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17932), .ZN(n17921) );
  OAI21_X1 U21047 ( .B1(n17965), .B2(n17922), .A(n17921), .ZN(n17923) );
  AOI211_X1 U21048 ( .C1(n18039), .C2(n18261), .A(n17924), .B(n17923), .ZN(
        n17925) );
  OAI221_X1 U21049 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17927), 
        .C1(n21233), .C2(n17926), .A(n17925), .ZN(P3_U2814) );
  NOR2_X1 U21050 ( .A1(n17950), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18266) );
  NAND2_X1 U21051 ( .A1(n9802), .A2(n18265), .ZN(n17943) );
  NAND2_X1 U21052 ( .A1(n18385), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18278) );
  INV_X1 U21053 ( .A(n18278), .ZN(n17931) );
  OAI22_X1 U21054 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17929), .B1(
        n17928), .B2(n17965), .ZN(n17930) );
  AOI211_X1 U21055 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17932), .A(
        n17931), .B(n17930), .ZN(n17942) );
  NOR2_X1 U21056 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17937) );
  INV_X1 U21057 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17985) );
  NOR2_X1 U21058 ( .A1(n17933), .A2(n17985), .ZN(n17958) );
  NOR2_X1 U21059 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17934), .ZN(
        n18011) );
  NAND3_X1 U21060 ( .A1(n17988), .A2(n18011), .A3(n17991), .ZN(n17956) );
  NOR2_X1 U21061 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17956), .ZN(
        n17952) );
  INV_X1 U21062 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18290) );
  INV_X1 U21063 ( .A(n18300), .ZN(n18312) );
  NOR4_X1 U21064 ( .A1(n18290), .A2(n18312), .A3(n18286), .A4(n17935), .ZN(
        n17936) );
  OAI22_X1 U21065 ( .A1(n17937), .A2(n17958), .B1(n17952), .B2(n17936), .ZN(
        n17938) );
  XOR2_X1 U21066 ( .A(n18274), .B(n17938), .Z(n18277) );
  AND2_X1 U21067 ( .A1(n18272), .A2(n18115), .ZN(n17940) );
  INV_X1 U21068 ( .A(n18283), .ZN(n18282) );
  NAND4_X1 U21069 ( .A1(n18282), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n17939), .ZN(n17944) );
  NAND2_X1 U21070 ( .A1(n18274), .A2(n17944), .ZN(n18276) );
  AOI22_X1 U21071 ( .A1(n18039), .A2(n18277), .B1(n17940), .B2(n18276), .ZN(
        n17941) );
  OAI211_X1 U21072 ( .C1(n18266), .C2(n17943), .A(n17942), .B(n17941), .ZN(
        P3_U2815) );
  NOR2_X1 U21073 ( .A1(n18324), .A2(n18283), .ZN(n18304) );
  OAI221_X1 U21074 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18304), .A(n17944), .ZN(
        n18298) );
  AOI221_X1 U21075 ( .B1(n18507), .B2(n17947), .C1(n17946), .C2(n17947), .A(
        n17945), .ZN(n17948) );
  NOR2_X1 U21076 ( .A1(n18384), .A2(n19023), .ZN(n18293) );
  AOI211_X1 U21077 ( .C1(n17949), .C2(n17902), .A(n17948), .B(n18293), .ZN(
        n17955) );
  NOR2_X1 U21078 ( .A1(n18322), .A2(n18283), .ZN(n18302) );
  INV_X1 U21079 ( .A(n18302), .ZN(n17951) );
  AOI221_X1 U21080 ( .B1(n18286), .B2(n18290), .C1(n17951), .C2(n18290), .A(
        n17950), .ZN(n18295) );
  AOI22_X1 U21081 ( .A1(n18010), .A2(n18285), .B1(n17952), .B2(n17985), .ZN(
        n17953) );
  XOR2_X1 U21082 ( .A(n18290), .B(n17953), .Z(n18294) );
  AOI22_X1 U21083 ( .A1(n9802), .A2(n18295), .B1(n18039), .B2(n18294), .ZN(
        n17954) );
  OAI211_X1 U21084 ( .C1(n18130), .C2(n18298), .A(n17955), .B(n17954), .ZN(
        P3_U2816) );
  INV_X1 U21085 ( .A(n17956), .ZN(n17974) );
  NOR2_X1 U21086 ( .A1(n18312), .A2(n17935), .ZN(n17957) );
  OAI22_X1 U21087 ( .A1(n17958), .A2(n17974), .B1(n17957), .B2(n17985), .ZN(
        n17959) );
  XOR2_X1 U21088 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17959), .Z(
        n18311) );
  OAI21_X1 U21089 ( .B1(n18030), .B2(n17977), .A(n18126), .ZN(n17960) );
  AOI21_X1 U21090 ( .B1(n17961), .B2(n17960), .A(n18079), .ZN(n17962) );
  INV_X1 U21091 ( .A(n17962), .ZN(n17980) );
  NOR2_X1 U21092 ( .A1(n18384), .A2(n19020), .ZN(n17970) );
  NOR2_X1 U21093 ( .A1(n17964), .A2(n17963), .ZN(n17968) );
  OAI211_X1 U21094 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17977), .B(n17976), .ZN(n17967) );
  OAI22_X1 U21095 ( .A1(n17968), .A2(n17967), .B1(n17966), .B2(n17965), .ZN(
        n17969) );
  AOI211_X1 U21096 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17980), .A(
        n17970), .B(n17969), .ZN(n17973) );
  OAI22_X1 U21097 ( .A1(n18304), .A2(n18130), .B1(n18302), .B2(n17971), .ZN(
        n17984) );
  NOR2_X1 U21098 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18283), .ZN(
        n18299) );
  AOI22_X1 U21099 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17984), .B1(
        n18299), .B2(n18020), .ZN(n17972) );
  OAI211_X1 U21100 ( .C1(n18024), .C2(n18311), .A(n17973), .B(n17972), .ZN(
        P3_U2817) );
  AOI21_X1 U21101 ( .B1(n18010), .B2(n18300), .A(n17974), .ZN(n17975) );
  XOR2_X1 U21102 ( .A(n17975), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18320) );
  NAND2_X1 U21103 ( .A1(n17977), .A2(n17976), .ZN(n17982) );
  AOI22_X1 U21104 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17980), .B1(
        n17979), .B2(n17978), .ZN(n17981) );
  NAND2_X1 U21105 ( .A1(n18385), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18318) );
  OAI211_X1 U21106 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17982), .A(
        n17981), .B(n18318), .ZN(n17983) );
  AOI21_X1 U21107 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17984), .A(
        n17983), .ZN(n17987) );
  NAND3_X1 U21108 ( .A1(n18300), .A2(n17985), .A3(n18020), .ZN(n17986) );
  OAI211_X1 U21109 ( .C1(n18320), .C2(n18024), .A(n17987), .B(n17986), .ZN(
        P3_U2818) );
  INV_X1 U21110 ( .A(n18329), .ZN(n17989) );
  AOI22_X1 U21111 ( .A1(n17989), .A2(n18010), .B1(n17988), .B2(n18011), .ZN(
        n17990) );
  XOR2_X1 U21112 ( .A(n17990), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18335) );
  NOR2_X1 U21113 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18329), .ZN(
        n18321) );
  AOI22_X1 U21114 ( .A1(n9802), .A2(n18322), .B1(n18115), .B2(n18324), .ZN(
        n18019) );
  NAND2_X1 U21115 ( .A1(n18329), .A2(n18020), .ZN(n18000) );
  AOI21_X1 U21116 ( .B1(n18019), .B2(n18000), .A(n17991), .ZN(n17997) );
  OR2_X1 U21117 ( .A1(n18507), .A2(n17992), .ZN(n17999) );
  OAI21_X1 U21118 ( .B1(n17992), .B2(n18507), .A(n18060), .ZN(n18008) );
  AOI22_X1 U21119 ( .A1(n18385), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17993), 
        .B2(n17902), .ZN(n17994) );
  OAI221_X1 U21120 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17999), .C1(
        n17995), .C2(n18008), .A(n17994), .ZN(n17996) );
  AOI211_X1 U21121 ( .C1(n18321), .C2(n18020), .A(n17997), .B(n17996), .ZN(
        n17998) );
  OAI21_X1 U21122 ( .B1(n18335), .B2(n18024), .A(n17998), .ZN(P3_U2819) );
  NAND3_X1 U21123 ( .A1(n18854), .A2(n18029), .A3(n18027), .ZN(n18015) );
  NOR2_X1 U21124 ( .A1(n18014), .A2(n18015), .ZN(n18013) );
  AOI22_X1 U21125 ( .A1(n18385), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18013), 
        .B2(n17999), .ZN(n18007) );
  OAI21_X1 U21126 ( .B1(n18019), .B2(n18339), .A(n18000), .ZN(n18004) );
  AOI22_X1 U21127 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18010), .B1(
        n18011), .B2(n18343), .ZN(n18001) );
  XOR2_X1 U21128 ( .A(n18001), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(
        n18342) );
  OAI22_X1 U21129 ( .A1(n18101), .A2(n18002), .B1(n18342), .B2(n18024), .ZN(
        n18003) );
  AOI21_X1 U21130 ( .B1(n18005), .B2(n18004), .A(n18003), .ZN(n18006) );
  OAI211_X1 U21131 ( .C1(n18009), .C2(n18008), .A(n18007), .B(n18006), .ZN(
        P3_U2820) );
  NOR2_X1 U21132 ( .A1(n18011), .A2(n18010), .ZN(n18012) );
  XOR2_X1 U21133 ( .A(n18012), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18353) );
  AOI211_X1 U21134 ( .C1(n18015), .C2(n18014), .A(n18122), .B(n18013), .ZN(
        n18017) );
  NOR2_X1 U21135 ( .A1(n18384), .A2(n19013), .ZN(n18016) );
  AOI211_X1 U21136 ( .C1(n18018), .C2(n17902), .A(n18017), .B(n18016), .ZN(
        n18023) );
  INV_X1 U21137 ( .A(n18019), .ZN(n18021) );
  AOI22_X1 U21138 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18021), .B1(
        n18020), .B2(n18343), .ZN(n18022) );
  OAI211_X1 U21139 ( .C1(n18353), .C2(n18024), .A(n18023), .B(n18022), .ZN(
        P3_U2821) );
  OAI21_X1 U21140 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18026), .A(
        n18025), .ZN(n18371) );
  NAND2_X1 U21141 ( .A1(n18029), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18028) );
  AOI211_X1 U21142 ( .C1(n18031), .C2(n18028), .A(n18027), .B(n18507), .ZN(
        n18035) );
  OAI21_X1 U21143 ( .B1(n18030), .B2(n18029), .A(n18125), .ZN(n18047) );
  INV_X1 U21144 ( .A(n18047), .ZN(n18032) );
  OAI22_X1 U21145 ( .A1(n18101), .A2(n18033), .B1(n18032), .B2(n18031), .ZN(
        n18034) );
  AOI211_X1 U21146 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n18385), .A(n18035), .B(
        n18034), .ZN(n18041) );
  OAI21_X1 U21147 ( .B1(n18038), .B2(n18036), .A(n18037), .ZN(n18366) );
  AOI22_X1 U21148 ( .A1(n9802), .A2(n18036), .B1(n18039), .B2(n18366), .ZN(
        n18040) );
  OAI211_X1 U21149 ( .C1(n18130), .C2(n18371), .A(n18041), .B(n18040), .ZN(
        P3_U2822) );
  OAI21_X1 U21150 ( .B1(n18044), .B2(n18043), .A(n18042), .ZN(n18045) );
  XOR2_X1 U21151 ( .A(n18045), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18382) );
  NOR2_X1 U21152 ( .A1(n18507), .A2(n18046), .ZN(n18049) );
  NOR2_X1 U21153 ( .A1(n18384), .A2(n19009), .ZN(n18373) );
  AOI221_X1 U21154 ( .B1(n18049), .B2(n18048), .C1(n18047), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18373), .ZN(n18054) );
  AOI21_X1 U21155 ( .B1(n18378), .B2(n18051), .A(n18050), .ZN(n18374) );
  AOI22_X1 U21156 ( .A1(n18118), .A2(n18374), .B1(n18052), .B2(n17902), .ZN(
        n18053) );
  OAI211_X1 U21157 ( .C1(n18130), .C2(n18382), .A(n18054), .B(n18053), .ZN(
        P3_U2823) );
  OAI21_X1 U21158 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18056), .A(
        n18055), .ZN(n18391) );
  NOR2_X1 U21159 ( .A1(n18507), .A2(n18061), .ZN(n18057) );
  AOI22_X1 U21160 ( .A1(n18385), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18057), 
        .B2(n18062), .ZN(n18066) );
  AOI21_X1 U21161 ( .B1(n9786), .B2(n18059), .A(n18058), .ZN(n18389) );
  OAI21_X1 U21162 ( .B1(n18061), .B2(n18507), .A(n18060), .ZN(n18074) );
  OAI22_X1 U21163 ( .A1(n18101), .A2(n18063), .B1(n18062), .B2(n18074), .ZN(
        n18064) );
  AOI21_X1 U21164 ( .B1(n18118), .B2(n18389), .A(n18064), .ZN(n18065) );
  OAI211_X1 U21165 ( .C1(n18130), .C2(n18391), .A(n18066), .B(n18065), .ZN(
        P3_U2824) );
  OAI21_X1 U21166 ( .B1(n18069), .B2(n18068), .A(n18067), .ZN(n18400) );
  AOI21_X1 U21167 ( .B1(n18072), .B2(n18071), .A(n18070), .ZN(n18397) );
  AOI21_X1 U21168 ( .B1(n18073), .B2(n18125), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18075) );
  OAI22_X1 U21169 ( .A1(n18101), .A2(n18076), .B1(n18075), .B2(n18074), .ZN(
        n18077) );
  AOI21_X1 U21170 ( .B1(n18118), .B2(n18397), .A(n18077), .ZN(n18078) );
  NAND2_X1 U21171 ( .A1(n18385), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18398) );
  OAI211_X1 U21172 ( .C1(n18130), .C2(n18400), .A(n18078), .B(n18398), .ZN(
        P3_U2825) );
  AOI21_X1 U21173 ( .B1(n18080), .B2(n18085), .A(n18079), .ZN(n18105) );
  AOI21_X1 U21174 ( .B1(n18083), .B2(n18082), .A(n18081), .ZN(n18084) );
  XOR2_X1 U21175 ( .A(n18084), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18402) );
  NOR2_X1 U21176 ( .A1(n18384), .A2(n19003), .ZN(n18401) );
  NOR3_X1 U21177 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18085), .A3(
        n18507), .ZN(n18086) );
  AOI211_X1 U21178 ( .C1(n18115), .C2(n18402), .A(n18401), .B(n18086), .ZN(
        n18092) );
  AOI21_X1 U21179 ( .B1(n18089), .B2(n18088), .A(n18087), .ZN(n18405) );
  AOI22_X1 U21180 ( .A1(n18118), .A2(n18405), .B1(n18090), .B2(n17902), .ZN(
        n18091) );
  OAI211_X1 U21181 ( .C1(n18093), .C2(n18105), .A(n18092), .B(n18091), .ZN(
        P3_U2826) );
  INV_X1 U21182 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18104) );
  NAND2_X1 U21183 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18125), .ZN(
        n18110) );
  AOI21_X1 U21184 ( .B1(n18096), .B2(n18095), .A(n18094), .ZN(n18415) );
  NOR2_X1 U21185 ( .A1(n18384), .A2(n19000), .ZN(n18414) );
  OAI21_X1 U21186 ( .B1(n18099), .B2(n18098), .A(n18097), .ZN(n18420) );
  OAI22_X1 U21187 ( .A1(n18101), .A2(n18100), .B1(n18130), .B2(n18420), .ZN(
        n18102) );
  AOI211_X1 U21188 ( .C1(n18118), .C2(n18415), .A(n18414), .B(n18102), .ZN(
        n18103) );
  OAI221_X1 U21189 ( .B1(n18105), .B2(n18104), .C1(n18105), .C2(n18110), .A(
        n18103), .ZN(P3_U2827) );
  AOI21_X1 U21190 ( .B1(n18108), .B2(n18107), .A(n18106), .ZN(n18436) );
  AOI22_X1 U21191 ( .A1(n18118), .A2(n18436), .B1(n18109), .B2(n17902), .ZN(
        n18113) );
  OAI21_X1 U21192 ( .B1(n18854), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n18110), .ZN(n18112) );
  NAND2_X1 U21193 ( .A1(n18385), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18437) );
  OAI211_X1 U21194 ( .C1(n18431), .C2(n18430), .A(n18115), .B(n18429), .ZN(
        n18111) );
  NAND4_X1 U21195 ( .A1(n18113), .A2(n18112), .A3(n18437), .A4(n18111), .ZN(
        P3_U2828) );
  NOR2_X1 U21196 ( .A1(n18124), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18114) );
  XNOR2_X1 U21197 ( .A(n18117), .B(n18114), .ZN(n18442) );
  AOI22_X1 U21198 ( .A1(n18115), .A2(n18442), .B1(n18385), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18120) );
  AOI21_X1 U21199 ( .B1(n18123), .B2(n18117), .A(n18116), .ZN(n18440) );
  AOI22_X1 U21200 ( .A1(n18118), .A2(n18440), .B1(n18121), .B2(n17902), .ZN(
        n18119) );
  OAI211_X1 U21201 ( .C1(n18122), .C2(n18121), .A(n18120), .B(n18119), .ZN(
        P3_U2829) );
  OAI21_X1 U21202 ( .B1(n18124), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18123), .ZN(n18456) );
  INV_X1 U21203 ( .A(n18456), .ZN(n18458) );
  NAND3_X1 U21204 ( .A1(n19075), .A2(n18126), .A3(n18125), .ZN(n18127) );
  AOI22_X1 U21205 ( .A1(n18385), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18127), .ZN(n18128) );
  OAI221_X1 U21206 ( .B1(n18458), .B2(n18130), .C1(n18456), .C2(n18129), .A(
        n18128), .ZN(P3_U2830) );
  AOI22_X1 U21207 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18445), .B1(
        n18385), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n18143) );
  INV_X1 U21208 ( .A(n18131), .ZN(n18137) );
  NAND2_X1 U21209 ( .A1(n18937), .A2(n18330), .ZN(n18421) );
  INV_X1 U21210 ( .A(n18421), .ZN(n18354) );
  NAND2_X1 U21211 ( .A1(n9660), .A2(n19091), .ZN(n18423) );
  INV_X1 U21212 ( .A(n18423), .ZN(n18358) );
  AOI21_X1 U21213 ( .B1(n18132), .B2(n18421), .A(n18358), .ZN(n18169) );
  OAI21_X1 U21214 ( .B1(n18133), .B2(n18354), .A(n18169), .ZN(n18153) );
  OAI21_X1 U21215 ( .B1(n18135), .B2(n18354), .A(n18134), .ZN(n18136) );
  AOI211_X1 U21216 ( .C1(n18906), .C2(n18137), .A(n18153), .B(n18136), .ZN(
        n18138) );
  OAI21_X1 U21217 ( .B1(n18139), .B2(n18301), .A(n18138), .ZN(n18148) );
  OAI221_X1 U21218 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18141), 
        .C1(n18140), .C2(n18148), .A(n18451), .ZN(n18142) );
  OAI211_X1 U21219 ( .C1(n18144), .C2(n18352), .A(n18143), .B(n18142), .ZN(
        P3_U2835) );
  INV_X1 U21220 ( .A(n18145), .ZN(n18198) );
  NAND2_X1 U21221 ( .A1(n18451), .A2(n18198), .ZN(n18203) );
  AOI21_X1 U21222 ( .B1(n18367), .B2(n18147), .A(n18146), .ZN(n18150) );
  OAI211_X1 U21223 ( .C1(n18433), .C2(n18148), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n18384), .ZN(n18149) );
  OAI211_X1 U21224 ( .C1(n18203), .C2(n18151), .A(n18150), .B(n18149), .ZN(
        P3_U2836) );
  NAND2_X1 U21225 ( .A1(n18155), .A2(n18152), .ZN(n18162) );
  NOR3_X1 U21226 ( .A1(n18154), .A2(n18155), .A3(n18153), .ZN(n18156) );
  INV_X1 U21227 ( .A(n18445), .ZN(n18439) );
  OAI22_X1 U21228 ( .A1(n18156), .A2(n18433), .B1(n18155), .B2(n18439), .ZN(
        n18161) );
  OAI22_X1 U21229 ( .A1(n18457), .A2(n18158), .B1(n18352), .B2(n18157), .ZN(
        n18159) );
  AOI211_X1 U21230 ( .C1(n18162), .C2(n18161), .A(n18160), .B(n18159), .ZN(
        n18163) );
  OAI21_X1 U21231 ( .B1(n18165), .B2(n18164), .A(n18163), .ZN(P3_U2837) );
  AOI22_X1 U21232 ( .A1(n18385), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18367), 
        .B2(n18166), .ZN(n18176) );
  AOI21_X1 U21233 ( .B1(n18323), .B2(n18167), .A(n18445), .ZN(n18168) );
  OAI211_X1 U21234 ( .C1(n18170), .C2(n18303), .A(n18169), .B(n18168), .ZN(
        n18174) );
  AOI211_X1 U21235 ( .C1(n18933), .C2(n18172), .A(n18171), .B(n18174), .ZN(
        n18173) );
  NOR2_X1 U21236 ( .A1(n18385), .A2(n18173), .ZN(n18181) );
  OAI211_X1 U21237 ( .C1(n18359), .C2(n18174), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18181), .ZN(n18175) );
  OAI211_X1 U21238 ( .C1(n18177), .C2(n18203), .A(n18176), .B(n18175), .ZN(
        P3_U2838) );
  AND3_X1 U21239 ( .A1(n18439), .A2(n18178), .A3(n18198), .ZN(n18180) );
  AOI221_X1 U21240 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18181), 
        .C1(n18180), .C2(n18181), .A(n18179), .ZN(n18182) );
  OAI21_X1 U21241 ( .B1(n18352), .B2(n18183), .A(n18182), .ZN(P3_U2839) );
  AOI22_X1 U21242 ( .A1(n18906), .A2(n18272), .B1(n18323), .B2(n18265), .ZN(
        n18206) );
  INV_X1 U21243 ( .A(n18206), .ZN(n18194) );
  OAI22_X1 U21244 ( .A1(n18937), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n18184), .B2(n18924), .ZN(n18193) );
  NAND2_X1 U21245 ( .A1(n18303), .A2(n18301), .ZN(n18328) );
  AOI21_X1 U21246 ( .B1(n18186), .B2(n18185), .A(n18937), .ZN(n18187) );
  AOI21_X1 U21247 ( .B1(n18933), .B2(n18188), .A(n18187), .ZN(n18219) );
  OAI21_X1 U21248 ( .B1(n18937), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n18219), .ZN(n18189) );
  AOI21_X1 U21249 ( .B1(n18190), .B2(n18328), .A(n18189), .ZN(n18210) );
  OAI211_X1 U21250 ( .C1(n18191), .C2(n18330), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18210), .ZN(n18192) );
  NOR3_X1 U21251 ( .A1(n18194), .A2(n18193), .A3(n18192), .ZN(n18196) );
  OAI22_X1 U21252 ( .A1(n18196), .A2(n18433), .B1(n18195), .B2(n18439), .ZN(
        n18197) );
  OAI221_X1 U21253 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18199), 
        .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18198), .A(n18197), .ZN(
        n18200) );
  OAI211_X1 U21254 ( .C1(n18202), .C2(n18352), .A(n18201), .B(n18200), .ZN(
        P3_U2840) );
  NOR2_X1 U21255 ( .A1(n18204), .A2(n18203), .ZN(n18229) );
  NAND2_X1 U21256 ( .A1(n18330), .A2(n18924), .ZN(n18444) );
  AND2_X1 U21257 ( .A1(n9660), .A2(n18205), .ZN(n18216) );
  NAND2_X1 U21258 ( .A1(n18451), .A2(n18206), .ZN(n18260) );
  AOI211_X1 U21259 ( .C1(n18444), .C2(n18207), .A(n18216), .B(n18260), .ZN(
        n18209) );
  AOI211_X1 U21260 ( .C1(n18210), .C2(n18209), .A(n18385), .B(n18208), .ZN(
        n18211) );
  AOI21_X1 U21261 ( .B1(n18212), .B2(n18229), .A(n18211), .ZN(n18214) );
  OAI211_X1 U21262 ( .C1(n18215), .C2(n18352), .A(n18214), .B(n18213), .ZN(
        P3_U2841) );
  NOR2_X1 U21263 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19123), .ZN(
        n18220) );
  AOI211_X1 U21264 ( .C1(n18217), .C2(n18328), .A(n18216), .B(n18260), .ZN(
        n18218) );
  AOI21_X1 U21265 ( .B1(n18219), .B2(n18218), .A(n18385), .ZN(n18230) );
  AOI21_X1 U21266 ( .B1(n18220), .B2(n18444), .A(n18230), .ZN(n18226) );
  NOR2_X1 U21267 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18228), .ZN(
        n18221) );
  AOI22_X1 U21268 ( .A1(n18367), .A2(n18222), .B1(n18229), .B2(n18221), .ZN(
        n18224) );
  OAI211_X1 U21269 ( .C1(n18226), .C2(n18225), .A(n18224), .B(n18223), .ZN(
        P3_U2842) );
  NOR2_X1 U21270 ( .A1(n18384), .A2(n19032), .ZN(n18227) );
  AOI221_X1 U21271 ( .B1(n18230), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), 
        .C1(n18229), .C2(n18228), .A(n18227), .ZN(n18231) );
  OAI21_X1 U21272 ( .B1(n18232), .B2(n18352), .A(n18231), .ZN(P3_U2843) );
  OAI22_X1 U21273 ( .A1(n18428), .A2(n18924), .B1(n18406), .B2(n18425), .ZN(
        n18417) );
  INV_X1 U21274 ( .A(n18417), .ZN(n18361) );
  NOR2_X1 U21275 ( .A1(n18233), .A2(n18361), .ZN(n18375) );
  NAND2_X1 U21276 ( .A1(n18234), .A2(n18375), .ZN(n18289) );
  INV_X1 U21277 ( .A(n18289), .ZN(n18236) );
  NOR2_X1 U21278 ( .A1(n18236), .A2(n18235), .ZN(n18313) );
  NAND2_X1 U21279 ( .A1(n18237), .A2(n18344), .ZN(n18264) );
  NOR3_X1 U21280 ( .A1(n18358), .A2(n18238), .A3(n21233), .ZN(n18239) );
  OAI22_X1 U21281 ( .A1(n18240), .A2(n18924), .B1(n18354), .B2(n18239), .ZN(
        n18241) );
  AOI211_X1 U21282 ( .C1(n18242), .C2(n18328), .A(n18260), .B(n18241), .ZN(
        n18248) );
  AOI221_X1 U21283 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18248), 
        .C1(n18354), .C2(n18248), .A(n18385), .ZN(n18244) );
  AOI22_X1 U21284 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18244), .B1(
        n18367), .B2(n18243), .ZN(n18246) );
  NAND2_X1 U21285 ( .A1(n18385), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18245) );
  OAI211_X1 U21286 ( .C1(n18247), .C2(n18264), .A(n18246), .B(n18245), .ZN(
        P3_U2844) );
  NOR2_X1 U21287 ( .A1(n18385), .A2(n18248), .ZN(n18251) );
  INV_X1 U21288 ( .A(n18264), .ZN(n18250) );
  AOI22_X1 U21289 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18251), .B1(
        n18250), .B2(n18249), .ZN(n18254) );
  INV_X1 U21290 ( .A(n18252), .ZN(n18253) );
  OAI211_X1 U21291 ( .C1(n18255), .C2(n18352), .A(n18254), .B(n18253), .ZN(
        P3_U2845) );
  INV_X1 U21292 ( .A(n18267), .ZN(n18259) );
  NAND2_X1 U21293 ( .A1(n18256), .A2(n18933), .ZN(n18345) );
  INV_X1 U21294 ( .A(n18345), .ZN(n18307) );
  AOI21_X1 U21295 ( .B1(n18921), .B2(n18281), .A(n18307), .ZN(n18326) );
  OAI21_X1 U21296 ( .B1(n18274), .B2(n9660), .A(n18257), .ZN(n18258) );
  OAI211_X1 U21297 ( .C1(n18337), .C2(n18259), .A(n18326), .B(n18258), .ZN(
        n18269) );
  OAI221_X1 U21298 ( .B1(n18260), .B2(n18359), .C1(n18260), .C2(n18269), .A(
        n18384), .ZN(n18263) );
  AOI22_X1 U21299 ( .A1(n18385), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18367), 
        .B2(n18261), .ZN(n18262) );
  OAI221_X1 U21300 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18264), 
        .C1(n21233), .C2(n18263), .A(n18262), .ZN(P3_U2846) );
  AND2_X1 U21301 ( .A1(n18265), .A2(n18323), .ZN(n18271) );
  INV_X1 U21302 ( .A(n18266), .ZN(n18270) );
  OAI21_X1 U21303 ( .B1(n18267), .B2(n18289), .A(n18274), .ZN(n18268) );
  AOI22_X1 U21304 ( .A1(n18271), .A2(n18270), .B1(n18269), .B2(n18268), .ZN(
        n18280) );
  NAND2_X1 U21305 ( .A1(n18906), .A2(n18272), .ZN(n18273) );
  OAI22_X1 U21306 ( .A1(n18274), .A2(n18439), .B1(n18433), .B2(n18273), .ZN(
        n18275) );
  AOI22_X1 U21307 ( .A1(n18367), .A2(n18277), .B1(n18276), .B2(n18275), .ZN(
        n18279) );
  OAI211_X1 U21308 ( .C1(n18280), .C2(n18433), .A(n18279), .B(n18278), .ZN(
        P3_U2847) );
  INV_X1 U21309 ( .A(n18285), .ZN(n18291) );
  AOI21_X1 U21310 ( .B1(n18921), .B2(n18281), .A(n9660), .ZN(n18346) );
  AOI21_X1 U21311 ( .B1(n18347), .B2(n18282), .A(n18346), .ZN(n18306) );
  AOI211_X1 U21312 ( .C1(n18933), .C2(n18283), .A(n18307), .B(n18306), .ZN(
        n18284) );
  OAI211_X1 U21313 ( .C1(n18937), .C2(n18285), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18284), .ZN(n18287) );
  OAI221_X1 U21314 ( .B1(n18287), .B2(n18286), .C1(n18287), .C2(n18444), .A(
        n18451), .ZN(n18288) );
  AOI221_X1 U21315 ( .B1(n18291), .B2(n18290), .C1(n18289), .C2(n18290), .A(
        n18288), .ZN(n18292) );
  AOI211_X1 U21316 ( .C1(n18445), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18293), .B(n18292), .ZN(n18297) );
  AOI22_X1 U21317 ( .A1(n18368), .A2(n18295), .B1(n18367), .B2(n18294), .ZN(
        n18296) );
  OAI211_X1 U21318 ( .C1(n18457), .C2(n18298), .A(n18297), .B(n18296), .ZN(
        P3_U2848) );
  AOI22_X1 U21319 ( .A1(n18385), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18344), 
        .B2(n18299), .ZN(n18310) );
  NOR2_X1 U21320 ( .A1(n18337), .A2(n18300), .ZN(n18332) );
  OAI22_X1 U21321 ( .A1(n18304), .A2(n18303), .B1(n18302), .B2(n18301), .ZN(
        n18305) );
  NOR4_X1 U21322 ( .A1(n18307), .A2(n18306), .A3(n18332), .A4(n18305), .ZN(
        n18314) );
  OAI211_X1 U21323 ( .C1(n18337), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18451), .B(n18314), .ZN(n18308) );
  NAND3_X1 U21324 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18384), .A3(
        n18308), .ZN(n18309) );
  OAI211_X1 U21325 ( .C1(n18352), .C2(n18311), .A(n18310), .B(n18309), .ZN(
        P3_U2849) );
  NOR2_X1 U21326 ( .A1(n18313), .A2(n18312), .ZN(n18316) );
  INV_X1 U21327 ( .A(n18314), .ZN(n18315) );
  MUX2_X1 U21328 ( .A(n18316), .B(n18315), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n18317) );
  AOI22_X1 U21329 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18445), .B1(
        n18451), .B2(n18317), .ZN(n18319) );
  OAI211_X1 U21330 ( .C1(n18320), .C2(n18352), .A(n18319), .B(n18318), .ZN(
        P3_U2850) );
  AOI22_X1 U21331 ( .A1(n18385), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18344), 
        .B2(n18321), .ZN(n18334) );
  AOI22_X1 U21332 ( .A1(n18906), .A2(n18324), .B1(n18323), .B2(n18322), .ZN(
        n18325) );
  NAND2_X1 U21333 ( .A1(n18451), .A2(n18325), .ZN(n18349) );
  OAI221_X1 U21334 ( .B1(n18330), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n18330), .C2(n18347), .A(n18326), .ZN(n18327) );
  AOI211_X1 U21335 ( .C1(n18329), .C2(n18328), .A(n18349), .B(n18327), .ZN(
        n18336) );
  OAI21_X1 U21336 ( .B1(n18330), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18336), .ZN(n18331) );
  OAI211_X1 U21337 ( .C1(n18332), .C2(n18331), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18384), .ZN(n18333) );
  OAI211_X1 U21338 ( .C1(n18335), .C2(n18352), .A(n18334), .B(n18333), .ZN(
        P3_U2851) );
  AOI221_X1 U21339 ( .B1(n18337), .B2(n18336), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18336), .A(n18339), .ZN(
        n18338) );
  AOI22_X1 U21340 ( .A1(n18385), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18338), 
        .B2(n18384), .ZN(n18341) );
  NAND3_X1 U21341 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18344), .A3(
        n18339), .ZN(n18340) );
  OAI211_X1 U21342 ( .C1(n18342), .C2(n18352), .A(n18341), .B(n18340), .ZN(
        P3_U2852) );
  AOI22_X1 U21343 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n18385), .B1(n18344), 
        .B2(n18343), .ZN(n18351) );
  OAI21_X1 U21344 ( .B1(n18347), .B2(n18346), .A(n18345), .ZN(n18348) );
  OAI211_X1 U21345 ( .C1(n18349), .C2(n18348), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n18384), .ZN(n18350) );
  OAI211_X1 U21346 ( .C1(n18353), .C2(n18352), .A(n18351), .B(n18350), .ZN(
        P3_U2853) );
  OAI22_X1 U21347 ( .A1(n18356), .A2(n18924), .B1(n18355), .B2(n18354), .ZN(
        n18357) );
  OR3_X1 U21348 ( .A1(n18358), .A2(n18433), .A3(n18357), .ZN(n18383) );
  AOI21_X1 U21349 ( .B1(n18359), .B2(n18362), .A(n18383), .ZN(n18376) );
  NOR2_X1 U21350 ( .A1(n18376), .A2(n18360), .ZN(n18365) );
  NOR3_X1 U21351 ( .A1(n18361), .A2(n18433), .A3(n18412), .ZN(n18404) );
  NAND3_X1 U21352 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n18404), .ZN(n18387) );
  NOR3_X1 U21353 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18362), .A3(
        n18387), .ZN(n18364) );
  NOR2_X1 U21354 ( .A1(n18384), .A2(n19012), .ZN(n18363) );
  AOI211_X1 U21355 ( .C1(n18365), .C2(n18408), .A(n18364), .B(n18363), .ZN(
        n18370) );
  AOI22_X1 U21356 ( .A1(n18036), .A2(n18368), .B1(n18367), .B2(n18366), .ZN(
        n18369) );
  OAI211_X1 U21357 ( .C1(n18457), .C2(n18371), .A(n18370), .B(n18369), .ZN(
        P3_U2854) );
  NAND2_X1 U21358 ( .A1(n18372), .A2(n18451), .ZN(n18455) );
  AOI21_X1 U21359 ( .B1(n18374), .B2(n18441), .A(n18373), .ZN(n18381) );
  INV_X1 U21360 ( .A(n18375), .ZN(n18377) );
  AOI221_X1 U21361 ( .B1(n21195), .B2(n18378), .C1(n18377), .C2(n18378), .A(
        n18376), .ZN(n18379) );
  OAI211_X1 U21362 ( .C1(n18451), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18384), .B(n18379), .ZN(n18380) );
  OAI211_X1 U21363 ( .C1(n18382), .C2(n18457), .A(n18381), .B(n18380), .ZN(
        P3_U2855) );
  NAND2_X1 U21364 ( .A1(n18384), .A2(n18383), .ZN(n18393) );
  NAND2_X1 U21365 ( .A1(n18385), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18386) );
  OAI221_X1 U21366 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18387), .C1(
        n21195), .C2(n18393), .A(n18386), .ZN(n18388) );
  AOI21_X1 U21367 ( .B1(n18441), .B2(n18389), .A(n18388), .ZN(n18390) );
  OAI21_X1 U21368 ( .B1(n18457), .B2(n18391), .A(n18390), .ZN(P3_U2856) );
  INV_X1 U21369 ( .A(n18404), .ZN(n18392) );
  NOR2_X1 U21370 ( .A1(n18403), .A2(n18392), .ZN(n18395) );
  INV_X1 U21371 ( .A(n18393), .ZN(n18394) );
  MUX2_X1 U21372 ( .A(n18395), .B(n18394), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18396) );
  AOI21_X1 U21373 ( .B1(n18441), .B2(n18397), .A(n18396), .ZN(n18399) );
  OAI211_X1 U21374 ( .C1(n18457), .C2(n18400), .A(n18399), .B(n18398), .ZN(
        P3_U2857) );
  AOI21_X1 U21375 ( .B1(n18443), .B2(n18402), .A(n18401), .ZN(n18411) );
  AOI22_X1 U21376 ( .A1(n18405), .A2(n18441), .B1(n18404), .B2(n18403), .ZN(
        n18410) );
  AOI22_X1 U21377 ( .A1(n18933), .A2(n18428), .B1(n18406), .B2(n18421), .ZN(
        n18407) );
  NAND3_X1 U21378 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18407), .A3(
        n18423), .ZN(n18416) );
  OAI211_X1 U21379 ( .C1(n18445), .C2(n18416), .A(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n18408), .ZN(n18409) );
  NAND3_X1 U21380 ( .A1(n18411), .A2(n18410), .A3(n18409), .ZN(P3_U2858) );
  NOR2_X1 U21381 ( .A1(n18412), .A2(n18439), .ZN(n18413) );
  AOI211_X1 U21382 ( .C1(n18441), .C2(n18415), .A(n18414), .B(n18413), .ZN(
        n18419) );
  OAI211_X1 U21383 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18417), .A(
        n18451), .B(n18416), .ZN(n18418) );
  OAI211_X1 U21384 ( .C1(n18420), .C2(n18457), .A(n18419), .B(n18418), .ZN(
        P3_U2859) );
  NOR2_X1 U21385 ( .A1(n19073), .A2(n19091), .ZN(n18422) );
  AOI22_X1 U21386 ( .A1(n18933), .A2(n18422), .B1(n19073), .B2(n18421), .ZN(
        n18424) );
  AOI21_X1 U21387 ( .B1(n18424), .B2(n18423), .A(n12274), .ZN(n18427) );
  NOR3_X1 U21388 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19073), .A3(
        n18425), .ZN(n18426) );
  AOI211_X1 U21389 ( .C1(n18428), .C2(n18933), .A(n18427), .B(n18426), .ZN(
        n18434) );
  OAI21_X1 U21390 ( .B1(n18431), .B2(n18430), .A(n18429), .ZN(n18432) );
  OAI22_X1 U21391 ( .A1(n18434), .A2(n18433), .B1(n18457), .B2(n18432), .ZN(
        n18435) );
  AOI21_X1 U21392 ( .B1(n18441), .B2(n18436), .A(n18435), .ZN(n18438) );
  OAI211_X1 U21393 ( .C1(n18439), .C2(n12274), .A(n18438), .B(n18437), .ZN(
        P3_U2860) );
  AOI22_X1 U21394 ( .A1(n18443), .A2(n18442), .B1(n18441), .B2(n18440), .ZN(
        n18450) );
  NAND2_X1 U21395 ( .A1(n18385), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18449) );
  AND3_X1 U21396 ( .A1(n19091), .A2(n18444), .A3(n18451), .ZN(n18452) );
  OAI21_X1 U21397 ( .B1(n18445), .B2(n18452), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18448) );
  OAI211_X1 U21398 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18921), .A(
        n18446), .B(n19073), .ZN(n18447) );
  NAND4_X1 U21399 ( .A1(n18450), .A2(n18449), .A3(n18448), .A4(n18447), .ZN(
        P3_U2861) );
  AOI21_X1 U21400 ( .B1(n18937), .B2(n18451), .A(n19091), .ZN(n18453) );
  AOI221_X1 U21401 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n18385), .C1(n18453), 
        .C2(n18384), .A(n18452), .ZN(n18454) );
  OAI221_X1 U21402 ( .B1(n18458), .B2(n18457), .C1(n18456), .C2(n18455), .A(
        n18454), .ZN(P3_U2862) );
  AOI211_X1 U21403 ( .C1(n18460), .C2(n18459), .A(n19123), .B(n19075), .ZN(
        n18961) );
  OAI21_X1 U21404 ( .B1(n18961), .B2(n18524), .A(n18470), .ZN(n18461) );
  OAI221_X1 U21405 ( .B1(n18940), .B2(n19106), .C1(n18940), .C2(n18470), .A(
        n18461), .ZN(P3_U2863) );
  AOI221_X1 U21406 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18942), .C1(n18463), 
        .C2(n18942), .A(n18462), .ZN(n18469) );
  NOR2_X1 U21407 ( .A1(n18464), .A2(n18942), .ZN(n18466) );
  OAI21_X1 U21408 ( .B1(n18466), .B2(n18465), .A(n18470), .ZN(n18467) );
  AOI22_X1 U21409 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18469), .B1(
        n18467), .B2(n18947), .ZN(P3_U2865) );
  INV_X1 U21410 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18950) );
  NAND2_X1 U21411 ( .A1(n18950), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18641) );
  INV_X1 U21412 ( .A(n18641), .ZN(n18665) );
  NAND2_X1 U21413 ( .A1(n18947), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18733) );
  INV_X1 U21414 ( .A(n18733), .ZN(n18710) );
  NOR2_X1 U21415 ( .A1(n18665), .A2(n18710), .ZN(n18468) );
  OAI22_X1 U21416 ( .A1(n18469), .A2(n18950), .B1(n18468), .B2(n18467), .ZN(
        P3_U2866) );
  NOR2_X1 U21417 ( .A1(n18951), .A2(n18470), .ZN(P3_U2867) );
  NOR3_X1 U21418 ( .A1(n18947), .A2(n18950), .A3(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18853) );
  NAND2_X1 U21419 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18853), .ZN(
        n18821) );
  INV_X1 U21420 ( .A(n18821), .ZN(n18898) );
  NOR3_X1 U21421 ( .A1(n18942), .A2(n18947), .A3(n18950), .ZN(n18852) );
  NAND2_X1 U21422 ( .A1(n18940), .A2(n18852), .ZN(n18847) );
  NOR2_X1 U21423 ( .A1(n18898), .A2(n18827), .ZN(n18822) );
  NAND2_X1 U21424 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18852), .ZN(
        n18905) );
  INV_X1 U21425 ( .A(n18905), .ZN(n18569) );
  NAND2_X1 U21426 ( .A1(n18942), .A2(n18940), .ZN(n18943) );
  NOR2_X1 U21427 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18576) );
  INV_X1 U21428 ( .A(n18576), .ZN(n18550) );
  NOR2_X1 U21429 ( .A1(n18943), .A2(n18550), .ZN(n18570) );
  CLKBUF_X1 U21430 ( .A(n18570), .Z(n18592) );
  NOR2_X1 U21431 ( .A1(n18569), .A2(n18592), .ZN(n18552) );
  INV_X1 U21432 ( .A(n18597), .ZN(n18826) );
  OAI21_X1 U21433 ( .B1(n18940), .B2(n19068), .A(n18826), .ZN(n18687) );
  OAI22_X1 U21434 ( .A1(n18822), .A2(n18507), .B1(n18552), .B2(n18687), .ZN(
        n18521) );
  AND2_X1 U21435 ( .A1(n18854), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18850) );
  NOR2_X2 U21436 ( .A1(n18597), .A2(n18471), .ZN(n18849) );
  NOR2_X1 U21437 ( .A1(n18971), .A2(n18552), .ZN(n18515) );
  AOI22_X1 U21438 ( .A1(n18827), .A2(n18850), .B1(n18849), .B2(n18515), .ZN(
        n18477) );
  INV_X1 U21439 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18472) );
  NOR2_X2 U21440 ( .A1(n18472), .A2(n18507), .ZN(n18855) );
  NAND2_X1 U21441 ( .A1(n18474), .A2(n18473), .ZN(n18517) );
  NOR2_X1 U21442 ( .A1(n18475), .A2(n18517), .ZN(n18523) );
  AOI22_X1 U21443 ( .A1(n18898), .A2(n18855), .B1(n18570), .B2(n18523), .ZN(
        n18476) );
  OAI211_X1 U21444 ( .C1(n18478), .C2(n18521), .A(n18477), .B(n18476), .ZN(
        P3_U2868) );
  INV_X1 U21445 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18479) );
  NOR2_X2 U21446 ( .A1(n18479), .A2(n18507), .ZN(n18859) );
  AND2_X1 U21447 ( .A1(n18826), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18860) );
  AOI22_X1 U21448 ( .A1(n18898), .A2(n18859), .B1(n18515), .B2(n18860), .ZN(
        n18481) );
  AND2_X1 U21449 ( .A1(n18854), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18861) );
  NOR2_X1 U21450 ( .A1(n19112), .A2(n18517), .ZN(n18527) );
  AOI22_X1 U21451 ( .A1(n18827), .A2(n18861), .B1(n18592), .B2(n18527), .ZN(
        n18480) );
  OAI211_X1 U21452 ( .C1(n18482), .C2(n18521), .A(n18481), .B(n18480), .ZN(
        P3_U2869) );
  AND2_X1 U21453 ( .A1(n18854), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18867) );
  NOR2_X2 U21454 ( .A1(n18597), .A2(n18483), .ZN(n18865) );
  AOI22_X1 U21455 ( .A1(n18827), .A2(n18867), .B1(n18515), .B2(n18865), .ZN(
        n18487) );
  INV_X1 U21456 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18484) );
  NOR2_X2 U21457 ( .A1(n18484), .A2(n18507), .ZN(n18866) );
  NOR2_X1 U21458 ( .A1(n18485), .A2(n18517), .ZN(n18530) );
  AOI22_X1 U21459 ( .A1(n18898), .A2(n18866), .B1(n18570), .B2(n18530), .ZN(
        n18486) );
  OAI211_X1 U21460 ( .C1(n18488), .C2(n18521), .A(n18487), .B(n18486), .ZN(
        P3_U2870) );
  NOR2_X2 U21461 ( .A1(n18507), .A2(n19543), .ZN(n18872) );
  NOR2_X2 U21462 ( .A1(n18597), .A2(n18489), .ZN(n18871) );
  AOI22_X1 U21463 ( .A1(n18827), .A2(n18872), .B1(n18515), .B2(n18871), .ZN(
        n18493) );
  INV_X1 U21464 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18490) );
  NOR2_X2 U21465 ( .A1(n18490), .A2(n18507), .ZN(n18873) );
  NOR2_X1 U21466 ( .A1(n18491), .A2(n18517), .ZN(n18533) );
  AOI22_X1 U21467 ( .A1(n18898), .A2(n18873), .B1(n18570), .B2(n18533), .ZN(
        n18492) );
  OAI211_X1 U21468 ( .C1(n18494), .C2(n18521), .A(n18493), .B(n18492), .ZN(
        P3_U2871) );
  AND2_X1 U21469 ( .A1(n18854), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18878) );
  NOR2_X2 U21470 ( .A1(n18597), .A2(n18495), .ZN(n18877) );
  AOI22_X1 U21471 ( .A1(n18827), .A2(n18878), .B1(n18515), .B2(n18877), .ZN(
        n18499) );
  NOR2_X2 U21472 ( .A1(n18496), .A2(n18507), .ZN(n18879) );
  NOR2_X1 U21473 ( .A1(n18497), .A2(n18517), .ZN(n18536) );
  AOI22_X1 U21474 ( .A1(n18898), .A2(n18879), .B1(n18570), .B2(n18536), .ZN(
        n18498) );
  OAI211_X1 U21475 ( .C1(n18500), .C2(n18521), .A(n18499), .B(n18498), .ZN(
        P3_U2872) );
  AND2_X1 U21476 ( .A1(n18854), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18884) );
  NOR2_X2 U21477 ( .A1(n18597), .A2(n18501), .ZN(n18883) );
  AOI22_X1 U21478 ( .A1(n18827), .A2(n18884), .B1(n18515), .B2(n18883), .ZN(
        n18505) );
  INV_X1 U21479 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18502) );
  NOR2_X2 U21480 ( .A1(n18502), .A2(n18507), .ZN(n18885) );
  NOR2_X1 U21481 ( .A1(n18503), .A2(n18517), .ZN(n18539) );
  AOI22_X1 U21482 ( .A1(n18898), .A2(n18885), .B1(n18570), .B2(n18539), .ZN(
        n18504) );
  OAI211_X1 U21483 ( .C1(n18506), .C2(n18521), .A(n18505), .B(n18504), .ZN(
        P3_U2873) );
  NOR2_X2 U21484 ( .A1(n18508), .A2(n18507), .ZN(n18891) );
  NOR2_X2 U21485 ( .A1(n18597), .A2(n18509), .ZN(n18889) );
  AOI22_X1 U21486 ( .A1(n18898), .A2(n18891), .B1(n18515), .B2(n18889), .ZN(
        n18512) );
  NOR2_X2 U21487 ( .A1(n18507), .A2(n19557), .ZN(n18890) );
  NOR2_X1 U21488 ( .A1(n18510), .A2(n18517), .ZN(n18542) );
  AOI22_X1 U21489 ( .A1(n18827), .A2(n18890), .B1(n18570), .B2(n18542), .ZN(
        n18511) );
  OAI211_X1 U21490 ( .C1(n18513), .C2(n18521), .A(n18512), .B(n18511), .ZN(
        P3_U2874) );
  AND2_X1 U21491 ( .A1(n18854), .A2(BUF2_REG_23__SCAN_IN), .ZN(n18897) );
  NOR2_X2 U21492 ( .A1(n18597), .A2(n18514), .ZN(n18896) );
  AOI22_X1 U21493 ( .A1(n18827), .A2(n18897), .B1(n18515), .B2(n18896), .ZN(
        n18520) );
  NOR2_X2 U21494 ( .A1(n18507), .A2(n18516), .ZN(n18900) );
  NOR2_X1 U21495 ( .A1(n18518), .A2(n18517), .ZN(n18545) );
  AOI22_X1 U21496 ( .A1(n18898), .A2(n18900), .B1(n18570), .B2(n18545), .ZN(
        n18519) );
  OAI211_X1 U21497 ( .C1(n18522), .C2(n18521), .A(n18520), .B(n18519), .ZN(
        P3_U2875) );
  NOR2_X1 U21498 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18940), .ZN(
        n18711) );
  NAND2_X1 U21499 ( .A1(n18576), .A2(n18711), .ZN(n18551) );
  NAND2_X1 U21500 ( .A1(n18942), .A2(n18964), .ZN(n18712) );
  NOR2_X1 U21501 ( .A1(n18550), .A2(n18712), .ZN(n18546) );
  AOI22_X1 U21502 ( .A1(n18827), .A2(n18855), .B1(n18849), .B2(n18546), .ZN(
        n18526) );
  NOR2_X1 U21503 ( .A1(n18597), .A2(n18524), .ZN(n18851) );
  INV_X1 U21504 ( .A(n18851), .ZN(n18575) );
  NOR2_X1 U21505 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18575), .ZN(
        n18620) );
  AOI22_X1 U21506 ( .A1(n18854), .A2(n18852), .B1(n18576), .B2(n18620), .ZN(
        n18547) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18547), .B1(
        n18569), .B2(n18850), .ZN(n18525) );
  OAI211_X1 U21508 ( .C1(n18858), .C2(n18551), .A(n18526), .B(n18525), .ZN(
        P3_U2876) );
  INV_X1 U21509 ( .A(n18527), .ZN(n18864) );
  AOI22_X1 U21510 ( .A1(n18569), .A2(n18861), .B1(n18860), .B2(n18546), .ZN(
        n18529) );
  AOI22_X1 U21511 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18547), .B1(
        n18827), .B2(n18859), .ZN(n18528) );
  OAI211_X1 U21512 ( .C1(n18864), .C2(n18551), .A(n18529), .B(n18528), .ZN(
        P3_U2877) );
  INV_X1 U21513 ( .A(n18530), .ZN(n18870) );
  AOI22_X1 U21514 ( .A1(n18569), .A2(n18867), .B1(n18865), .B2(n18546), .ZN(
        n18532) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18547), .B1(
        n18827), .B2(n18866), .ZN(n18531) );
  OAI211_X1 U21516 ( .C1(n18870), .C2(n18551), .A(n18532), .B(n18531), .ZN(
        P3_U2878) );
  INV_X1 U21517 ( .A(n18533), .ZN(n18876) );
  AOI22_X1 U21518 ( .A1(n18827), .A2(n18873), .B1(n18871), .B2(n18546), .ZN(
        n18535) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18547), .B1(
        n18569), .B2(n18872), .ZN(n18534) );
  OAI211_X1 U21520 ( .C1(n18876), .C2(n18551), .A(n18535), .B(n18534), .ZN(
        P3_U2879) );
  INV_X1 U21521 ( .A(n18536), .ZN(n18882) );
  AOI22_X1 U21522 ( .A1(n18827), .A2(n18879), .B1(n18877), .B2(n18546), .ZN(
        n18538) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18547), .B1(
        n18569), .B2(n18878), .ZN(n18537) );
  OAI211_X1 U21524 ( .C1(n18882), .C2(n18551), .A(n18538), .B(n18537), .ZN(
        P3_U2880) );
  AOI22_X1 U21525 ( .A1(n18569), .A2(n18884), .B1(n18883), .B2(n18546), .ZN(
        n18541) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18547), .B1(
        n18827), .B2(n18885), .ZN(n18540) );
  OAI211_X1 U21527 ( .C1(n18888), .C2(n18551), .A(n18541), .B(n18540), .ZN(
        P3_U2881) );
  INV_X1 U21528 ( .A(n18542), .ZN(n18894) );
  AOI22_X1 U21529 ( .A1(n18827), .A2(n18891), .B1(n18889), .B2(n18546), .ZN(
        n18544) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18547), .B1(
        n18569), .B2(n18890), .ZN(n18543) );
  OAI211_X1 U21531 ( .C1(n18894), .C2(n18551), .A(n18544), .B(n18543), .ZN(
        P3_U2882) );
  INV_X1 U21532 ( .A(n18545), .ZN(n18904) );
  AOI22_X1 U21533 ( .A1(n18827), .A2(n18900), .B1(n18896), .B2(n18546), .ZN(
        n18549) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18547), .B1(
        n18569), .B2(n18897), .ZN(n18548) );
  OAI211_X1 U21535 ( .C1(n18904), .C2(n18551), .A(n18549), .B(n18548), .ZN(
        P3_U2883) );
  NOR2_X1 U21536 ( .A1(n18942), .A2(n18550), .ZN(n18621) );
  NAND2_X1 U21537 ( .A1(n18621), .A2(n18940), .ZN(n18574) );
  INV_X1 U21538 ( .A(n18551), .ZN(n18615) );
  NOR2_X1 U21539 ( .A1(n18615), .A2(n18637), .ZN(n18598) );
  NOR2_X1 U21540 ( .A1(n18971), .A2(n18598), .ZN(n18568) );
  AOI22_X1 U21541 ( .A1(n18569), .A2(n18855), .B1(n18849), .B2(n18568), .ZN(
        n18555) );
  AOI221_X1 U21542 ( .B1(n18598), .B2(n18823), .C1(n18598), .C2(n18552), .A(
        n18687), .ZN(n18553) );
  INV_X1 U21543 ( .A(n18553), .ZN(n18571) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18571), .B1(
        n18570), .B2(n18850), .ZN(n18554) );
  OAI211_X1 U21545 ( .C1(n18858), .C2(n18574), .A(n18555), .B(n18554), .ZN(
        P3_U2884) );
  AOI22_X1 U21546 ( .A1(n18569), .A2(n18859), .B1(n18860), .B2(n18568), .ZN(
        n18557) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18571), .B1(
        n18570), .B2(n18861), .ZN(n18556) );
  OAI211_X1 U21548 ( .C1(n18864), .C2(n18574), .A(n18557), .B(n18556), .ZN(
        P3_U2885) );
  AOI22_X1 U21549 ( .A1(n18569), .A2(n18866), .B1(n18865), .B2(n18568), .ZN(
        n18559) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18571), .B1(
        n18570), .B2(n18867), .ZN(n18558) );
  OAI211_X1 U21551 ( .C1(n18870), .C2(n18574), .A(n18559), .B(n18558), .ZN(
        P3_U2886) );
  AOI22_X1 U21552 ( .A1(n18592), .A2(n18872), .B1(n18871), .B2(n18568), .ZN(
        n18561) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18571), .B1(
        n18569), .B2(n18873), .ZN(n18560) );
  OAI211_X1 U21554 ( .C1(n18876), .C2(n18574), .A(n18561), .B(n18560), .ZN(
        P3_U2887) );
  AOI22_X1 U21555 ( .A1(n18592), .A2(n18878), .B1(n18877), .B2(n18568), .ZN(
        n18563) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18571), .B1(
        n18569), .B2(n18879), .ZN(n18562) );
  OAI211_X1 U21557 ( .C1(n18882), .C2(n18574), .A(n18563), .B(n18562), .ZN(
        P3_U2888) );
  AOI22_X1 U21558 ( .A1(n18592), .A2(n18884), .B1(n18883), .B2(n18568), .ZN(
        n18565) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18571), .B1(
        n18569), .B2(n18885), .ZN(n18564) );
  OAI211_X1 U21560 ( .C1(n18888), .C2(n18574), .A(n18565), .B(n18564), .ZN(
        P3_U2889) );
  AOI22_X1 U21561 ( .A1(n18592), .A2(n18890), .B1(n18889), .B2(n18568), .ZN(
        n18567) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18571), .B1(
        n18569), .B2(n18891), .ZN(n18566) );
  OAI211_X1 U21563 ( .C1(n18894), .C2(n18574), .A(n18567), .B(n18566), .ZN(
        P3_U2890) );
  AOI22_X1 U21564 ( .A1(n18569), .A2(n18900), .B1(n18896), .B2(n18568), .ZN(
        n18573) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18571), .B1(
        n18570), .B2(n18897), .ZN(n18572) );
  OAI211_X1 U21566 ( .C1(n18904), .C2(n18574), .A(n18573), .B(n18572), .ZN(
        P3_U2891) );
  NAND2_X1 U21567 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18621), .ZN(
        n18596) );
  AND2_X1 U21568 ( .A1(n18964), .A2(n18621), .ZN(n18591) );
  AOI22_X1 U21569 ( .A1(n18592), .A2(n18855), .B1(n18849), .B2(n18591), .ZN(
        n18578) );
  AOI21_X1 U21570 ( .B1(n18942), .B2(n18823), .A(n18575), .ZN(n18666) );
  NAND2_X1 U21571 ( .A1(n18576), .A2(n18666), .ZN(n18593) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18593), .B1(
        n18850), .B2(n18615), .ZN(n18577) );
  OAI211_X1 U21573 ( .C1(n18858), .C2(n18596), .A(n18578), .B(n18577), .ZN(
        P3_U2892) );
  AOI22_X1 U21574 ( .A1(n18861), .A2(n18615), .B1(n18860), .B2(n18591), .ZN(
        n18580) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18593), .B1(
        n18592), .B2(n18859), .ZN(n18579) );
  OAI211_X1 U21576 ( .C1(n18864), .C2(n18596), .A(n18580), .B(n18579), .ZN(
        P3_U2893) );
  AOI22_X1 U21577 ( .A1(n18592), .A2(n18866), .B1(n18865), .B2(n18591), .ZN(
        n18582) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18593), .B1(
        n18867), .B2(n18615), .ZN(n18581) );
  OAI211_X1 U21579 ( .C1(n18870), .C2(n18596), .A(n18582), .B(n18581), .ZN(
        P3_U2894) );
  AOI22_X1 U21580 ( .A1(n18592), .A2(n18873), .B1(n18871), .B2(n18591), .ZN(
        n18584) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18593), .B1(
        n18872), .B2(n18615), .ZN(n18583) );
  OAI211_X1 U21582 ( .C1(n18876), .C2(n18596), .A(n18584), .B(n18583), .ZN(
        P3_U2895) );
  AOI22_X1 U21583 ( .A1(n18878), .A2(n18615), .B1(n18877), .B2(n18591), .ZN(
        n18586) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18593), .B1(
        n18592), .B2(n18879), .ZN(n18585) );
  OAI211_X1 U21585 ( .C1(n18882), .C2(n18596), .A(n18586), .B(n18585), .ZN(
        P3_U2896) );
  AOI22_X1 U21586 ( .A1(n18592), .A2(n18885), .B1(n18883), .B2(n18591), .ZN(
        n18588) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18593), .B1(
        n18884), .B2(n18615), .ZN(n18587) );
  OAI211_X1 U21588 ( .C1(n18888), .C2(n18596), .A(n18588), .B(n18587), .ZN(
        P3_U2897) );
  AOI22_X1 U21589 ( .A1(n18890), .A2(n18615), .B1(n18889), .B2(n18591), .ZN(
        n18590) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18593), .B1(
        n18592), .B2(n18891), .ZN(n18589) );
  OAI211_X1 U21591 ( .C1(n18894), .C2(n18596), .A(n18590), .B(n18589), .ZN(
        P3_U2898) );
  AOI22_X1 U21592 ( .A1(n18592), .A2(n18900), .B1(n18896), .B2(n18591), .ZN(
        n18595) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18593), .B1(
        n18897), .B2(n18615), .ZN(n18594) );
  OAI211_X1 U21594 ( .C1(n18904), .C2(n18596), .A(n18595), .B(n18594), .ZN(
        P3_U2899) );
  NOR2_X2 U21595 ( .A1(n18943), .A2(n18641), .ZN(n18682) );
  INV_X1 U21596 ( .A(n18682), .ZN(n18619) );
  INV_X1 U21597 ( .A(n18596), .ZN(n18660) );
  NOR2_X1 U21598 ( .A1(n18660), .A2(n18682), .ZN(n18643) );
  NOR2_X1 U21599 ( .A1(n18971), .A2(n18643), .ZN(n18614) );
  AOI22_X1 U21600 ( .A1(n18855), .A2(n18615), .B1(n18849), .B2(n18614), .ZN(
        n18601) );
  OAI22_X1 U21601 ( .A1(n18598), .A2(n18507), .B1(n18643), .B2(n18597), .ZN(
        n18599) );
  OAI21_X1 U21602 ( .B1(n18682), .B2(n19068), .A(n18599), .ZN(n18616) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18616), .B1(
        n18850), .B2(n18637), .ZN(n18600) );
  OAI211_X1 U21604 ( .C1(n18858), .C2(n18619), .A(n18601), .B(n18600), .ZN(
        P3_U2900) );
  AOI22_X1 U21605 ( .A1(n18861), .A2(n18637), .B1(n18860), .B2(n18614), .ZN(
        n18603) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18616), .B1(
        n18859), .B2(n18615), .ZN(n18602) );
  OAI211_X1 U21607 ( .C1(n18864), .C2(n18619), .A(n18603), .B(n18602), .ZN(
        P3_U2901) );
  AOI22_X1 U21608 ( .A1(n18867), .A2(n18637), .B1(n18865), .B2(n18614), .ZN(
        n18605) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18616), .B1(
        n18866), .B2(n18615), .ZN(n18604) );
  OAI211_X1 U21610 ( .C1(n18870), .C2(n18619), .A(n18605), .B(n18604), .ZN(
        P3_U2902) );
  AOI22_X1 U21611 ( .A1(n18873), .A2(n18615), .B1(n18871), .B2(n18614), .ZN(
        n18607) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18616), .B1(
        n18872), .B2(n18637), .ZN(n18606) );
  OAI211_X1 U21613 ( .C1(n18876), .C2(n18619), .A(n18607), .B(n18606), .ZN(
        P3_U2903) );
  AOI22_X1 U21614 ( .A1(n18879), .A2(n18615), .B1(n18877), .B2(n18614), .ZN(
        n18609) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18616), .B1(
        n18878), .B2(n18637), .ZN(n18608) );
  OAI211_X1 U21616 ( .C1(n18882), .C2(n18619), .A(n18609), .B(n18608), .ZN(
        P3_U2904) );
  AOI22_X1 U21617 ( .A1(n18885), .A2(n18615), .B1(n18883), .B2(n18614), .ZN(
        n18611) );
  AOI22_X1 U21618 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18616), .B1(
        n18884), .B2(n18637), .ZN(n18610) );
  OAI211_X1 U21619 ( .C1(n18888), .C2(n18619), .A(n18611), .B(n18610), .ZN(
        P3_U2905) );
  AOI22_X1 U21620 ( .A1(n18890), .A2(n18637), .B1(n18889), .B2(n18614), .ZN(
        n18613) );
  AOI22_X1 U21621 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18616), .B1(
        n18891), .B2(n18615), .ZN(n18612) );
  OAI211_X1 U21622 ( .C1(n18894), .C2(n18619), .A(n18613), .B(n18612), .ZN(
        P3_U2906) );
  AOI22_X1 U21623 ( .A1(n18900), .A2(n18615), .B1(n18896), .B2(n18614), .ZN(
        n18618) );
  AOI22_X1 U21624 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18616), .B1(
        n18897), .B2(n18637), .ZN(n18617) );
  OAI211_X1 U21625 ( .C1(n18904), .C2(n18619), .A(n18618), .B(n18617), .ZN(
        P3_U2907) );
  NAND2_X1 U21626 ( .A1(n18711), .A2(n18665), .ZN(n18642) );
  NOR2_X1 U21627 ( .A1(n18712), .A2(n18641), .ZN(n18636) );
  AOI22_X1 U21628 ( .A1(n18850), .A2(n18660), .B1(n18849), .B2(n18636), .ZN(
        n18623) );
  AOI22_X1 U21629 ( .A1(n18854), .A2(n18621), .B1(n18620), .B2(n18665), .ZN(
        n18638) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18638), .B1(
        n18855), .B2(n18637), .ZN(n18622) );
  OAI211_X1 U21631 ( .C1(n18858), .C2(n18642), .A(n18623), .B(n18622), .ZN(
        P3_U2908) );
  AOI22_X1 U21632 ( .A1(n18860), .A2(n18636), .B1(n18859), .B2(n18637), .ZN(
        n18625) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18638), .B1(
        n18861), .B2(n18660), .ZN(n18624) );
  OAI211_X1 U21634 ( .C1(n18864), .C2(n18642), .A(n18625), .B(n18624), .ZN(
        P3_U2909) );
  AOI22_X1 U21635 ( .A1(n18866), .A2(n18637), .B1(n18865), .B2(n18636), .ZN(
        n18627) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18638), .B1(
        n18867), .B2(n18660), .ZN(n18626) );
  OAI211_X1 U21637 ( .C1(n18870), .C2(n18642), .A(n18627), .B(n18626), .ZN(
        P3_U2910) );
  AOI22_X1 U21638 ( .A1(n18872), .A2(n18660), .B1(n18871), .B2(n18636), .ZN(
        n18629) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18638), .B1(
        n18873), .B2(n18637), .ZN(n18628) );
  OAI211_X1 U21640 ( .C1(n18876), .C2(n18642), .A(n18629), .B(n18628), .ZN(
        P3_U2911) );
  AOI22_X1 U21641 ( .A1(n18879), .A2(n18637), .B1(n18877), .B2(n18636), .ZN(
        n18631) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18638), .B1(
        n18878), .B2(n18660), .ZN(n18630) );
  OAI211_X1 U21643 ( .C1(n18882), .C2(n18642), .A(n18631), .B(n18630), .ZN(
        P3_U2912) );
  AOI22_X1 U21644 ( .A1(n18884), .A2(n18660), .B1(n18883), .B2(n18636), .ZN(
        n18633) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18638), .B1(
        n18885), .B2(n18637), .ZN(n18632) );
  OAI211_X1 U21646 ( .C1(n18888), .C2(n18642), .A(n18633), .B(n18632), .ZN(
        P3_U2913) );
  AOI22_X1 U21647 ( .A1(n18890), .A2(n18660), .B1(n18889), .B2(n18636), .ZN(
        n18635) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18638), .B1(
        n18891), .B2(n18637), .ZN(n18634) );
  OAI211_X1 U21649 ( .C1(n18894), .C2(n18642), .A(n18635), .B(n18634), .ZN(
        P3_U2914) );
  AOI22_X1 U21650 ( .A1(n18897), .A2(n18660), .B1(n18896), .B2(n18636), .ZN(
        n18640) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18638), .B1(
        n18900), .B2(n18637), .ZN(n18639) );
  OAI211_X1 U21652 ( .C1(n18904), .C2(n18642), .A(n18640), .B(n18639), .ZN(
        P3_U2915) );
  NOR2_X1 U21653 ( .A1(n18942), .A2(n18641), .ZN(n18713) );
  NAND2_X1 U21654 ( .A1(n18713), .A2(n18940), .ZN(n18664) );
  INV_X1 U21655 ( .A(n18642), .ZN(n18705) );
  NOR2_X1 U21656 ( .A1(n18705), .A2(n18729), .ZN(n18688) );
  NOR2_X1 U21657 ( .A1(n18971), .A2(n18688), .ZN(n18659) );
  AOI22_X1 U21658 ( .A1(n18855), .A2(n18660), .B1(n18849), .B2(n18659), .ZN(
        n18646) );
  OAI21_X1 U21659 ( .B1(n18643), .B2(n18823), .A(n18688), .ZN(n18644) );
  OAI211_X1 U21660 ( .C1(n18729), .C2(n19068), .A(n18826), .B(n18644), .ZN(
        n18661) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18661), .B1(
        n18850), .B2(n18682), .ZN(n18645) );
  OAI211_X1 U21662 ( .C1(n18858), .C2(n18664), .A(n18646), .B(n18645), .ZN(
        P3_U2916) );
  AOI22_X1 U21663 ( .A1(n18861), .A2(n18682), .B1(n18860), .B2(n18659), .ZN(
        n18648) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18661), .B1(
        n18859), .B2(n18660), .ZN(n18647) );
  OAI211_X1 U21665 ( .C1(n18864), .C2(n18664), .A(n18648), .B(n18647), .ZN(
        P3_U2917) );
  AOI22_X1 U21666 ( .A1(n18866), .A2(n18660), .B1(n18865), .B2(n18659), .ZN(
        n18650) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18661), .B1(
        n18867), .B2(n18682), .ZN(n18649) );
  OAI211_X1 U21668 ( .C1(n18870), .C2(n18664), .A(n18650), .B(n18649), .ZN(
        P3_U2918) );
  AOI22_X1 U21669 ( .A1(n18872), .A2(n18682), .B1(n18871), .B2(n18659), .ZN(
        n18652) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18661), .B1(
        n18873), .B2(n18660), .ZN(n18651) );
  OAI211_X1 U21671 ( .C1(n18876), .C2(n18664), .A(n18652), .B(n18651), .ZN(
        P3_U2919) );
  AOI22_X1 U21672 ( .A1(n18879), .A2(n18660), .B1(n18877), .B2(n18659), .ZN(
        n18654) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18661), .B1(
        n18878), .B2(n18682), .ZN(n18653) );
  OAI211_X1 U21674 ( .C1(n18882), .C2(n18664), .A(n18654), .B(n18653), .ZN(
        P3_U2920) );
  AOI22_X1 U21675 ( .A1(n18885), .A2(n18660), .B1(n18883), .B2(n18659), .ZN(
        n18656) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18661), .B1(
        n18884), .B2(n18682), .ZN(n18655) );
  OAI211_X1 U21677 ( .C1(n18888), .C2(n18664), .A(n18656), .B(n18655), .ZN(
        P3_U2921) );
  AOI22_X1 U21678 ( .A1(n18890), .A2(n18682), .B1(n18889), .B2(n18659), .ZN(
        n18658) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18661), .B1(
        n18891), .B2(n18660), .ZN(n18657) );
  OAI211_X1 U21680 ( .C1(n18894), .C2(n18664), .A(n18658), .B(n18657), .ZN(
        P3_U2922) );
  AOI22_X1 U21681 ( .A1(n18900), .A2(n18660), .B1(n18896), .B2(n18659), .ZN(
        n18663) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18661), .B1(
        n18897), .B2(n18682), .ZN(n18662) );
  OAI211_X1 U21683 ( .C1(n18904), .C2(n18664), .A(n18663), .B(n18662), .ZN(
        P3_U2923) );
  NAND2_X1 U21684 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18713), .ZN(
        n18686) );
  AND2_X1 U21685 ( .A1(n18964), .A2(n18713), .ZN(n18681) );
  AOI22_X1 U21686 ( .A1(n18855), .A2(n18682), .B1(n18849), .B2(n18681), .ZN(
        n18668) );
  NAND2_X1 U21687 ( .A1(n18666), .A2(n18665), .ZN(n18683) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18683), .B1(
        n18850), .B2(n18705), .ZN(n18667) );
  OAI211_X1 U21689 ( .C1(n18858), .C2(n18686), .A(n18668), .B(n18667), .ZN(
        P3_U2924) );
  AOI22_X1 U21690 ( .A1(n18860), .A2(n18681), .B1(n18859), .B2(n18682), .ZN(
        n18670) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18683), .B1(
        n18861), .B2(n18705), .ZN(n18669) );
  OAI211_X1 U21692 ( .C1(n18864), .C2(n18686), .A(n18670), .B(n18669), .ZN(
        P3_U2925) );
  AOI22_X1 U21693 ( .A1(n18866), .A2(n18682), .B1(n18865), .B2(n18681), .ZN(
        n18672) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18683), .B1(
        n18867), .B2(n18705), .ZN(n18671) );
  OAI211_X1 U21695 ( .C1(n18870), .C2(n18686), .A(n18672), .B(n18671), .ZN(
        P3_U2926) );
  AOI22_X1 U21696 ( .A1(n18872), .A2(n18705), .B1(n18871), .B2(n18681), .ZN(
        n18674) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18683), .B1(
        n18873), .B2(n18682), .ZN(n18673) );
  OAI211_X1 U21698 ( .C1(n18876), .C2(n18686), .A(n18674), .B(n18673), .ZN(
        P3_U2927) );
  AOI22_X1 U21699 ( .A1(n18879), .A2(n18682), .B1(n18877), .B2(n18681), .ZN(
        n18676) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18683), .B1(
        n18878), .B2(n18705), .ZN(n18675) );
  OAI211_X1 U21701 ( .C1(n18882), .C2(n18686), .A(n18676), .B(n18675), .ZN(
        P3_U2928) );
  AOI22_X1 U21702 ( .A1(n18884), .A2(n18705), .B1(n18883), .B2(n18681), .ZN(
        n18678) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18683), .B1(
        n18885), .B2(n18682), .ZN(n18677) );
  OAI211_X1 U21704 ( .C1(n18888), .C2(n18686), .A(n18678), .B(n18677), .ZN(
        P3_U2929) );
  AOI22_X1 U21705 ( .A1(n18890), .A2(n18705), .B1(n18889), .B2(n18681), .ZN(
        n18680) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18683), .B1(
        n18891), .B2(n18682), .ZN(n18679) );
  OAI211_X1 U21707 ( .C1(n18894), .C2(n18686), .A(n18680), .B(n18679), .ZN(
        P3_U2930) );
  AOI22_X1 U21708 ( .A1(n18900), .A2(n18682), .B1(n18896), .B2(n18681), .ZN(
        n18685) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18683), .B1(
        n18897), .B2(n18705), .ZN(n18684) );
  OAI211_X1 U21710 ( .C1(n18904), .C2(n18686), .A(n18685), .B(n18684), .ZN(
        P3_U2931) );
  NOR2_X2 U21711 ( .A1(n18943), .A2(n18733), .ZN(n18773) );
  INV_X1 U21712 ( .A(n18773), .ZN(n18709) );
  INV_X1 U21713 ( .A(n18686), .ZN(n18752) );
  NOR2_X1 U21714 ( .A1(n18752), .A2(n18773), .ZN(n18735) );
  NOR2_X1 U21715 ( .A1(n18971), .A2(n18735), .ZN(n18704) );
  AOI22_X1 U21716 ( .A1(n18855), .A2(n18705), .B1(n18849), .B2(n18704), .ZN(
        n18691) );
  AOI221_X1 U21717 ( .B1(n18735), .B2(n18823), .C1(n18735), .C2(n18688), .A(
        n18687), .ZN(n18689) );
  INV_X1 U21718 ( .A(n18689), .ZN(n18706) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18706), .B1(
        n18850), .B2(n18729), .ZN(n18690) );
  OAI211_X1 U21720 ( .C1(n18858), .C2(n18709), .A(n18691), .B(n18690), .ZN(
        P3_U2932) );
  AOI22_X1 U21721 ( .A1(n18860), .A2(n18704), .B1(n18859), .B2(n18705), .ZN(
        n18693) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18706), .B1(
        n18861), .B2(n18729), .ZN(n18692) );
  OAI211_X1 U21723 ( .C1(n18864), .C2(n18709), .A(n18693), .B(n18692), .ZN(
        P3_U2933) );
  AOI22_X1 U21724 ( .A1(n18866), .A2(n18705), .B1(n18865), .B2(n18704), .ZN(
        n18695) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18706), .B1(
        n18867), .B2(n18729), .ZN(n18694) );
  OAI211_X1 U21726 ( .C1(n18870), .C2(n18709), .A(n18695), .B(n18694), .ZN(
        P3_U2934) );
  AOI22_X1 U21727 ( .A1(n18872), .A2(n18729), .B1(n18871), .B2(n18704), .ZN(
        n18697) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18706), .B1(
        n18873), .B2(n18705), .ZN(n18696) );
  OAI211_X1 U21729 ( .C1(n18876), .C2(n18709), .A(n18697), .B(n18696), .ZN(
        P3_U2935) );
  AOI22_X1 U21730 ( .A1(n18878), .A2(n18729), .B1(n18877), .B2(n18704), .ZN(
        n18699) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18706), .B1(
        n18879), .B2(n18705), .ZN(n18698) );
  OAI211_X1 U21732 ( .C1(n18882), .C2(n18709), .A(n18699), .B(n18698), .ZN(
        P3_U2936) );
  AOI22_X1 U21733 ( .A1(n18884), .A2(n18729), .B1(n18883), .B2(n18704), .ZN(
        n18701) );
  AOI22_X1 U21734 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18706), .B1(
        n18885), .B2(n18705), .ZN(n18700) );
  OAI211_X1 U21735 ( .C1(n18888), .C2(n18709), .A(n18701), .B(n18700), .ZN(
        P3_U2937) );
  AOI22_X1 U21736 ( .A1(n18889), .A2(n18704), .B1(n18891), .B2(n18705), .ZN(
        n18703) );
  AOI22_X1 U21737 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18706), .B1(
        n18890), .B2(n18729), .ZN(n18702) );
  OAI211_X1 U21738 ( .C1(n18894), .C2(n18709), .A(n18703), .B(n18702), .ZN(
        P3_U2938) );
  AOI22_X1 U21739 ( .A1(n18900), .A2(n18705), .B1(n18896), .B2(n18704), .ZN(
        n18708) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18706), .B1(
        n18897), .B2(n18729), .ZN(n18707) );
  OAI211_X1 U21741 ( .C1(n18904), .C2(n18709), .A(n18708), .B(n18707), .ZN(
        P3_U2939) );
  NAND2_X1 U21742 ( .A1(n18711), .A2(n18710), .ZN(n18734) );
  NOR2_X1 U21743 ( .A1(n18712), .A2(n18733), .ZN(n18728) );
  AOI22_X1 U21744 ( .A1(n18850), .A2(n18752), .B1(n18849), .B2(n18728), .ZN(
        n18715) );
  NOR2_X1 U21745 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18733), .ZN(
        n18757) );
  AOI22_X1 U21746 ( .A1(n18854), .A2(n18713), .B1(n18851), .B2(n18757), .ZN(
        n18730) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18730), .B1(
        n18855), .B2(n18729), .ZN(n18714) );
  OAI211_X1 U21748 ( .C1(n18858), .C2(n18734), .A(n18715), .B(n18714), .ZN(
        P3_U2940) );
  AOI22_X1 U21749 ( .A1(n18860), .A2(n18728), .B1(n18859), .B2(n18729), .ZN(
        n18717) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18730), .B1(
        n18861), .B2(n18752), .ZN(n18716) );
  OAI211_X1 U21751 ( .C1(n18864), .C2(n18734), .A(n18717), .B(n18716), .ZN(
        P3_U2941) );
  AOI22_X1 U21752 ( .A1(n18866), .A2(n18729), .B1(n18865), .B2(n18728), .ZN(
        n18719) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18730), .B1(
        n18867), .B2(n18752), .ZN(n18718) );
  OAI211_X1 U21754 ( .C1(n18870), .C2(n18734), .A(n18719), .B(n18718), .ZN(
        P3_U2942) );
  AOI22_X1 U21755 ( .A1(n18873), .A2(n18729), .B1(n18871), .B2(n18728), .ZN(
        n18721) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18730), .B1(
        n18872), .B2(n18752), .ZN(n18720) );
  OAI211_X1 U21757 ( .C1(n18876), .C2(n18734), .A(n18721), .B(n18720), .ZN(
        P3_U2943) );
  AOI22_X1 U21758 ( .A1(n18879), .A2(n18729), .B1(n18877), .B2(n18728), .ZN(
        n18723) );
  AOI22_X1 U21759 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18730), .B1(
        n18878), .B2(n18752), .ZN(n18722) );
  OAI211_X1 U21760 ( .C1(n18882), .C2(n18734), .A(n18723), .B(n18722), .ZN(
        P3_U2944) );
  AOI22_X1 U21761 ( .A1(n18884), .A2(n18752), .B1(n18883), .B2(n18728), .ZN(
        n18725) );
  AOI22_X1 U21762 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18730), .B1(
        n18885), .B2(n18729), .ZN(n18724) );
  OAI211_X1 U21763 ( .C1(n18888), .C2(n18734), .A(n18725), .B(n18724), .ZN(
        P3_U2945) );
  AOI22_X1 U21764 ( .A1(n18890), .A2(n18752), .B1(n18889), .B2(n18728), .ZN(
        n18727) );
  AOI22_X1 U21765 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18730), .B1(
        n18891), .B2(n18729), .ZN(n18726) );
  OAI211_X1 U21766 ( .C1(n18894), .C2(n18734), .A(n18727), .B(n18726), .ZN(
        P3_U2946) );
  AOI22_X1 U21767 ( .A1(n18900), .A2(n18729), .B1(n18896), .B2(n18728), .ZN(
        n18732) );
  AOI22_X1 U21768 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18730), .B1(
        n18897), .B2(n18752), .ZN(n18731) );
  OAI211_X1 U21769 ( .C1(n18904), .C2(n18734), .A(n18732), .B(n18731), .ZN(
        P3_U2947) );
  NOR2_X1 U21770 ( .A1(n18942), .A2(n18733), .ZN(n18801) );
  NAND2_X1 U21771 ( .A1(n18801), .A2(n18940), .ZN(n18756) );
  INV_X1 U21772 ( .A(n18734), .ZN(n18795) );
  NOR2_X1 U21773 ( .A1(n18795), .A2(n18817), .ZN(n18778) );
  NOR2_X1 U21774 ( .A1(n18971), .A2(n18778), .ZN(n18751) );
  AOI22_X1 U21775 ( .A1(n18850), .A2(n18773), .B1(n18849), .B2(n18751), .ZN(
        n18738) );
  OAI21_X1 U21776 ( .B1(n18735), .B2(n18823), .A(n18778), .ZN(n18736) );
  OAI211_X1 U21777 ( .C1(n18817), .C2(n19068), .A(n18826), .B(n18736), .ZN(
        n18753) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18753), .B1(
        n18855), .B2(n18752), .ZN(n18737) );
  OAI211_X1 U21779 ( .C1(n18858), .C2(n18756), .A(n18738), .B(n18737), .ZN(
        P3_U2948) );
  AOI22_X1 U21780 ( .A1(n18860), .A2(n18751), .B1(n18859), .B2(n18752), .ZN(
        n18740) );
  AOI22_X1 U21781 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18753), .B1(
        n18861), .B2(n18773), .ZN(n18739) );
  OAI211_X1 U21782 ( .C1(n18864), .C2(n18756), .A(n18740), .B(n18739), .ZN(
        P3_U2949) );
  AOI22_X1 U21783 ( .A1(n18867), .A2(n18773), .B1(n18865), .B2(n18751), .ZN(
        n18742) );
  AOI22_X1 U21784 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18753), .B1(
        n18866), .B2(n18752), .ZN(n18741) );
  OAI211_X1 U21785 ( .C1(n18870), .C2(n18756), .A(n18742), .B(n18741), .ZN(
        P3_U2950) );
  AOI22_X1 U21786 ( .A1(n18873), .A2(n18752), .B1(n18871), .B2(n18751), .ZN(
        n18744) );
  AOI22_X1 U21787 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18753), .B1(
        n18872), .B2(n18773), .ZN(n18743) );
  OAI211_X1 U21788 ( .C1(n18876), .C2(n18756), .A(n18744), .B(n18743), .ZN(
        P3_U2951) );
  AOI22_X1 U21789 ( .A1(n18879), .A2(n18752), .B1(n18877), .B2(n18751), .ZN(
        n18746) );
  AOI22_X1 U21790 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18753), .B1(
        n18878), .B2(n18773), .ZN(n18745) );
  OAI211_X1 U21791 ( .C1(n18882), .C2(n18756), .A(n18746), .B(n18745), .ZN(
        P3_U2952) );
  AOI22_X1 U21792 ( .A1(n18884), .A2(n18773), .B1(n18883), .B2(n18751), .ZN(
        n18748) );
  AOI22_X1 U21793 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18753), .B1(
        n18885), .B2(n18752), .ZN(n18747) );
  OAI211_X1 U21794 ( .C1(n18888), .C2(n18756), .A(n18748), .B(n18747), .ZN(
        P3_U2953) );
  AOI22_X1 U21795 ( .A1(n18889), .A2(n18751), .B1(n18891), .B2(n18752), .ZN(
        n18750) );
  AOI22_X1 U21796 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18753), .B1(
        n18890), .B2(n18773), .ZN(n18749) );
  OAI211_X1 U21797 ( .C1(n18894), .C2(n18756), .A(n18750), .B(n18749), .ZN(
        P3_U2954) );
  AOI22_X1 U21798 ( .A1(n18897), .A2(n18773), .B1(n18896), .B2(n18751), .ZN(
        n18755) );
  AOI22_X1 U21799 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18753), .B1(
        n18900), .B2(n18752), .ZN(n18754) );
  OAI211_X1 U21800 ( .C1(n18904), .C2(n18756), .A(n18755), .B(n18754), .ZN(
        P3_U2955) );
  NAND2_X1 U21801 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18801), .ZN(
        n18777) );
  AND2_X1 U21802 ( .A1(n18964), .A2(n18801), .ZN(n18772) );
  AOI22_X1 U21803 ( .A1(n18850), .A2(n18795), .B1(n18849), .B2(n18772), .ZN(
        n18759) );
  AOI22_X1 U21804 ( .A1(n18854), .A2(n18757), .B1(n18851), .B2(n18801), .ZN(
        n18774) );
  AOI22_X1 U21805 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18774), .B1(
        n18855), .B2(n18773), .ZN(n18758) );
  OAI211_X1 U21806 ( .C1(n18858), .C2(n18777), .A(n18759), .B(n18758), .ZN(
        P3_U2956) );
  AOI22_X1 U21807 ( .A1(n18861), .A2(n18795), .B1(n18860), .B2(n18772), .ZN(
        n18761) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18774), .B1(
        n18859), .B2(n18773), .ZN(n18760) );
  OAI211_X1 U21809 ( .C1(n18864), .C2(n18777), .A(n18761), .B(n18760), .ZN(
        P3_U2957) );
  AOI22_X1 U21810 ( .A1(n18866), .A2(n18773), .B1(n18865), .B2(n18772), .ZN(
        n18763) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18774), .B1(
        n18867), .B2(n18795), .ZN(n18762) );
  OAI211_X1 U21812 ( .C1(n18870), .C2(n18777), .A(n18763), .B(n18762), .ZN(
        P3_U2958) );
  AOI22_X1 U21813 ( .A1(n18872), .A2(n18795), .B1(n18871), .B2(n18772), .ZN(
        n18765) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18774), .B1(
        n18873), .B2(n18773), .ZN(n18764) );
  OAI211_X1 U21815 ( .C1(n18876), .C2(n18777), .A(n18765), .B(n18764), .ZN(
        P3_U2959) );
  AOI22_X1 U21816 ( .A1(n18879), .A2(n18773), .B1(n18877), .B2(n18772), .ZN(
        n18767) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18774), .B1(
        n18878), .B2(n18795), .ZN(n18766) );
  OAI211_X1 U21818 ( .C1(n18882), .C2(n18777), .A(n18767), .B(n18766), .ZN(
        P3_U2960) );
  AOI22_X1 U21819 ( .A1(n18885), .A2(n18773), .B1(n18883), .B2(n18772), .ZN(
        n18769) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18774), .B1(
        n18884), .B2(n18795), .ZN(n18768) );
  OAI211_X1 U21821 ( .C1(n18888), .C2(n18777), .A(n18769), .B(n18768), .ZN(
        P3_U2961) );
  AOI22_X1 U21822 ( .A1(n18890), .A2(n18795), .B1(n18889), .B2(n18772), .ZN(
        n18771) );
  AOI22_X1 U21823 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18774), .B1(
        n18891), .B2(n18773), .ZN(n18770) );
  OAI211_X1 U21824 ( .C1(n18894), .C2(n18777), .A(n18771), .B(n18770), .ZN(
        P3_U2962) );
  AOI22_X1 U21825 ( .A1(n18897), .A2(n18795), .B1(n18896), .B2(n18772), .ZN(
        n18776) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18774), .B1(
        n18900), .B2(n18773), .ZN(n18775) );
  OAI211_X1 U21827 ( .C1(n18904), .C2(n18777), .A(n18776), .B(n18775), .ZN(
        P3_U2963) );
  INV_X1 U21828 ( .A(n18853), .ZN(n18800) );
  NOR2_X2 U21829 ( .A1(n18800), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18899) );
  INV_X1 U21830 ( .A(n18899), .ZN(n18799) );
  INV_X1 U21831 ( .A(n18777), .ZN(n18843) );
  NOR2_X1 U21832 ( .A1(n18843), .A2(n18899), .ZN(n18824) );
  NOR2_X1 U21833 ( .A1(n18971), .A2(n18824), .ZN(n18794) );
  AOI22_X1 U21834 ( .A1(n18850), .A2(n18817), .B1(n18849), .B2(n18794), .ZN(
        n18781) );
  OAI21_X1 U21835 ( .B1(n18778), .B2(n18823), .A(n18824), .ZN(n18779) );
  OAI211_X1 U21836 ( .C1(n18899), .C2(n19068), .A(n18826), .B(n18779), .ZN(
        n18796) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18796), .B1(
        n18855), .B2(n18795), .ZN(n18780) );
  OAI211_X1 U21838 ( .C1(n18858), .C2(n18799), .A(n18781), .B(n18780), .ZN(
        P3_U2964) );
  AOI22_X1 U21839 ( .A1(n18861), .A2(n18817), .B1(n18860), .B2(n18794), .ZN(
        n18783) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18796), .B1(
        n18859), .B2(n18795), .ZN(n18782) );
  OAI211_X1 U21841 ( .C1(n18864), .C2(n18799), .A(n18783), .B(n18782), .ZN(
        P3_U2965) );
  AOI22_X1 U21842 ( .A1(n18866), .A2(n18795), .B1(n18865), .B2(n18794), .ZN(
        n18785) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18796), .B1(
        n18867), .B2(n18817), .ZN(n18784) );
  OAI211_X1 U21844 ( .C1(n18870), .C2(n18799), .A(n18785), .B(n18784), .ZN(
        P3_U2966) );
  AOI22_X1 U21845 ( .A1(n18873), .A2(n18795), .B1(n18871), .B2(n18794), .ZN(
        n18787) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18796), .B1(
        n18872), .B2(n18817), .ZN(n18786) );
  OAI211_X1 U21847 ( .C1(n18876), .C2(n18799), .A(n18787), .B(n18786), .ZN(
        P3_U2967) );
  AOI22_X1 U21848 ( .A1(n18879), .A2(n18795), .B1(n18877), .B2(n18794), .ZN(
        n18789) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18796), .B1(
        n18878), .B2(n18817), .ZN(n18788) );
  OAI211_X1 U21850 ( .C1(n18882), .C2(n18799), .A(n18789), .B(n18788), .ZN(
        P3_U2968) );
  AOI22_X1 U21851 ( .A1(n18884), .A2(n18817), .B1(n18883), .B2(n18794), .ZN(
        n18791) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18796), .B1(
        n18885), .B2(n18795), .ZN(n18790) );
  OAI211_X1 U21853 ( .C1(n18888), .C2(n18799), .A(n18791), .B(n18790), .ZN(
        P3_U2969) );
  AOI22_X1 U21854 ( .A1(n18890), .A2(n18817), .B1(n18889), .B2(n18794), .ZN(
        n18793) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18796), .B1(
        n18891), .B2(n18795), .ZN(n18792) );
  OAI211_X1 U21856 ( .C1(n18894), .C2(n18799), .A(n18793), .B(n18792), .ZN(
        P3_U2970) );
  AOI22_X1 U21857 ( .A1(n18900), .A2(n18795), .B1(n18896), .B2(n18794), .ZN(
        n18798) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18796), .B1(
        n18897), .B2(n18817), .ZN(n18797) );
  OAI211_X1 U21859 ( .C1(n18904), .C2(n18799), .A(n18798), .B(n18797), .ZN(
        P3_U2971) );
  NOR2_X1 U21860 ( .A1(n18971), .A2(n18800), .ZN(n18816) );
  AOI22_X1 U21861 ( .A1(n18855), .A2(n18817), .B1(n18849), .B2(n18816), .ZN(
        n18803) );
  AOI22_X1 U21862 ( .A1(n18854), .A2(n18801), .B1(n18853), .B2(n18851), .ZN(
        n18818) );
  AOI22_X1 U21863 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18818), .B1(
        n18850), .B2(n18843), .ZN(n18802) );
  OAI211_X1 U21864 ( .C1(n18821), .C2(n18858), .A(n18803), .B(n18802), .ZN(
        P3_U2972) );
  AOI22_X1 U21865 ( .A1(n18860), .A2(n18816), .B1(n18859), .B2(n18817), .ZN(
        n18805) );
  AOI22_X1 U21866 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18818), .B1(
        n18861), .B2(n18843), .ZN(n18804) );
  OAI211_X1 U21867 ( .C1(n18821), .C2(n18864), .A(n18805), .B(n18804), .ZN(
        P3_U2973) );
  AOI22_X1 U21868 ( .A1(n18867), .A2(n18843), .B1(n18865), .B2(n18816), .ZN(
        n18807) );
  AOI22_X1 U21869 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18818), .B1(
        n18866), .B2(n18817), .ZN(n18806) );
  OAI211_X1 U21870 ( .C1(n18821), .C2(n18870), .A(n18807), .B(n18806), .ZN(
        P3_U2974) );
  AOI22_X1 U21871 ( .A1(n18872), .A2(n18843), .B1(n18871), .B2(n18816), .ZN(
        n18809) );
  AOI22_X1 U21872 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18818), .B1(
        n18873), .B2(n18817), .ZN(n18808) );
  OAI211_X1 U21873 ( .C1(n18821), .C2(n18876), .A(n18809), .B(n18808), .ZN(
        P3_U2975) );
  AOI22_X1 U21874 ( .A1(n18879), .A2(n18817), .B1(n18877), .B2(n18816), .ZN(
        n18811) );
  AOI22_X1 U21875 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18818), .B1(
        n18878), .B2(n18843), .ZN(n18810) );
  OAI211_X1 U21876 ( .C1(n18821), .C2(n18882), .A(n18811), .B(n18810), .ZN(
        P3_U2976) );
  AOI22_X1 U21877 ( .A1(n18885), .A2(n18817), .B1(n18883), .B2(n18816), .ZN(
        n18813) );
  AOI22_X1 U21878 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18818), .B1(
        n18884), .B2(n18843), .ZN(n18812) );
  OAI211_X1 U21879 ( .C1(n18821), .C2(n18888), .A(n18813), .B(n18812), .ZN(
        P3_U2977) );
  AOI22_X1 U21880 ( .A1(n18889), .A2(n18816), .B1(n18891), .B2(n18817), .ZN(
        n18815) );
  AOI22_X1 U21881 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18818), .B1(
        n18890), .B2(n18843), .ZN(n18814) );
  OAI211_X1 U21882 ( .C1(n18821), .C2(n18894), .A(n18815), .B(n18814), .ZN(
        P3_U2978) );
  AOI22_X1 U21883 ( .A1(n18900), .A2(n18817), .B1(n18896), .B2(n18816), .ZN(
        n18820) );
  AOI22_X1 U21884 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18818), .B1(
        n18897), .B2(n18843), .ZN(n18819) );
  OAI211_X1 U21885 ( .C1(n18821), .C2(n18904), .A(n18820), .B(n18819), .ZN(
        P3_U2979) );
  NOR2_X1 U21886 ( .A1(n18971), .A2(n18822), .ZN(n18842) );
  AOI22_X1 U21887 ( .A1(n18850), .A2(n18899), .B1(n18849), .B2(n18842), .ZN(
        n18829) );
  OAI21_X1 U21888 ( .B1(n18824), .B2(n18823), .A(n18822), .ZN(n18825) );
  OAI211_X1 U21889 ( .C1(n18827), .C2(n19068), .A(n18826), .B(n18825), .ZN(
        n18844) );
  AOI22_X1 U21890 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18844), .B1(
        n18855), .B2(n18843), .ZN(n18828) );
  OAI211_X1 U21891 ( .C1(n18847), .C2(n18858), .A(n18829), .B(n18828), .ZN(
        P3_U2980) );
  AOI22_X1 U21892 ( .A1(n18861), .A2(n18899), .B1(n18860), .B2(n18842), .ZN(
        n18831) );
  AOI22_X1 U21893 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18844), .B1(
        n18859), .B2(n18843), .ZN(n18830) );
  OAI211_X1 U21894 ( .C1(n18847), .C2(n18864), .A(n18831), .B(n18830), .ZN(
        P3_U2981) );
  AOI22_X1 U21895 ( .A1(n18866), .A2(n18843), .B1(n18865), .B2(n18842), .ZN(
        n18833) );
  AOI22_X1 U21896 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18844), .B1(
        n18867), .B2(n18899), .ZN(n18832) );
  OAI211_X1 U21897 ( .C1(n18847), .C2(n18870), .A(n18833), .B(n18832), .ZN(
        P3_U2982) );
  AOI22_X1 U21898 ( .A1(n18872), .A2(n18899), .B1(n18871), .B2(n18842), .ZN(
        n18835) );
  AOI22_X1 U21899 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18844), .B1(
        n18873), .B2(n18843), .ZN(n18834) );
  OAI211_X1 U21900 ( .C1(n18847), .C2(n18876), .A(n18835), .B(n18834), .ZN(
        P3_U2983) );
  AOI22_X1 U21901 ( .A1(n18878), .A2(n18899), .B1(n18877), .B2(n18842), .ZN(
        n18837) );
  AOI22_X1 U21902 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18844), .B1(
        n18879), .B2(n18843), .ZN(n18836) );
  OAI211_X1 U21903 ( .C1(n18847), .C2(n18882), .A(n18837), .B(n18836), .ZN(
        P3_U2984) );
  AOI22_X1 U21904 ( .A1(n18885), .A2(n18843), .B1(n18883), .B2(n18842), .ZN(
        n18839) );
  AOI22_X1 U21905 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18844), .B1(
        n18884), .B2(n18899), .ZN(n18838) );
  OAI211_X1 U21906 ( .C1(n18847), .C2(n18888), .A(n18839), .B(n18838), .ZN(
        P3_U2985) );
  AOI22_X1 U21907 ( .A1(n18889), .A2(n18842), .B1(n18891), .B2(n18843), .ZN(
        n18841) );
  AOI22_X1 U21908 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18844), .B1(
        n18890), .B2(n18899), .ZN(n18840) );
  OAI211_X1 U21909 ( .C1(n18847), .C2(n18894), .A(n18841), .B(n18840), .ZN(
        P3_U2986) );
  AOI22_X1 U21910 ( .A1(n18897), .A2(n18899), .B1(n18896), .B2(n18842), .ZN(
        n18846) );
  AOI22_X1 U21911 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18844), .B1(
        n18900), .B2(n18843), .ZN(n18845) );
  OAI211_X1 U21912 ( .C1(n18847), .C2(n18904), .A(n18846), .B(n18845), .ZN(
        P3_U2987) );
  INV_X1 U21913 ( .A(n18852), .ZN(n18848) );
  NOR2_X1 U21914 ( .A1(n18971), .A2(n18848), .ZN(n18895) );
  AOI22_X1 U21915 ( .A1(n18898), .A2(n18850), .B1(n18849), .B2(n18895), .ZN(
        n18857) );
  AOI22_X1 U21916 ( .A1(n18854), .A2(n18853), .B1(n18852), .B2(n18851), .ZN(
        n18901) );
  AOI22_X1 U21917 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18901), .B1(
        n18855), .B2(n18899), .ZN(n18856) );
  OAI211_X1 U21918 ( .C1(n18905), .C2(n18858), .A(n18857), .B(n18856), .ZN(
        P3_U2988) );
  AOI22_X1 U21919 ( .A1(n18860), .A2(n18895), .B1(n18859), .B2(n18899), .ZN(
        n18863) );
  AOI22_X1 U21920 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18901), .B1(
        n18898), .B2(n18861), .ZN(n18862) );
  OAI211_X1 U21921 ( .C1(n18905), .C2(n18864), .A(n18863), .B(n18862), .ZN(
        P3_U2989) );
  AOI22_X1 U21922 ( .A1(n18866), .A2(n18899), .B1(n18865), .B2(n18895), .ZN(
        n18869) );
  AOI22_X1 U21923 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18901), .B1(
        n18898), .B2(n18867), .ZN(n18868) );
  OAI211_X1 U21924 ( .C1(n18905), .C2(n18870), .A(n18869), .B(n18868), .ZN(
        P3_U2990) );
  AOI22_X1 U21925 ( .A1(n18898), .A2(n18872), .B1(n18871), .B2(n18895), .ZN(
        n18875) );
  AOI22_X1 U21926 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18901), .B1(
        n18873), .B2(n18899), .ZN(n18874) );
  OAI211_X1 U21927 ( .C1(n18905), .C2(n18876), .A(n18875), .B(n18874), .ZN(
        P3_U2991) );
  AOI22_X1 U21928 ( .A1(n18898), .A2(n18878), .B1(n18877), .B2(n18895), .ZN(
        n18881) );
  AOI22_X1 U21929 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18901), .B1(
        n18879), .B2(n18899), .ZN(n18880) );
  OAI211_X1 U21930 ( .C1(n18905), .C2(n18882), .A(n18881), .B(n18880), .ZN(
        P3_U2992) );
  AOI22_X1 U21931 ( .A1(n18898), .A2(n18884), .B1(n18883), .B2(n18895), .ZN(
        n18887) );
  AOI22_X1 U21932 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18901), .B1(
        n18885), .B2(n18899), .ZN(n18886) );
  OAI211_X1 U21933 ( .C1(n18905), .C2(n18888), .A(n18887), .B(n18886), .ZN(
        P3_U2993) );
  AOI22_X1 U21934 ( .A1(n18898), .A2(n18890), .B1(n18889), .B2(n18895), .ZN(
        n18893) );
  AOI22_X1 U21935 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18901), .B1(
        n18891), .B2(n18899), .ZN(n18892) );
  OAI211_X1 U21936 ( .C1(n18905), .C2(n18894), .A(n18893), .B(n18892), .ZN(
        P3_U2994) );
  AOI22_X1 U21937 ( .A1(n18898), .A2(n18897), .B1(n18896), .B2(n18895), .ZN(
        n18903) );
  AOI22_X1 U21938 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18901), .B1(
        n18900), .B2(n18899), .ZN(n18902) );
  OAI211_X1 U21939 ( .C1(n18905), .C2(n18904), .A(n18903), .B(n18902), .ZN(
        P3_U2995) );
  NOR2_X1 U21940 ( .A1(n18933), .A2(n18906), .ZN(n18908) );
  OAI222_X1 U21941 ( .A1(n18912), .A2(n18911), .B1(n18910), .B2(n18909), .C1(
        n18908), .C2(n18907), .ZN(n19105) );
  OAI21_X1 U21942 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18913), .ZN(n18915) );
  OAI211_X1 U21943 ( .C1(n18934), .C2(n18916), .A(n18915), .B(n18914), .ZN(
        n18956) );
  INV_X1 U21944 ( .A(n18934), .ZN(n18945) );
  NAND3_X1 U21945 ( .A1(n18918), .A2(n18917), .A3(n18937), .ZN(n18928) );
  AOI211_X1 U21946 ( .C1(n18928), .C2(n18922), .A(n18923), .B(n19072), .ZN(
        n18927) );
  OAI21_X1 U21947 ( .B1(n18919), .B2(n18918), .A(n18917), .ZN(n18920) );
  NAND2_X1 U21948 ( .A1(n17147), .A2(n18920), .ZN(n18930) );
  AOI21_X1 U21949 ( .B1(n9660), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n18921), .ZN(n18938) );
  OAI22_X1 U21950 ( .A1(n18924), .A2(n18923), .B1(n18922), .B2(n18938), .ZN(
        n18925) );
  INV_X1 U21951 ( .A(n18925), .ZN(n18926) );
  AOI22_X1 U21952 ( .A1(n18927), .A2(n18930), .B1(n18926), .B2(n19072), .ZN(
        n19070) );
  AOI22_X1 U21953 ( .A1(n18945), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19070), .B2(n18934), .ZN(n18954) );
  NOR3_X1 U21954 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18938), .A3(
        n12318), .ZN(n18932) );
  INV_X1 U21955 ( .A(n18928), .ZN(n18929) );
  AOI211_X1 U21956 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n18930), .A(
        n18929), .B(n12320), .ZN(n18931) );
  AOI211_X1 U21957 ( .C1(n18933), .C2(n19076), .A(n18932), .B(n18931), .ZN(
        n19079) );
  AOI22_X1 U21958 ( .A1(n18945), .A2(n12320), .B1(n19079), .B2(n18934), .ZN(
        n18949) );
  NOR2_X1 U21959 ( .A1(n18936), .A2(n9660), .ZN(n18939) );
  AOI22_X1 U21960 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18937), .B1(
        n18939), .B2(n17147), .ZN(n19090) );
  OAI22_X1 U21961 ( .A1(n18939), .A2(n19083), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18938), .ZN(n19087) );
  OR3_X1 U21962 ( .A1(n19090), .A2(n18942), .A3(n18940), .ZN(n18941) );
  AOI22_X1 U21963 ( .A1(n19090), .A2(n18942), .B1(n19087), .B2(n18941), .ZN(
        n18944) );
  OAI21_X1 U21964 ( .B1(n18945), .B2(n18944), .A(n18943), .ZN(n18948) );
  AND2_X1 U21965 ( .A1(n18949), .A2(n18948), .ZN(n18946) );
  OAI221_X1 U21966 ( .B1(n18949), .B2(n18948), .C1(n18947), .C2(n18946), .A(
        n18951), .ZN(n18953) );
  AOI21_X1 U21967 ( .B1(n18951), .B2(n18950), .A(n18949), .ZN(n18952) );
  AOI222_X1 U21968 ( .A1(n18954), .A2(n18953), .B1(n18954), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18953), .C2(n18952), .ZN(
        n18955) );
  NOR4_X1 U21969 ( .A1(n18957), .A2(n19105), .A3(n18956), .A4(n18955), .ZN(
        n18968) );
  INV_X1 U21970 ( .A(n19077), .ZN(n19089) );
  NAND2_X1 U21971 ( .A1(n19075), .A2(n19123), .ZN(n18977) );
  INV_X1 U21972 ( .A(n18977), .ZN(n19115) );
  AOI22_X1 U21973 ( .A1(n19089), .A2(n19115), .B1(n18988), .B2(n19109), .ZN(
        n18958) );
  INV_X1 U21974 ( .A(n18958), .ZN(n18963) );
  OAI211_X1 U21975 ( .C1(n18960), .C2(n18959), .A(n19107), .B(n18968), .ZN(
        n19067) );
  OAI21_X1 U21976 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19113), .A(n19067), 
        .ZN(n18969) );
  NOR2_X1 U21977 ( .A1(n18961), .A2(n18969), .ZN(n18962) );
  MUX2_X1 U21978 ( .A(n18963), .B(n18962), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18966) );
  OR2_X1 U21979 ( .A1(n18970), .A2(n18964), .ZN(n18965) );
  OAI211_X1 U21980 ( .C1(n18968), .C2(n18967), .A(n18966), .B(n18965), .ZN(
        P3_U2996) );
  NAND2_X1 U21981 ( .A1(n18988), .A2(n19109), .ZN(n18973) );
  NAND4_X1 U21982 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n18988), .A4(n19123), .ZN(n18975) );
  OR3_X1 U21983 ( .A1(n18971), .A2(n18970), .A3(n18969), .ZN(n18972) );
  NAND4_X1 U21984 ( .A1(n18974), .A2(n18973), .A3(n18975), .A4(n18972), .ZN(
        P3_U2997) );
  AND4_X1 U21985 ( .A1(n18977), .A2(n18976), .A3(n18975), .A4(n19066), .ZN(
        P3_U2998) );
  AND2_X1 U21986 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18978), .ZN(
        P3_U2999) );
  AND2_X1 U21987 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18978), .ZN(
        P3_U3000) );
  AND2_X1 U21988 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18978), .ZN(
        P3_U3001) );
  AND2_X1 U21989 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18978), .ZN(
        P3_U3002) );
  AND2_X1 U21990 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18978), .ZN(
        P3_U3003) );
  AND2_X1 U21991 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18978), .ZN(
        P3_U3004) );
  AND2_X1 U21992 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18978), .ZN(
        P3_U3005) );
  AND2_X1 U21993 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18978), .ZN(
        P3_U3006) );
  AND2_X1 U21994 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18978), .ZN(
        P3_U3007) );
  AND2_X1 U21995 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18978), .ZN(
        P3_U3008) );
  AND2_X1 U21996 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18978), .ZN(
        P3_U3009) );
  INV_X1 U21997 ( .A(n19065), .ZN(n18979) );
  AND2_X1 U21998 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18979), .ZN(
        P3_U3010) );
  AND2_X1 U21999 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18979), .ZN(
        P3_U3011) );
  AND2_X1 U22000 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18979), .ZN(
        P3_U3012) );
  AND2_X1 U22001 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18979), .ZN(
        P3_U3013) );
  INV_X1 U22002 ( .A(P3_DATAWIDTH_REG_16__SCAN_IN), .ZN(n21092) );
  NOR2_X1 U22003 ( .A1(n21092), .A2(n19065), .ZN(P3_U3014) );
  AND2_X1 U22004 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18979), .ZN(
        P3_U3015) );
  AND2_X1 U22005 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18979), .ZN(
        P3_U3016) );
  AND2_X1 U22006 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18979), .ZN(
        P3_U3017) );
  AND2_X1 U22007 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18979), .ZN(
        P3_U3018) );
  AND2_X1 U22008 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18979), .ZN(
        P3_U3019) );
  AND2_X1 U22009 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18979), .ZN(
        P3_U3020) );
  AND2_X1 U22010 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18979), .ZN(P3_U3021) );
  AND2_X1 U22011 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18979), .ZN(P3_U3022) );
  AND2_X1 U22012 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18978), .ZN(P3_U3023) );
  AND2_X1 U22013 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18979), .ZN(P3_U3024) );
  AND2_X1 U22014 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18978), .ZN(P3_U3025) );
  AND2_X1 U22015 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18979), .ZN(P3_U3026) );
  AND2_X1 U22016 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18979), .ZN(P3_U3027) );
  AND2_X1 U22017 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18979), .ZN(P3_U3028) );
  INV_X1 U22018 ( .A(n18985), .ZN(n18984) );
  OAI21_X1 U22019 ( .B1(n18980), .B2(n20110), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18981) );
  AOI22_X1 U22020 ( .A1(n18994), .A2(n18996), .B1(n19120), .B2(n18981), .ZN(
        n18983) );
  NAND3_X1 U22021 ( .A1(NA), .A2(n18994), .A3(n18982), .ZN(n18987) );
  OAI211_X1 U22022 ( .C1(n19113), .C2(n18984), .A(n18983), .B(n18987), .ZN(
        P3_U3029) );
  NAND2_X1 U22023 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n18989) );
  AOI22_X1 U22024 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18989), .B1(HOLD), 
        .B2(n18985), .ZN(n18986) );
  NAND2_X1 U22025 ( .A1(n18988), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18990) );
  OAI211_X1 U22026 ( .C1(n18986), .C2(n18994), .A(n18990), .B(n19110), .ZN(
        P3_U3030) );
  AOI22_X1 U22027 ( .A1(n18988), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n18994), 
        .B2(n18987), .ZN(n18995) );
  INV_X1 U22028 ( .A(n18989), .ZN(n18992) );
  OAI22_X1 U22029 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18990), .ZN(n18991) );
  OAI22_X1 U22030 ( .A1(n18992), .A2(n18991), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18993) );
  OAI22_X1 U22031 ( .A1(n18995), .A2(n18996), .B1(n18994), .B2(n18993), .ZN(
        P3_U3031) );
  OAI222_X1 U22032 ( .A1(n19095), .A2(n9664), .B1(n18997), .B2(n19055), .C1(
        n18998), .C2(n19044), .ZN(P3_U3032) );
  OAI222_X1 U22033 ( .A1(n19044), .A2(n19000), .B1(n18999), .B2(n19121), .C1(
        n18998), .C2(n9664), .ZN(P3_U3033) );
  OAI222_X1 U22034 ( .A1(n19044), .A2(n19003), .B1(n19001), .B2(n19055), .C1(
        n19000), .C2(n9664), .ZN(P3_U3034) );
  OAI222_X1 U22035 ( .A1(n19044), .A2(n19005), .B1(n19004), .B2(n19121), .C1(
        n19003), .C2(n9664), .ZN(P3_U3035) );
  OAI222_X1 U22036 ( .A1(n19044), .A2(n19007), .B1(n19006), .B2(n19055), .C1(
        n19005), .C2(n9664), .ZN(P3_U3036) );
  OAI222_X1 U22037 ( .A1(n19044), .A2(n19009), .B1(n19008), .B2(n19121), .C1(
        n19007), .C2(n9664), .ZN(P3_U3037) );
  OAI222_X1 U22038 ( .A1(n19044), .A2(n19012), .B1(n19010), .B2(n19121), .C1(
        n19009), .C2(n9664), .ZN(P3_U3038) );
  OAI222_X1 U22039 ( .A1(n19012), .A2(n9664), .B1(n19011), .B2(n19121), .C1(
        n19013), .C2(n19044), .ZN(P3_U3039) );
  OAI222_X1 U22040 ( .A1(n19044), .A2(n21188), .B1(n19014), .B2(n19121), .C1(
        n19013), .C2(n9664), .ZN(P3_U3040) );
  INV_X1 U22041 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19016) );
  OAI222_X1 U22042 ( .A1(n19044), .A2(n19016), .B1(n19015), .B2(n19121), .C1(
        n21188), .C2(n9664), .ZN(P3_U3041) );
  OAI222_X1 U22043 ( .A1(n19044), .A2(n19018), .B1(n19017), .B2(n19121), .C1(
        n19016), .C2(n9664), .ZN(P3_U3042) );
  OAI222_X1 U22044 ( .A1(n19044), .A2(n19020), .B1(n19019), .B2(n19121), .C1(
        n19018), .C2(n9664), .ZN(P3_U3043) );
  OAI222_X1 U22045 ( .A1(n19044), .A2(n19023), .B1(n19021), .B2(n19121), .C1(
        n19020), .C2(n9664), .ZN(P3_U3044) );
  OAI222_X1 U22046 ( .A1(n19023), .A2(n9664), .B1(n19022), .B2(n19121), .C1(
        n19024), .C2(n19044), .ZN(P3_U3045) );
  OAI222_X1 U22047 ( .A1(n19044), .A2(n19026), .B1(n19025), .B2(n19121), .C1(
        n19024), .C2(n9664), .ZN(P3_U3046) );
  OAI222_X1 U22048 ( .A1(n19044), .A2(n19028), .B1(n19027), .B2(n19121), .C1(
        n19026), .C2(n9664), .ZN(P3_U3047) );
  OAI222_X1 U22049 ( .A1(n19044), .A2(n19030), .B1(n19029), .B2(n19121), .C1(
        n19028), .C2(n9664), .ZN(P3_U3048) );
  OAI222_X1 U22050 ( .A1(n19044), .A2(n19032), .B1(n19031), .B2(n19121), .C1(
        n19030), .C2(n9664), .ZN(P3_U3049) );
  OAI222_X1 U22051 ( .A1(n19044), .A2(n19034), .B1(n19033), .B2(n19121), .C1(
        n19032), .C2(n9664), .ZN(P3_U3050) );
  OAI222_X1 U22052 ( .A1(n19044), .A2(n19036), .B1(n19035), .B2(n19121), .C1(
        n19034), .C2(n9664), .ZN(P3_U3051) );
  OAI222_X1 U22053 ( .A1(n19044), .A2(n19038), .B1(n19037), .B2(n19121), .C1(
        n19036), .C2(n9664), .ZN(P3_U3052) );
  OAI222_X1 U22054 ( .A1(n19044), .A2(n19040), .B1(n19039), .B2(n19121), .C1(
        n19038), .C2(n9664), .ZN(P3_U3053) );
  OAI222_X1 U22055 ( .A1(n19044), .A2(n19042), .B1(n19041), .B2(n19121), .C1(
        n19040), .C2(n9664), .ZN(P3_U3054) );
  OAI222_X1 U22056 ( .A1(n19044), .A2(n19045), .B1(n19043), .B2(n19055), .C1(
        n19042), .C2(n9664), .ZN(P3_U3055) );
  OAI222_X1 U22057 ( .A1(n19044), .A2(n19047), .B1(n19046), .B2(n19055), .C1(
        n19045), .C2(n9664), .ZN(P3_U3056) );
  OAI222_X1 U22058 ( .A1(n19044), .A2(n19049), .B1(n19048), .B2(n19055), .C1(
        n19047), .C2(n9664), .ZN(P3_U3057) );
  INV_X1 U22059 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21069) );
  OAI222_X1 U22060 ( .A1(n19044), .A2(n21069), .B1(n19050), .B2(n19055), .C1(
        n19049), .C2(n9664), .ZN(P3_U3058) );
  INV_X1 U22061 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19052) );
  OAI222_X1 U22062 ( .A1(n21069), .A2(n9664), .B1(n19051), .B2(n19055), .C1(
        n19052), .C2(n19044), .ZN(P3_U3059) );
  OAI222_X1 U22063 ( .A1(n19044), .A2(n19057), .B1(n19053), .B2(n19055), .C1(
        n19052), .C2(n9664), .ZN(P3_U3060) );
  OAI222_X1 U22064 ( .A1(n9664), .A2(n19057), .B1(n19056), .B2(n19055), .C1(
        n19054), .C2(n19044), .ZN(P3_U3061) );
  OAI22_X1 U22065 ( .A1(n19120), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19121), .ZN(n19058) );
  INV_X1 U22066 ( .A(n19058), .ZN(P3_U3274) );
  OAI22_X1 U22067 ( .A1(n19120), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19121), .ZN(n19059) );
  INV_X1 U22068 ( .A(n19059), .ZN(P3_U3275) );
  OAI22_X1 U22069 ( .A1(n19120), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19121), .ZN(n19060) );
  INV_X1 U22070 ( .A(n19060), .ZN(P3_U3276) );
  OAI22_X1 U22071 ( .A1(n19120), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19121), .ZN(n19061) );
  INV_X1 U22072 ( .A(n19061), .ZN(P3_U3277) );
  OAI21_X1 U22073 ( .B1(n19065), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19063), 
        .ZN(n19062) );
  INV_X1 U22074 ( .A(n19062), .ZN(P3_U3280) );
  OAI21_X1 U22075 ( .B1(n19065), .B2(n19064), .A(n19063), .ZN(P3_U3281) );
  OAI221_X1 U22076 ( .B1(n19068), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19068), 
        .C2(n19067), .A(n19066), .ZN(P3_U3282) );
  INV_X1 U22077 ( .A(n19078), .ZN(n19124) );
  AOI22_X1 U22078 ( .A1(n19124), .A2(n19070), .B1(n19089), .B2(n19069), .ZN(
        n19071) );
  INV_X1 U22079 ( .A(n19094), .ZN(n19092) );
  AOI22_X1 U22080 ( .A1(n19094), .A2(n19072), .B1(n19071), .B2(n19092), .ZN(
        P3_U3285) );
  OAI22_X1 U22081 ( .A1(n19074), .A2(n19073), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19085) );
  INV_X1 U22082 ( .A(n19085), .ZN(n19081) );
  NOR2_X1 U22083 ( .A1(n19075), .A2(n19091), .ZN(n19084) );
  OAI22_X1 U22084 ( .A1(n19079), .A2(n19078), .B1(n19077), .B2(n19076), .ZN(
        n19080) );
  AOI21_X1 U22085 ( .B1(n19081), .B2(n19084), .A(n19080), .ZN(n19082) );
  AOI22_X1 U22086 ( .A1(n19094), .A2(n12320), .B1(n19082), .B2(n19092), .ZN(
        P3_U3288) );
  INV_X1 U22087 ( .A(n19083), .ZN(n19086) );
  AOI222_X1 U22088 ( .A1(n19087), .A2(n19124), .B1(n19089), .B2(n19086), .C1(
        n19085), .C2(n19084), .ZN(n19088) );
  AOI22_X1 U22089 ( .A1(n19094), .A2(n12318), .B1(n19088), .B2(n19092), .ZN(
        P3_U3289) );
  AOI222_X1 U22090 ( .A1(n19091), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19124), 
        .B2(n19090), .C1(n17147), .C2(n19089), .ZN(n19093) );
  AOI22_X1 U22091 ( .A1(n19094), .A2(n17147), .B1(n19093), .B2(n19092), .ZN(
        P3_U3290) );
  AOI21_X1 U22092 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19096) );
  AOI22_X1 U22093 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19096), .B2(n19095), .ZN(n19099) );
  INV_X1 U22094 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19098) );
  AOI22_X1 U22095 ( .A1(n19102), .A2(n19099), .B1(n19098), .B2(n19097), .ZN(
        P3_U3292) );
  INV_X1 U22096 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19101) );
  OAI21_X1 U22097 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19102), .ZN(n19100) );
  OAI21_X1 U22098 ( .B1(n19102), .B2(n19101), .A(n19100), .ZN(P3_U3293) );
  INV_X1 U22099 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19103) );
  AOI22_X1 U22100 ( .A1(n19121), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19103), 
        .B2(n19120), .ZN(P3_U3294) );
  MUX2_X1 U22101 ( .A(P3_MORE_REG_SCAN_IN), .B(n19105), .S(n19104), .Z(
        P3_U3295) );
  OAI21_X1 U22102 ( .B1(n19107), .B2(n19106), .A(n19126), .ZN(n19108) );
  AOI21_X1 U22103 ( .B1(n19109), .B2(n19113), .A(n19108), .ZN(n19119) );
  AOI21_X1 U22104 ( .B1(n19112), .B2(n19111), .A(n19110), .ZN(n19114) );
  OAI211_X1 U22105 ( .C1(n19125), .C2(n19114), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19113), .ZN(n19116) );
  AOI21_X1 U22106 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19116), .A(n19115), 
        .ZN(n19118) );
  NAND2_X1 U22107 ( .A1(n19119), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19117) );
  OAI21_X1 U22108 ( .B1(n19119), .B2(n19118), .A(n19117), .ZN(P3_U3296) );
  INV_X1 U22109 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19130) );
  AOI22_X1 U22110 ( .A1(n19121), .A2(n19130), .B1(n21206), .B2(n19120), .ZN(
        P3_U3297) );
  AOI21_X1 U22111 ( .B1(n19124), .B2(n19123), .A(n19122), .ZN(n19131) );
  INV_X1 U22112 ( .A(n19131), .ZN(n19127) );
  OAI22_X1 U22113 ( .A1(n19127), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19126), 
        .B2(n19125), .ZN(n19128) );
  INV_X1 U22114 ( .A(n19128), .ZN(P3_U3298) );
  AOI21_X1 U22115 ( .B1(n19131), .B2(n19130), .A(n19129), .ZN(P3_U3299) );
  NAND2_X1 U22116 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20120), .ZN(n20109) );
  AOI22_X1 U22117 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20109), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n20103), .ZN(n20173) );
  AOI21_X1 U22118 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20173), .ZN(n19132) );
  INV_X1 U22119 ( .A(n19132), .ZN(P2_U2815) );
  INV_X1 U22120 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19134) );
  OAI22_X1 U22121 ( .A1(n20221), .A2(n19134), .B1(n19133), .B2(n20183), .ZN(
        P2_U2816) );
  NAND2_X1 U22122 ( .A1(n20103), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20235) );
  INV_X2 U22123 ( .A(n20235), .ZN(n20163) );
  NAND2_X1 U22124 ( .A1(n19136), .A2(n20235), .ZN(n20106) );
  AOI21_X1 U22125 ( .B1(n20103), .B2(n20106), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19135) );
  AOI21_X1 U22126 ( .B1(n20163), .B2(P2_CODEFETCH_REG_SCAN_IN), .A(n19135), 
        .ZN(P2_U2817) );
  INV_X1 U22127 ( .A(n19136), .ZN(n20112) );
  OAI21_X1 U22128 ( .B1(n20112), .B2(BS16), .A(n20173), .ZN(n20171) );
  OAI21_X1 U22129 ( .B1(n20173), .B2(n20228), .A(n20171), .ZN(P2_U2818) );
  NOR4_X1 U22130 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19140) );
  NOR4_X1 U22131 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19139) );
  NOR4_X1 U22132 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19138) );
  NOR4_X1 U22133 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19137) );
  NAND4_X1 U22134 ( .A1(n19140), .A2(n19139), .A3(n19138), .A4(n19137), .ZN(
        n19146) );
  NOR4_X1 U22135 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19144) );
  AOI211_X1 U22136 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19143) );
  NOR4_X1 U22137 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19142) );
  NOR4_X1 U22138 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19141) );
  NAND4_X1 U22139 ( .A1(n19144), .A2(n19143), .A3(n19142), .A4(n19141), .ZN(
        n19145) );
  NOR2_X1 U22140 ( .A1(n19146), .A2(n19145), .ZN(n19156) );
  INV_X1 U22141 ( .A(n19156), .ZN(n19154) );
  NOR2_X1 U22142 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19154), .ZN(n19149) );
  INV_X1 U22143 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19147) );
  AOI22_X1 U22144 ( .A1(n19149), .A2(n19315), .B1(n19154), .B2(n19147), .ZN(
        P2_U2820) );
  OR3_X1 U22145 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19153) );
  INV_X1 U22146 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19148) );
  AOI22_X1 U22147 ( .A1(n19149), .A2(n19153), .B1(n19154), .B2(n19148), .ZN(
        P2_U2821) );
  INV_X1 U22148 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20172) );
  NAND2_X1 U22149 ( .A1(n19149), .A2(n20172), .ZN(n19152) );
  OAI21_X1 U22150 ( .B1(n20121), .B2(n19315), .A(n19156), .ZN(n19150) );
  OAI21_X1 U22151 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19156), .A(n19150), 
        .ZN(n19151) );
  OAI221_X1 U22152 ( .B1(n19152), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19152), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19151), .ZN(P2_U2822) );
  INV_X1 U22153 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19155) );
  OAI221_X1 U22154 ( .B1(n19156), .B2(n19155), .C1(n19154), .C2(n19153), .A(
        n19152), .ZN(P2_U2823) );
  AOI211_X1 U22155 ( .C1(n19159), .C2(n19157), .A(n19158), .B(n20099), .ZN(
        n19160) );
  INV_X1 U22156 ( .A(n19160), .ZN(n19170) );
  AOI22_X1 U22157 ( .A1(n19320), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n19318), .ZN(n19169) );
  OAI22_X1 U22158 ( .A1(n19161), .A2(n19300), .B1(n19326), .B2(n10763), .ZN(
        n19162) );
  INV_X1 U22159 ( .A(n19162), .ZN(n19168) );
  INV_X1 U22160 ( .A(n19163), .ZN(n19164) );
  OAI22_X1 U22161 ( .A1(n19165), .A2(n19292), .B1(n19312), .B2(n19164), .ZN(
        n19166) );
  INV_X1 U22162 ( .A(n19166), .ZN(n19167) );
  NAND4_X1 U22163 ( .A1(n19170), .A2(n19169), .A3(n19168), .A4(n19167), .ZN(
        P2_U2834) );
  INV_X1 U22164 ( .A(n19171), .ZN(n19172) );
  AOI22_X1 U22165 ( .A1(n19173), .A2(n19313), .B1(n19319), .B2(n19172), .ZN(
        n19182) );
  AOI211_X1 U22166 ( .C1(n19176), .C2(n19175), .A(n19174), .B(n20099), .ZN(
        n19180) );
  AOI22_X1 U22167 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19318), .ZN(n19177) );
  OAI21_X1 U22168 ( .B1(n19178), .B2(n19300), .A(n19177), .ZN(n19179) );
  AOI211_X1 U22169 ( .C1(P2_EBX_REG_20__SCAN_IN), .C2(n19320), .A(n19180), .B(
        n19179), .ZN(n19181) );
  NAND2_X1 U22170 ( .A1(n19182), .A2(n19181), .ZN(P2_U2835) );
  INV_X1 U22171 ( .A(n19183), .ZN(n19184) );
  NOR2_X1 U22172 ( .A1(n19186), .A2(n19184), .ZN(n19185) );
  AOI211_X1 U22173 ( .C1(n19186), .C2(n19184), .A(n19185), .B(n20099), .ZN(
        n19195) );
  OAI22_X1 U22174 ( .A1(n19188), .A2(n19300), .B1(n19326), .B2(n19187), .ZN(
        n19189) );
  AOI211_X1 U22175 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19320), .A(n19303), .B(
        n19189), .ZN(n19190) );
  OAI21_X1 U22176 ( .B1(n10759), .B2(n19260), .A(n19190), .ZN(n19191) );
  INV_X1 U22177 ( .A(n19191), .ZN(n19192) );
  OAI21_X1 U22178 ( .B1(n19193), .B2(n19292), .A(n19192), .ZN(n19194) );
  NOR2_X1 U22179 ( .A1(n19195), .A2(n19194), .ZN(n19196) );
  OAI21_X1 U22180 ( .B1(n19197), .B2(n19312), .A(n19196), .ZN(P2_U2836) );
  AOI211_X1 U22181 ( .C1(n19200), .C2(n19199), .A(n19198), .B(n20099), .ZN(
        n19209) );
  NAND2_X1 U22182 ( .A1(n19201), .A2(n19317), .ZN(n19207) );
  NAND2_X1 U22183 ( .A1(n19318), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n19203) );
  AOI22_X1 U22184 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n19320), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19298), .ZN(n19202) );
  NAND3_X1 U22185 ( .A1(n19203), .A2(n19202), .A3(n19277), .ZN(n19204) );
  AOI21_X1 U22186 ( .B1(n19205), .B2(n19313), .A(n19204), .ZN(n19206) );
  NAND2_X1 U22187 ( .A1(n19207), .A2(n19206), .ZN(n19208) );
  NOR2_X1 U22188 ( .A1(n19209), .A2(n19208), .ZN(n19210) );
  OAI21_X1 U22189 ( .B1(n19211), .B2(n19312), .A(n19210), .ZN(P2_U2837) );
  OAI22_X1 U22190 ( .A1(n19213), .A2(n19292), .B1(n19312), .B2(n19212), .ZN(
        n19214) );
  INV_X1 U22191 ( .A(n19214), .ZN(n19224) );
  INV_X1 U22192 ( .A(n19325), .ZN(n19245) );
  AOI211_X1 U22193 ( .C1(n19222), .C2(n19216), .A(n19215), .B(n19331), .ZN(
        n19221) );
  OAI22_X1 U22194 ( .A1(n15817), .A2(n19326), .B1(n20143), .B2(n19260), .ZN(
        n19217) );
  AOI211_X1 U22195 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19320), .A(n19303), .B(
        n19217), .ZN(n19218) );
  OAI21_X1 U22196 ( .B1(n19219), .B2(n19300), .A(n19218), .ZN(n19220) );
  AOI211_X1 U22197 ( .C1(n19222), .C2(n19245), .A(n19221), .B(n19220), .ZN(
        n19223) );
  NAND2_X1 U22198 ( .A1(n19224), .A2(n19223), .ZN(P2_U2838) );
  NOR2_X1 U22199 ( .A1(n19289), .A2(n19237), .ZN(n19226) );
  XOR2_X1 U22200 ( .A(n19226), .B(n19225), .Z(n19236) );
  INV_X1 U22201 ( .A(n19227), .ZN(n19229) );
  AOI22_X1 U22202 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19318), .ZN(n19228) );
  OAI21_X1 U22203 ( .B1(n19229), .B2(n19300), .A(n19228), .ZN(n19230) );
  AOI211_X1 U22204 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n19320), .A(n19303), .B(
        n19230), .ZN(n19235) );
  INV_X1 U22205 ( .A(n19231), .ZN(n19352) );
  OAI22_X1 U22206 ( .A1(n19232), .A2(n19292), .B1(n19312), .B2(n19352), .ZN(
        n19233) );
  INV_X1 U22207 ( .A(n19233), .ZN(n19234) );
  OAI211_X1 U22208 ( .C1(n20099), .C2(n19236), .A(n19235), .B(n19234), .ZN(
        P2_U2841) );
  AOI211_X1 U22209 ( .C1(n19246), .C2(n19238), .A(n19237), .B(n19331), .ZN(
        n19244) );
  NAND2_X1 U22210 ( .A1(n19239), .A2(n19317), .ZN(n19242) );
  AOI22_X1 U22211 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n19320), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19298), .ZN(n19241) );
  NAND2_X1 U22212 ( .A1(n19318), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n19240) );
  NAND4_X1 U22213 ( .A1(n19242), .A2(n19241), .A3(n19277), .A4(n19240), .ZN(
        n19243) );
  NOR2_X1 U22214 ( .A1(n19244), .A2(n19243), .ZN(n19249) );
  AOI22_X1 U22215 ( .A1(n19247), .A2(n19313), .B1(n19246), .B2(n19245), .ZN(
        n19248) );
  OAI211_X1 U22216 ( .C1(n19312), .C2(n19354), .A(n19249), .B(n19248), .ZN(
        P2_U2842) );
  XNOR2_X1 U22217 ( .A(n19251), .B(n19250), .ZN(n19259) );
  INV_X1 U22218 ( .A(n19252), .ZN(n19253) );
  AOI22_X1 U22219 ( .A1(n19253), .A2(n19317), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19298), .ZN(n19254) );
  OAI211_X1 U22220 ( .C1(n20136), .C2(n19260), .A(n19254), .B(n19277), .ZN(
        n19257) );
  OAI22_X1 U22221 ( .A1(n19357), .A2(n19312), .B1(n19292), .B2(n19255), .ZN(
        n19256) );
  AOI211_X1 U22222 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n19320), .A(n19257), .B(
        n19256), .ZN(n19258) );
  OAI21_X1 U22223 ( .B1(n20099), .B2(n19259), .A(n19258), .ZN(P2_U2843) );
  OAI21_X1 U22224 ( .B1(n20132), .B2(n19260), .A(n19277), .ZN(n19265) );
  INV_X1 U22225 ( .A(n19261), .ZN(n19263) );
  OAI22_X1 U22226 ( .A1(n19263), .A2(n19300), .B1(n19326), .B2(n19262), .ZN(
        n19264) );
  AOI211_X1 U22227 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19320), .A(n19265), .B(
        n19264), .ZN(n19272) );
  NAND2_X1 U22228 ( .A1(n12811), .A2(n19266), .ZN(n19267) );
  XNOR2_X1 U22229 ( .A(n19268), .B(n19267), .ZN(n19270) );
  AOI22_X1 U22230 ( .A1(n19270), .A2(n19308), .B1(n19313), .B2(n19269), .ZN(
        n19271) );
  OAI211_X1 U22231 ( .C1(n19312), .C2(n19364), .A(n19272), .B(n19271), .ZN(
        P2_U2846) );
  NAND2_X1 U22232 ( .A1(n12811), .A2(n19273), .ZN(n19275) );
  XOR2_X1 U22233 ( .A(n19275), .B(n19274), .Z(n19283) );
  AOI22_X1 U22234 ( .A1(n19276), .A2(n19317), .B1(n19318), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n19278) );
  OAI211_X1 U22235 ( .C1(n19285), .C2(n10813), .A(n19278), .B(n19277), .ZN(
        n19281) );
  OAI22_X1 U22236 ( .A1(n19279), .A2(n19292), .B1(n19312), .B2(n19369), .ZN(
        n19280) );
  AOI211_X1 U22237 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19298), .A(
        n19281), .B(n19280), .ZN(n19282) );
  OAI21_X1 U22238 ( .B1(n19283), .B2(n20099), .A(n19282), .ZN(P2_U2848) );
  OAI22_X1 U22239 ( .A1(n19286), .A2(n19300), .B1(n19285), .B2(n19284), .ZN(
        n19287) );
  AOI211_X1 U22240 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n19318), .A(n19303), .B(
        n19287), .ZN(n19297) );
  NOR2_X1 U22241 ( .A1(n19289), .A2(n19288), .ZN(n19290) );
  XNOR2_X1 U22242 ( .A(n19291), .B(n19290), .ZN(n19295) );
  OAI22_X1 U22243 ( .A1(n19293), .A2(n19292), .B1(n19312), .B2(n19370), .ZN(
        n19294) );
  AOI21_X1 U22244 ( .B1(n19295), .B2(n19308), .A(n19294), .ZN(n19296) );
  OAI211_X1 U22245 ( .C1(n10723), .C2(n19326), .A(n19297), .B(n19296), .ZN(
        P2_U2849) );
  AOI22_X1 U22246 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n19318), .ZN(n19299) );
  OAI21_X1 U22247 ( .B1(n19301), .B2(n19300), .A(n19299), .ZN(n19302) );
  AOI211_X1 U22248 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n19320), .A(n19303), .B(
        n19302), .ZN(n19311) );
  NAND2_X1 U22249 ( .A1(n12811), .A2(n19304), .ZN(n19305) );
  XNOR2_X1 U22250 ( .A(n19306), .B(n19305), .ZN(n19309) );
  AOI22_X1 U22251 ( .A1(n19309), .A2(n19308), .B1(n19313), .B2(n19307), .ZN(
        n19310) );
  OAI211_X1 U22252 ( .C1(n19312), .C2(n19378), .A(n19311), .B(n19310), .ZN(
        P2_U2850) );
  NAND2_X1 U22253 ( .A1(n19314), .A2(n19313), .ZN(n19323) );
  AOI22_X1 U22254 ( .A1(n19318), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19317), 
        .B2(n19316), .ZN(n19322) );
  AOI22_X1 U22255 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(n19320), .B1(n19319), .B2(
        n19373), .ZN(n19321) );
  NAND3_X1 U22256 ( .A1(n19323), .A2(n19322), .A3(n19321), .ZN(n19328) );
  INV_X1 U22257 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19324) );
  AOI21_X1 U22258 ( .B1(n19326), .B2(n19325), .A(n19324), .ZN(n19327) );
  AOI211_X1 U22259 ( .C1(n19329), .C2(n19784), .A(n19328), .B(n19327), .ZN(
        n19330) );
  OAI21_X1 U22260 ( .B1(n19332), .B2(n19331), .A(n19330), .ZN(P2_U2855) );
  INV_X1 U22261 ( .A(n19333), .ZN(n19334) );
  AOI22_X1 U22262 ( .A1(n19334), .A2(n19400), .B1(n19340), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19336) );
  AOI22_X1 U22263 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19399), .B1(n19339), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19335) );
  NAND2_X1 U22264 ( .A1(n19336), .A2(n19335), .ZN(P2_U2888) );
  AOI22_X1 U22265 ( .A1(n19338), .A2(n19337), .B1(n19399), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19347) );
  AOI22_X1 U22266 ( .A1(n19340), .A2(BUF2_REG_16__SCAN_IN), .B1(n19339), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19346) );
  NOR2_X1 U22267 ( .A1(n19342), .A2(n19341), .ZN(n19343) );
  AOI21_X1 U22268 ( .B1(n19344), .B2(n19404), .A(n19343), .ZN(n19345) );
  NAND3_X1 U22269 ( .A1(n19347), .A2(n19346), .A3(n19345), .ZN(P2_U2903) );
  OAI222_X1 U22270 ( .A1(n19349), .A2(n19379), .B1(n12945), .B2(n19371), .C1(
        n19348), .C2(n19408), .ZN(P2_U2904) );
  AOI22_X1 U22271 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19399), .B1(n19350), 
        .B2(n19365), .ZN(n19351) );
  OAI21_X1 U22272 ( .B1(n19379), .B2(n19352), .A(n19351), .ZN(P2_U2905) );
  INV_X1 U22273 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19452) );
  OAI222_X1 U22274 ( .A1(n19354), .A2(n19379), .B1(n19452), .B2(n19371), .C1(
        n19408), .C2(n19353), .ZN(P2_U2906) );
  AOI22_X1 U22275 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19399), .B1(n19355), 
        .B2(n19365), .ZN(n19356) );
  OAI21_X1 U22276 ( .B1(n19379), .B2(n19357), .A(n19356), .ZN(P2_U2907) );
  OAI222_X1 U22277 ( .A1(n19359), .A2(n19379), .B1(n12856), .B2(n19371), .C1(
        n19408), .C2(n19358), .ZN(P2_U2908) );
  AOI22_X1 U22278 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19399), .B1(n19360), 
        .B2(n19365), .ZN(n19361) );
  OAI21_X1 U22279 ( .B1(n19379), .B2(n19362), .A(n19361), .ZN(P2_U2909) );
  OAI222_X1 U22280 ( .A1(n19364), .A2(n19379), .B1(n12892), .B2(n19371), .C1(
        n19408), .C2(n19363), .ZN(P2_U2910) );
  AOI22_X1 U22281 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19399), .B1(n19366), .B2(
        n19365), .ZN(n19367) );
  OAI21_X1 U22282 ( .B1(n19379), .B2(n19368), .A(n19367), .ZN(P2_U2911) );
  INV_X1 U22283 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19464) );
  OAI222_X1 U22284 ( .A1(n19369), .A2(n19379), .B1(n19464), .B2(n19371), .C1(
        n19408), .C2(n19567), .ZN(P2_U2912) );
  INV_X1 U22285 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19466) );
  OAI222_X1 U22286 ( .A1(n19370), .A2(n19379), .B1(n19466), .B2(n19371), .C1(
        n19408), .C2(n19560), .ZN(P2_U2913) );
  INV_X1 U22287 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19468) );
  OAI22_X1 U22288 ( .A1(n19468), .A2(n19371), .B1(n19553), .B2(n19408), .ZN(
        n19372) );
  INV_X1 U22289 ( .A(n19372), .ZN(n19377) );
  XNOR2_X1 U22290 ( .A(n19520), .B(n20188), .ZN(n19395) );
  XNOR2_X1 U22291 ( .A(n19657), .B(n20197), .ZN(n19403) );
  NAND2_X1 U22292 ( .A1(n19784), .A2(n19373), .ZN(n19402) );
  NAND2_X1 U22293 ( .A1(n19403), .A2(n19402), .ZN(n19401) );
  OAI21_X1 U22294 ( .B1(n20197), .B2(n20193), .A(n19401), .ZN(n19394) );
  NAND2_X1 U22295 ( .A1(n19395), .A2(n19394), .ZN(n19393) );
  OAI21_X1 U22296 ( .B1(n20184), .B2(n20188), .A(n19393), .ZN(n19388) );
  XNOR2_X1 U22297 ( .A(n20177), .B(n20180), .ZN(n19389) );
  NAND2_X1 U22298 ( .A1(n19388), .A2(n19389), .ZN(n19387) );
  OAI21_X1 U22299 ( .B1(n20180), .B2(n19521), .A(n19387), .ZN(n19374) );
  NAND2_X1 U22300 ( .A1(n19374), .A2(n19380), .ZN(n19383) );
  INV_X1 U22301 ( .A(n19382), .ZN(n19375) );
  NAND3_X1 U22302 ( .A1(n19383), .A2(n19375), .A3(n19404), .ZN(n19376) );
  OAI211_X1 U22303 ( .C1(n19379), .C2(n19378), .A(n19377), .B(n19376), .ZN(
        P2_U2914) );
  INV_X1 U22304 ( .A(n19380), .ZN(n19381) );
  AOI22_X1 U22305 ( .A1(n19400), .A2(n19381), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19399), .ZN(n19386) );
  XNOR2_X1 U22306 ( .A(n19383), .B(n19382), .ZN(n19384) );
  NAND2_X1 U22307 ( .A1(n19384), .A2(n19404), .ZN(n19385) );
  OAI211_X1 U22308 ( .C1(n19550), .C2(n19408), .A(n19386), .B(n19385), .ZN(
        P2_U2915) );
  AOI22_X1 U22309 ( .A1(n19400), .A2(n20180), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19399), .ZN(n19392) );
  OAI21_X1 U22310 ( .B1(n19389), .B2(n19388), .A(n19387), .ZN(n19390) );
  NAND2_X1 U22311 ( .A1(n19390), .A2(n19404), .ZN(n19391) );
  OAI211_X1 U22312 ( .C1(n19546), .C2(n19408), .A(n19392), .B(n19391), .ZN(
        P2_U2916) );
  AOI22_X1 U22313 ( .A1(n19400), .A2(n20188), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19399), .ZN(n19398) );
  OAI21_X1 U22314 ( .B1(n19395), .B2(n19394), .A(n19393), .ZN(n19396) );
  NAND2_X1 U22315 ( .A1(n19396), .A2(n19404), .ZN(n19397) );
  OAI211_X1 U22316 ( .C1(n19540), .C2(n19408), .A(n19398), .B(n19397), .ZN(
        P2_U2917) );
  AOI22_X1 U22317 ( .A1(n19400), .A2(n20197), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19399), .ZN(n19407) );
  OAI21_X1 U22318 ( .B1(n19403), .B2(n19402), .A(n19401), .ZN(n19405) );
  NAND2_X1 U22319 ( .A1(n19405), .A2(n19404), .ZN(n19406) );
  OAI211_X1 U22320 ( .C1(n19536), .C2(n19408), .A(n19407), .B(n19406), .ZN(
        P2_U2918) );
  NAND2_X1 U22321 ( .A1(n19409), .A2(n20095), .ZN(n19411) );
  OAI21_X1 U22322 ( .B1(n19412), .B2(n19411), .A(n19410), .ZN(n19414) );
  INV_X1 U22323 ( .A(n20227), .ZN(n19413) );
  NOR2_X1 U22324 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20200), .ZN(n19440) );
  CLKBUF_X1 U22325 ( .A(n19440), .Z(n20223) );
  NOR2_X1 U22326 ( .A1(n19459), .A2(n19415), .ZN(P2_U2920) );
  NAND2_X1 U22327 ( .A1(n19456), .A2(n19416), .ZN(n19446) );
  INV_X2 U22328 ( .A(n19459), .ZN(n19476) );
  AOI22_X1 U22329 ( .A1(n20223), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n19417) );
  OAI21_X1 U22330 ( .B1(n19418), .B2(n19446), .A(n19417), .ZN(P2_U2921) );
  AOI22_X1 U22331 ( .A1(n20223), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19419) );
  OAI21_X1 U22332 ( .B1(n19420), .B2(n19446), .A(n19419), .ZN(P2_U2922) );
  AOI22_X1 U22333 ( .A1(n20223), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19421) );
  OAI21_X1 U22334 ( .B1(n21198), .B2(n19446), .A(n19421), .ZN(P2_U2923) );
  AOI22_X1 U22335 ( .A1(n19440), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19422) );
  OAI21_X1 U22336 ( .B1(n19423), .B2(n19446), .A(n19422), .ZN(P2_U2924) );
  AOI22_X1 U22337 ( .A1(n19440), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19424) );
  OAI21_X1 U22338 ( .B1(n19425), .B2(n19446), .A(n19424), .ZN(P2_U2925) );
  AOI22_X1 U22339 ( .A1(n19440), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19426) );
  OAI21_X1 U22340 ( .B1(n19427), .B2(n19446), .A(n19426), .ZN(P2_U2926) );
  AOI22_X1 U22341 ( .A1(n19440), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19428) );
  OAI21_X1 U22342 ( .B1(n19429), .B2(n19446), .A(n19428), .ZN(P2_U2927) );
  INV_X1 U22343 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19431) );
  AOI22_X1 U22344 ( .A1(n19440), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19430) );
  OAI21_X1 U22345 ( .B1(n19431), .B2(n19446), .A(n19430), .ZN(P2_U2928) );
  INV_X1 U22346 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19433) );
  AOI22_X1 U22347 ( .A1(n19440), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19432) );
  OAI21_X1 U22348 ( .B1(n19433), .B2(n19446), .A(n19432), .ZN(P2_U2929) );
  AOI22_X1 U22349 ( .A1(n19440), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19434) );
  OAI21_X1 U22350 ( .B1(n19435), .B2(n19446), .A(n19434), .ZN(P2_U2930) );
  INV_X1 U22351 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19437) );
  AOI22_X1 U22352 ( .A1(n19440), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19436) );
  OAI21_X1 U22353 ( .B1(n19437), .B2(n19446), .A(n19436), .ZN(P2_U2931) );
  INV_X1 U22354 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19439) );
  AOI22_X1 U22355 ( .A1(n19440), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19438) );
  OAI21_X1 U22356 ( .B1(n19439), .B2(n19446), .A(n19438), .ZN(P2_U2932) );
  INV_X1 U22357 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19442) );
  AOI22_X1 U22358 ( .A1(n19440), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19441) );
  OAI21_X1 U22359 ( .B1(n19442), .B2(n19446), .A(n19441), .ZN(P2_U2933) );
  AOI22_X1 U22360 ( .A1(n20223), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19443) );
  OAI21_X1 U22361 ( .B1(n19444), .B2(n19446), .A(n19443), .ZN(P2_U2934) );
  INV_X1 U22362 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19447) );
  AOI22_X1 U22363 ( .A1(n20223), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19445) );
  OAI21_X1 U22364 ( .B1(n19447), .B2(n19446), .A(n19445), .ZN(P2_U2935) );
  AOI22_X1 U22365 ( .A1(n20223), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19448) );
  OAI21_X1 U22366 ( .B1(n12945), .B2(n19478), .A(n19448), .ZN(P2_U2936) );
  AOI22_X1 U22367 ( .A1(n20223), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19449) );
  OAI21_X1 U22368 ( .B1(n19450), .B2(n19478), .A(n19449), .ZN(P2_U2937) );
  AOI22_X1 U22369 ( .A1(n20223), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19451) );
  OAI21_X1 U22370 ( .B1(n19452), .B2(n19478), .A(n19451), .ZN(P2_U2938) );
  AOI22_X1 U22371 ( .A1(n20223), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19453) );
  OAI21_X1 U22372 ( .B1(n19454), .B2(n19478), .A(n19453), .ZN(P2_U2939) );
  AOI22_X1 U22373 ( .A1(n20223), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19455) );
  OAI21_X1 U22374 ( .B1(n12856), .B2(n19478), .A(n19455), .ZN(P2_U2940) );
  AOI22_X1 U22375 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19456), .B1(n20223), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n19457) );
  OAI21_X1 U22376 ( .B1(n19459), .B2(n19458), .A(n19457), .ZN(P2_U2941) );
  AOI22_X1 U22377 ( .A1(n20223), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19460) );
  OAI21_X1 U22378 ( .B1(n12892), .B2(n19478), .A(n19460), .ZN(P2_U2942) );
  AOI22_X1 U22379 ( .A1(n20223), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19461) );
  OAI21_X1 U22380 ( .B1(n19462), .B2(n19478), .A(n19461), .ZN(P2_U2943) );
  AOI22_X1 U22381 ( .A1(n20223), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19463) );
  OAI21_X1 U22382 ( .B1(n19464), .B2(n19478), .A(n19463), .ZN(P2_U2944) );
  AOI22_X1 U22383 ( .A1(n20223), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19465) );
  OAI21_X1 U22384 ( .B1(n19466), .B2(n19478), .A(n19465), .ZN(P2_U2945) );
  AOI22_X1 U22385 ( .A1(n20223), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19467) );
  OAI21_X1 U22386 ( .B1(n19468), .B2(n19478), .A(n19467), .ZN(P2_U2946) );
  INV_X1 U22387 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19470) );
  AOI22_X1 U22388 ( .A1(n20223), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19469) );
  OAI21_X1 U22389 ( .B1(n19470), .B2(n19478), .A(n19469), .ZN(P2_U2947) );
  INV_X1 U22390 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19472) );
  AOI22_X1 U22391 ( .A1(n20223), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19471) );
  OAI21_X1 U22392 ( .B1(n19472), .B2(n19478), .A(n19471), .ZN(P2_U2948) );
  INV_X1 U22393 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19474) );
  AOI22_X1 U22394 ( .A1(n20223), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19473) );
  OAI21_X1 U22395 ( .B1(n19474), .B2(n19478), .A(n19473), .ZN(P2_U2949) );
  AOI22_X1 U22396 ( .A1(n20223), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19475) );
  OAI21_X1 U22397 ( .B1(n12895), .B2(n19478), .A(n19475), .ZN(P2_U2950) );
  INV_X1 U22398 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19479) );
  AOI22_X1 U22399 ( .A1(n20223), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19476), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19477) );
  OAI21_X1 U22400 ( .B1(n19479), .B2(n19478), .A(n19477), .ZN(P2_U2951) );
  AOI22_X1 U22401 ( .A1(n19481), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19480), 
        .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n19483) );
  NAND2_X1 U22402 ( .A1(n19483), .A2(n19482), .ZN(P2_U2977) );
  AOI22_X1 U22403 ( .A1(n19484), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19303), .ZN(n19494) );
  NAND2_X1 U22404 ( .A1(n19485), .A2(n10990), .ZN(n19489) );
  NAND2_X1 U22405 ( .A1(n19487), .A2(n19486), .ZN(n19488) );
  OAI211_X1 U22406 ( .C1(n19491), .C2(n19490), .A(n19489), .B(n19488), .ZN(
        n19492) );
  INV_X1 U22407 ( .A(n19492), .ZN(n19493) );
  OAI211_X1 U22408 ( .C1(n19496), .C2(n19495), .A(n19494), .B(n19493), .ZN(
        P2_U3010) );
  AOI22_X1 U22409 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19500), .B2(n19497), .ZN(
        n19498) );
  NAND2_X1 U22410 ( .A1(n19499), .A2(n19498), .ZN(n19512) );
  OAI22_X1 U22411 ( .A1(n19503), .A2(n19502), .B1(n19501), .B2(n19500), .ZN(
        n19504) );
  INV_X1 U22412 ( .A(n19504), .ZN(n19511) );
  NAND2_X1 U22413 ( .A1(n19506), .A2(n19505), .ZN(n19510) );
  INV_X1 U22414 ( .A(n20197), .ZN(n19507) );
  OR2_X1 U22415 ( .A1(n19508), .A2(n19507), .ZN(n19509) );
  AND4_X1 U22416 ( .A1(n19512), .A2(n19511), .A3(n19510), .A4(n19509), .ZN(
        n19514) );
  OAI211_X1 U22417 ( .C1(n19516), .C2(n19515), .A(n19514), .B(n19513), .ZN(
        P2_U3045) );
  AOI22_X1 U22418 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19563), .ZN(n20001) );
  AOI22_X1 U22419 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19563), .ZN(n20045) );
  NOR2_X2 U22420 ( .A1(n13056), .A2(n19565), .ZN(n20033) );
  NAND3_X1 U22421 ( .A1(n20199), .A2(n20208), .A3(n19626), .ZN(n19524) );
  INV_X1 U22422 ( .A(n19524), .ZN(n19566) );
  AOI22_X1 U22423 ( .A1(n19988), .A2(n20061), .B1(n20033), .B2(n19566), .ZN(
        n19533) );
  INV_X1 U22424 ( .A(n19597), .ZN(n19522) );
  OAI21_X1 U22425 ( .B1(n20061), .B2(n19522), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19523) );
  NAND2_X1 U22426 ( .A1(n19523), .A2(n19989), .ZN(n19531) );
  NOR2_X1 U22427 ( .A1(n20085), .A2(n19566), .ZN(n19530) );
  INV_X1 U22428 ( .A(n19530), .ZN(n19526) );
  OAI211_X1 U22429 ( .C1(n10551), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19524), 
        .B(n20183), .ZN(n19525) );
  OAI211_X1 U22430 ( .C1(n19531), .C2(n19526), .A(n20039), .B(n19525), .ZN(
        n19569) );
  NOR2_X2 U22431 ( .A1(n19527), .A2(n19956), .ZN(n20034) );
  INV_X1 U22432 ( .A(n10551), .ZN(n19528) );
  OAI21_X1 U22433 ( .B1(n19528), .B2(n19566), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19529) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19569), .B1(
        n20034), .B2(n19568), .ZN(n19532) );
  OAI211_X1 U22435 ( .C1(n20001), .C2(n19597), .A(n19533), .B(n19532), .ZN(
        P2_U3048) );
  AOI22_X1 U22436 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19563), .ZN(n19935) );
  AOI22_X1 U22437 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19563), .ZN(n20051) );
  INV_X1 U22438 ( .A(n19565), .ZN(n19534) );
  AND2_X1 U22439 ( .A1(n9676), .A2(n19534), .ZN(n20046) );
  AOI22_X1 U22440 ( .A1(n19932), .A2(n20061), .B1(n20046), .B2(n19566), .ZN(
        n19538) );
  NOR2_X2 U22441 ( .A1(n19536), .A2(n19956), .ZN(n20047) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19569), .B1(
        n20047), .B2(n19568), .ZN(n19537) );
  OAI211_X1 U22443 ( .C1(n19935), .C2(n19597), .A(n19538), .B(n19537), .ZN(
        P2_U3049) );
  AOI22_X1 U22444 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19563), .ZN(n20007) );
  AOI22_X1 U22445 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19563), .ZN(n20057) );
  NOR2_X2 U22446 ( .A1(n19539), .A2(n19565), .ZN(n20052) );
  AOI22_X1 U22447 ( .A1(n20004), .A2(n20061), .B1(n20052), .B2(n19566), .ZN(
        n19542) );
  NOR2_X2 U22448 ( .A1(n19540), .A2(n19956), .ZN(n20053) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19569), .B1(
        n20053), .B2(n19568), .ZN(n19541) );
  OAI211_X1 U22450 ( .C1(n20007), .C2(n19597), .A(n19542), .B(n19541), .ZN(
        P2_U3050) );
  INV_X1 U22451 ( .A(n19564), .ZN(n19558) );
  INV_X1 U22452 ( .A(n19563), .ZN(n19556) );
  INV_X1 U22453 ( .A(n20060), .ZN(n20011) );
  AOI22_X1 U22454 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19563), .ZN(n20065) );
  NOR2_X2 U22455 ( .A1(n19545), .A2(n19565), .ZN(n20058) );
  AOI22_X1 U22456 ( .A1(n20008), .A2(n20061), .B1(n20058), .B2(n19566), .ZN(
        n19548) );
  NOR2_X2 U22457 ( .A1(n19546), .A2(n19956), .ZN(n20059) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19569), .B1(
        n20059), .B2(n19568), .ZN(n19547) );
  OAI211_X1 U22459 ( .C1(n20011), .C2(n19597), .A(n19548), .B(n19547), .ZN(
        P2_U3051) );
  AOI22_X1 U22460 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19563), .ZN(n20071) );
  AOI22_X1 U22461 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19563), .ZN(n19974) );
  NOR2_X2 U22462 ( .A1(n19549), .A2(n19565), .ZN(n20066) );
  AOI22_X1 U22463 ( .A1(n20068), .A2(n20061), .B1(n20066), .B2(n19566), .ZN(
        n19552) );
  NOR2_X2 U22464 ( .A1(n19550), .A2(n19956), .ZN(n20067) );
  AOI22_X1 U22465 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19569), .B1(
        n20067), .B2(n19568), .ZN(n19551) );
  OAI211_X1 U22466 ( .C1(n20071), .C2(n19597), .A(n19552), .B(n19551), .ZN(
        P2_U3052) );
  AOI22_X1 U22467 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19563), .ZN(n19978) );
  NOR2_X2 U22468 ( .A1(n10812), .A2(n19565), .ZN(n20072) );
  AOI22_X1 U22469 ( .A1(n20061), .A2(n20074), .B1(n20072), .B2(n19566), .ZN(
        n19555) );
  NOR2_X2 U22470 ( .A1(n19553), .A2(n19956), .ZN(n20073) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19569), .B1(
        n20073), .B2(n19568), .ZN(n19554) );
  OAI211_X1 U22472 ( .C1(n20077), .C2(n19597), .A(n19555), .B(n19554), .ZN(
        P2_U3053) );
  INV_X1 U22473 ( .A(n20017), .ZN(n20083) );
  AOI22_X1 U22474 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19563), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19564), .ZN(n20020) );
  NOR2_X2 U22475 ( .A1(n10300), .A2(n19565), .ZN(n20078) );
  AOI22_X1 U22476 ( .A1(n20080), .A2(n20061), .B1(n20078), .B2(n19566), .ZN(
        n19562) );
  NOR2_X2 U22477 ( .A1(n19560), .A2(n19956), .ZN(n20079) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19569), .B1(
        n20079), .B2(n19568), .ZN(n19561) );
  OAI211_X1 U22479 ( .C1(n20083), .C2(n19597), .A(n19562), .B(n19561), .ZN(
        P2_U3054) );
  AOI22_X1 U22480 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19563), .ZN(n20094) );
  AOI22_X1 U22481 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19564), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19563), .ZN(n20028) );
  NOR2_X2 U22482 ( .A1(n10322), .A2(n19565), .ZN(n20084) );
  AOI22_X1 U22483 ( .A1(n20088), .A2(n20061), .B1(n20084), .B2(n19566), .ZN(
        n19571) );
  NOR2_X2 U22484 ( .A1(n19567), .A2(n19956), .ZN(n20086) );
  AOI22_X1 U22485 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19569), .B1(
        n20086), .B2(n19568), .ZN(n19570) );
  OAI211_X1 U22486 ( .C1(n20094), .C2(n19597), .A(n19571), .B(n19570), .ZN(
        P2_U3055) );
  NAND2_X1 U22487 ( .A1(n19626), .A2(n20199), .ZN(n19575) );
  INV_X1 U22488 ( .A(n19572), .ZN(n19573) );
  NAND2_X1 U22489 ( .A1(n20199), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19824) );
  NOR2_X1 U22490 ( .A1(n19824), .A2(n19625), .ZN(n19592) );
  NOR3_X1 U22491 ( .A1(n19573), .A2(n19592), .A3(n19953), .ZN(n19574) );
  AOI211_X2 U22492 ( .C1(n19575), .C2(n19953), .A(n19758), .B(n19574), .ZN(
        n19593) );
  AOI22_X1 U22493 ( .A1(n19593), .A2(n20034), .B1(n20033), .B2(n19592), .ZN(
        n19579) );
  INV_X1 U22494 ( .A(n19831), .ZN(n19822) );
  NAND2_X1 U22495 ( .A1(n19822), .A2(n19749), .ZN(n19576) );
  AOI21_X1 U22496 ( .B1(n19576), .B2(n19575), .A(n19574), .ZN(n19577) );
  OAI211_X1 U22497 ( .C1(n19592), .C2(n20041), .A(n19577), .B(n20039), .ZN(
        n19594) );
  NOR2_X2 U22498 ( .A1(n19831), .A2(n19760), .ZN(n19621) );
  INV_X1 U22499 ( .A(n20001), .ZN(n20042) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19594), .B1(
        n19621), .B2(n20042), .ZN(n19578) );
  OAI211_X1 U22501 ( .C1(n20045), .C2(n19597), .A(n19579), .B(n19578), .ZN(
        P2_U3056) );
  AOI22_X1 U22502 ( .A1(n19593), .A2(n20047), .B1(n20046), .B2(n19592), .ZN(
        n19581) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19594), .B1(
        n19621), .B2(n20048), .ZN(n19580) );
  OAI211_X1 U22504 ( .C1(n20051), .C2(n19597), .A(n19581), .B(n19580), .ZN(
        P2_U3057) );
  AOI22_X1 U22505 ( .A1(n19593), .A2(n20053), .B1(n20052), .B2(n19592), .ZN(
        n19583) );
  INV_X1 U22506 ( .A(n20007), .ZN(n20054) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19594), .B1(
        n19621), .B2(n20054), .ZN(n19582) );
  OAI211_X1 U22508 ( .C1(n20057), .C2(n19597), .A(n19583), .B(n19582), .ZN(
        P2_U3058) );
  AOI22_X1 U22509 ( .A1(n19593), .A2(n20059), .B1(n20058), .B2(n19592), .ZN(
        n19585) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19594), .B1(
        n19621), .B2(n20060), .ZN(n19584) );
  OAI211_X1 U22511 ( .C1(n20065), .C2(n19597), .A(n19585), .B(n19584), .ZN(
        P2_U3059) );
  AOI22_X1 U22512 ( .A1(n19593), .A2(n20067), .B1(n20066), .B2(n19592), .ZN(
        n19587) );
  INV_X1 U22513 ( .A(n20071), .ZN(n19971) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19594), .B1(
        n19621), .B2(n19971), .ZN(n19586) );
  OAI211_X1 U22515 ( .C1(n19974), .C2(n19597), .A(n19587), .B(n19586), .ZN(
        P2_U3060) );
  AOI22_X1 U22516 ( .A1(n19593), .A2(n20073), .B1(n20072), .B2(n19592), .ZN(
        n19589) );
  INV_X1 U22517 ( .A(n20077), .ZN(n19975) );
  AOI22_X1 U22518 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19594), .B1(
        n19621), .B2(n19975), .ZN(n19588) );
  OAI211_X1 U22519 ( .C1(n19978), .C2(n19597), .A(n19589), .B(n19588), .ZN(
        P2_U3061) );
  AOI22_X1 U22520 ( .A1(n19593), .A2(n20079), .B1(n20078), .B2(n19592), .ZN(
        n19591) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19594), .B1(
        n19621), .B2(n20017), .ZN(n19590) );
  OAI211_X1 U22522 ( .C1(n20020), .C2(n19597), .A(n19591), .B(n19590), .ZN(
        P2_U3062) );
  AOI22_X1 U22523 ( .A1(n19593), .A2(n20086), .B1(n20084), .B2(n19592), .ZN(
        n19596) );
  INV_X1 U22524 ( .A(n20094), .ZN(n20022) );
  AOI22_X1 U22525 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19594), .B1(
        n19621), .B2(n20022), .ZN(n19595) );
  OAI211_X1 U22526 ( .C1(n20028), .C2(n19597), .A(n19596), .B(n19595), .ZN(
        P2_U3063) );
  OR2_X1 U22527 ( .A1(n19625), .A2(n19659), .ZN(n19602) );
  INV_X1 U22528 ( .A(n19600), .ZN(n19598) );
  NAND2_X1 U22529 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20208), .ZN(
        n19858) );
  NOR2_X1 U22530 ( .A1(n19858), .A2(n19625), .ZN(n19619) );
  OAI21_X1 U22531 ( .B1(n19598), .B2(n19619), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19599) );
  OAI21_X1 U22532 ( .B1(n19602), .B2(n20183), .A(n19599), .ZN(n19620) );
  AOI22_X1 U22533 ( .A1(n19620), .A2(n20034), .B1(n20033), .B2(n19619), .ZN(
        n19606) );
  AOI21_X1 U22534 ( .B1(n19600), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19604) );
  OAI21_X1 U22535 ( .B1(n19621), .B2(n19647), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19601) );
  NAND2_X1 U22536 ( .A1(n19602), .A2(n19601), .ZN(n19603) );
  OAI211_X1 U22537 ( .C1(n19619), .C2(n19604), .A(n19603), .B(n20039), .ZN(
        n19622) );
  AOI22_X1 U22538 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19622), .B1(
        n19621), .B2(n19988), .ZN(n19605) );
  OAI211_X1 U22539 ( .C1(n20001), .C2(n19656), .A(n19606), .B(n19605), .ZN(
        P2_U3064) );
  AOI22_X1 U22540 ( .A1(n19620), .A2(n20047), .B1(n20046), .B2(n19619), .ZN(
        n19608) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19622), .B1(
        n19621), .B2(n19932), .ZN(n19607) );
  OAI211_X1 U22542 ( .C1(n19935), .C2(n19656), .A(n19608), .B(n19607), .ZN(
        P2_U3065) );
  AOI22_X1 U22543 ( .A1(n19620), .A2(n20053), .B1(n20052), .B2(n19619), .ZN(
        n19610) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19622), .B1(
        n19621), .B2(n20004), .ZN(n19609) );
  OAI211_X1 U22545 ( .C1(n20007), .C2(n19656), .A(n19610), .B(n19609), .ZN(
        P2_U3066) );
  AOI22_X1 U22546 ( .A1(n19620), .A2(n20059), .B1(n20058), .B2(n19619), .ZN(
        n19612) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19622), .B1(
        n19621), .B2(n20008), .ZN(n19611) );
  OAI211_X1 U22548 ( .C1(n20011), .C2(n19656), .A(n19612), .B(n19611), .ZN(
        P2_U3067) );
  AOI22_X1 U22549 ( .A1(n19620), .A2(n20067), .B1(n20066), .B2(n19619), .ZN(
        n19614) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19622), .B1(
        n19621), .B2(n20068), .ZN(n19613) );
  OAI211_X1 U22551 ( .C1(n20071), .C2(n19656), .A(n19614), .B(n19613), .ZN(
        P2_U3068) );
  AOI22_X1 U22552 ( .A1(n19620), .A2(n20073), .B1(n20072), .B2(n19619), .ZN(
        n19616) );
  AOI22_X1 U22553 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19622), .B1(
        n19621), .B2(n20074), .ZN(n19615) );
  OAI211_X1 U22554 ( .C1(n20077), .C2(n19656), .A(n19616), .B(n19615), .ZN(
        P2_U3069) );
  AOI22_X1 U22555 ( .A1(n19620), .A2(n20079), .B1(n20078), .B2(n19619), .ZN(
        n19618) );
  AOI22_X1 U22556 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19622), .B1(
        n19621), .B2(n20080), .ZN(n19617) );
  OAI211_X1 U22557 ( .C1(n20083), .C2(n19656), .A(n19618), .B(n19617), .ZN(
        P2_U3070) );
  AOI22_X1 U22558 ( .A1(n19620), .A2(n20086), .B1(n20084), .B2(n19619), .ZN(
        n19624) );
  AOI22_X1 U22559 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19622), .B1(
        n19621), .B2(n20088), .ZN(n19623) );
  OAI211_X1 U22560 ( .C1(n20094), .C2(n19656), .A(n19624), .B(n19623), .ZN(
        P2_U3071) );
  NOR2_X2 U22561 ( .A1(n19886), .A2(n19760), .ZN(n19683) );
  NOR2_X1 U22562 ( .A1(n19625), .A2(n19888), .ZN(n19651) );
  AOI22_X1 U22563 ( .A1(n20042), .A2(n19683), .B1(n19651), .B2(n20033), .ZN(
        n19636) );
  INV_X1 U22564 ( .A(n19749), .ZN(n19687) );
  OAI21_X1 U22565 ( .B1(n19687), .B2(n19886), .A(n19989), .ZN(n19634) );
  NAND2_X1 U22566 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19626), .ZN(
        n19633) );
  INV_X1 U22567 ( .A(n19633), .ZN(n19629) );
  INV_X1 U22568 ( .A(n19651), .ZN(n19627) );
  OAI211_X1 U22569 ( .C1(n19630), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19627), 
        .B(n20183), .ZN(n19628) );
  OAI211_X1 U22570 ( .C1(n19634), .C2(n19629), .A(n20039), .B(n19628), .ZN(
        n19653) );
  INV_X1 U22571 ( .A(n19630), .ZN(n19631) );
  OAI21_X1 U22572 ( .B1(n19631), .B2(n19651), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19632) );
  OAI21_X1 U22573 ( .B1(n19634), .B2(n19633), .A(n19632), .ZN(n19652) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19653), .B1(
        n20034), .B2(n19652), .ZN(n19635) );
  OAI211_X1 U22575 ( .C1(n20045), .C2(n19656), .A(n19636), .B(n19635), .ZN(
        P2_U3072) );
  INV_X1 U22576 ( .A(n19683), .ZN(n19650) );
  AOI22_X1 U22577 ( .A1(n19647), .A2(n19932), .B1(n19651), .B2(n20046), .ZN(
        n19638) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19653), .B1(
        n20047), .B2(n19652), .ZN(n19637) );
  OAI211_X1 U22579 ( .C1(n19935), .C2(n19650), .A(n19638), .B(n19637), .ZN(
        P2_U3073) );
  AOI22_X1 U22580 ( .A1(n20054), .A2(n19683), .B1(n19651), .B2(n20052), .ZN(
        n19640) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19653), .B1(
        n20053), .B2(n19652), .ZN(n19639) );
  OAI211_X1 U22582 ( .C1(n20057), .C2(n19656), .A(n19640), .B(n19639), .ZN(
        P2_U3074) );
  AOI22_X1 U22583 ( .A1(n20060), .A2(n19683), .B1(n19651), .B2(n20058), .ZN(
        n19642) );
  AOI22_X1 U22584 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19653), .B1(
        n20059), .B2(n19652), .ZN(n19641) );
  OAI211_X1 U22585 ( .C1(n20065), .C2(n19656), .A(n19642), .B(n19641), .ZN(
        P2_U3075) );
  AOI22_X1 U22586 ( .A1(n19971), .A2(n19683), .B1(n19651), .B2(n20066), .ZN(
        n19644) );
  AOI22_X1 U22587 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19653), .B1(
        n20067), .B2(n19652), .ZN(n19643) );
  OAI211_X1 U22588 ( .C1(n19974), .C2(n19656), .A(n19644), .B(n19643), .ZN(
        P2_U3076) );
  AOI22_X1 U22589 ( .A1(n19647), .A2(n20074), .B1(n19651), .B2(n20072), .ZN(
        n19646) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19653), .B1(
        n20073), .B2(n19652), .ZN(n19645) );
  OAI211_X1 U22591 ( .C1(n20077), .C2(n19650), .A(n19646), .B(n19645), .ZN(
        P2_U3077) );
  AOI22_X1 U22592 ( .A1(n19647), .A2(n20080), .B1(n19651), .B2(n20078), .ZN(
        n19649) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19653), .B1(
        n20079), .B2(n19652), .ZN(n19648) );
  OAI211_X1 U22594 ( .C1(n20083), .C2(n19650), .A(n19649), .B(n19648), .ZN(
        P2_U3078) );
  AOI22_X1 U22595 ( .A1(n20022), .A2(n19683), .B1(n19651), .B2(n20084), .ZN(
        n19655) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19653), .B1(
        n20086), .B2(n19652), .ZN(n19654) );
  OAI211_X1 U22597 ( .C1(n20028), .C2(n19656), .A(n19655), .B(n19654), .ZN(
        P2_U3079) );
  INV_X1 U22598 ( .A(n19659), .ZN(n19661) );
  NOR2_X1 U22599 ( .A1(n19661), .A2(n19660), .ZN(n19928) );
  NAND2_X1 U22600 ( .A1(n19928), .A2(n20182), .ZN(n19665) );
  NAND3_X1 U22601 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20182), .A3(
        n20199), .ZN(n19693) );
  NOR2_X1 U22602 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19693), .ZN(
        n19681) );
  OAI21_X1 U22603 ( .B1(n10564), .B2(n19681), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19662) );
  OAI21_X1 U22604 ( .B1(n19665), .B2(n20183), .A(n19662), .ZN(n19682) );
  AOI22_X1 U22605 ( .A1(n19682), .A2(n20034), .B1(n20033), .B2(n19681), .ZN(
        n19668) );
  OAI21_X1 U22606 ( .B1(n19683), .B2(n19705), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19664) );
  AOI211_X1 U22607 ( .C1(n10564), .C2(n20041), .A(n19681), .B(n19989), .ZN(
        n19663) );
  AOI211_X1 U22608 ( .C1(n19665), .C2(n19664), .A(n19956), .B(n19663), .ZN(
        n19666) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n19988), .ZN(n19667) );
  OAI211_X1 U22610 ( .C1(n20001), .C2(n19714), .A(n19668), .B(n19667), .ZN(
        P2_U3080) );
  AOI22_X1 U22611 ( .A1(n19682), .A2(n20047), .B1(n20046), .B2(n19681), .ZN(
        n19670) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n19932), .ZN(n19669) );
  OAI211_X1 U22613 ( .C1(n19935), .C2(n19714), .A(n19670), .B(n19669), .ZN(
        P2_U3081) );
  AOI22_X1 U22614 ( .A1(n19682), .A2(n20053), .B1(n20052), .B2(n19681), .ZN(
        n19672) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n20004), .ZN(n19671) );
  OAI211_X1 U22616 ( .C1(n20007), .C2(n19714), .A(n19672), .B(n19671), .ZN(
        P2_U3082) );
  AOI22_X1 U22617 ( .A1(n19682), .A2(n20059), .B1(n20058), .B2(n19681), .ZN(
        n19674) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n20008), .ZN(n19673) );
  OAI211_X1 U22619 ( .C1(n20011), .C2(n19714), .A(n19674), .B(n19673), .ZN(
        P2_U3083) );
  AOI22_X1 U22620 ( .A1(n19682), .A2(n20067), .B1(n20066), .B2(n19681), .ZN(
        n19676) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n20068), .ZN(n19675) );
  OAI211_X1 U22622 ( .C1(n20071), .C2(n19714), .A(n19676), .B(n19675), .ZN(
        P2_U3084) );
  AOI22_X1 U22623 ( .A1(n19682), .A2(n20073), .B1(n20072), .B2(n19681), .ZN(
        n19678) );
  AOI22_X1 U22624 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n20074), .ZN(n19677) );
  OAI211_X1 U22625 ( .C1(n20077), .C2(n19714), .A(n19678), .B(n19677), .ZN(
        P2_U3085) );
  AOI22_X1 U22626 ( .A1(n19682), .A2(n20079), .B1(n20078), .B2(n19681), .ZN(
        n19680) );
  AOI22_X1 U22627 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n20080), .ZN(n19679) );
  OAI211_X1 U22628 ( .C1(n20083), .C2(n19714), .A(n19680), .B(n19679), .ZN(
        P2_U3086) );
  AOI22_X1 U22629 ( .A1(n19682), .A2(n20086), .B1(n20084), .B2(n19681), .ZN(
        n19686) );
  AOI22_X1 U22630 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19684), .B1(
        n19683), .B2(n20088), .ZN(n19685) );
  OAI211_X1 U22631 ( .C1(n20094), .C2(n19714), .A(n19686), .B(n19685), .ZN(
        P2_U3087) );
  NOR2_X1 U22632 ( .A1(n20208), .A2(n19693), .ZN(n19718) );
  AOI22_X1 U22633 ( .A1(n20042), .A2(n19745), .B1(n19718), .B2(n20033), .ZN(
        n19696) );
  OAI21_X1 U22634 ( .B1(n19687), .B2(n19961), .A(n19989), .ZN(n19694) );
  INV_X1 U22635 ( .A(n19693), .ZN(n19690) );
  INV_X1 U22636 ( .A(n19718), .ZN(n19688) );
  OAI211_X1 U22637 ( .C1(n10546), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19688), 
        .B(n20183), .ZN(n19689) );
  OAI211_X1 U22638 ( .C1(n19694), .C2(n19690), .A(n20039), .B(n19689), .ZN(
        n19711) );
  INV_X1 U22639 ( .A(n10546), .ZN(n19691) );
  OAI21_X1 U22640 ( .B1(n19691), .B2(n19718), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19692) );
  OAI21_X1 U22641 ( .B1(n19694), .B2(n19693), .A(n19692), .ZN(n19710) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19711), .B1(
        n20034), .B2(n19710), .ZN(n19695) );
  OAI211_X1 U22643 ( .C1(n20045), .C2(n19714), .A(n19696), .B(n19695), .ZN(
        P2_U3088) );
  AOI22_X1 U22644 ( .A1(n20048), .A2(n19745), .B1(n19718), .B2(n20046), .ZN(
        n19698) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19711), .B1(
        n20047), .B2(n19710), .ZN(n19697) );
  OAI211_X1 U22646 ( .C1(n20051), .C2(n19714), .A(n19698), .B(n19697), .ZN(
        P2_U3089) );
  AOI22_X1 U22647 ( .A1(n20054), .A2(n19745), .B1(n19718), .B2(n20052), .ZN(
        n19700) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19711), .B1(
        n20053), .B2(n19710), .ZN(n19699) );
  OAI211_X1 U22649 ( .C1(n20057), .C2(n19714), .A(n19700), .B(n19699), .ZN(
        P2_U3090) );
  AOI22_X1 U22650 ( .A1(n20060), .A2(n19745), .B1(n19718), .B2(n20058), .ZN(
        n19702) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19711), .B1(
        n20059), .B2(n19710), .ZN(n19701) );
  OAI211_X1 U22652 ( .C1(n20065), .C2(n19714), .A(n19702), .B(n19701), .ZN(
        P2_U3091) );
  AOI22_X1 U22653 ( .A1(n19705), .A2(n20068), .B1(n20066), .B2(n19718), .ZN(
        n19704) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19711), .B1(
        n20067), .B2(n19710), .ZN(n19703) );
  OAI211_X1 U22655 ( .C1(n20071), .C2(n19738), .A(n19704), .B(n19703), .ZN(
        P2_U3092) );
  AOI22_X1 U22656 ( .A1(n19705), .A2(n20074), .B1(n19718), .B2(n20072), .ZN(
        n19707) );
  AOI22_X1 U22657 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19711), .B1(
        n20073), .B2(n19710), .ZN(n19706) );
  OAI211_X1 U22658 ( .C1(n20077), .C2(n19738), .A(n19707), .B(n19706), .ZN(
        P2_U3093) );
  AOI22_X1 U22659 ( .A1(n20017), .A2(n19745), .B1(n19718), .B2(n20078), .ZN(
        n19709) );
  AOI22_X1 U22660 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19711), .B1(
        n20079), .B2(n19710), .ZN(n19708) );
  OAI211_X1 U22661 ( .C1(n20020), .C2(n19714), .A(n19709), .B(n19708), .ZN(
        P2_U3094) );
  AOI22_X1 U22662 ( .A1(n20022), .A2(n19745), .B1(n19718), .B2(n20084), .ZN(
        n19713) );
  AOI22_X1 U22663 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19711), .B1(
        n20086), .B2(n19710), .ZN(n19712) );
  OAI211_X1 U22664 ( .C1(n20028), .C2(n19714), .A(n19713), .B(n19712), .ZN(
        P2_U3095) );
  NAND2_X1 U22665 ( .A1(n10563), .A2(n20041), .ZN(n19717) );
  NAND2_X1 U22666 ( .A1(n19987), .A2(n20182), .ZN(n19759) );
  NOR2_X1 U22667 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19759), .ZN(
        n19743) );
  INV_X1 U22668 ( .A(n19743), .ZN(n19715) );
  AND2_X1 U22669 ( .A1(n20183), .A2(n19715), .ZN(n19716) );
  NAND2_X1 U22670 ( .A1(n19717), .A2(n19716), .ZN(n19723) );
  NOR2_X1 U22671 ( .A1(n19718), .A2(n19743), .ZN(n19725) );
  OAI21_X1 U22672 ( .B1(n19745), .B2(n19765), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19720) );
  AND2_X1 U22673 ( .A1(n19725), .A2(n19720), .ZN(n19721) );
  NOR2_X1 U22674 ( .A1(n19956), .A2(n19721), .ZN(n19722) );
  OAI21_X1 U22675 ( .B1(n10563), .B2(n19743), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19724) );
  OAI21_X1 U22676 ( .B1(n19725), .B2(n20183), .A(n19724), .ZN(n19744) );
  AOI22_X1 U22677 ( .A1(n19744), .A2(n20034), .B1(n20033), .B2(n19743), .ZN(
        n19727) );
  AOI22_X1 U22678 ( .A1(n19745), .A2(n19988), .B1(n19765), .B2(n20042), .ZN(
        n19726) );
  OAI211_X1 U22679 ( .C1(n19729), .C2(n19728), .A(n19727), .B(n19726), .ZN(
        P2_U3096) );
  AOI22_X1 U22680 ( .A1(n19744), .A2(n20047), .B1(n20046), .B2(n19743), .ZN(
        n19731) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19746), .B1(
        n19765), .B2(n20048), .ZN(n19730) );
  OAI211_X1 U22682 ( .C1(n20051), .C2(n19738), .A(n19731), .B(n19730), .ZN(
        P2_U3097) );
  AOI22_X1 U22683 ( .A1(n19744), .A2(n20053), .B1(n20052), .B2(n19743), .ZN(
        n19733) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19746), .B1(
        n19765), .B2(n20054), .ZN(n19732) );
  OAI211_X1 U22685 ( .C1(n20057), .C2(n19738), .A(n19733), .B(n19732), .ZN(
        P2_U3098) );
  AOI22_X1 U22686 ( .A1(n19744), .A2(n20059), .B1(n20058), .B2(n19743), .ZN(
        n19735) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19746), .B1(
        n19765), .B2(n20060), .ZN(n19734) );
  OAI211_X1 U22688 ( .C1(n20065), .C2(n19738), .A(n19735), .B(n19734), .ZN(
        P2_U3099) );
  AOI22_X1 U22689 ( .A1(n19744), .A2(n20067), .B1(n20066), .B2(n19743), .ZN(
        n19737) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19746), .B1(
        n19765), .B2(n19971), .ZN(n19736) );
  OAI211_X1 U22691 ( .C1(n19974), .C2(n19738), .A(n19737), .B(n19736), .ZN(
        P2_U3100) );
  AOI22_X1 U22692 ( .A1(n19744), .A2(n20073), .B1(n20072), .B2(n19743), .ZN(
        n19740) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n20074), .ZN(n19739) );
  OAI211_X1 U22694 ( .C1(n20077), .C2(n19783), .A(n19740), .B(n19739), .ZN(
        P2_U3101) );
  AOI22_X1 U22695 ( .A1(n19744), .A2(n20079), .B1(n20078), .B2(n19743), .ZN(
        n19742) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n20080), .ZN(n19741) );
  OAI211_X1 U22697 ( .C1(n20083), .C2(n19783), .A(n19742), .B(n19741), .ZN(
        P2_U3102) );
  AOI22_X1 U22698 ( .A1(n19744), .A2(n20086), .B1(n20084), .B2(n19743), .ZN(
        n19748) );
  AOI22_X1 U22699 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n20088), .ZN(n19747) );
  OAI211_X1 U22700 ( .C1(n20094), .C2(n19783), .A(n19748), .B(n19747), .ZN(
        P2_U3103) );
  NAND2_X1 U22701 ( .A1(n19749), .A2(n20174), .ZN(n20178) );
  NAND2_X1 U22702 ( .A1(n20178), .A2(n19759), .ZN(n19755) );
  NOR2_X1 U22703 ( .A1(n20208), .A2(n19759), .ZN(n19788) );
  INV_X1 U22704 ( .A(n19788), .ZN(n19750) );
  AND2_X1 U22705 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19750), .ZN(n19751) );
  NAND2_X1 U22706 ( .A1(n19752), .A2(n19751), .ZN(n19756) );
  OAI211_X1 U22707 ( .C1(n19788), .C2(n20041), .A(n19756), .B(n20039), .ZN(
        n19753) );
  INV_X1 U22708 ( .A(n19753), .ZN(n19754) );
  INV_X1 U22709 ( .A(n19756), .ZN(n19757) );
  AOI211_X2 U22710 ( .C1(n19759), .C2(n19953), .A(n19758), .B(n19757), .ZN(
        n19779) );
  AOI22_X1 U22711 ( .A1(n19779), .A2(n20034), .B1(n20033), .B2(n19788), .ZN(
        n19763) );
  AOI22_X1 U22712 ( .A1(n19765), .A2(n19988), .B1(n19816), .B2(n20042), .ZN(
        n19762) );
  OAI211_X1 U22713 ( .C1(n19768), .C2(n19764), .A(n19763), .B(n19762), .ZN(
        P2_U3104) );
  AOI22_X1 U22714 ( .A1(n19779), .A2(n20047), .B1(n20046), .B2(n19788), .ZN(
        n19767) );
  AOI22_X1 U22715 ( .A1(n19765), .A2(n19932), .B1(n19816), .B2(n20048), .ZN(
        n19766) );
  OAI211_X1 U22716 ( .C1(n19768), .C2(n21236), .A(n19767), .B(n19766), .ZN(
        P2_U3105) );
  AOI22_X1 U22717 ( .A1(n19779), .A2(n20053), .B1(n20052), .B2(n19788), .ZN(
        n19770) );
  INV_X1 U22718 ( .A(n19768), .ZN(n19780) );
  AOI22_X1 U22719 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19780), .B1(
        n19816), .B2(n20054), .ZN(n19769) );
  OAI211_X1 U22720 ( .C1(n20057), .C2(n19783), .A(n19770), .B(n19769), .ZN(
        P2_U3106) );
  AOI22_X1 U22721 ( .A1(n19779), .A2(n20059), .B1(n20058), .B2(n19788), .ZN(
        n19772) );
  AOI22_X1 U22722 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19780), .B1(
        n19816), .B2(n20060), .ZN(n19771) );
  OAI211_X1 U22723 ( .C1(n20065), .C2(n19783), .A(n19772), .B(n19771), .ZN(
        P2_U3107) );
  AOI22_X1 U22724 ( .A1(n19779), .A2(n20067), .B1(n20066), .B2(n19788), .ZN(
        n19774) );
  AOI22_X1 U22725 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19780), .B1(
        n19816), .B2(n19971), .ZN(n19773) );
  OAI211_X1 U22726 ( .C1(n19974), .C2(n19783), .A(n19774), .B(n19773), .ZN(
        P2_U3108) );
  AOI22_X1 U22727 ( .A1(n19779), .A2(n20073), .B1(n20072), .B2(n19788), .ZN(
        n19776) );
  AOI22_X1 U22728 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19780), .B1(
        n19816), .B2(n19975), .ZN(n19775) );
  OAI211_X1 U22729 ( .C1(n19978), .C2(n19783), .A(n19776), .B(n19775), .ZN(
        P2_U3109) );
  AOI22_X1 U22730 ( .A1(n19779), .A2(n20079), .B1(n20078), .B2(n19788), .ZN(
        n19778) );
  AOI22_X1 U22731 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19780), .B1(
        n19816), .B2(n20017), .ZN(n19777) );
  OAI211_X1 U22732 ( .C1(n20020), .C2(n19783), .A(n19778), .B(n19777), .ZN(
        P2_U3110) );
  AOI22_X1 U22733 ( .A1(n19779), .A2(n20086), .B1(n20084), .B2(n19788), .ZN(
        n19782) );
  AOI22_X1 U22734 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19780), .B1(
        n19816), .B2(n20022), .ZN(n19781) );
  OAI211_X1 U22735 ( .C1(n20028), .C2(n19783), .A(n19782), .B(n19781), .ZN(
        P2_U3111) );
  INV_X1 U22736 ( .A(n19851), .ZN(n19786) );
  INV_X1 U22737 ( .A(n19816), .ZN(n19785) );
  AOI21_X1 U22738 ( .B1(n19786), .B2(n19785), .A(n20228), .ZN(n19787) );
  NOR2_X1 U22739 ( .A1(n19787), .A2(n20183), .ZN(n19790) );
  NAND2_X1 U22740 ( .A1(n20190), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19889) );
  OR2_X1 U22741 ( .A1(n19889), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19829) );
  NOR2_X1 U22742 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19829), .ZN(
        n19815) );
  NOR2_X1 U22743 ( .A1(n19815), .A2(n19788), .ZN(n19791) );
  AOI211_X1 U22744 ( .C1(n10560), .C2(n20041), .A(n19815), .B(n19989), .ZN(
        n19789) );
  INV_X1 U22745 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n19796) );
  AOI22_X1 U22746 ( .A1(n19851), .A2(n20042), .B1(n20033), .B2(n19815), .ZN(
        n19795) );
  INV_X1 U22747 ( .A(n19790), .ZN(n19793) );
  OAI21_X1 U22748 ( .B1(n10560), .B2(n19815), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19792) );
  AOI22_X1 U22749 ( .A1(n20034), .A2(n19817), .B1(n19816), .B2(n19988), .ZN(
        n19794) );
  OAI211_X1 U22750 ( .C1(n19821), .C2(n19796), .A(n19795), .B(n19794), .ZN(
        P2_U3112) );
  INV_X1 U22751 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n19799) );
  AOI22_X1 U22752 ( .A1(n19851), .A2(n20048), .B1(n20046), .B2(n19815), .ZN(
        n19798) );
  AOI22_X1 U22753 ( .A1(n20047), .A2(n19817), .B1(n19816), .B2(n19932), .ZN(
        n19797) );
  OAI211_X1 U22754 ( .C1(n19821), .C2(n19799), .A(n19798), .B(n19797), .ZN(
        P2_U3113) );
  INV_X1 U22755 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n19802) );
  AOI22_X1 U22756 ( .A1(n19851), .A2(n20054), .B1(n20052), .B2(n19815), .ZN(
        n19801) );
  AOI22_X1 U22757 ( .A1(n20053), .A2(n19817), .B1(n19816), .B2(n20004), .ZN(
        n19800) );
  OAI211_X1 U22758 ( .C1(n19821), .C2(n19802), .A(n19801), .B(n19800), .ZN(
        P2_U3114) );
  INV_X1 U22759 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n19805) );
  AOI22_X1 U22760 ( .A1(n19851), .A2(n20060), .B1(n20058), .B2(n19815), .ZN(
        n19804) );
  AOI22_X1 U22761 ( .A1(n20059), .A2(n19817), .B1(n19816), .B2(n20008), .ZN(
        n19803) );
  OAI211_X1 U22762 ( .C1(n19821), .C2(n19805), .A(n19804), .B(n19803), .ZN(
        P2_U3115) );
  AOI22_X1 U22763 ( .A1(n19851), .A2(n19971), .B1(n20066), .B2(n19815), .ZN(
        n19807) );
  AOI22_X1 U22764 ( .A1(n20067), .A2(n19817), .B1(n19816), .B2(n20068), .ZN(
        n19806) );
  OAI211_X1 U22765 ( .C1(n19821), .C2(n19808), .A(n19807), .B(n19806), .ZN(
        P2_U3116) );
  INV_X1 U22766 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n19811) );
  AOI22_X1 U22767 ( .A1(n19851), .A2(n19975), .B1(n20072), .B2(n19815), .ZN(
        n19810) );
  AOI22_X1 U22768 ( .A1(n20073), .A2(n19817), .B1(n19816), .B2(n20074), .ZN(
        n19809) );
  OAI211_X1 U22769 ( .C1(n19821), .C2(n19811), .A(n19810), .B(n19809), .ZN(
        P2_U3117) );
  INV_X1 U22770 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n19814) );
  AOI22_X1 U22771 ( .A1(n19851), .A2(n20017), .B1(n20078), .B2(n19815), .ZN(
        n19813) );
  AOI22_X1 U22772 ( .A1(n20079), .A2(n19817), .B1(n19816), .B2(n20080), .ZN(
        n19812) );
  OAI211_X1 U22773 ( .C1(n19821), .C2(n19814), .A(n19813), .B(n19812), .ZN(
        P2_U3118) );
  INV_X1 U22774 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n19820) );
  AOI22_X1 U22775 ( .A1(n19851), .A2(n20022), .B1(n20084), .B2(n19815), .ZN(
        n19819) );
  AOI22_X1 U22776 ( .A1(n20086), .A2(n19817), .B1(n19816), .B2(n20088), .ZN(
        n19818) );
  OAI211_X1 U22777 ( .C1(n19821), .C2(n19820), .A(n19819), .B(n19818), .ZN(
        P2_U3119) );
  NOR2_X1 U22778 ( .A1(n20177), .A2(n20228), .ZN(n20035) );
  AOI21_X1 U22779 ( .B1(n20035), .B2(n19822), .A(n20183), .ZN(n19827) );
  INV_X1 U22780 ( .A(n10543), .ZN(n19823) );
  AOI21_X1 U22781 ( .B1(n19823), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19825) );
  NOR2_X1 U22782 ( .A1(n19824), .A2(n19889), .ZN(n19861) );
  OAI21_X1 U22783 ( .B1(n19825), .B2(n19861), .A(n20039), .ZN(n19826) );
  INV_X1 U22784 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19834) );
  AOI22_X1 U22785 ( .A1(n19851), .A2(n19988), .B1(n20033), .B2(n19861), .ZN(
        n19833) );
  INV_X1 U22786 ( .A(n19827), .ZN(n19830) );
  OAI21_X1 U22787 ( .B1(n10543), .B2(n19861), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19828) );
  OAI21_X1 U22788 ( .B1(n19830), .B2(n19829), .A(n19828), .ZN(n19852) );
  NOR2_X2 U22789 ( .A1(n19962), .A2(n19831), .ZN(n19882) );
  AOI22_X1 U22790 ( .A1(n20034), .A2(n19852), .B1(n19882), .B2(n20042), .ZN(
        n19832) );
  OAI211_X1 U22791 ( .C1(n19855), .C2(n19834), .A(n19833), .B(n19832), .ZN(
        P2_U3120) );
  INV_X1 U22792 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n19837) );
  AOI22_X1 U22793 ( .A1(n20048), .A2(n19882), .B1(n20046), .B2(n19861), .ZN(
        n19836) );
  AOI22_X1 U22794 ( .A1(n20047), .A2(n19852), .B1(n19851), .B2(n19932), .ZN(
        n19835) );
  OAI211_X1 U22795 ( .C1(n19855), .C2(n19837), .A(n19836), .B(n19835), .ZN(
        P2_U3121) );
  AOI22_X1 U22796 ( .A1(n20054), .A2(n19882), .B1(n20052), .B2(n19861), .ZN(
        n19839) );
  AOI22_X1 U22797 ( .A1(n20053), .A2(n19852), .B1(n19851), .B2(n20004), .ZN(
        n19838) );
  OAI211_X1 U22798 ( .C1(n19855), .C2(n10488), .A(n19839), .B(n19838), .ZN(
        P2_U3122) );
  AOI22_X1 U22799 ( .A1(n20060), .A2(n19882), .B1(n20058), .B2(n19861), .ZN(
        n19841) );
  AOI22_X1 U22800 ( .A1(n20059), .A2(n19852), .B1(n19851), .B2(n20008), .ZN(
        n19840) );
  OAI211_X1 U22801 ( .C1(n19855), .C2(n19842), .A(n19841), .B(n19840), .ZN(
        P2_U3123) );
  AOI22_X1 U22802 ( .A1(n19971), .A2(n19882), .B1(n20066), .B2(n19861), .ZN(
        n19844) );
  AOI22_X1 U22803 ( .A1(n20067), .A2(n19852), .B1(n19851), .B2(n20068), .ZN(
        n19843) );
  OAI211_X1 U22804 ( .C1(n19855), .C2(n21197), .A(n19844), .B(n19843), .ZN(
        P2_U3124) );
  INV_X1 U22805 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n19847) );
  AOI22_X1 U22806 ( .A1(n19851), .A2(n20074), .B1(n20072), .B2(n19861), .ZN(
        n19846) );
  AOI22_X1 U22807 ( .A1(n20073), .A2(n19852), .B1(n19882), .B2(n19975), .ZN(
        n19845) );
  OAI211_X1 U22808 ( .C1(n19855), .C2(n19847), .A(n19846), .B(n19845), .ZN(
        P2_U3125) );
  INV_X1 U22809 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n19850) );
  AOI22_X1 U22810 ( .A1(n20017), .A2(n19882), .B1(n20078), .B2(n19861), .ZN(
        n19849) );
  AOI22_X1 U22811 ( .A1(n20079), .A2(n19852), .B1(n19851), .B2(n20080), .ZN(
        n19848) );
  OAI211_X1 U22812 ( .C1(n19855), .C2(n19850), .A(n19849), .B(n19848), .ZN(
        P2_U3126) );
  AOI22_X1 U22813 ( .A1(n19851), .A2(n20088), .B1(n20084), .B2(n19861), .ZN(
        n19854) );
  AOI22_X1 U22814 ( .A1(n20086), .A2(n19852), .B1(n19882), .B2(n20022), .ZN(
        n19853) );
  OAI211_X1 U22815 ( .C1(n19855), .C2(n10652), .A(n19854), .B(n19853), .ZN(
        P2_U3127) );
  INV_X1 U22816 ( .A(n19857), .ZN(n19860) );
  NOR2_X1 U22817 ( .A1(n19858), .A2(n19889), .ZN(n19880) );
  OAI21_X1 U22818 ( .B1(n10562), .B2(n19880), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19859) );
  OAI21_X1 U22819 ( .B1(n19889), .B2(n19860), .A(n19859), .ZN(n19881) );
  AOI22_X1 U22820 ( .A1(n19881), .A2(n20034), .B1(n20033), .B2(n19880), .ZN(
        n19867) );
  OAI21_X1 U22821 ( .B1(n19882), .B2(n19910), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19864) );
  INV_X1 U22822 ( .A(n19861), .ZN(n19863) );
  OAI21_X1 U22823 ( .B1(n10562), .B2(n19953), .A(n20041), .ZN(n19862) );
  AOI21_X1 U22824 ( .B1(n19864), .B2(n19863), .A(n19862), .ZN(n19865) );
  OAI21_X1 U22825 ( .B1(n19865), .B2(n19880), .A(n20039), .ZN(n19883) );
  AOI22_X1 U22826 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n19988), .ZN(n19866) );
  OAI211_X1 U22827 ( .C1(n20001), .C2(n19920), .A(n19867), .B(n19866), .ZN(
        P2_U3128) );
  AOI22_X1 U22828 ( .A1(n19881), .A2(n20047), .B1(n20046), .B2(n19880), .ZN(
        n19869) );
  AOI22_X1 U22829 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n19932), .ZN(n19868) );
  OAI211_X1 U22830 ( .C1(n19935), .C2(n19920), .A(n19869), .B(n19868), .ZN(
        P2_U3129) );
  AOI22_X1 U22831 ( .A1(n19881), .A2(n20053), .B1(n20052), .B2(n19880), .ZN(
        n19871) );
  AOI22_X1 U22832 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n20004), .ZN(n19870) );
  OAI211_X1 U22833 ( .C1(n20007), .C2(n19920), .A(n19871), .B(n19870), .ZN(
        P2_U3130) );
  AOI22_X1 U22834 ( .A1(n19881), .A2(n20059), .B1(n20058), .B2(n19880), .ZN(
        n19873) );
  AOI22_X1 U22835 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n20008), .ZN(n19872) );
  OAI211_X1 U22836 ( .C1(n20011), .C2(n19920), .A(n19873), .B(n19872), .ZN(
        P2_U3131) );
  AOI22_X1 U22837 ( .A1(n19881), .A2(n20067), .B1(n20066), .B2(n19880), .ZN(
        n19875) );
  AOI22_X1 U22838 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n20068), .ZN(n19874) );
  OAI211_X1 U22839 ( .C1(n20071), .C2(n19920), .A(n19875), .B(n19874), .ZN(
        P2_U3132) );
  AOI22_X1 U22840 ( .A1(n19881), .A2(n20073), .B1(n20072), .B2(n19880), .ZN(
        n19877) );
  AOI22_X1 U22841 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n20074), .ZN(n19876) );
  OAI211_X1 U22842 ( .C1(n20077), .C2(n19920), .A(n19877), .B(n19876), .ZN(
        P2_U3133) );
  AOI22_X1 U22843 ( .A1(n19881), .A2(n20079), .B1(n20078), .B2(n19880), .ZN(
        n19879) );
  AOI22_X1 U22844 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n20080), .ZN(n19878) );
  OAI211_X1 U22845 ( .C1(n20083), .C2(n19920), .A(n19879), .B(n19878), .ZN(
        P2_U3134) );
  AOI22_X1 U22846 ( .A1(n19881), .A2(n20086), .B1(n20084), .B2(n19880), .ZN(
        n19885) );
  AOI22_X1 U22847 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19883), .B1(
        n19882), .B2(n20088), .ZN(n19884) );
  OAI211_X1 U22848 ( .C1(n20094), .C2(n19920), .A(n19885), .B(n19884), .ZN(
        P2_U3135) );
  NOR2_X2 U22849 ( .A1(n19962), .A2(n19886), .ZN(n19948) );
  NOR2_X1 U22850 ( .A1(n20199), .A2(n19889), .ZN(n19899) );
  INV_X1 U22851 ( .A(n19899), .ZN(n19887) );
  OR2_X1 U22852 ( .A1(n19887), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19893) );
  INV_X1 U22853 ( .A(n19888), .ZN(n19891) );
  INV_X1 U22854 ( .A(n19889), .ZN(n19890) );
  NAND2_X1 U22855 ( .A1(n19891), .A2(n19890), .ZN(n19894) );
  NAND2_X1 U22856 ( .A1(n19894), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19892) );
  NOR2_X1 U22857 ( .A1(n10542), .A2(n19892), .ZN(n19896) );
  AOI21_X1 U22858 ( .B1(n19953), .B2(n19893), .A(n19896), .ZN(n19916) );
  INV_X1 U22859 ( .A(n19894), .ZN(n19915) );
  AOI22_X1 U22860 ( .A1(n19916), .A2(n20034), .B1(n20033), .B2(n19915), .ZN(
        n19901) );
  AND2_X1 U22861 ( .A1(n19894), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19895) );
  NOR3_X1 U22862 ( .A1(n19896), .A2(n19956), .A3(n19895), .ZN(n19897) );
  OAI221_X1 U22863 ( .B1(n19899), .B2(n19898), .C1(n19899), .C2(n20035), .A(
        n19897), .ZN(n19917) );
  AOI22_X1 U22864 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19917), .B1(
        n19910), .B2(n19988), .ZN(n19900) );
  OAI211_X1 U22865 ( .C1(n20001), .C2(n19925), .A(n19901), .B(n19900), .ZN(
        P2_U3136) );
  AOI22_X1 U22866 ( .A1(n19916), .A2(n20047), .B1(n20046), .B2(n19915), .ZN(
        n19903) );
  AOI22_X1 U22867 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19917), .B1(
        n19948), .B2(n20048), .ZN(n19902) );
  OAI211_X1 U22868 ( .C1(n20051), .C2(n19920), .A(n19903), .B(n19902), .ZN(
        P2_U3137) );
  AOI22_X1 U22869 ( .A1(n19916), .A2(n20053), .B1(n20052), .B2(n19915), .ZN(
        n19905) );
  AOI22_X1 U22870 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19917), .B1(
        n19910), .B2(n20004), .ZN(n19904) );
  OAI211_X1 U22871 ( .C1(n20007), .C2(n19925), .A(n19905), .B(n19904), .ZN(
        P2_U3138) );
  AOI22_X1 U22872 ( .A1(n19916), .A2(n20059), .B1(n20058), .B2(n19915), .ZN(
        n19907) );
  AOI22_X1 U22873 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19917), .B1(
        n19910), .B2(n20008), .ZN(n19906) );
  OAI211_X1 U22874 ( .C1(n20011), .C2(n19925), .A(n19907), .B(n19906), .ZN(
        P2_U3139) );
  AOI22_X1 U22875 ( .A1(n19916), .A2(n20067), .B1(n20066), .B2(n19915), .ZN(
        n19909) );
  AOI22_X1 U22876 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19917), .B1(
        n19948), .B2(n19971), .ZN(n19908) );
  OAI211_X1 U22877 ( .C1(n19974), .C2(n19920), .A(n19909), .B(n19908), .ZN(
        P2_U3140) );
  AOI22_X1 U22878 ( .A1(n19916), .A2(n20073), .B1(n20072), .B2(n19915), .ZN(
        n19912) );
  AOI22_X1 U22879 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19917), .B1(
        n19910), .B2(n20074), .ZN(n19911) );
  OAI211_X1 U22880 ( .C1(n20077), .C2(n19925), .A(n19912), .B(n19911), .ZN(
        P2_U3141) );
  AOI22_X1 U22881 ( .A1(n19916), .A2(n20079), .B1(n20078), .B2(n19915), .ZN(
        n19914) );
  AOI22_X1 U22882 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19917), .B1(
        n19948), .B2(n20017), .ZN(n19913) );
  OAI211_X1 U22883 ( .C1(n20020), .C2(n19920), .A(n19914), .B(n19913), .ZN(
        P2_U3142) );
  AOI22_X1 U22884 ( .A1(n19916), .A2(n20086), .B1(n20084), .B2(n19915), .ZN(
        n19919) );
  AOI22_X1 U22885 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19917), .B1(
        n19948), .B2(n20022), .ZN(n19918) );
  OAI211_X1 U22886 ( .C1(n20028), .C2(n19920), .A(n19919), .B(n19918), .ZN(
        P2_U3143) );
  INV_X1 U22887 ( .A(n19921), .ZN(n19924) );
  INV_X1 U22888 ( .A(n19928), .ZN(n19923) );
  NAND3_X1 U22889 ( .A1(n20199), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19952) );
  INV_X1 U22890 ( .A(n19952), .ZN(n19960) );
  AND2_X1 U22891 ( .A1(n20208), .A2(n19960), .ZN(n19946) );
  OAI21_X1 U22892 ( .B1(n10561), .B2(n19946), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19922) );
  OAI21_X1 U22893 ( .B1(n19924), .B2(n19923), .A(n19922), .ZN(n19947) );
  AOI22_X1 U22894 ( .A1(n19947), .A2(n20034), .B1(n20033), .B2(n19946), .ZN(
        n19931) );
  AOI21_X1 U22895 ( .B1(n19985), .B2(n19925), .A(n20228), .ZN(n19929) );
  AOI211_X1 U22896 ( .C1(n10561), .C2(n20041), .A(n19989), .B(n19946), .ZN(
        n19926) );
  NOR2_X1 U22897 ( .A1(n19926), .A2(n19956), .ZN(n19927) );
  OAI211_X1 U22898 ( .C1(n19929), .C2(n19928), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19927), .ZN(n19949) );
  AOI22_X1 U22899 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19949), .B1(
        n19948), .B2(n19988), .ZN(n19930) );
  OAI211_X1 U22900 ( .C1(n20001), .C2(n19985), .A(n19931), .B(n19930), .ZN(
        P2_U3144) );
  AOI22_X1 U22901 ( .A1(n19947), .A2(n20047), .B1(n20046), .B2(n19946), .ZN(
        n19934) );
  AOI22_X1 U22902 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19949), .B1(
        n19948), .B2(n19932), .ZN(n19933) );
  OAI211_X1 U22903 ( .C1(n19935), .C2(n19985), .A(n19934), .B(n19933), .ZN(
        P2_U3145) );
  AOI22_X1 U22904 ( .A1(n19947), .A2(n20053), .B1(n20052), .B2(n19946), .ZN(
        n19937) );
  AOI22_X1 U22905 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19949), .B1(
        n19948), .B2(n20004), .ZN(n19936) );
  OAI211_X1 U22906 ( .C1(n20007), .C2(n19985), .A(n19937), .B(n19936), .ZN(
        P2_U3146) );
  AOI22_X1 U22907 ( .A1(n19947), .A2(n20059), .B1(n20058), .B2(n19946), .ZN(
        n19939) );
  AOI22_X1 U22908 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19949), .B1(
        n19948), .B2(n20008), .ZN(n19938) );
  OAI211_X1 U22909 ( .C1(n20011), .C2(n19985), .A(n19939), .B(n19938), .ZN(
        P2_U3147) );
  AOI22_X1 U22910 ( .A1(n19947), .A2(n20067), .B1(n20066), .B2(n19946), .ZN(
        n19941) );
  AOI22_X1 U22911 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19949), .B1(
        n19948), .B2(n20068), .ZN(n19940) );
  OAI211_X1 U22912 ( .C1(n20071), .C2(n19985), .A(n19941), .B(n19940), .ZN(
        P2_U3148) );
  AOI22_X1 U22913 ( .A1(n19947), .A2(n20073), .B1(n20072), .B2(n19946), .ZN(
        n19943) );
  AOI22_X1 U22914 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19949), .B1(
        n19948), .B2(n20074), .ZN(n19942) );
  OAI211_X1 U22915 ( .C1(n20077), .C2(n19985), .A(n19943), .B(n19942), .ZN(
        P2_U3149) );
  AOI22_X1 U22916 ( .A1(n19947), .A2(n20079), .B1(n20078), .B2(n19946), .ZN(
        n19945) );
  AOI22_X1 U22917 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19949), .B1(
        n19948), .B2(n20080), .ZN(n19944) );
  OAI211_X1 U22918 ( .C1(n20083), .C2(n19985), .A(n19945), .B(n19944), .ZN(
        P2_U3150) );
  AOI22_X1 U22919 ( .A1(n19947), .A2(n20086), .B1(n20084), .B2(n19946), .ZN(
        n19951) );
  AOI22_X1 U22920 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19949), .B1(
        n19948), .B2(n20088), .ZN(n19950) );
  OAI211_X1 U22921 ( .C1(n20094), .C2(n19985), .A(n19951), .B(n19950), .ZN(
        P2_U3151) );
  NOR2_X1 U22922 ( .A1(n20208), .A2(n19952), .ZN(n19991) );
  NOR3_X1 U22923 ( .A1(n10540), .A2(n19991), .A3(n19953), .ZN(n19955) );
  AOI21_X1 U22924 ( .B1(n20041), .B2(n19960), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19954) );
  NOR2_X1 U22925 ( .A1(n19955), .A2(n19954), .ZN(n19981) );
  AOI22_X1 U22926 ( .A1(n19981), .A2(n20034), .B1(n20033), .B2(n19991), .ZN(
        n19964) );
  INV_X1 U22927 ( .A(n19991), .ZN(n19957) );
  AOI211_X1 U22928 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19957), .A(n19956), 
        .B(n19955), .ZN(n19958) );
  OAI221_X1 U22929 ( .B1(n19960), .B2(n19959), .C1(n19960), .C2(n20035), .A(
        n19958), .ZN(n19982) );
  AOI22_X1 U22930 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19982), .B1(
        n20014), .B2(n20042), .ZN(n19963) );
  OAI211_X1 U22931 ( .C1(n20045), .C2(n19985), .A(n19964), .B(n19963), .ZN(
        P2_U3152) );
  AOI22_X1 U22932 ( .A1(n19981), .A2(n20047), .B1(n20046), .B2(n19991), .ZN(
        n19966) );
  AOI22_X1 U22933 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19982), .B1(
        n20014), .B2(n20048), .ZN(n19965) );
  OAI211_X1 U22934 ( .C1(n20051), .C2(n19985), .A(n19966), .B(n19965), .ZN(
        P2_U3153) );
  AOI22_X1 U22935 ( .A1(n19981), .A2(n20053), .B1(n20052), .B2(n19991), .ZN(
        n19968) );
  AOI22_X1 U22936 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19982), .B1(
        n20014), .B2(n20054), .ZN(n19967) );
  OAI211_X1 U22937 ( .C1(n20057), .C2(n19985), .A(n19968), .B(n19967), .ZN(
        P2_U3154) );
  AOI22_X1 U22938 ( .A1(n19981), .A2(n20059), .B1(n20058), .B2(n19991), .ZN(
        n19970) );
  AOI22_X1 U22939 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19982), .B1(
        n20014), .B2(n20060), .ZN(n19969) );
  OAI211_X1 U22940 ( .C1(n20065), .C2(n19985), .A(n19970), .B(n19969), .ZN(
        P2_U3155) );
  AOI22_X1 U22941 ( .A1(n19981), .A2(n20067), .B1(n20066), .B2(n19991), .ZN(
        n19973) );
  AOI22_X1 U22942 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19982), .B1(
        n20014), .B2(n19971), .ZN(n19972) );
  OAI211_X1 U22943 ( .C1(n19974), .C2(n19985), .A(n19973), .B(n19972), .ZN(
        P2_U3156) );
  AOI22_X1 U22944 ( .A1(n19981), .A2(n20073), .B1(n20072), .B2(n19991), .ZN(
        n19977) );
  AOI22_X1 U22945 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19982), .B1(
        n20014), .B2(n19975), .ZN(n19976) );
  OAI211_X1 U22946 ( .C1(n19978), .C2(n19985), .A(n19977), .B(n19976), .ZN(
        P2_U3157) );
  AOI22_X1 U22947 ( .A1(n19981), .A2(n20079), .B1(n20078), .B2(n19991), .ZN(
        n19980) );
  AOI22_X1 U22948 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19982), .B1(
        n20014), .B2(n20017), .ZN(n19979) );
  OAI211_X1 U22949 ( .C1(n20020), .C2(n19985), .A(n19980), .B(n19979), .ZN(
        P2_U3158) );
  AOI22_X1 U22950 ( .A1(n19981), .A2(n20086), .B1(n20084), .B2(n19991), .ZN(
        n19984) );
  AOI22_X1 U22951 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19982), .B1(
        n20014), .B2(n20022), .ZN(n19983) );
  OAI211_X1 U22952 ( .C1(n20028), .C2(n19985), .A(n19984), .B(n19983), .ZN(
        P2_U3159) );
  NAND2_X1 U22953 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19987), .ZN(
        n20037) );
  NOR2_X1 U22954 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20037), .ZN(
        n20021) );
  AOI22_X1 U22955 ( .A1(n19988), .A2(n20014), .B1(n20033), .B2(n20021), .ZN(
        n20000) );
  OAI21_X1 U22956 ( .B1(n20014), .B2(n20089), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19990) );
  NAND2_X1 U22957 ( .A1(n19990), .A2(n19989), .ZN(n19998) );
  NOR2_X1 U22958 ( .A1(n20021), .A2(n19991), .ZN(n19997) );
  INV_X1 U22959 ( .A(n19997), .ZN(n19995) );
  INV_X1 U22960 ( .A(n20021), .ZN(n19992) );
  OAI211_X1 U22961 ( .C1(n19993), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19992), 
        .B(n20183), .ZN(n19994) );
  OAI211_X1 U22962 ( .C1(n19998), .C2(n19995), .A(n20039), .B(n19994), .ZN(
        n20024) );
  OAI21_X1 U22963 ( .B1(n10559), .B2(n20021), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19996) );
  AOI22_X1 U22964 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20024), .B1(
        n20034), .B2(n20023), .ZN(n19999) );
  OAI211_X1 U22965 ( .C1(n20001), .C2(n20064), .A(n20000), .B(n19999), .ZN(
        P2_U3160) );
  AOI22_X1 U22966 ( .A1(n20048), .A2(n20089), .B1(n20046), .B2(n20021), .ZN(
        n20003) );
  AOI22_X1 U22967 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20024), .B1(
        n20047), .B2(n20023), .ZN(n20002) );
  OAI211_X1 U22968 ( .C1(n20051), .C2(n20027), .A(n20003), .B(n20002), .ZN(
        P2_U3161) );
  AOI22_X1 U22969 ( .A1(n20004), .A2(n20014), .B1(n20052), .B2(n20021), .ZN(
        n20006) );
  AOI22_X1 U22970 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20024), .B1(
        n20053), .B2(n20023), .ZN(n20005) );
  OAI211_X1 U22971 ( .C1(n20007), .C2(n20064), .A(n20006), .B(n20005), .ZN(
        P2_U3162) );
  AOI22_X1 U22972 ( .A1(n20008), .A2(n20014), .B1(n20058), .B2(n20021), .ZN(
        n20010) );
  AOI22_X1 U22973 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20024), .B1(
        n20059), .B2(n20023), .ZN(n20009) );
  OAI211_X1 U22974 ( .C1(n20011), .C2(n20064), .A(n20010), .B(n20009), .ZN(
        P2_U3163) );
  AOI22_X1 U22975 ( .A1(n20068), .A2(n20014), .B1(n20066), .B2(n20021), .ZN(
        n20013) );
  AOI22_X1 U22976 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20024), .B1(
        n20067), .B2(n20023), .ZN(n20012) );
  OAI211_X1 U22977 ( .C1(n20071), .C2(n20064), .A(n20013), .B(n20012), .ZN(
        P2_U3164) );
  AOI22_X1 U22978 ( .A1(n20014), .A2(n20074), .B1(n20072), .B2(n20021), .ZN(
        n20016) );
  AOI22_X1 U22979 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20024), .B1(
        n20073), .B2(n20023), .ZN(n20015) );
  OAI211_X1 U22980 ( .C1(n20077), .C2(n20064), .A(n20016), .B(n20015), .ZN(
        P2_U3165) );
  AOI22_X1 U22981 ( .A1(n20017), .A2(n20089), .B1(n20078), .B2(n20021), .ZN(
        n20019) );
  AOI22_X1 U22982 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20024), .B1(
        n20079), .B2(n20023), .ZN(n20018) );
  OAI211_X1 U22983 ( .C1(n20020), .C2(n20027), .A(n20019), .B(n20018), .ZN(
        P2_U3166) );
  AOI22_X1 U22984 ( .A1(n20022), .A2(n20089), .B1(n20084), .B2(n20021), .ZN(
        n20026) );
  AOI22_X1 U22985 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20024), .B1(
        n20086), .B2(n20023), .ZN(n20025) );
  OAI211_X1 U22986 ( .C1(n20028), .C2(n20027), .A(n20026), .B(n20025), .ZN(
        P2_U3167) );
  NAND2_X1 U22987 ( .A1(n20029), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20030) );
  NOR2_X1 U22988 ( .A1(n10541), .A2(n20030), .ZN(n20036) );
  INV_X1 U22989 ( .A(n20037), .ZN(n20031) );
  AOI21_X1 U22990 ( .B1(n20041), .B2(n20031), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20032) );
  NOR2_X1 U22991 ( .A1(n20036), .A2(n20032), .ZN(n20087) );
  AOI22_X1 U22992 ( .A1(n20087), .A2(n20034), .B1(n20085), .B2(n20033), .ZN(
        n20044) );
  NAND2_X1 U22993 ( .A1(n20035), .A2(n20174), .ZN(n20038) );
  AOI21_X1 U22994 ( .B1(n20038), .B2(n20037), .A(n20036), .ZN(n20040) );
  OAI211_X1 U22995 ( .C1(n20085), .C2(n20041), .A(n20040), .B(n20039), .ZN(
        n20090) );
  AOI22_X1 U22996 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20090), .B1(
        n20061), .B2(n20042), .ZN(n20043) );
  OAI211_X1 U22997 ( .C1(n20045), .C2(n20064), .A(n20044), .B(n20043), .ZN(
        P2_U3168) );
  AOI22_X1 U22998 ( .A1(n20087), .A2(n20047), .B1(n20085), .B2(n20046), .ZN(
        n20050) );
  AOI22_X1 U22999 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20090), .B1(
        n20061), .B2(n20048), .ZN(n20049) );
  OAI211_X1 U23000 ( .C1(n20051), .C2(n20064), .A(n20050), .B(n20049), .ZN(
        P2_U3169) );
  AOI22_X1 U23001 ( .A1(n20087), .A2(n20053), .B1(n20085), .B2(n20052), .ZN(
        n20056) );
  AOI22_X1 U23002 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20090), .B1(
        n20061), .B2(n20054), .ZN(n20055) );
  OAI211_X1 U23003 ( .C1(n20057), .C2(n20064), .A(n20056), .B(n20055), .ZN(
        P2_U3170) );
  AOI22_X1 U23004 ( .A1(n20087), .A2(n20059), .B1(n20085), .B2(n20058), .ZN(
        n20063) );
  AOI22_X1 U23005 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20090), .B1(
        n20061), .B2(n20060), .ZN(n20062) );
  OAI211_X1 U23006 ( .C1(n20065), .C2(n20064), .A(n20063), .B(n20062), .ZN(
        P2_U3171) );
  AOI22_X1 U23007 ( .A1(n20087), .A2(n20067), .B1(n20085), .B2(n20066), .ZN(
        n20070) );
  AOI22_X1 U23008 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20090), .B1(
        n20089), .B2(n20068), .ZN(n20069) );
  OAI211_X1 U23009 ( .C1(n20071), .C2(n20093), .A(n20070), .B(n20069), .ZN(
        P2_U3172) );
  AOI22_X1 U23010 ( .A1(n20087), .A2(n20073), .B1(n20085), .B2(n20072), .ZN(
        n20076) );
  AOI22_X1 U23011 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20090), .B1(
        n20089), .B2(n20074), .ZN(n20075) );
  OAI211_X1 U23012 ( .C1(n20077), .C2(n20093), .A(n20076), .B(n20075), .ZN(
        P2_U3173) );
  AOI22_X1 U23013 ( .A1(n20087), .A2(n20079), .B1(n20085), .B2(n20078), .ZN(
        n20082) );
  AOI22_X1 U23014 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20090), .B1(
        n20089), .B2(n20080), .ZN(n20081) );
  OAI211_X1 U23015 ( .C1(n20083), .C2(n20093), .A(n20082), .B(n20081), .ZN(
        P2_U3174) );
  AOI22_X1 U23016 ( .A1(n20087), .A2(n20086), .B1(n20085), .B2(n20084), .ZN(
        n20092) );
  AOI22_X1 U23017 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20090), .B1(
        n20089), .B2(n20088), .ZN(n20091) );
  OAI211_X1 U23018 ( .C1(n20094), .C2(n20093), .A(n20092), .B(n20091), .ZN(
        P2_U3175) );
  AOI21_X1 U23019 ( .B1(n20176), .B2(n20096), .A(n20095), .ZN(n20100) );
  NOR2_X1 U23020 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n9681), .ZN(n20097) );
  OAI211_X1 U23021 ( .C1(n20101), .C2(n20097), .A(n20114), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20098) );
  OAI211_X1 U23022 ( .C1(n20101), .C2(n20100), .A(n20099), .B(n20098), .ZN(
        P2_U3177) );
  INV_X1 U23023 ( .A(n20173), .ZN(n20102) );
  AND2_X1 U23024 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20102), .ZN(
        P2_U3179) );
  AND2_X1 U23025 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20102), .ZN(
        P2_U3180) );
  AND2_X1 U23026 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20102), .ZN(
        P2_U3181) );
  AND2_X1 U23027 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20102), .ZN(
        P2_U3182) );
  AND2_X1 U23028 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20102), .ZN(
        P2_U3183) );
  AND2_X1 U23029 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20102), .ZN(
        P2_U3184) );
  AND2_X1 U23030 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20102), .ZN(
        P2_U3185) );
  AND2_X1 U23031 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20102), .ZN(
        P2_U3186) );
  AND2_X1 U23032 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20102), .ZN(
        P2_U3187) );
  AND2_X1 U23033 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20102), .ZN(
        P2_U3188) );
  AND2_X1 U23034 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20102), .ZN(
        P2_U3189) );
  AND2_X1 U23035 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20102), .ZN(
        P2_U3190) );
  AND2_X1 U23036 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20102), .ZN(
        P2_U3191) );
  AND2_X1 U23037 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20102), .ZN(
        P2_U3192) );
  AND2_X1 U23038 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20102), .ZN(
        P2_U3193) );
  AND2_X1 U23039 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20102), .ZN(
        P2_U3194) );
  AND2_X1 U23040 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20102), .ZN(
        P2_U3195) );
  AND2_X1 U23041 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20102), .ZN(
        P2_U3196) );
  AND2_X1 U23042 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20102), .ZN(
        P2_U3197) );
  AND2_X1 U23043 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20102), .ZN(
        P2_U3198) );
  AND2_X1 U23044 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20102), .ZN(
        P2_U3199) );
  AND2_X1 U23045 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20102), .ZN(
        P2_U3200) );
  AND2_X1 U23046 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20102), .ZN(P2_U3201) );
  AND2_X1 U23047 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20102), .ZN(P2_U3202) );
  AND2_X1 U23048 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20102), .ZN(P2_U3203) );
  AND2_X1 U23049 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20102), .ZN(P2_U3204) );
  AND2_X1 U23050 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20102), .ZN(P2_U3205) );
  AND2_X1 U23051 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20102), .ZN(P2_U3206) );
  AND2_X1 U23052 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20102), .ZN(P2_U3207) );
  AND2_X1 U23053 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20102), .ZN(P2_U3208) );
  INV_X1 U23054 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20233) );
  NOR2_X1 U23055 ( .A1(n20226), .A2(n21221), .ZN(n20111) );
  OR3_X1 U23056 ( .A1(n20233), .A2(n20103), .A3(n20111), .ZN(n20104) );
  INV_X1 U23057 ( .A(NA), .ZN(n20975) );
  NOR3_X1 U23058 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n20975), .ZN(n20117) );
  AOI21_X1 U23059 ( .B1(n20120), .B2(n20104), .A(n20117), .ZN(n20105) );
  OAI221_X1 U23060 ( .B1(n20106), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20106), .C2(n20110), .A(n20105), .ZN(P2_U3209) );
  AOI21_X1 U23061 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20110), .A(n20120), 
        .ZN(n20113) );
  NOR3_X1 U23062 ( .A1(n20113), .A2(n20233), .A3(n20103), .ZN(n20107) );
  NOR2_X1 U23063 ( .A1(n20107), .A2(n20111), .ZN(n20108) );
  OAI211_X1 U23064 ( .C1(n20110), .C2(n20109), .A(n20108), .B(n20227), .ZN(
        P2_U3210) );
  AOI22_X1 U23065 ( .A1(n20112), .A2(n20233), .B1(n20111), .B2(n20975), .ZN(
        n20119) );
  OAI21_X1 U23066 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n20118) );
  NOR2_X1 U23067 ( .A1(n21221), .A2(n20120), .ZN(n20115) );
  AOI21_X1 U23068 ( .B1(n20115), .B2(n20114), .A(n20113), .ZN(n20116) );
  OAI22_X1 U23069 ( .A1(n20119), .A2(n20118), .B1(n20117), .B2(n20116), .ZN(
        P2_U3211) );
  OAI222_X1 U23070 ( .A1(n20166), .A2(n21208), .B1(n20122), .B2(n20163), .C1(
        n20121), .C2(n20162), .ZN(P2_U3212) );
  OAI222_X1 U23071 ( .A1(n20166), .A2(n13609), .B1(n20123), .B2(n20163), .C1(
        n21208), .C2(n20162), .ZN(P2_U3213) );
  OAI222_X1 U23072 ( .A1(n20166), .A2(n12536), .B1(n20124), .B2(n20163), .C1(
        n13609), .C2(n20162), .ZN(P2_U3214) );
  OAI222_X1 U23073 ( .A1(n20166), .A2(n12527), .B1(n20125), .B2(n20163), .C1(
        n12536), .C2(n20162), .ZN(P2_U3215) );
  OAI222_X1 U23074 ( .A1(n20166), .A2(n20127), .B1(n20126), .B2(n20163), .C1(
        n12527), .C2(n20162), .ZN(P2_U3216) );
  OAI222_X1 U23075 ( .A1(n20166), .A2(n20129), .B1(n20128), .B2(n20163), .C1(
        n20127), .C2(n20162), .ZN(P2_U3217) );
  OAI222_X1 U23076 ( .A1(n20166), .A2(n12590), .B1(n20130), .B2(n20163), .C1(
        n20129), .C2(n20162), .ZN(P2_U3218) );
  OAI222_X1 U23077 ( .A1(n20166), .A2(n20132), .B1(n20131), .B2(n20163), .C1(
        n12590), .C2(n20162), .ZN(P2_U3219) );
  OAI222_X1 U23078 ( .A1(n20166), .A2(n12635), .B1(n20133), .B2(n20163), .C1(
        n20132), .C2(n20162), .ZN(P2_U3220) );
  OAI222_X1 U23079 ( .A1(n20166), .A2(n10738), .B1(n20134), .B2(n20163), .C1(
        n12635), .C2(n20162), .ZN(P2_U3221) );
  OAI222_X1 U23080 ( .A1(n20166), .A2(n20136), .B1(n20135), .B2(n20163), .C1(
        n10738), .C2(n20162), .ZN(P2_U3222) );
  OAI222_X1 U23081 ( .A1(n20166), .A2(n16109), .B1(n20137), .B2(n20163), .C1(
        n20136), .C2(n20162), .ZN(P2_U3223) );
  OAI222_X1 U23082 ( .A1(n20166), .A2(n12721), .B1(n20138), .B2(n20163), .C1(
        n16109), .C2(n20162), .ZN(P2_U3224) );
  OAI222_X1 U23083 ( .A1(n20166), .A2(n15841), .B1(n20139), .B2(n20163), .C1(
        n12721), .C2(n20162), .ZN(P2_U3225) );
  OAI222_X1 U23084 ( .A1(n20166), .A2(n20141), .B1(n20140), .B2(n20163), .C1(
        n15841), .C2(n20162), .ZN(P2_U3226) );
  OAI222_X1 U23085 ( .A1(n20166), .A2(n20143), .B1(n20142), .B2(n20163), .C1(
        n20141), .C2(n20162), .ZN(P2_U3227) );
  OAI222_X1 U23086 ( .A1(n20166), .A2(n10756), .B1(n20144), .B2(n20163), .C1(
        n20143), .C2(n20162), .ZN(P2_U3228) );
  OAI222_X1 U23087 ( .A1(n20166), .A2(n10759), .B1(n20145), .B2(n20163), .C1(
        n10756), .C2(n20162), .ZN(P2_U3229) );
  OAI222_X1 U23088 ( .A1(n20166), .A2(n12749), .B1(n20146), .B2(n20163), .C1(
        n10759), .C2(n20162), .ZN(P2_U3230) );
  OAI222_X1 U23089 ( .A1(n20166), .A2(n20148), .B1(n20147), .B2(n20163), .C1(
        n12749), .C2(n20162), .ZN(P2_U3231) );
  OAI222_X1 U23090 ( .A1(n20166), .A2(n10767), .B1(n20149), .B2(n20163), .C1(
        n20148), .C2(n20162), .ZN(P2_U3232) );
  OAI222_X1 U23091 ( .A1(n20166), .A2(n10770), .B1(n20150), .B2(n20163), .C1(
        n10767), .C2(n20162), .ZN(P2_U3233) );
  INV_X1 U23092 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20152) );
  OAI222_X1 U23093 ( .A1(n20166), .A2(n20152), .B1(n20151), .B2(n20163), .C1(
        n10770), .C2(n20162), .ZN(P2_U3234) );
  INV_X1 U23094 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20154) );
  OAI222_X1 U23095 ( .A1(n20166), .A2(n20154), .B1(n20153), .B2(n20163), .C1(
        n20152), .C2(n20162), .ZN(P2_U3235) );
  OAI222_X1 U23096 ( .A1(n20166), .A2(n16455), .B1(n21237), .B2(n20163), .C1(
        n20154), .C2(n20162), .ZN(P2_U3236) );
  OAI222_X1 U23097 ( .A1(n20166), .A2(n20157), .B1(n20155), .B2(n20163), .C1(
        n16455), .C2(n20162), .ZN(P2_U3237) );
  INV_X1 U23098 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20158) );
  OAI222_X1 U23099 ( .A1(n20162), .A2(n20157), .B1(n20156), .B2(n20163), .C1(
        n20158), .C2(n20166), .ZN(P2_U3238) );
  OAI222_X1 U23100 ( .A1(n20166), .A2(n20160), .B1(n20159), .B2(n20163), .C1(
        n20158), .C2(n20162), .ZN(P2_U3239) );
  OAI222_X1 U23101 ( .A1(n20166), .A2(n12787), .B1(n20161), .B2(n20163), .C1(
        n20160), .C2(n20162), .ZN(P2_U3240) );
  OAI222_X1 U23102 ( .A1(n20166), .A2(n20165), .B1(n20164), .B2(n20163), .C1(
        n12787), .C2(n20162), .ZN(P2_U3241) );
  OAI22_X1 U23103 ( .A1(n20235), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20163), .ZN(n20167) );
  INV_X1 U23104 ( .A(n20167), .ZN(P2_U3585) );
  MUX2_X1 U23105 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20235), .Z(P2_U3586) );
  OAI22_X1 U23106 ( .A1(n20235), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20163), .ZN(n20168) );
  INV_X1 U23107 ( .A(n20168), .ZN(P2_U3587) );
  OAI22_X1 U23108 ( .A1(n20235), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20163), .ZN(n20169) );
  INV_X1 U23109 ( .A(n20169), .ZN(P2_U3588) );
  OAI21_X1 U23110 ( .B1(n20173), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20171), 
        .ZN(n20170) );
  INV_X1 U23111 ( .A(n20170), .ZN(P2_U3591) );
  OAI21_X1 U23112 ( .B1(n20173), .B2(n20172), .A(n20171), .ZN(P2_U3592) );
  INV_X1 U23113 ( .A(n20207), .ZN(n20206) );
  NAND2_X1 U23114 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20174), .ZN(n20175) );
  OAI21_X1 U23115 ( .B1(n20176), .B2(n20175), .A(n20191), .ZN(n20185) );
  OAI22_X1 U23116 ( .A1(n20178), .A2(n20183), .B1(n20177), .B2(n20185), .ZN(
        n20179) );
  AOI21_X1 U23117 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20180), .A(n20179), 
        .ZN(n20181) );
  AOI22_X1 U23118 ( .A1(n20206), .A2(n20182), .B1(n20181), .B2(n20207), .ZN(
        P2_U3602) );
  NOR2_X1 U23119 ( .A1(n20183), .A2(n20228), .ZN(n20195) );
  AOI21_X1 U23120 ( .B1(n20195), .B2(n20193), .A(n20184), .ZN(n20186) );
  NOR2_X1 U23121 ( .A1(n20186), .A2(n20185), .ZN(n20187) );
  AOI21_X1 U23122 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20188), .A(n20187), 
        .ZN(n20189) );
  AOI22_X1 U23123 ( .A1(n20206), .A2(n20190), .B1(n20189), .B2(n20207), .ZN(
        P2_U3603) );
  INV_X1 U23124 ( .A(n20191), .ZN(n20202) );
  NOR2_X1 U23125 ( .A1(n20202), .A2(n20192), .ZN(n20194) );
  MUX2_X1 U23126 ( .A(n20195), .B(n20194), .S(n20193), .Z(n20196) );
  AOI21_X1 U23127 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20197), .A(n20196), 
        .ZN(n20198) );
  AOI22_X1 U23128 ( .A1(n20206), .A2(n20199), .B1(n20198), .B2(n20207), .ZN(
        P2_U3604) );
  OAI22_X1 U23129 ( .A1(n20203), .A2(n20202), .B1(n20201), .B2(n20200), .ZN(
        n20204) );
  AOI21_X1 U23130 ( .B1(n20208), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20204), 
        .ZN(n20205) );
  OAI22_X1 U23131 ( .A1(n20208), .A2(n20207), .B1(n20206), .B2(n20205), .ZN(
        P2_U3605) );
  INV_X1 U23132 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20209) );
  AOI22_X1 U23133 ( .A1(n20163), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20209), 
        .B2(n20235), .ZN(P2_U3608) );
  INV_X1 U23134 ( .A(n20210), .ZN(n20216) );
  INV_X1 U23135 ( .A(n20211), .ZN(n20215) );
  NAND2_X1 U23136 ( .A1(n20213), .A2(n20212), .ZN(n20214) );
  OAI211_X1 U23137 ( .C1(n20217), .C2(n20216), .A(n20215), .B(n20214), .ZN(
        n20219) );
  MUX2_X1 U23138 ( .A(P2_MORE_REG_SCAN_IN), .B(n20219), .S(n20218), .Z(
        P2_U3609) );
  AOI21_X1 U23139 ( .B1(n20220), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20222) );
  AOI211_X1 U23140 ( .C1(n20226), .C2(n20223), .A(n20222), .B(n20221), .ZN(
        n20224) );
  INV_X1 U23141 ( .A(n20224), .ZN(n20234) );
  AOI21_X1 U23142 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20226), .A(n20225), 
        .ZN(n20231) );
  AOI21_X1 U23143 ( .B1(n10292), .B2(n20228), .A(n20227), .ZN(n20229) );
  NOR3_X1 U23144 ( .A1(n12840), .A2(n20229), .A3(n16267), .ZN(n20230) );
  OAI21_X1 U23145 ( .B1(n20231), .B2(n20230), .A(n20234), .ZN(n20232) );
  OAI21_X1 U23146 ( .B1(n20234), .B2(n20233), .A(n20232), .ZN(P2_U3610) );
  OAI22_X1 U23147 ( .A1(n20235), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20163), .ZN(n20236) );
  INV_X1 U23148 ( .A(n20236), .ZN(P2_U3611) );
  AOI21_X1 U23149 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20982), .A(n20969), 
        .ZN(n20243) );
  INV_X1 U23150 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20237) );
  AND2_X1 U23151 ( .A1(n20969), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21046) );
  AOI21_X1 U23152 ( .B1(n20243), .B2(n20237), .A(n21046), .ZN(P1_U2802) );
  OAI21_X1 U23153 ( .B1(n20239), .B2(n20238), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20240) );
  OAI21_X1 U23154 ( .B1(n20241), .B2(n20963), .A(n20240), .ZN(P1_U2803) );
  INV_X2 U23155 ( .A(n21046), .ZN(n21059) );
  NOR2_X1 U23156 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20244) );
  OAI21_X1 U23157 ( .B1(n20244), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21059), .ZN(
        n20242) );
  OAI21_X1 U23158 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21059), .A(n20242), 
        .ZN(P1_U2804) );
  NOR2_X1 U23159 ( .A1(n21046), .A2(n20243), .ZN(n21036) );
  OAI21_X1 U23160 ( .B1(BS16), .B2(n20244), .A(n21036), .ZN(n21034) );
  OAI21_X1 U23161 ( .B1(n21036), .B2(n20852), .A(n21034), .ZN(P1_U2805) );
  OAI21_X1 U23162 ( .B1(n20245), .B2(n21176), .A(n20363), .ZN(P1_U2806) );
  NOR4_X1 U23163 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20249) );
  NOR4_X1 U23164 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20248) );
  NOR4_X1 U23165 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20247) );
  NOR4_X1 U23166 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20246) );
  NAND4_X1 U23167 ( .A1(n20249), .A2(n20248), .A3(n20247), .A4(n20246), .ZN(
        n20255) );
  NOR4_X1 U23168 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20253) );
  AOI211_X1 U23169 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20252) );
  NOR4_X1 U23170 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20251) );
  NOR4_X1 U23171 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20250) );
  NAND4_X1 U23172 ( .A1(n20253), .A2(n20252), .A3(n20251), .A4(n20250), .ZN(
        n20254) );
  NOR2_X1 U23173 ( .A1(n20255), .A2(n20254), .ZN(n21044) );
  INV_X1 U23174 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20257) );
  NOR3_X1 U23175 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20258) );
  OAI21_X1 U23176 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20258), .A(n21044), .ZN(
        n20256) );
  OAI21_X1 U23177 ( .B1(n21044), .B2(n20257), .A(n20256), .ZN(P1_U2807) );
  INV_X1 U23178 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21035) );
  AOI21_X1 U23179 ( .B1(n21037), .B2(n21035), .A(n20258), .ZN(n20260) );
  INV_X1 U23180 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20259) );
  INV_X1 U23181 ( .A(n21044), .ZN(n21039) );
  AOI22_X1 U23182 ( .A1(n21044), .A2(n20260), .B1(n20259), .B2(n21039), .ZN(
        P1_U2808) );
  NAND2_X1 U23183 ( .A1(n20262), .A2(n20261), .ZN(n20293) );
  OAI21_X1 U23184 ( .B1(n20263), .B2(n20293), .A(n20292), .ZN(n20291) );
  INV_X1 U23185 ( .A(n20264), .ZN(n20268) );
  NAND2_X1 U23186 ( .A1(n20340), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n20265) );
  OAI211_X1 U23187 ( .C1(n20308), .C2(n20266), .A(n20322), .B(n20265), .ZN(
        n20267) );
  AOI21_X1 U23188 ( .B1(n20268), .B2(n20334), .A(n20267), .ZN(n20269) );
  OAI21_X1 U23189 ( .B1(n20270), .B2(P1_REIP_REG_9__SCAN_IN), .A(n20269), .ZN(
        n20271) );
  INV_X1 U23190 ( .A(n20271), .ZN(n20276) );
  INV_X1 U23191 ( .A(n20272), .ZN(n20274) );
  AOI22_X1 U23192 ( .A1(n20274), .A2(n20317), .B1(n20339), .B2(n20273), .ZN(
        n20275) );
  OAI211_X1 U23193 ( .C1(n20291), .C2(n20277), .A(n20276), .B(n20275), .ZN(
        P1_U2831) );
  NAND2_X1 U23194 ( .A1(n20335), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n20278) );
  OAI211_X1 U23195 ( .C1(n20279), .C2(n21209), .A(n20278), .B(n20322), .ZN(
        n20283) );
  NAND3_X1 U23196 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n20281) );
  NOR3_X1 U23197 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20281), .A3(n20280), .ZN(
        n20282) );
  AOI211_X1 U23198 ( .C1(n20334), .C2(n20284), .A(n20283), .B(n20282), .ZN(
        n20285) );
  OAI21_X1 U23199 ( .B1(n20287), .B2(n20286), .A(n20285), .ZN(n20288) );
  AOI21_X1 U23200 ( .B1(n20289), .B2(n20339), .A(n20288), .ZN(n20290) );
  OAI21_X1 U23201 ( .B1(n20291), .B2(n14099), .A(n20290), .ZN(P1_U2832) );
  INV_X1 U23202 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20992) );
  NAND2_X1 U23203 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20320), .ZN(n20314) );
  NOR2_X1 U23204 ( .A1(n20992), .A2(n20314), .ZN(n20296) );
  NAND2_X1 U23205 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20294) );
  OAI21_X1 U23206 ( .B1(n20294), .B2(n20293), .A(n20292), .ZN(n20313) );
  INV_X1 U23207 ( .A(n20313), .ZN(n20295) );
  MUX2_X1 U23208 ( .A(n20296), .B(n20295), .S(P1_REIP_REG_7__SCAN_IN), .Z(
        n20305) );
  AND2_X1 U23209 ( .A1(n20297), .A2(n20317), .ZN(n20304) );
  INV_X1 U23210 ( .A(n20298), .ZN(n20299) );
  NAND2_X1 U23211 ( .A1(n20299), .A2(n20334), .ZN(n20302) );
  NAND2_X1 U23212 ( .A1(n20335), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n20301) );
  NAND2_X1 U23213 ( .A1(n20340), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n20300) );
  NAND4_X1 U23214 ( .A1(n20302), .A2(n20301), .A3(n20322), .A4(n20300), .ZN(
        n20303) );
  NOR3_X1 U23215 ( .A1(n20305), .A2(n20304), .A3(n20303), .ZN(n20306) );
  OAI21_X1 U23216 ( .B1(n20307), .B2(n20330), .A(n20306), .ZN(P1_U2833) );
  INV_X1 U23217 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20355) );
  NOR2_X1 U23218 ( .A1(n20308), .A2(n20355), .ZN(n20309) );
  AOI211_X1 U23219 ( .C1(n20340), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20310), .B(n20309), .ZN(n20311) );
  OAI21_X1 U23220 ( .B1(n20325), .B2(n20312), .A(n20311), .ZN(n20316) );
  AOI21_X1 U23221 ( .B1(n20992), .B2(n20314), .A(n20313), .ZN(n20315) );
  AOI211_X1 U23222 ( .C1(n20353), .C2(n20317), .A(n20316), .B(n20315), .ZN(
        n20318) );
  OAI21_X1 U23223 ( .B1(n20319), .B2(n20330), .A(n20318), .ZN(P1_U2834) );
  INV_X1 U23224 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20989) );
  AOI22_X1 U23225 ( .A1(n20320), .A2(n20989), .B1(n20335), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n20329) );
  AOI22_X1 U23226 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20340), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20321), .ZN(n20323) );
  OAI211_X1 U23227 ( .C1(n20325), .C2(n20324), .A(n20323), .B(n20322), .ZN(
        n20326) );
  AOI21_X1 U23228 ( .B1(n20327), .B2(n20345), .A(n20326), .ZN(n20328) );
  OAI211_X1 U23229 ( .C1(n20331), .C2(n20330), .A(n20329), .B(n20328), .ZN(
        P1_U2835) );
  AOI21_X1 U23230 ( .B1(n20333), .B2(n21037), .A(n20332), .ZN(n20349) );
  AOI22_X1 U23231 ( .A1(n20335), .A2(P1_EBX_REG_2__SCAN_IN), .B1(n20334), .B2(
        n20396), .ZN(n20348) );
  NOR2_X1 U23232 ( .A1(n20336), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20344) );
  INV_X1 U23233 ( .A(n20337), .ZN(n20338) );
  AOI22_X1 U23234 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20340), .B1(
        n20339), .B2(n20338), .ZN(n20341) );
  OAI21_X1 U23235 ( .B1(n13223), .B2(n20342), .A(n20341), .ZN(n20343) );
  AOI211_X1 U23236 ( .C1(n20346), .C2(n20345), .A(n20344), .B(n20343), .ZN(
        n20347) );
  OAI211_X1 U23237 ( .C1(n20349), .C2(n20392), .A(n20348), .B(n20347), .ZN(
        P1_U2838) );
  AOI22_X1 U23238 ( .A1(n20353), .A2(n20352), .B1(n20351), .B2(n20350), .ZN(
        n20354) );
  OAI21_X1 U23239 ( .B1(n20356), .B2(n20355), .A(n20354), .ZN(P1_U2866) );
  AOI22_X1 U23240 ( .A1(n20357), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20407), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20366) );
  OR2_X1 U23241 ( .A1(n20359), .A2(n20358), .ZN(n20360) );
  NAND2_X1 U23242 ( .A1(n20361), .A2(n20360), .ZN(n20376) );
  OAI22_X1 U23243 ( .A1(n20376), .A2(n20363), .B1(n20422), .B2(n20362), .ZN(
        n20364) );
  INV_X1 U23244 ( .A(n20364), .ZN(n20365) );
  OAI211_X1 U23245 ( .C1(n20368), .C2(n20367), .A(n20366), .B(n20365), .ZN(
        P1_U2995) );
  NOR2_X1 U23246 ( .A1(n20370), .A2(n20369), .ZN(n20395) );
  OAI21_X1 U23247 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20372), .A(
        n20371), .ZN(n20389) );
  AOI211_X1 U23248 ( .C1(n20403), .C2(n20373), .A(n20395), .B(n20389), .ZN(
        n20386) );
  AOI22_X1 U23249 ( .A1(n20407), .A2(P1_REIP_REG_4__SCAN_IN), .B1(n20406), 
        .B2(n20374), .ZN(n20380) );
  AOI211_X1 U23250 ( .C1(n20381), .C2(n20387), .A(n20388), .B(n20375), .ZN(
        n20378) );
  NOR2_X1 U23251 ( .A1(n20376), .A2(n20408), .ZN(n20377) );
  NOR2_X1 U23252 ( .A1(n20378), .A2(n20377), .ZN(n20379) );
  OAI211_X1 U23253 ( .C1(n20386), .C2(n20381), .A(n20380), .B(n20379), .ZN(
        P1_U3027) );
  INV_X1 U23254 ( .A(n20382), .ZN(n20383) );
  AOI222_X1 U23255 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n20407), .B1(n20406), 
        .B2(n20384), .C1(n20399), .C2(n20383), .ZN(n20385) );
  OAI221_X1 U23256 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20388), .C1(
        n20387), .C2(n20386), .A(n20385), .ZN(P1_U3028) );
  INV_X1 U23257 ( .A(n20389), .ZN(n20404) );
  NAND2_X1 U23258 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20391) );
  NAND2_X1 U23259 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20390), .ZN(
        n20410) );
  OAI22_X1 U23260 ( .A1(n20393), .A2(n20392), .B1(n20391), .B2(n20410), .ZN(
        n20394) );
  AOI211_X1 U23261 ( .C1(n20406), .C2(n20396), .A(n20395), .B(n20394), .ZN(
        n20402) );
  INV_X1 U23262 ( .A(n20397), .ZN(n20400) );
  AOI22_X1 U23263 ( .A1(n20400), .A2(n20399), .B1(n20398), .B2(n20403), .ZN(
        n20401) );
  OAI211_X1 U23264 ( .C1(n20404), .C2(n20403), .A(n20402), .B(n20401), .ZN(
        P1_U3029) );
  AOI22_X1 U23265 ( .A1(n20407), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n20406), 
        .B2(n20405), .ZN(n20415) );
  NOR2_X1 U23266 ( .A1(n20409), .A2(n20408), .ZN(n20413) );
  AOI21_X1 U23267 ( .B1(n20411), .B2(n20410), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20412) );
  AOI21_X1 U23268 ( .B1(n20413), .B2(n13656), .A(n20412), .ZN(n20414) );
  OAI211_X1 U23269 ( .C1(n20416), .C2(n9877), .A(n20415), .B(n20414), .ZN(
        P1_U3030) );
  NOR2_X1 U23270 ( .A1(n20418), .A2(n20417), .ZN(P1_U3032) );
  NOR2_X2 U23271 ( .A1(n20422), .A2(n20421), .ZN(n20459) );
  AOI22_X1 U23272 ( .A1(DATAI_16_), .A2(n20420), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20459), .ZN(n20914) );
  NOR2_X2 U23273 ( .A1(n20458), .A2(n11170), .ZN(n20901) );
  NOR3_X1 U23274 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20471) );
  INV_X1 U23275 ( .A(n20471), .ZN(n20468) );
  NOR2_X1 U23276 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20468), .ZN(
        n20461) );
  NAND2_X1 U23277 ( .A1(n9702), .A2(n20784), .ZN(n20760) );
  AOI22_X1 U23278 ( .A1(DATAI_24_), .A2(n20420), .B1(BUF1_REG_24__SCAN_IN), 
        .B2(n20459), .ZN(n20863) );
  INV_X1 U23279 ( .A(n20863), .ZN(n20911) );
  AOI22_X1 U23280 ( .A1(n20901), .A2(n20461), .B1(n20460), .B2(n20911), .ZN(
        n20434) );
  NAND2_X1 U23281 ( .A1(n20430), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20846) );
  INV_X1 U23282 ( .A(n20846), .ZN(n20424) );
  AOI21_X1 U23283 ( .B1(n20492), .B2(n20960), .A(n20852), .ZN(n20425) );
  NOR2_X1 U23284 ( .A1(n20425), .A2(n20903), .ZN(n20429) );
  INV_X1 U23285 ( .A(n13223), .ZN(n20666) );
  OR2_X1 U23286 ( .A1(n20426), .A2(n20666), .ZN(n20494) );
  INV_X1 U23287 ( .A(n9697), .ZN(n20854) );
  OR2_X1 U23288 ( .A1(n20494), .A2(n20854), .ZN(n20431) );
  NAND2_X1 U23289 ( .A1(n20725), .A2(n20668), .ZN(n20554) );
  AOI22_X1 U23290 ( .A1(n20429), .A2(n20431), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20554), .ZN(n20427) );
  OAI211_X1 U23291 ( .C1(n20461), .C2(n20674), .A(n20727), .B(n20427), .ZN(
        n20464) );
  NOR2_X2 U23292 ( .A1(n20428), .A2(n20557), .ZN(n20900) );
  INV_X1 U23293 ( .A(n20429), .ZN(n20432) );
  NOR2_X1 U23294 ( .A1(n20430), .A2(n20966), .ZN(n20558) );
  INV_X1 U23295 ( .A(n20558), .ZN(n20729) );
  OAI22_X1 U23296 ( .A1(n20432), .A2(n20431), .B1(n20729), .B2(n20554), .ZN(
        n20463) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20464), .B1(
        n20900), .B2(n20463), .ZN(n20433) );
  OAI211_X1 U23298 ( .C1(n20914), .C2(n20492), .A(n20434), .B(n20433), .ZN(
        P1_U3033) );
  NOR2_X2 U23299 ( .A1(n20458), .A2(n11968), .ZN(n20916) );
  AOI22_X1 U23300 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20459), .B1(DATAI_25_), 
        .B2(n20420), .ZN(n20867) );
  INV_X1 U23301 ( .A(n20867), .ZN(n20917) );
  AOI22_X1 U23302 ( .A1(n20916), .A2(n20461), .B1(n20460), .B2(n20917), .ZN(
        n20437) );
  NOR2_X2 U23303 ( .A1(n20435), .A2(n20557), .ZN(n20915) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20464), .B1(
        n20915), .B2(n20463), .ZN(n20436) );
  OAI211_X1 U23305 ( .C1(n20920), .C2(n20492), .A(n20437), .B(n20436), .ZN(
        P1_U3034) );
  AOI22_X1 U23306 ( .A1(DATAI_18_), .A2(n20420), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20459), .ZN(n20926) );
  NOR2_X2 U23307 ( .A1(n20458), .A2(n20438), .ZN(n20922) );
  AOI22_X1 U23308 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20459), .B1(DATAI_26_), 
        .B2(n20420), .ZN(n20871) );
  INV_X1 U23309 ( .A(n20871), .ZN(n20923) );
  AOI22_X1 U23310 ( .A1(n20922), .A2(n20461), .B1(n20460), .B2(n20923), .ZN(
        n20441) );
  NOR2_X2 U23311 ( .A1(n20439), .A2(n20557), .ZN(n20921) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20464), .B1(
        n20921), .B2(n20463), .ZN(n20440) );
  OAI211_X1 U23313 ( .C1(n20926), .C2(n20492), .A(n20441), .B(n20440), .ZN(
        P1_U3035) );
  AOI22_X1 U23314 ( .A1(DATAI_19_), .A2(n20420), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20459), .ZN(n20932) );
  NOR2_X2 U23315 ( .A1(n20458), .A2(n20442), .ZN(n20928) );
  AOI22_X1 U23316 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20459), .B1(DATAI_27_), 
        .B2(n20420), .ZN(n20875) );
  INV_X1 U23317 ( .A(n20875), .ZN(n20929) );
  AOI22_X1 U23318 ( .A1(n20928), .A2(n20461), .B1(n20460), .B2(n20929), .ZN(
        n20445) );
  NOR2_X2 U23319 ( .A1(n20443), .A2(n20557), .ZN(n20927) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20464), .B1(
        n20927), .B2(n20463), .ZN(n20444) );
  OAI211_X1 U23321 ( .C1(n20932), .C2(n20492), .A(n20445), .B(n20444), .ZN(
        P1_U3036) );
  AOI22_X1 U23322 ( .A1(DATAI_20_), .A2(n20420), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20459), .ZN(n20938) );
  NOR2_X2 U23323 ( .A1(n20458), .A2(n20446), .ZN(n20934) );
  AOI22_X1 U23324 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20459), .B1(DATAI_28_), 
        .B2(n20420), .ZN(n20879) );
  INV_X1 U23325 ( .A(n20879), .ZN(n20935) );
  AOI22_X1 U23326 ( .A1(n20934), .A2(n20461), .B1(n20460), .B2(n20935), .ZN(
        n20449) );
  NOR2_X2 U23327 ( .A1(n20447), .A2(n20557), .ZN(n20933) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20464), .B1(
        n20933), .B2(n20463), .ZN(n20448) );
  OAI211_X1 U23329 ( .C1(n20938), .C2(n20492), .A(n20449), .B(n20448), .ZN(
        P1_U3037) );
  AOI22_X1 U23330 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20459), .B1(DATAI_21_), 
        .B2(n20420), .ZN(n20944) );
  NOR2_X2 U23331 ( .A1(n20458), .A2(n20450), .ZN(n20939) );
  AOI22_X1 U23332 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20459), .B1(DATAI_29_), 
        .B2(n20420), .ZN(n20883) );
  INV_X1 U23333 ( .A(n20883), .ZN(n20941) );
  AOI22_X1 U23334 ( .A1(n20939), .A2(n20461), .B1(n20460), .B2(n20941), .ZN(
        n20453) );
  NOR2_X2 U23335 ( .A1(n20557), .A2(n20451), .ZN(n20940) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20464), .B1(
        n20940), .B2(n20463), .ZN(n20452) );
  OAI211_X1 U23337 ( .C1(n20944), .C2(n20492), .A(n20453), .B(n20452), .ZN(
        P1_U3038) );
  AOI22_X1 U23338 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20459), .B1(DATAI_22_), 
        .B2(n20420), .ZN(n20950) );
  NOR2_X2 U23339 ( .A1(n20458), .A2(n10038), .ZN(n20945) );
  AOI22_X1 U23340 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20459), .B1(DATAI_30_), 
        .B2(n20420), .ZN(n20887) );
  INV_X1 U23341 ( .A(n20887), .ZN(n20947) );
  AOI22_X1 U23342 ( .A1(n20945), .A2(n20461), .B1(n20460), .B2(n20947), .ZN(
        n20456) );
  NOR2_X2 U23343 ( .A1(n20557), .A2(n20454), .ZN(n20946) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20464), .B1(
        n20946), .B2(n20463), .ZN(n20455) );
  OAI211_X1 U23345 ( .C1(n20950), .C2(n20492), .A(n20456), .B(n20455), .ZN(
        P1_U3039) );
  AOI22_X1 U23346 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20459), .B1(DATAI_23_), 
        .B2(n20420), .ZN(n20961) );
  NOR2_X2 U23347 ( .A1(n20458), .A2(n20457), .ZN(n20952) );
  AOI22_X1 U23348 ( .A1(DATAI_31_), .A2(n20420), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20459), .ZN(n20895) );
  INV_X1 U23349 ( .A(n20895), .ZN(n20955) );
  AOI22_X1 U23350 ( .A1(n20952), .A2(n20461), .B1(n20460), .B2(n20955), .ZN(
        n20466) );
  NOR2_X2 U23351 ( .A1(n20557), .A2(n20462), .ZN(n20954) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20464), .B1(
        n20954), .B2(n20463), .ZN(n20465) );
  OAI211_X1 U23353 ( .C1(n20961), .C2(n20492), .A(n20466), .B(n20465), .ZN(
        P1_U3040) );
  NOR2_X1 U23354 ( .A1(n20820), .A2(n20468), .ZN(n20487) );
  INV_X1 U23355 ( .A(n20494), .ZN(n20524) );
  INV_X1 U23356 ( .A(n20467), .ZN(n20821) );
  AOI21_X1 U23357 ( .B1(n20524), .B2(n20821), .A(n20487), .ZN(n20469) );
  OAI22_X1 U23358 ( .A1(n20469), .A2(n20903), .B1(n20468), .B2(n20966), .ZN(
        n20488) );
  AOI22_X1 U23359 ( .A1(n20901), .A2(n20487), .B1(n20900), .B2(n20488), .ZN(
        n20473) );
  OAI211_X1 U23360 ( .C1(n20526), .C2(n20852), .A(n20909), .B(n20469), .ZN(
        n20470) );
  OAI211_X1 U23361 ( .C1(n20909), .C2(n20471), .A(n20908), .B(n20470), .ZN(
        n20489) );
  INV_X1 U23362 ( .A(n20914), .ZN(n20860) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20489), .B1(
        n20517), .B2(n20860), .ZN(n20472) );
  OAI211_X1 U23364 ( .C1(n20863), .C2(n20492), .A(n20473), .B(n20472), .ZN(
        P1_U3041) );
  AOI22_X1 U23365 ( .A1(n20916), .A2(n20487), .B1(n20915), .B2(n20488), .ZN(
        n20475) );
  INV_X1 U23366 ( .A(n20492), .ZN(n20476) );
  AOI22_X1 U23367 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20489), .B1(
        n20476), .B2(n20917), .ZN(n20474) );
  OAI211_X1 U23368 ( .C1(n20920), .C2(n20513), .A(n20475), .B(n20474), .ZN(
        P1_U3042) );
  AOI22_X1 U23369 ( .A1(n20922), .A2(n20487), .B1(n20921), .B2(n20488), .ZN(
        n20478) );
  AOI22_X1 U23370 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20489), .B1(
        n20476), .B2(n20923), .ZN(n20477) );
  OAI211_X1 U23371 ( .C1(n20926), .C2(n20513), .A(n20478), .B(n20477), .ZN(
        P1_U3043) );
  AOI22_X1 U23372 ( .A1(n20928), .A2(n20487), .B1(n20927), .B2(n20488), .ZN(
        n20480) );
  INV_X1 U23373 ( .A(n20932), .ZN(n20872) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20489), .B1(
        n20517), .B2(n20872), .ZN(n20479) );
  OAI211_X1 U23375 ( .C1(n20875), .C2(n20492), .A(n20480), .B(n20479), .ZN(
        P1_U3044) );
  AOI22_X1 U23376 ( .A1(n20934), .A2(n20487), .B1(n20933), .B2(n20488), .ZN(
        n20482) );
  INV_X1 U23377 ( .A(n20938), .ZN(n20876) );
  AOI22_X1 U23378 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20489), .B1(
        n20517), .B2(n20876), .ZN(n20481) );
  OAI211_X1 U23379 ( .C1(n20879), .C2(n20492), .A(n20482), .B(n20481), .ZN(
        P1_U3045) );
  AOI22_X1 U23380 ( .A1(n20940), .A2(n20488), .B1(n20939), .B2(n20487), .ZN(
        n20484) );
  INV_X1 U23381 ( .A(n20944), .ZN(n20880) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20489), .B1(
        n20517), .B2(n20880), .ZN(n20483) );
  OAI211_X1 U23383 ( .C1(n20883), .C2(n20492), .A(n20484), .B(n20483), .ZN(
        P1_U3046) );
  AOI22_X1 U23384 ( .A1(n20946), .A2(n20488), .B1(n20945), .B2(n20487), .ZN(
        n20486) );
  INV_X1 U23385 ( .A(n20950), .ZN(n20884) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20489), .B1(
        n20517), .B2(n20884), .ZN(n20485) );
  OAI211_X1 U23387 ( .C1(n20887), .C2(n20492), .A(n20486), .B(n20485), .ZN(
        P1_U3047) );
  AOI22_X1 U23388 ( .A1(n20954), .A2(n20488), .B1(n20952), .B2(n20487), .ZN(
        n20491) );
  INV_X1 U23389 ( .A(n20961), .ZN(n20890) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20489), .B1(
        n20517), .B2(n20890), .ZN(n20490) );
  OAI211_X1 U23391 ( .C1(n20895), .C2(n20492), .A(n20491), .B(n20490), .ZN(
        P1_U3048) );
  NAND3_X1 U23392 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20786), .A3(
        n20787), .ZN(n20529) );
  NOR2_X1 U23393 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20529), .ZN(
        n20516) );
  AOI22_X1 U23394 ( .A1(n20517), .A2(n20911), .B1(n20901), .B2(n20516), .ZN(
        n20502) );
  OAI21_X1 U23395 ( .B1(n20547), .B2(n20517), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20493) );
  NAND2_X1 U23396 ( .A1(n20493), .A2(n20909), .ZN(n20500) );
  INV_X1 U23397 ( .A(n20500), .ZN(n20496) );
  OR2_X1 U23398 ( .A1(n20494), .A2(n9697), .ZN(n20499) );
  INV_X1 U23399 ( .A(n20516), .ZN(n20495) );
  AOI22_X1 U23400 ( .A1(n20496), .A2(n20499), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20495), .ZN(n20497) );
  OAI21_X1 U23401 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20725), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20609) );
  NAND3_X1 U23402 ( .A1(n20727), .A2(n20497), .A3(n20609), .ZN(n20519) );
  INV_X1 U23403 ( .A(n20725), .ZN(n20498) );
  NAND2_X1 U23404 ( .A1(n20498), .A2(n20786), .ZN(n20612) );
  OAI22_X1 U23405 ( .A1(n20500), .A2(n20499), .B1(n20729), .B2(n20612), .ZN(
        n20518) );
  AOI22_X1 U23406 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20519), .B1(
        n20900), .B2(n20518), .ZN(n20501) );
  OAI211_X1 U23407 ( .C1(n20914), .C2(n20546), .A(n20502), .B(n20501), .ZN(
        P1_U3049) );
  AOI22_X1 U23408 ( .A1(n20517), .A2(n20917), .B1(n20916), .B2(n20516), .ZN(
        n20504) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20519), .B1(
        n20915), .B2(n20518), .ZN(n20503) );
  OAI211_X1 U23410 ( .C1(n20920), .C2(n20546), .A(n20504), .B(n20503), .ZN(
        P1_U3050) );
  INV_X1 U23411 ( .A(n20926), .ZN(n20868) );
  AOI22_X1 U23412 ( .A1(n20547), .A2(n20868), .B1(n20922), .B2(n20516), .ZN(
        n20506) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20519), .B1(
        n20921), .B2(n20518), .ZN(n20505) );
  OAI211_X1 U23414 ( .C1(n20871), .C2(n20513), .A(n20506), .B(n20505), .ZN(
        P1_U3051) );
  AOI22_X1 U23415 ( .A1(n20547), .A2(n20872), .B1(n20928), .B2(n20516), .ZN(
        n20508) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20519), .B1(
        n20927), .B2(n20518), .ZN(n20507) );
  OAI211_X1 U23417 ( .C1(n20875), .C2(n20513), .A(n20508), .B(n20507), .ZN(
        P1_U3052) );
  AOI22_X1 U23418 ( .A1(n20547), .A2(n20876), .B1(n20934), .B2(n20516), .ZN(
        n20510) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20519), .B1(
        n20933), .B2(n20518), .ZN(n20509) );
  OAI211_X1 U23420 ( .C1(n20879), .C2(n20513), .A(n20510), .B(n20509), .ZN(
        P1_U3053) );
  AOI22_X1 U23421 ( .A1(n20547), .A2(n20880), .B1(n20939), .B2(n20516), .ZN(
        n20512) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20519), .B1(
        n20940), .B2(n20518), .ZN(n20511) );
  OAI211_X1 U23423 ( .C1(n20883), .C2(n20513), .A(n20512), .B(n20511), .ZN(
        P1_U3054) );
  AOI22_X1 U23424 ( .A1(n20517), .A2(n20947), .B1(n20945), .B2(n20516), .ZN(
        n20515) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20519), .B1(
        n20946), .B2(n20518), .ZN(n20514) );
  OAI211_X1 U23426 ( .C1(n20950), .C2(n20546), .A(n20515), .B(n20514), .ZN(
        P1_U3055) );
  AOI22_X1 U23427 ( .A1(n20517), .A2(n20955), .B1(n20952), .B2(n20516), .ZN(
        n20521) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20519), .B1(
        n20954), .B2(n20518), .ZN(n20520) );
  OAI211_X1 U23429 ( .C1(n20961), .C2(n20546), .A(n20521), .B(n20520), .ZN(
        P1_U3056) );
  AOI22_X1 U23430 ( .A1(n20547), .A2(n20911), .B1(n20901), .B2(n10186), .ZN(
        n20533) );
  NOR2_X1 U23431 ( .A1(n20523), .A2(n20522), .ZN(n20897) );
  AOI21_X1 U23432 ( .B1(n20524), .B2(n20897), .A(n10186), .ZN(n20530) );
  AOI21_X1 U23433 ( .B1(n20526), .B2(n20909), .A(n20525), .ZN(n20531) );
  INV_X1 U23434 ( .A(n20531), .ZN(n20527) );
  AOI22_X1 U23435 ( .A1(n20530), .A2(n20527), .B1(n20903), .B2(n20529), .ZN(
        n20528) );
  NAND2_X1 U23436 ( .A1(n20908), .A2(n20528), .ZN(n20549) );
  OAI22_X1 U23437 ( .A1(n20531), .A2(n20530), .B1(n20966), .B2(n20529), .ZN(
        n20548) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20549), .B1(
        n20900), .B2(n20548), .ZN(n20532) );
  OAI211_X1 U23439 ( .C1(n20914), .C2(n20572), .A(n20533), .B(n20532), .ZN(
        P1_U3057) );
  AOI22_X1 U23440 ( .A1(n20547), .A2(n20917), .B1(n20916), .B2(n10186), .ZN(
        n20535) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20549), .B1(
        n20915), .B2(n20548), .ZN(n20534) );
  OAI211_X1 U23442 ( .C1(n20920), .C2(n20572), .A(n20535), .B(n20534), .ZN(
        P1_U3058) );
  AOI22_X1 U23443 ( .A1(n20577), .A2(n20868), .B1(n20922), .B2(n10186), .ZN(
        n20537) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20549), .B1(
        n20921), .B2(n20548), .ZN(n20536) );
  OAI211_X1 U23445 ( .C1(n20871), .C2(n20546), .A(n20537), .B(n20536), .ZN(
        P1_U3059) );
  AOI22_X1 U23446 ( .A1(n20577), .A2(n20872), .B1(n20928), .B2(n10186), .ZN(
        n20539) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20549), .B1(
        n20927), .B2(n20548), .ZN(n20538) );
  OAI211_X1 U23448 ( .C1(n20875), .C2(n20546), .A(n20539), .B(n20538), .ZN(
        P1_U3060) );
  AOI22_X1 U23449 ( .A1(n20577), .A2(n20876), .B1(n20934), .B2(n10186), .ZN(
        n20541) );
  AOI22_X1 U23450 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20549), .B1(
        n20933), .B2(n20548), .ZN(n20540) );
  OAI211_X1 U23451 ( .C1(n20879), .C2(n20546), .A(n20541), .B(n20540), .ZN(
        P1_U3061) );
  AOI22_X1 U23452 ( .A1(n20547), .A2(n20941), .B1(n20939), .B2(n10186), .ZN(
        n20543) );
  AOI22_X1 U23453 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20549), .B1(
        n20940), .B2(n20548), .ZN(n20542) );
  OAI211_X1 U23454 ( .C1(n20944), .C2(n20572), .A(n20543), .B(n20542), .ZN(
        P1_U3062) );
  AOI22_X1 U23455 ( .A1(n20577), .A2(n20884), .B1(n20945), .B2(n10186), .ZN(
        n20545) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20549), .B1(
        n20946), .B2(n20548), .ZN(n20544) );
  OAI211_X1 U23457 ( .C1(n20887), .C2(n20546), .A(n20545), .B(n20544), .ZN(
        P1_U3063) );
  AOI22_X1 U23458 ( .A1(n20547), .A2(n20955), .B1(n20952), .B2(n10186), .ZN(
        n20551) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20549), .B1(
        n20954), .B2(n20548), .ZN(n20550) );
  OAI211_X1 U23460 ( .C1(n20961), .C2(n20572), .A(n20551), .B(n20550), .ZN(
        P1_U3064) );
  NOR3_X1 U23461 ( .A1(n20787), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20585) );
  INV_X1 U23462 ( .A(n20585), .ZN(n20581) );
  NOR2_X1 U23463 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20581), .ZN(
        n20575) );
  NOR2_X1 U23464 ( .A1(n13223), .A2(n20552), .ZN(n20637) );
  NAND3_X1 U23465 ( .A1(n20637), .A2(n20909), .A3(n9697), .ZN(n20553) );
  OAI21_X1 U23466 ( .B1(n20846), .B2(n20554), .A(n20553), .ZN(n20576) );
  AOI22_X1 U23467 ( .A1(n20901), .A2(n20575), .B1(n20900), .B2(n20576), .ZN(
        n20561) );
  INV_X1 U23468 ( .A(n20637), .ZN(n20556) );
  OAI21_X1 U23469 ( .B1(n20577), .B2(n20603), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20555) );
  OAI21_X1 U23470 ( .B1(n20854), .B2(n20556), .A(n20555), .ZN(n20559) );
  OAI221_X1 U23471 ( .B1(n20575), .B2(n20674), .C1(n20575), .C2(n20559), .A(
        n20857), .ZN(n20578) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20911), .ZN(n20560) );
  OAI211_X1 U23473 ( .C1(n20914), .C2(n20600), .A(n20561), .B(n20560), .ZN(
        P1_U3065) );
  AOI22_X1 U23474 ( .A1(n20916), .A2(n20575), .B1(n20915), .B2(n20576), .ZN(
        n20563) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20917), .ZN(n20562) );
  OAI211_X1 U23476 ( .C1(n20920), .C2(n20600), .A(n20563), .B(n20562), .ZN(
        P1_U3066) );
  AOI22_X1 U23477 ( .A1(n20922), .A2(n20575), .B1(n20921), .B2(n20576), .ZN(
        n20565) );
  AOI22_X1 U23478 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20578), .B1(
        n20603), .B2(n20868), .ZN(n20564) );
  OAI211_X1 U23479 ( .C1(n20871), .C2(n20572), .A(n20565), .B(n20564), .ZN(
        P1_U3067) );
  AOI22_X1 U23480 ( .A1(n20928), .A2(n20575), .B1(n20927), .B2(n20576), .ZN(
        n20567) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20578), .B1(
        n20603), .B2(n20872), .ZN(n20566) );
  OAI211_X1 U23482 ( .C1(n20875), .C2(n20572), .A(n20567), .B(n20566), .ZN(
        P1_U3068) );
  AOI22_X1 U23483 ( .A1(n20934), .A2(n20575), .B1(n20933), .B2(n20576), .ZN(
        n20569) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20578), .B1(
        n20603), .B2(n20876), .ZN(n20568) );
  OAI211_X1 U23485 ( .C1(n20879), .C2(n20572), .A(n20569), .B(n20568), .ZN(
        P1_U3069) );
  AOI22_X1 U23486 ( .A1(n20940), .A2(n20576), .B1(n20939), .B2(n20575), .ZN(
        n20571) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20578), .B1(
        n20603), .B2(n20880), .ZN(n20570) );
  OAI211_X1 U23488 ( .C1(n20883), .C2(n20572), .A(n20571), .B(n20570), .ZN(
        P1_U3070) );
  AOI22_X1 U23489 ( .A1(n20946), .A2(n20576), .B1(n20945), .B2(n20575), .ZN(
        n20574) );
  AOI22_X1 U23490 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20947), .ZN(n20573) );
  OAI211_X1 U23491 ( .C1(n20950), .C2(n20600), .A(n20574), .B(n20573), .ZN(
        P1_U3071) );
  AOI22_X1 U23492 ( .A1(n20954), .A2(n20576), .B1(n20952), .B2(n20575), .ZN(
        n20580) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20955), .ZN(n20579) );
  OAI211_X1 U23494 ( .C1(n20961), .C2(n20600), .A(n20580), .B(n20579), .ZN(
        P1_U3072) );
  NOR2_X1 U23495 ( .A1(n20820), .A2(n20581), .ZN(n20601) );
  AOI21_X1 U23496 ( .B1(n20637), .B2(n20821), .A(n20601), .ZN(n20582) );
  OAI22_X1 U23497 ( .A1(n20582), .A2(n20903), .B1(n20581), .B2(n20966), .ZN(
        n20602) );
  AOI22_X1 U23498 ( .A1(n20901), .A2(n20601), .B1(n20900), .B2(n20602), .ZN(
        n20587) );
  INV_X1 U23499 ( .A(n20789), .ZN(n20583) );
  OAI21_X1 U23500 ( .B1(n20641), .B2(n20583), .A(n20582), .ZN(n20584) );
  OAI211_X1 U23501 ( .C1(n20909), .C2(n20585), .A(n20908), .B(n20584), .ZN(
        n20604) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20604), .B1(
        n20603), .B2(n20911), .ZN(n20586) );
  OAI211_X1 U23503 ( .C1(n20914), .C2(n20629), .A(n20587), .B(n20586), .ZN(
        P1_U3073) );
  AOI22_X1 U23504 ( .A1(n20916), .A2(n20601), .B1(n20915), .B2(n20602), .ZN(
        n20589) );
  INV_X1 U23505 ( .A(n20920), .ZN(n20864) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20604), .B1(
        n20630), .B2(n20864), .ZN(n20588) );
  OAI211_X1 U23507 ( .C1(n20867), .C2(n20600), .A(n20589), .B(n20588), .ZN(
        P1_U3074) );
  AOI22_X1 U23508 ( .A1(n20922), .A2(n20601), .B1(n20921), .B2(n20602), .ZN(
        n20591) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20604), .B1(
        n20630), .B2(n20868), .ZN(n20590) );
  OAI211_X1 U23510 ( .C1(n20871), .C2(n20600), .A(n20591), .B(n20590), .ZN(
        P1_U3075) );
  AOI22_X1 U23511 ( .A1(n20928), .A2(n20601), .B1(n20927), .B2(n20602), .ZN(
        n20593) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20604), .B1(
        n20630), .B2(n20872), .ZN(n20592) );
  OAI211_X1 U23513 ( .C1(n20875), .C2(n20600), .A(n20593), .B(n20592), .ZN(
        P1_U3076) );
  AOI22_X1 U23514 ( .A1(n20934), .A2(n20601), .B1(n20933), .B2(n20602), .ZN(
        n20595) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20604), .B1(
        n20603), .B2(n20935), .ZN(n20594) );
  OAI211_X1 U23516 ( .C1(n20938), .C2(n20629), .A(n20595), .B(n20594), .ZN(
        P1_U3077) );
  AOI22_X1 U23517 ( .A1(n20940), .A2(n20602), .B1(n20939), .B2(n20601), .ZN(
        n20597) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20604), .B1(
        n20603), .B2(n20941), .ZN(n20596) );
  OAI211_X1 U23519 ( .C1(n20944), .C2(n20629), .A(n20597), .B(n20596), .ZN(
        P1_U3078) );
  AOI22_X1 U23520 ( .A1(n20946), .A2(n20602), .B1(n20945), .B2(n20601), .ZN(
        n20599) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20604), .B1(
        n20630), .B2(n20884), .ZN(n20598) );
  OAI211_X1 U23522 ( .C1(n20887), .C2(n20600), .A(n20599), .B(n20598), .ZN(
        P1_U3079) );
  AOI22_X1 U23523 ( .A1(n20954), .A2(n20602), .B1(n20952), .B2(n20601), .ZN(
        n20606) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20604), .B1(
        n20603), .B2(n20955), .ZN(n20605) );
  OAI211_X1 U23525 ( .C1(n20961), .C2(n20629), .A(n20606), .B(n20605), .ZN(
        P1_U3080) );
  NAND2_X1 U23526 ( .A1(n20820), .A2(n11329), .ZN(n20608) );
  INV_X1 U23527 ( .A(n20608), .ZN(n20631) );
  AOI22_X1 U23528 ( .A1(n20901), .A2(n20631), .B1(n20654), .B2(n20860), .ZN(
        n20616) );
  NAND2_X1 U23529 ( .A1(n20663), .A2(n20629), .ZN(n20607) );
  AOI21_X1 U23530 ( .B1(n20607), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20903), 
        .ZN(n20611) );
  NAND2_X1 U23531 ( .A1(n20637), .A2(n20854), .ZN(n20613) );
  AOI22_X1 U23532 ( .A1(n20611), .A2(n20613), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20608), .ZN(n20610) );
  NAND3_X1 U23533 ( .A1(n20857), .A2(n20610), .A3(n20609), .ZN(n20633) );
  INV_X1 U23534 ( .A(n20611), .ZN(n20614) );
  OAI22_X1 U23535 ( .A1(n20614), .A2(n20613), .B1(n20612), .B2(n20846), .ZN(
        n20632) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20633), .B1(
        n20900), .B2(n20632), .ZN(n20615) );
  OAI211_X1 U23537 ( .C1(n20863), .C2(n20629), .A(n20616), .B(n20615), .ZN(
        P1_U3081) );
  AOI22_X1 U23538 ( .A1(n20916), .A2(n20631), .B1(n20630), .B2(n20917), .ZN(
        n20618) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20633), .B1(
        n20915), .B2(n20632), .ZN(n20617) );
  OAI211_X1 U23540 ( .C1(n20920), .C2(n20663), .A(n20618), .B(n20617), .ZN(
        P1_U3082) );
  AOI22_X1 U23541 ( .A1(n20922), .A2(n20631), .B1(n20654), .B2(n20868), .ZN(
        n20620) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20633), .B1(
        n20921), .B2(n20632), .ZN(n20619) );
  OAI211_X1 U23543 ( .C1(n20871), .C2(n20629), .A(n20620), .B(n20619), .ZN(
        P1_U3083) );
  AOI22_X1 U23544 ( .A1(n20928), .A2(n20631), .B1(n20630), .B2(n20929), .ZN(
        n20622) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20633), .B1(
        n20927), .B2(n20632), .ZN(n20621) );
  OAI211_X1 U23546 ( .C1(n20932), .C2(n20663), .A(n20622), .B(n20621), .ZN(
        P1_U3084) );
  AOI22_X1 U23547 ( .A1(n20934), .A2(n20631), .B1(n20630), .B2(n20935), .ZN(
        n20624) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20633), .B1(
        n20933), .B2(n20632), .ZN(n20623) );
  OAI211_X1 U23549 ( .C1(n20938), .C2(n20663), .A(n20624), .B(n20623), .ZN(
        P1_U3085) );
  AOI22_X1 U23550 ( .A1(n20939), .A2(n20631), .B1(n20630), .B2(n20941), .ZN(
        n20626) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20633), .B1(
        n20940), .B2(n20632), .ZN(n20625) );
  OAI211_X1 U23552 ( .C1(n20944), .C2(n20663), .A(n20626), .B(n20625), .ZN(
        P1_U3086) );
  AOI22_X1 U23553 ( .A1(n20945), .A2(n20631), .B1(n20654), .B2(n20884), .ZN(
        n20628) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20633), .B1(
        n20946), .B2(n20632), .ZN(n20627) );
  OAI211_X1 U23555 ( .C1(n20887), .C2(n20629), .A(n20628), .B(n20627), .ZN(
        P1_U3087) );
  AOI22_X1 U23556 ( .A1(n20952), .A2(n20631), .B1(n20630), .B2(n20955), .ZN(
        n20635) );
  AOI22_X1 U23557 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20633), .B1(
        n20954), .B2(n20632), .ZN(n20634) );
  OAI211_X1 U23558 ( .C1(n20961), .C2(n20663), .A(n20635), .B(n20634), .ZN(
        P1_U3088) );
  INV_X1 U23559 ( .A(n20636), .ZN(n20658) );
  AOI21_X1 U23560 ( .B1(n20637), .B2(n20897), .A(n20658), .ZN(n20639) );
  OAI22_X1 U23561 ( .A1(n20639), .A2(n20903), .B1(n20638), .B2(n20966), .ZN(
        n20659) );
  AOI22_X1 U23562 ( .A1(n20901), .A2(n20658), .B1(n20900), .B2(n20659), .ZN(
        n20643) );
  OAI21_X1 U23563 ( .B1(n11329), .B2(n20640), .A(n20908), .ZN(n20660) );
  OR2_X1 U23564 ( .A1(n20641), .A2(n20760), .ZN(n20657) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20660), .B1(
        n20691), .B2(n20860), .ZN(n20642) );
  OAI211_X1 U23566 ( .C1(n20863), .C2(n20663), .A(n20643), .B(n20642), .ZN(
        P1_U3089) );
  AOI22_X1 U23567 ( .A1(n20916), .A2(n20658), .B1(n20915), .B2(n20659), .ZN(
        n20645) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20660), .B1(
        n20654), .B2(n20917), .ZN(n20644) );
  OAI211_X1 U23569 ( .C1(n20920), .C2(n20657), .A(n20645), .B(n20644), .ZN(
        P1_U3090) );
  AOI22_X1 U23570 ( .A1(n20922), .A2(n20658), .B1(n20921), .B2(n20659), .ZN(
        n20647) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20660), .B1(
        n20691), .B2(n20868), .ZN(n20646) );
  OAI211_X1 U23572 ( .C1(n20871), .C2(n20663), .A(n20647), .B(n20646), .ZN(
        P1_U3091) );
  AOI22_X1 U23573 ( .A1(n20928), .A2(n20658), .B1(n20927), .B2(n20659), .ZN(
        n20649) );
  AOI22_X1 U23574 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20660), .B1(
        n20654), .B2(n20929), .ZN(n20648) );
  OAI211_X1 U23575 ( .C1(n20932), .C2(n20657), .A(n20649), .B(n20648), .ZN(
        P1_U3092) );
  AOI22_X1 U23576 ( .A1(n20934), .A2(n20658), .B1(n20933), .B2(n20659), .ZN(
        n20651) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20660), .B1(
        n20691), .B2(n20876), .ZN(n20650) );
  OAI211_X1 U23578 ( .C1(n20879), .C2(n20663), .A(n20651), .B(n20650), .ZN(
        P1_U3093) );
  AOI22_X1 U23579 ( .A1(n20940), .A2(n20659), .B1(n20939), .B2(n20658), .ZN(
        n20653) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20660), .B1(
        n20691), .B2(n20880), .ZN(n20652) );
  OAI211_X1 U23581 ( .C1(n20883), .C2(n20663), .A(n20653), .B(n20652), .ZN(
        P1_U3094) );
  AOI22_X1 U23582 ( .A1(n20946), .A2(n20659), .B1(n20945), .B2(n20658), .ZN(
        n20656) );
  AOI22_X1 U23583 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20660), .B1(
        n20654), .B2(n20947), .ZN(n20655) );
  OAI211_X1 U23584 ( .C1(n20950), .C2(n20657), .A(n20656), .B(n20655), .ZN(
        P1_U3095) );
  AOI22_X1 U23585 ( .A1(n20954), .A2(n20659), .B1(n20952), .B2(n20658), .ZN(
        n20662) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20660), .B1(
        n20691), .B2(n20890), .ZN(n20661) );
  OAI211_X1 U23587 ( .C1(n20895), .C2(n20663), .A(n20662), .B(n20661), .ZN(
        P1_U3096) );
  INV_X1 U23588 ( .A(n20664), .ZN(n20665) );
  NOR3_X1 U23589 ( .A1(n20786), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20699) );
  INV_X1 U23590 ( .A(n20699), .ZN(n20695) );
  NOR2_X1 U23591 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20695), .ZN(
        n20689) );
  AOI21_X1 U23592 ( .B1(n20754), .B2(n9697), .A(n20689), .ZN(n20671) );
  INV_X1 U23593 ( .A(n20668), .ZN(n20669) );
  NAND2_X1 U23594 ( .A1(n20669), .A2(n20725), .ZN(n20796) );
  OAI22_X1 U23595 ( .A1(n20671), .A2(n20903), .B1(n20729), .B2(n20796), .ZN(
        n20690) );
  AOI22_X1 U23596 ( .A1(n20901), .A2(n20689), .B1(n20900), .B2(n20690), .ZN(
        n20676) );
  INV_X1 U23597 ( .A(n20720), .ZN(n20670) );
  OAI21_X1 U23598 ( .B1(n20670), .B2(n20691), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20672) );
  NAND2_X1 U23599 ( .A1(n20672), .A2(n20671), .ZN(n20673) );
  AOI22_X1 U23600 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20692), .B1(
        n20691), .B2(n20911), .ZN(n20675) );
  OAI211_X1 U23601 ( .C1(n20914), .C2(n20720), .A(n20676), .B(n20675), .ZN(
        P1_U3097) );
  AOI22_X1 U23602 ( .A1(n20916), .A2(n20689), .B1(n20915), .B2(n20690), .ZN(
        n20678) );
  AOI22_X1 U23603 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20692), .B1(
        n20691), .B2(n20917), .ZN(n20677) );
  OAI211_X1 U23604 ( .C1(n20920), .C2(n20720), .A(n20678), .B(n20677), .ZN(
        P1_U3098) );
  AOI22_X1 U23605 ( .A1(n20922), .A2(n20689), .B1(n20921), .B2(n20690), .ZN(
        n20680) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20692), .B1(
        n20691), .B2(n20923), .ZN(n20679) );
  OAI211_X1 U23607 ( .C1(n20926), .C2(n20720), .A(n20680), .B(n20679), .ZN(
        P1_U3099) );
  AOI22_X1 U23608 ( .A1(n20928), .A2(n20689), .B1(n20927), .B2(n20690), .ZN(
        n20682) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20692), .B1(
        n20691), .B2(n20929), .ZN(n20681) );
  OAI211_X1 U23610 ( .C1(n20932), .C2(n20720), .A(n20682), .B(n20681), .ZN(
        P1_U3100) );
  AOI22_X1 U23611 ( .A1(n20934), .A2(n20689), .B1(n20933), .B2(n20690), .ZN(
        n20684) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20692), .B1(
        n20691), .B2(n20935), .ZN(n20683) );
  OAI211_X1 U23613 ( .C1(n20938), .C2(n20720), .A(n20684), .B(n20683), .ZN(
        P1_U3101) );
  AOI22_X1 U23614 ( .A1(n20940), .A2(n20690), .B1(n20939), .B2(n20689), .ZN(
        n20686) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20692), .B1(
        n20691), .B2(n20941), .ZN(n20685) );
  OAI211_X1 U23616 ( .C1(n20944), .C2(n20720), .A(n20686), .B(n20685), .ZN(
        P1_U3102) );
  AOI22_X1 U23617 ( .A1(n20946), .A2(n20690), .B1(n20945), .B2(n20689), .ZN(
        n20688) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20692), .B1(
        n20691), .B2(n20947), .ZN(n20687) );
  OAI211_X1 U23619 ( .C1(n20950), .C2(n20720), .A(n20688), .B(n20687), .ZN(
        P1_U3103) );
  AOI22_X1 U23620 ( .A1(n20954), .A2(n20690), .B1(n20952), .B2(n20689), .ZN(
        n20694) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20692), .B1(
        n20691), .B2(n20955), .ZN(n20693) );
  OAI211_X1 U23622 ( .C1(n20961), .C2(n20720), .A(n20694), .B(n20693), .ZN(
        P1_U3104) );
  NOR2_X1 U23623 ( .A1(n20820), .A2(n20695), .ZN(n20715) );
  AOI21_X1 U23624 ( .B1(n20754), .B2(n20821), .A(n20715), .ZN(n20696) );
  OAI22_X1 U23625 ( .A1(n20696), .A2(n20903), .B1(n20695), .B2(n20966), .ZN(
        n20716) );
  AOI22_X1 U23626 ( .A1(n20901), .A2(n20715), .B1(n20900), .B2(n20716), .ZN(
        n20702) );
  OAI211_X1 U23627 ( .C1(n20697), .C2(n20852), .A(n20909), .B(n20696), .ZN(
        n20698) );
  OAI211_X1 U23628 ( .C1(n20909), .C2(n20699), .A(n20908), .B(n20698), .ZN(
        n20717) );
  NAND2_X1 U23629 ( .A1(n20762), .A2(n20819), .ZN(n20752) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20717), .B1(
        n20744), .B2(n20860), .ZN(n20701) );
  OAI211_X1 U23631 ( .C1(n20863), .C2(n20720), .A(n20702), .B(n20701), .ZN(
        P1_U3105) );
  AOI22_X1 U23632 ( .A1(n20916), .A2(n20715), .B1(n20915), .B2(n20716), .ZN(
        n20704) );
  AOI22_X1 U23633 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20717), .B1(
        n20744), .B2(n20864), .ZN(n20703) );
  OAI211_X1 U23634 ( .C1(n20867), .C2(n20720), .A(n20704), .B(n20703), .ZN(
        P1_U3106) );
  AOI22_X1 U23635 ( .A1(n20922), .A2(n20715), .B1(n20921), .B2(n20716), .ZN(
        n20706) );
  AOI22_X1 U23636 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20717), .B1(
        n20744), .B2(n20868), .ZN(n20705) );
  OAI211_X1 U23637 ( .C1(n20871), .C2(n20720), .A(n20706), .B(n20705), .ZN(
        P1_U3107) );
  AOI22_X1 U23638 ( .A1(n20928), .A2(n20715), .B1(n20927), .B2(n20716), .ZN(
        n20708) );
  AOI22_X1 U23639 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20717), .B1(
        n20744), .B2(n20872), .ZN(n20707) );
  OAI211_X1 U23640 ( .C1(n20875), .C2(n20720), .A(n20708), .B(n20707), .ZN(
        P1_U3108) );
  AOI22_X1 U23641 ( .A1(n20934), .A2(n20715), .B1(n20933), .B2(n20716), .ZN(
        n20710) );
  AOI22_X1 U23642 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20717), .B1(
        n20744), .B2(n20876), .ZN(n20709) );
  OAI211_X1 U23643 ( .C1(n20879), .C2(n20720), .A(n20710), .B(n20709), .ZN(
        P1_U3109) );
  AOI22_X1 U23644 ( .A1(n20940), .A2(n20716), .B1(n20939), .B2(n20715), .ZN(
        n20712) );
  AOI22_X1 U23645 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20717), .B1(
        n20744), .B2(n20880), .ZN(n20711) );
  OAI211_X1 U23646 ( .C1(n20883), .C2(n20720), .A(n20712), .B(n20711), .ZN(
        P1_U3110) );
  AOI22_X1 U23647 ( .A1(n20946), .A2(n20716), .B1(n20945), .B2(n20715), .ZN(
        n20714) );
  AOI22_X1 U23648 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20717), .B1(
        n20744), .B2(n20884), .ZN(n20713) );
  OAI211_X1 U23649 ( .C1(n20887), .C2(n20720), .A(n20714), .B(n20713), .ZN(
        P1_U3111) );
  AOI22_X1 U23650 ( .A1(n20954), .A2(n20716), .B1(n20952), .B2(n20715), .ZN(
        n20719) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20717), .B1(
        n20744), .B2(n20890), .ZN(n20718) );
  OAI211_X1 U23652 ( .C1(n20895), .C2(n20720), .A(n20719), .B(n20718), .ZN(
        P1_U3112) );
  NOR3_X1 U23653 ( .A1(n20786), .A2(n20722), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20759) );
  NAND2_X1 U23654 ( .A1(n20820), .A2(n20759), .ZN(n20724) );
  INV_X1 U23655 ( .A(n20724), .ZN(n20747) );
  AOI22_X1 U23656 ( .A1(n20744), .A2(n20911), .B1(n20901), .B2(n20747), .ZN(
        n20733) );
  NAND2_X1 U23657 ( .A1(n20783), .A2(n20752), .ZN(n20723) );
  AOI21_X1 U23658 ( .B1(n20723), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20903), 
        .ZN(n20728) );
  NAND2_X1 U23659 ( .A1(n20754), .A2(n20854), .ZN(n20730) );
  AOI22_X1 U23660 ( .A1(n20728), .A2(n20730), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20724), .ZN(n20726) );
  OR2_X1 U23661 ( .A1(n20725), .A2(n20786), .ZN(n20847) );
  NAND2_X1 U23662 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20847), .ZN(n20856) );
  NAND3_X1 U23663 ( .A1(n20727), .A2(n20726), .A3(n20856), .ZN(n20749) );
  INV_X1 U23664 ( .A(n20728), .ZN(n20731) );
  AOI22_X1 U23665 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20749), .B1(
        n20900), .B2(n20748), .ZN(n20732) );
  OAI211_X1 U23666 ( .C1(n20914), .C2(n20783), .A(n20733), .B(n20732), .ZN(
        P1_U3113) );
  AOI22_X1 U23667 ( .A1(n20744), .A2(n20917), .B1(n20916), .B2(n20747), .ZN(
        n20735) );
  AOI22_X1 U23668 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20749), .B1(
        n20915), .B2(n20748), .ZN(n20734) );
  OAI211_X1 U23669 ( .C1(n20920), .C2(n20783), .A(n20735), .B(n20734), .ZN(
        P1_U3114) );
  INV_X1 U23670 ( .A(n20783), .ZN(n20771) );
  AOI22_X1 U23671 ( .A1(n20771), .A2(n20868), .B1(n20922), .B2(n20747), .ZN(
        n20737) );
  AOI22_X1 U23672 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20749), .B1(
        n20921), .B2(n20748), .ZN(n20736) );
  OAI211_X1 U23673 ( .C1(n20871), .C2(n20752), .A(n20737), .B(n20736), .ZN(
        P1_U3115) );
  AOI22_X1 U23674 ( .A1(n20744), .A2(n20929), .B1(n20928), .B2(n20747), .ZN(
        n20739) );
  AOI22_X1 U23675 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20749), .B1(
        n20927), .B2(n20748), .ZN(n20738) );
  OAI211_X1 U23676 ( .C1(n20932), .C2(n20783), .A(n20739), .B(n20738), .ZN(
        P1_U3116) );
  AOI22_X1 U23677 ( .A1(n20744), .A2(n20935), .B1(n20934), .B2(n20747), .ZN(
        n20741) );
  AOI22_X1 U23678 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20749), .B1(
        n20933), .B2(n20748), .ZN(n20740) );
  OAI211_X1 U23679 ( .C1(n20938), .C2(n20783), .A(n20741), .B(n20740), .ZN(
        P1_U3117) );
  AOI22_X1 U23680 ( .A1(n20744), .A2(n20941), .B1(n20939), .B2(n20747), .ZN(
        n20743) );
  AOI22_X1 U23681 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20749), .B1(
        n20940), .B2(n20748), .ZN(n20742) );
  OAI211_X1 U23682 ( .C1(n20944), .C2(n20783), .A(n20743), .B(n20742), .ZN(
        P1_U3118) );
  AOI22_X1 U23683 ( .A1(n20744), .A2(n20947), .B1(n20945), .B2(n20747), .ZN(
        n20746) );
  AOI22_X1 U23684 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20749), .B1(
        n20946), .B2(n20748), .ZN(n20745) );
  OAI211_X1 U23685 ( .C1(n20950), .C2(n20783), .A(n20746), .B(n20745), .ZN(
        P1_U3119) );
  AOI22_X1 U23686 ( .A1(n20771), .A2(n20890), .B1(n20952), .B2(n20747), .ZN(
        n20751) );
  AOI22_X1 U23687 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20749), .B1(
        n20954), .B2(n20748), .ZN(n20750) );
  OAI211_X1 U23688 ( .C1(n20895), .C2(n20752), .A(n20751), .B(n20750), .ZN(
        P1_U3120) );
  AOI21_X1 U23689 ( .B1(n20754), .B2(n20897), .A(n10170), .ZN(n20756) );
  INV_X1 U23690 ( .A(n20759), .ZN(n20755) );
  OAI22_X1 U23691 ( .A1(n20756), .A2(n20903), .B1(n20755), .B2(n20966), .ZN(
        n20778) );
  AOI22_X1 U23692 ( .A1(n20901), .A2(n10170), .B1(n20900), .B2(n20778), .ZN(
        n20764) );
  OAI21_X1 U23693 ( .B1(n20762), .B2(n20903), .A(n20902), .ZN(n20757) );
  NAND2_X1 U23694 ( .A1(n20757), .A2(n20756), .ZN(n20758) );
  OAI211_X1 U23695 ( .C1(n20909), .C2(n20759), .A(n20908), .B(n20758), .ZN(
        n20780) );
  INV_X1 U23696 ( .A(n20760), .ZN(n20761) );
  AOI22_X1 U23697 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20780), .B1(
        n20779), .B2(n20860), .ZN(n20763) );
  OAI211_X1 U23698 ( .C1(n20863), .C2(n20783), .A(n20764), .B(n20763), .ZN(
        P1_U3121) );
  AOI22_X1 U23699 ( .A1(n20916), .A2(n10170), .B1(n20915), .B2(n20778), .ZN(
        n20766) );
  AOI22_X1 U23700 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20780), .B1(
        n20779), .B2(n20864), .ZN(n20765) );
  OAI211_X1 U23701 ( .C1(n20867), .C2(n20783), .A(n20766), .B(n20765), .ZN(
        P1_U3122) );
  AOI22_X1 U23702 ( .A1(n20922), .A2(n10170), .B1(n20921), .B2(n20778), .ZN(
        n20768) );
  AOI22_X1 U23703 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20780), .B1(
        n20771), .B2(n20923), .ZN(n20767) );
  OAI211_X1 U23704 ( .C1(n20926), .C2(n20818), .A(n20768), .B(n20767), .ZN(
        P1_U3123) );
  AOI22_X1 U23705 ( .A1(n20928), .A2(n10170), .B1(n20927), .B2(n20778), .ZN(
        n20770) );
  AOI22_X1 U23706 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20780), .B1(
        n20779), .B2(n20872), .ZN(n20769) );
  OAI211_X1 U23707 ( .C1(n20875), .C2(n20783), .A(n20770), .B(n20769), .ZN(
        P1_U3124) );
  AOI22_X1 U23708 ( .A1(n20934), .A2(n10170), .B1(n20933), .B2(n20778), .ZN(
        n20773) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20780), .B1(
        n20771), .B2(n20935), .ZN(n20772) );
  OAI211_X1 U23710 ( .C1(n20938), .C2(n20818), .A(n20773), .B(n20772), .ZN(
        P1_U3125) );
  AOI22_X1 U23711 ( .A1(n20940), .A2(n20778), .B1(n20939), .B2(n10170), .ZN(
        n20775) );
  AOI22_X1 U23712 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20780), .B1(
        n20779), .B2(n20880), .ZN(n20774) );
  OAI211_X1 U23713 ( .C1(n20883), .C2(n20783), .A(n20775), .B(n20774), .ZN(
        P1_U3126) );
  AOI22_X1 U23714 ( .A1(n20946), .A2(n20778), .B1(n20945), .B2(n10170), .ZN(
        n20777) );
  AOI22_X1 U23715 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20780), .B1(
        n20779), .B2(n20884), .ZN(n20776) );
  OAI211_X1 U23716 ( .C1(n20887), .C2(n20783), .A(n20777), .B(n20776), .ZN(
        P1_U3127) );
  AOI22_X1 U23717 ( .A1(n20954), .A2(n20778), .B1(n20952), .B2(n10170), .ZN(
        n20782) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20780), .B1(
        n20779), .B2(n20890), .ZN(n20781) );
  OAI211_X1 U23719 ( .C1(n20895), .C2(n20783), .A(n20782), .B(n20781), .ZN(
        P1_U3128) );
  NOR3_X1 U23720 ( .A1(n20787), .A2(n20786), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20825) );
  NAND2_X1 U23721 ( .A1(n20820), .A2(n20825), .ZN(n20792) );
  INV_X1 U23722 ( .A(n20792), .ZN(n20813) );
  AOI22_X1 U23723 ( .A1(n20842), .A2(n20860), .B1(n20901), .B2(n20813), .ZN(
        n20800) );
  INV_X1 U23724 ( .A(n20796), .ZN(n20794) );
  INV_X1 U23725 ( .A(n20842), .ZN(n20788) );
  NAND3_X1 U23726 ( .A1(n20788), .A2(n20909), .A3(n20818), .ZN(n20790) );
  NAND2_X1 U23727 ( .A1(n20790), .A2(n20789), .ZN(n20795) );
  OR2_X1 U23728 ( .A1(n13223), .A2(n20791), .ZN(n20849) );
  OR2_X1 U23729 ( .A1(n20849), .A2(n20854), .ZN(n20797) );
  AOI22_X1 U23730 ( .A1(n20795), .A2(n20797), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20792), .ZN(n20793) );
  OAI211_X1 U23731 ( .C1(n20794), .C2(n20966), .A(n20857), .B(n20793), .ZN(
        n20815) );
  INV_X1 U23732 ( .A(n20795), .ZN(n20798) );
  AOI22_X1 U23733 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20815), .B1(
        n20900), .B2(n20814), .ZN(n20799) );
  OAI211_X1 U23734 ( .C1(n20863), .C2(n20818), .A(n20800), .B(n20799), .ZN(
        P1_U3129) );
  AOI22_X1 U23735 ( .A1(n20842), .A2(n20864), .B1(n20916), .B2(n20813), .ZN(
        n20802) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20815), .B1(
        n20915), .B2(n20814), .ZN(n20801) );
  OAI211_X1 U23737 ( .C1(n20867), .C2(n20818), .A(n20802), .B(n20801), .ZN(
        P1_U3130) );
  AOI22_X1 U23738 ( .A1(n20842), .A2(n20868), .B1(n20922), .B2(n20813), .ZN(
        n20804) );
  AOI22_X1 U23739 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20815), .B1(
        n20921), .B2(n20814), .ZN(n20803) );
  OAI211_X1 U23740 ( .C1(n20871), .C2(n20818), .A(n20804), .B(n20803), .ZN(
        P1_U3131) );
  AOI22_X1 U23741 ( .A1(n20842), .A2(n20872), .B1(n20928), .B2(n20813), .ZN(
        n20806) );
  AOI22_X1 U23742 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20815), .B1(
        n20927), .B2(n20814), .ZN(n20805) );
  OAI211_X1 U23743 ( .C1(n20875), .C2(n20818), .A(n20806), .B(n20805), .ZN(
        P1_U3132) );
  AOI22_X1 U23744 ( .A1(n20842), .A2(n20876), .B1(n20934), .B2(n20813), .ZN(
        n20808) );
  AOI22_X1 U23745 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20815), .B1(
        n20933), .B2(n20814), .ZN(n20807) );
  OAI211_X1 U23746 ( .C1(n20879), .C2(n20818), .A(n20808), .B(n20807), .ZN(
        P1_U3133) );
  AOI22_X1 U23747 ( .A1(n20842), .A2(n20880), .B1(n20939), .B2(n20813), .ZN(
        n20810) );
  AOI22_X1 U23748 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20815), .B1(
        n20940), .B2(n20814), .ZN(n20809) );
  OAI211_X1 U23749 ( .C1(n20883), .C2(n20818), .A(n20810), .B(n20809), .ZN(
        P1_U3134) );
  AOI22_X1 U23750 ( .A1(n20842), .A2(n20884), .B1(n20945), .B2(n20813), .ZN(
        n20812) );
  AOI22_X1 U23751 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20815), .B1(
        n20946), .B2(n20814), .ZN(n20811) );
  OAI211_X1 U23752 ( .C1(n20887), .C2(n20818), .A(n20812), .B(n20811), .ZN(
        P1_U3135) );
  AOI22_X1 U23753 ( .A1(n20842), .A2(n20890), .B1(n20952), .B2(n20813), .ZN(
        n20817) );
  AOI22_X1 U23754 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20815), .B1(
        n20954), .B2(n20814), .ZN(n20816) );
  OAI211_X1 U23755 ( .C1(n20895), .C2(n20818), .A(n20817), .B(n20816), .ZN(
        P1_U3136) );
  INV_X1 U23756 ( .A(n20851), .ZN(n20904) );
  INV_X1 U23757 ( .A(n20825), .ZN(n20822) );
  NOR2_X1 U23758 ( .A1(n20820), .A2(n20822), .ZN(n20840) );
  INV_X1 U23759 ( .A(n20849), .ZN(n20898) );
  AOI21_X1 U23760 ( .B1(n20898), .B2(n20821), .A(n20840), .ZN(n20823) );
  OAI22_X1 U23761 ( .A1(n20823), .A2(n20903), .B1(n20822), .B2(n20966), .ZN(
        n20841) );
  AOI22_X1 U23762 ( .A1(n20901), .A2(n20840), .B1(n20900), .B2(n20841), .ZN(
        n20827) );
  OAI211_X1 U23763 ( .C1(n20851), .C2(n20852), .A(n20909), .B(n20823), .ZN(
        n20824) );
  OAI211_X1 U23764 ( .C1(n20909), .C2(n20825), .A(n20908), .B(n20824), .ZN(
        n20843) );
  AOI22_X1 U23765 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20911), .ZN(n20826) );
  OAI211_X1 U23766 ( .C1(n20914), .C2(n20894), .A(n20827), .B(n20826), .ZN(
        P1_U3137) );
  AOI22_X1 U23767 ( .A1(n20916), .A2(n20840), .B1(n20915), .B2(n20841), .ZN(
        n20829) );
  AOI22_X1 U23768 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20917), .ZN(n20828) );
  OAI211_X1 U23769 ( .C1(n20920), .C2(n20894), .A(n20829), .B(n20828), .ZN(
        P1_U3138) );
  AOI22_X1 U23770 ( .A1(n20922), .A2(n20840), .B1(n20921), .B2(n20841), .ZN(
        n20831) );
  AOI22_X1 U23771 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20923), .ZN(n20830) );
  OAI211_X1 U23772 ( .C1(n20926), .C2(n20894), .A(n20831), .B(n20830), .ZN(
        P1_U3139) );
  AOI22_X1 U23773 ( .A1(n20928), .A2(n20840), .B1(n20927), .B2(n20841), .ZN(
        n20833) );
  AOI22_X1 U23774 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20929), .ZN(n20832) );
  OAI211_X1 U23775 ( .C1(n20932), .C2(n20894), .A(n20833), .B(n20832), .ZN(
        P1_U3140) );
  AOI22_X1 U23776 ( .A1(n20934), .A2(n20840), .B1(n20933), .B2(n20841), .ZN(
        n20835) );
  AOI22_X1 U23777 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20935), .ZN(n20834) );
  OAI211_X1 U23778 ( .C1(n20938), .C2(n20894), .A(n20835), .B(n20834), .ZN(
        P1_U3141) );
  AOI22_X1 U23779 ( .A1(n20940), .A2(n20841), .B1(n20939), .B2(n20840), .ZN(
        n20837) );
  AOI22_X1 U23780 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20941), .ZN(n20836) );
  OAI211_X1 U23781 ( .C1(n20944), .C2(n20894), .A(n20837), .B(n20836), .ZN(
        P1_U3142) );
  AOI22_X1 U23782 ( .A1(n20946), .A2(n20841), .B1(n20945), .B2(n20840), .ZN(
        n20839) );
  AOI22_X1 U23783 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20947), .ZN(n20838) );
  OAI211_X1 U23784 ( .C1(n20950), .C2(n20894), .A(n20839), .B(n20838), .ZN(
        P1_U3143) );
  AOI22_X1 U23785 ( .A1(n20954), .A2(n20841), .B1(n20952), .B2(n20840), .ZN(
        n20845) );
  AOI22_X1 U23786 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20843), .B1(
        n20842), .B2(n20955), .ZN(n20844) );
  OAI211_X1 U23787 ( .C1(n20961), .C2(n20894), .A(n20845), .B(n20844), .ZN(
        P1_U3144) );
  INV_X1 U23788 ( .A(n20910), .ZN(n20899) );
  NOR2_X1 U23789 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20899), .ZN(
        n20888) );
  NAND2_X1 U23790 ( .A1(n20854), .A2(n20909), .ZN(n20848) );
  OAI22_X1 U23791 ( .A1(n20849), .A2(n20848), .B1(n20847), .B2(n20846), .ZN(
        n20889) );
  AOI22_X1 U23792 ( .A1(n20901), .A2(n20888), .B1(n20900), .B2(n20889), .ZN(
        n20862) );
  AOI21_X1 U23793 ( .B1(n20894), .B2(n20859), .A(n20852), .ZN(n20853) );
  AOI21_X1 U23794 ( .B1(n20898), .B2(n20854), .A(n20853), .ZN(n20855) );
  NOR2_X1 U23795 ( .A1(n20855), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20858) );
  AOI22_X1 U23796 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20891), .B1(
        n20956), .B2(n20860), .ZN(n20861) );
  OAI211_X1 U23797 ( .C1(n20863), .C2(n20894), .A(n20862), .B(n20861), .ZN(
        P1_U3145) );
  AOI22_X1 U23798 ( .A1(n20916), .A2(n20888), .B1(n20915), .B2(n20889), .ZN(
        n20866) );
  AOI22_X1 U23799 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20891), .B1(
        n20956), .B2(n20864), .ZN(n20865) );
  OAI211_X1 U23800 ( .C1(n20867), .C2(n20894), .A(n20866), .B(n20865), .ZN(
        P1_U3146) );
  AOI22_X1 U23801 ( .A1(n20922), .A2(n20888), .B1(n20921), .B2(n20889), .ZN(
        n20870) );
  AOI22_X1 U23802 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20891), .B1(
        n20956), .B2(n20868), .ZN(n20869) );
  OAI211_X1 U23803 ( .C1(n20871), .C2(n20894), .A(n20870), .B(n20869), .ZN(
        P1_U3147) );
  AOI22_X1 U23804 ( .A1(n20928), .A2(n20888), .B1(n20927), .B2(n20889), .ZN(
        n20874) );
  AOI22_X1 U23805 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20891), .B1(
        n20956), .B2(n20872), .ZN(n20873) );
  OAI211_X1 U23806 ( .C1(n20875), .C2(n20894), .A(n20874), .B(n20873), .ZN(
        P1_U3148) );
  AOI22_X1 U23807 ( .A1(n20934), .A2(n20888), .B1(n20933), .B2(n20889), .ZN(
        n20878) );
  AOI22_X1 U23808 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20891), .B1(
        n20956), .B2(n20876), .ZN(n20877) );
  OAI211_X1 U23809 ( .C1(n20879), .C2(n20894), .A(n20878), .B(n20877), .ZN(
        P1_U3149) );
  AOI22_X1 U23810 ( .A1(n20940), .A2(n20889), .B1(n20939), .B2(n20888), .ZN(
        n20882) );
  AOI22_X1 U23811 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20891), .B1(
        n20956), .B2(n20880), .ZN(n20881) );
  OAI211_X1 U23812 ( .C1(n20883), .C2(n20894), .A(n20882), .B(n20881), .ZN(
        P1_U3150) );
  AOI22_X1 U23813 ( .A1(n20946), .A2(n20889), .B1(n20945), .B2(n20888), .ZN(
        n20886) );
  AOI22_X1 U23814 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20891), .B1(
        n20956), .B2(n20884), .ZN(n20885) );
  OAI211_X1 U23815 ( .C1(n20887), .C2(n20894), .A(n20886), .B(n20885), .ZN(
        P1_U3151) );
  AOI22_X1 U23816 ( .A1(n20954), .A2(n20889), .B1(n20952), .B2(n20888), .ZN(
        n20893) );
  AOI22_X1 U23817 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20891), .B1(
        n20956), .B2(n20890), .ZN(n20892) );
  OAI211_X1 U23818 ( .C1(n20895), .C2(n20894), .A(n20893), .B(n20892), .ZN(
        P1_U3152) );
  INV_X1 U23819 ( .A(n20896), .ZN(n20951) );
  AOI21_X1 U23820 ( .B1(n20898), .B2(n20897), .A(n20951), .ZN(n20905) );
  OAI22_X1 U23821 ( .A1(n20905), .A2(n20903), .B1(n20966), .B2(n20899), .ZN(
        n20953) );
  AOI22_X1 U23822 ( .A1(n20901), .A2(n20951), .B1(n20900), .B2(n20953), .ZN(
        n20913) );
  OAI21_X1 U23823 ( .B1(n20904), .B2(n20903), .A(n20902), .ZN(n20906) );
  NAND2_X1 U23824 ( .A1(n20906), .A2(n20905), .ZN(n20907) );
  OAI211_X1 U23825 ( .C1(n20910), .C2(n20909), .A(n20908), .B(n20907), .ZN(
        n20957) );
  AOI22_X1 U23826 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20957), .B1(
        n20956), .B2(n20911), .ZN(n20912) );
  OAI211_X1 U23827 ( .C1(n20914), .C2(n20960), .A(n20913), .B(n20912), .ZN(
        P1_U3153) );
  AOI22_X1 U23828 ( .A1(n20916), .A2(n20951), .B1(n20915), .B2(n20953), .ZN(
        n20919) );
  AOI22_X1 U23829 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20957), .B1(
        n20956), .B2(n20917), .ZN(n20918) );
  OAI211_X1 U23830 ( .C1(n20920), .C2(n20960), .A(n20919), .B(n20918), .ZN(
        P1_U3154) );
  AOI22_X1 U23831 ( .A1(n20922), .A2(n20951), .B1(n20921), .B2(n20953), .ZN(
        n20925) );
  AOI22_X1 U23832 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20957), .B1(
        n20956), .B2(n20923), .ZN(n20924) );
  OAI211_X1 U23833 ( .C1(n20926), .C2(n20960), .A(n20925), .B(n20924), .ZN(
        P1_U3155) );
  AOI22_X1 U23834 ( .A1(n20928), .A2(n20951), .B1(n20927), .B2(n20953), .ZN(
        n20931) );
  AOI22_X1 U23835 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20957), .B1(
        n20956), .B2(n20929), .ZN(n20930) );
  OAI211_X1 U23836 ( .C1(n20932), .C2(n20960), .A(n20931), .B(n20930), .ZN(
        P1_U3156) );
  AOI22_X1 U23837 ( .A1(n20934), .A2(n20951), .B1(n20933), .B2(n20953), .ZN(
        n20937) );
  AOI22_X1 U23838 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20957), .B1(
        n20956), .B2(n20935), .ZN(n20936) );
  OAI211_X1 U23839 ( .C1(n20938), .C2(n20960), .A(n20937), .B(n20936), .ZN(
        P1_U3157) );
  AOI22_X1 U23840 ( .A1(n20940), .A2(n20953), .B1(n20939), .B2(n20951), .ZN(
        n20943) );
  AOI22_X1 U23841 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20957), .B1(
        n20956), .B2(n20941), .ZN(n20942) );
  OAI211_X1 U23842 ( .C1(n20944), .C2(n20960), .A(n20943), .B(n20942), .ZN(
        P1_U3158) );
  AOI22_X1 U23843 ( .A1(n20946), .A2(n20953), .B1(n20945), .B2(n20951), .ZN(
        n20949) );
  AOI22_X1 U23844 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20957), .B1(
        n20956), .B2(n20947), .ZN(n20948) );
  OAI211_X1 U23845 ( .C1(n20950), .C2(n20960), .A(n20949), .B(n20948), .ZN(
        P1_U3159) );
  AOI22_X1 U23846 ( .A1(n20954), .A2(n20953), .B1(n20952), .B2(n20951), .ZN(
        n20959) );
  AOI22_X1 U23847 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20957), .B1(
        n20956), .B2(n20955), .ZN(n20958) );
  OAI211_X1 U23848 ( .C1(n20961), .C2(n20960), .A(n20959), .B(n20958), .ZN(
        P1_U3160) );
  NOR2_X1 U23849 ( .A1(n20963), .A2(n20962), .ZN(n20967) );
  INV_X1 U23850 ( .A(n20964), .ZN(n20965) );
  OAI21_X1 U23851 ( .B1(n20967), .B2(n20966), .A(n20965), .ZN(P1_U3163) );
  AND2_X1 U23852 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20968), .ZN(
        P1_U3164) );
  AND2_X1 U23853 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20968), .ZN(
        P1_U3165) );
  AND2_X1 U23854 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20968), .ZN(
        P1_U3166) );
  AND2_X1 U23855 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20968), .ZN(
        P1_U3167) );
  AND2_X1 U23856 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20968), .ZN(
        P1_U3168) );
  AND2_X1 U23857 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20968), .ZN(
        P1_U3169) );
  AND2_X1 U23858 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20968), .ZN(
        P1_U3170) );
  AND2_X1 U23859 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20968), .ZN(
        P1_U3171) );
  AND2_X1 U23860 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20968), .ZN(
        P1_U3172) );
  AND2_X1 U23861 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20968), .ZN(
        P1_U3173) );
  AND2_X1 U23862 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20968), .ZN(
        P1_U3174) );
  AND2_X1 U23863 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20968), .ZN(
        P1_U3175) );
  AND2_X1 U23864 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20968), .ZN(
        P1_U3176) );
  AND2_X1 U23865 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20968), .ZN(
        P1_U3177) );
  AND2_X1 U23866 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20968), .ZN(
        P1_U3178) );
  AND2_X1 U23867 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20968), .ZN(
        P1_U3179) );
  AND2_X1 U23868 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20968), .ZN(
        P1_U3180) );
  AND2_X1 U23869 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20968), .ZN(
        P1_U3181) );
  AND2_X1 U23870 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20968), .ZN(
        P1_U3182) );
  AND2_X1 U23871 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20968), .ZN(
        P1_U3183) );
  AND2_X1 U23872 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20968), .ZN(
        P1_U3184) );
  AND2_X1 U23873 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20968), .ZN(
        P1_U3185) );
  AND2_X1 U23874 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20968), .ZN(P1_U3186) );
  AND2_X1 U23875 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20968), .ZN(P1_U3187) );
  AND2_X1 U23876 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20968), .ZN(P1_U3188) );
  AND2_X1 U23877 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20968), .ZN(P1_U3189) );
  AND2_X1 U23878 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20968), .ZN(P1_U3190) );
  AND2_X1 U23879 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20968), .ZN(P1_U3191) );
  AND2_X1 U23880 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20968), .ZN(P1_U3192) );
  AND2_X1 U23881 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20968), .ZN(P1_U3193) );
  AOI21_X1 U23882 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20976), .A(n20969), 
        .ZN(n20981) );
  OAI21_X1 U23883 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20975), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20970) );
  AOI211_X1 U23884 ( .C1(HOLD), .C2(P1_STATE_REG_2__SCAN_IN), .A(n20971), .B(
        n20970), .ZN(n20972) );
  OAI22_X1 U23885 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20981), .B1(n21046), 
        .B2(n20972), .ZN(P1_U3194) );
  NOR2_X1 U23886 ( .A1(NA), .A2(n20973), .ZN(n20974) );
  OAI22_X1 U23887 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20974), .B1(
        P1_STATE_REG_1__SCAN_IN), .B2(n20975), .ZN(n20980) );
  NAND2_X1 U23888 ( .A1(n20976), .A2(n20975), .ZN(n20977) );
  OAI221_X1 U23889 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(
        P1_STATE_REG_1__SCAN_IN), .C1(P1_REQUESTPENDING_REG_SCAN_IN), .C2(
        n20977), .A(n20982), .ZN(n20978) );
  NAND3_X1 U23890 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(HOLD), .A3(n20978), .ZN(
        n20979) );
  OAI21_X1 U23891 ( .B1(n20981), .B2(n20980), .A(n20979), .ZN(P1_U3196) );
  OR2_X1 U23892 ( .A1(n21059), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21011) );
  AOI222_X1 U23893 ( .A1(n21026), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n9652), .ZN(n20983) );
  INV_X1 U23894 ( .A(n20983), .ZN(P1_U3197) );
  AOI222_X1 U23895 ( .A1(n9652), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n21026), .ZN(n20984) );
  INV_X1 U23896 ( .A(n20984), .ZN(P1_U3198) );
  INV_X1 U23897 ( .A(n9652), .ZN(n21024) );
  AOI22_X1 U23898 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(n21059), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(n21026), .ZN(n20985) );
  OAI21_X1 U23899 ( .B1(n20986), .B2(n21024), .A(n20985), .ZN(P1_U3199) );
  OAI222_X1 U23900 ( .A1(n21011), .A2(n20989), .B1(n20988), .B2(n21046), .C1(
        n20987), .C2(n21024), .ZN(P1_U3200) );
  AOI222_X1 U23901 ( .A1(n9652), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n21026), .ZN(n20990) );
  INV_X1 U23902 ( .A(n20990), .ZN(P1_U3201) );
  INV_X1 U23903 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21177) );
  OAI222_X1 U23904 ( .A1(n21024), .A2(n20992), .B1(n21177), .B2(n21046), .C1(
        n20991), .C2(n21011), .ZN(P1_U3202) );
  AOI222_X1 U23905 ( .A1(n9652), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n21026), .ZN(n20993) );
  INV_X1 U23906 ( .A(n20993), .ZN(P1_U3203) );
  AOI222_X1 U23907 ( .A1(n21026), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n9652), .ZN(n20994) );
  INV_X1 U23908 ( .A(n20994), .ZN(P1_U3204) );
  AOI222_X1 U23909 ( .A1(n9652), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21026), .ZN(n20995) );
  INV_X1 U23910 ( .A(n20995), .ZN(P1_U3205) );
  AOI222_X1 U23911 ( .A1(n21026), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n9652), .ZN(n20996) );
  INV_X1 U23912 ( .A(n20996), .ZN(P1_U3206) );
  AOI22_X1 U23913 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21059), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21026), .ZN(n20997) );
  OAI21_X1 U23914 ( .B1(n20998), .B2(n21024), .A(n20997), .ZN(P1_U3207) );
  AOI22_X1 U23915 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n21059), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n9652), .ZN(n20999) );
  OAI21_X1 U23916 ( .B1(n21001), .B2(n21011), .A(n20999), .ZN(P1_U3208) );
  AOI22_X1 U23917 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n21059), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n21026), .ZN(n21000) );
  OAI21_X1 U23918 ( .B1(n21001), .B2(n21024), .A(n21000), .ZN(P1_U3209) );
  AOI22_X1 U23919 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n21059), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n9652), .ZN(n21002) );
  OAI21_X1 U23920 ( .B1(n21003), .B2(n21011), .A(n21002), .ZN(P1_U3210) );
  AOI222_X1 U23921 ( .A1(n9652), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n21026), .ZN(n21004) );
  INV_X1 U23922 ( .A(n21004), .ZN(P1_U3211) );
  INV_X1 U23923 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21006) );
  AOI22_X1 U23924 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21059), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21026), .ZN(n21005) );
  OAI21_X1 U23925 ( .B1(n21006), .B2(n21024), .A(n21005), .ZN(P1_U3212) );
  AOI22_X1 U23926 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21059), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n9652), .ZN(n21007) );
  OAI21_X1 U23927 ( .B1(n21009), .B2(n21011), .A(n21007), .ZN(P1_U3213) );
  AOI22_X1 U23928 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21059), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21026), .ZN(n21008) );
  OAI21_X1 U23929 ( .B1(n21009), .B2(n21024), .A(n21008), .ZN(P1_U3214) );
  AOI22_X1 U23930 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21059), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n9652), .ZN(n21010) );
  OAI21_X1 U23931 ( .B1(n21012), .B2(n21011), .A(n21010), .ZN(P1_U3215) );
  AOI222_X1 U23932 ( .A1(n9652), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n21026), .ZN(n21013) );
  INV_X1 U23933 ( .A(n21013), .ZN(P1_U3216) );
  AOI222_X1 U23934 ( .A1(n9652), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n21026), .ZN(n21014) );
  INV_X1 U23935 ( .A(n21014), .ZN(P1_U3217) );
  AOI222_X1 U23936 ( .A1(n9652), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n21026), .ZN(n21015) );
  INV_X1 U23937 ( .A(n21015), .ZN(P1_U3218) );
  AOI222_X1 U23938 ( .A1(n9652), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n21026), .ZN(n21016) );
  INV_X1 U23939 ( .A(n21016), .ZN(P1_U3219) );
  AOI222_X1 U23940 ( .A1(n9652), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n21026), .ZN(n21017) );
  INV_X1 U23941 ( .A(n21017), .ZN(P1_U3220) );
  AOI222_X1 U23942 ( .A1(n9652), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n21026), .ZN(n21018) );
  INV_X1 U23943 ( .A(n21018), .ZN(P1_U3221) );
  AOI222_X1 U23944 ( .A1(n9652), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n21026), .ZN(n21019) );
  INV_X1 U23945 ( .A(n21019), .ZN(P1_U3222) );
  AOI22_X1 U23946 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n21026), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21059), .ZN(n21020) );
  OAI21_X1 U23947 ( .B1(n21021), .B2(n21024), .A(n21020), .ZN(P1_U3223) );
  AOI222_X1 U23948 ( .A1(n9652), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21026), .ZN(n21022) );
  INV_X1 U23949 ( .A(n21022), .ZN(P1_U3224) );
  AOI22_X1 U23950 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n21026), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21059), .ZN(n21023) );
  OAI21_X1 U23951 ( .B1(n21025), .B2(n21024), .A(n21023), .ZN(P1_U3225) );
  AOI222_X1 U23952 ( .A1(n9652), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21059), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n21026), .ZN(n21028) );
  INV_X1 U23953 ( .A(n21028), .ZN(P1_U3226) );
  OAI22_X1 U23954 ( .A1(n21059), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21046), .ZN(n21029) );
  INV_X1 U23955 ( .A(n21029), .ZN(P1_U3458) );
  OAI22_X1 U23956 ( .A1(n21059), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21046), .ZN(n21030) );
  INV_X1 U23957 ( .A(n21030), .ZN(P1_U3459) );
  OAI22_X1 U23958 ( .A1(n21059), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21046), .ZN(n21031) );
  INV_X1 U23959 ( .A(n21031), .ZN(P1_U3460) );
  OAI22_X1 U23960 ( .A1(n21059), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21046), .ZN(n21032) );
  INV_X1 U23961 ( .A(n21032), .ZN(P1_U3461) );
  OAI21_X1 U23962 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21036), .A(n21034), 
        .ZN(n21033) );
  INV_X1 U23963 ( .A(n21033), .ZN(P1_U3464) );
  OAI21_X1 U23964 ( .B1(n21036), .B2(n21035), .A(n21034), .ZN(P1_U3465) );
  AOI21_X1 U23965 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21038) );
  AOI22_X1 U23966 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21038), .B2(n21037), .ZN(n21041) );
  INV_X1 U23967 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21040) );
  AOI22_X1 U23968 ( .A1(n21044), .A2(n21041), .B1(n21040), .B2(n21039), .ZN(
        P1_U3481) );
  INV_X1 U23969 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21043) );
  OAI21_X1 U23970 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21044), .ZN(n21042) );
  OAI21_X1 U23971 ( .B1(n21044), .B2(n21043), .A(n21042), .ZN(P1_U3482) );
  AOI22_X1 U23972 ( .A1(n21046), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21045), 
        .B2(n21059), .ZN(P1_U3483) );
  INV_X1 U23973 ( .A(n21047), .ZN(n21048) );
  AOI211_X1 U23974 ( .C1(n21051), .C2(n21050), .A(n21049), .B(n21048), .ZN(
        n21058) );
  NAND3_X1 U23975 ( .A1(n21053), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n21052), 
        .ZN(n21055) );
  AOI21_X1 U23976 ( .B1(n21055), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n21054), 
        .ZN(n21057) );
  NAND2_X1 U23977 ( .A1(n21058), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21056) );
  OAI21_X1 U23978 ( .B1(n21058), .B2(n21057), .A(n21056), .ZN(P1_U3485) );
  MUX2_X1 U23979 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n21059), .Z(P1_U3486) );
  AOI22_X1 U23980 ( .A1(n21177), .A2(keyinput81), .B1(n21203), .B2(keyinput65), 
        .ZN(n21060) );
  OAI221_X1 U23981 ( .B1(n21177), .B2(keyinput81), .C1(n21203), .C2(keyinput65), .A(n21060), .ZN(n21067) );
  AOI22_X1 U23982 ( .A1(n14042), .A2(keyinput95), .B1(keyinput73), .B2(n21218), 
        .ZN(n21061) );
  OAI221_X1 U23983 ( .B1(n14042), .B2(keyinput95), .C1(n21218), .C2(keyinput73), .A(n21061), .ZN(n21066) );
  INV_X1 U23984 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n21189) );
  AOI22_X1 U23985 ( .A1(n21189), .A2(keyinput121), .B1(n21197), .B2(keyinput97), .ZN(n21062) );
  OAI221_X1 U23986 ( .B1(n21189), .B2(keyinput121), .C1(n21197), .C2(
        keyinput97), .A(n21062), .ZN(n21065) );
  AOI22_X1 U23987 ( .A1(n21237), .A2(keyinput84), .B1(n21236), .B2(keyinput96), 
        .ZN(n21063) );
  OAI221_X1 U23988 ( .B1(n21237), .B2(keyinput84), .C1(n21236), .C2(keyinput96), .A(n21063), .ZN(n21064) );
  NOR4_X1 U23989 ( .A1(n21067), .A2(n21066), .A3(n21065), .A4(n21064), .ZN(
        n21107) );
  AOI22_X1 U23990 ( .A1(n21070), .A2(keyinput103), .B1(keyinput94), .B2(n21069), .ZN(n21068) );
  OAI221_X1 U23991 ( .B1(n21070), .B2(keyinput103), .C1(n21069), .C2(
        keyinput94), .A(n21068), .ZN(n21079) );
  INV_X1 U23992 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n21072) );
  INV_X1 U23993 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21240) );
  AOI22_X1 U23994 ( .A1(n21072), .A2(keyinput79), .B1(keyinput93), .B2(n21240), 
        .ZN(n21071) );
  OAI221_X1 U23995 ( .B1(n21072), .B2(keyinput79), .C1(n21240), .C2(keyinput93), .A(n21071), .ZN(n21078) );
  AOI22_X1 U23996 ( .A1(n21239), .A2(keyinput112), .B1(keyinput78), .B2(n13523), .ZN(n21073) );
  OAI221_X1 U23997 ( .B1(n21239), .B2(keyinput112), .C1(n13523), .C2(
        keyinput78), .A(n21073), .ZN(n21077) );
  AOI22_X1 U23998 ( .A1(n21075), .A2(keyinput102), .B1(keyinput124), .B2(
        n12941), .ZN(n21074) );
  OAI221_X1 U23999 ( .B1(n21075), .B2(keyinput102), .C1(n12941), .C2(
        keyinput124), .A(n21074), .ZN(n21076) );
  NOR4_X1 U24000 ( .A1(n21079), .A2(n21078), .A3(n21077), .A4(n21076), .ZN(
        n21106) );
  INV_X1 U24001 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n21081) );
  AOI22_X1 U24002 ( .A1(n21081), .A2(keyinput114), .B1(keyinput77), .B2(n21176), .ZN(n21080) );
  OAI221_X1 U24003 ( .B1(n21081), .B2(keyinput114), .C1(n21176), .C2(
        keyinput77), .A(n21080), .ZN(n21090) );
  INV_X1 U24004 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n21222) );
  AOI22_X1 U24005 ( .A1(n21222), .A2(keyinput119), .B1(n21083), .B2(
        keyinput118), .ZN(n21082) );
  OAI221_X1 U24006 ( .B1(n21222), .B2(keyinput119), .C1(n21083), .C2(
        keyinput118), .A(n21082), .ZN(n21089) );
  AOI22_X1 U24007 ( .A1(n21085), .A2(keyinput70), .B1(n14390), .B2(keyinput89), 
        .ZN(n21084) );
  OAI221_X1 U24008 ( .B1(n21085), .B2(keyinput70), .C1(n14390), .C2(keyinput89), .A(n21084), .ZN(n21088) );
  AOI22_X1 U24009 ( .A1(n21194), .A2(keyinput91), .B1(n12624), .B2(keyinput90), 
        .ZN(n21086) );
  OAI221_X1 U24010 ( .B1(n21194), .B2(keyinput91), .C1(n12624), .C2(keyinput90), .A(n21086), .ZN(n21087) );
  NOR4_X1 U24011 ( .A1(n21090), .A2(n21089), .A3(n21088), .A4(n21087), .ZN(
        n21105) );
  AOI22_X1 U24012 ( .A1(n21092), .A2(keyinput105), .B1(n21211), .B2(keyinput88), .ZN(n21091) );
  OAI221_X1 U24013 ( .B1(n21092), .B2(keyinput105), .C1(n21211), .C2(
        keyinput88), .A(n21091), .ZN(n21103) );
  AOI22_X1 U24014 ( .A1(n21208), .A2(keyinput75), .B1(keyinput106), .B2(n21094), .ZN(n21093) );
  OAI221_X1 U24015 ( .B1(n21208), .B2(keyinput75), .C1(n21094), .C2(
        keyinput106), .A(n21093), .ZN(n21102) );
  INV_X1 U24016 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n21096) );
  AOI22_X1 U24017 ( .A1(n21212), .A2(keyinput123), .B1(keyinput85), .B2(n21096), .ZN(n21095) );
  OAI221_X1 U24018 ( .B1(n21212), .B2(keyinput123), .C1(n21096), .C2(
        keyinput85), .A(n21095), .ZN(n21101) );
  AOI22_X1 U24019 ( .A1(n21099), .A2(keyinput117), .B1(n21098), .B2(
        keyinput127), .ZN(n21097) );
  OAI221_X1 U24020 ( .B1(n21099), .B2(keyinput117), .C1(n21098), .C2(
        keyinput127), .A(n21097), .ZN(n21100) );
  NOR4_X1 U24021 ( .A1(n21103), .A2(n21102), .A3(n21101), .A4(n21100), .ZN(
        n21104) );
  AND4_X1 U24022 ( .A1(n21107), .A2(n21106), .A3(n21105), .A4(n21104), .ZN(
        n21254) );
  OAI22_X1 U24023 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(keyinput126), 
        .B1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(keyinput113), .ZN(n21108) );
  AOI221_X1 U24024 ( .B1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(keyinput126), 
        .C1(keyinput113), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(n21108), 
        .ZN(n21115) );
  OAI22_X1 U24025 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(keyinput120), 
        .B1(keyinput116), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n21109) );
  AOI221_X1 U24026 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput120), 
        .C1(P3_EBX_REG_13__SCAN_IN), .C2(keyinput116), .A(n21109), .ZN(n21114)
         );
  OAI22_X1 U24027 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(keyinput71), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(keyinput115), .ZN(n21110) );
  AOI221_X1 U24028 ( .B1(P2_EBX_REG_31__SCAN_IN), .B2(keyinput71), .C1(
        keyinput115), .C2(P2_STATE_REG_1__SCAN_IN), .A(n21110), .ZN(n21113) );
  OAI22_X1 U24029 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(keyinput99), 
        .B1(keyinput107), .B2(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n21111) );
  AOI221_X1 U24030 ( .B1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B2(keyinput99), 
        .C1(P1_ADDRESS_REG_0__SCAN_IN), .C2(keyinput107), .A(n21111), .ZN(
        n21112) );
  NAND4_X1 U24031 ( .A1(n21115), .A2(n21114), .A3(n21113), .A4(n21112), .ZN(
        n21147) );
  OAI22_X1 U24032 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(keyinput98), .B1(
        keyinput111), .B2(P1_EAX_REG_8__SCAN_IN), .ZN(n21116) );
  AOI221_X1 U24033 ( .B1(P2_EAX_REG_28__SCAN_IN), .B2(keyinput98), .C1(
        P1_EAX_REG_8__SCAN_IN), .C2(keyinput111), .A(n21116), .ZN(n21123) );
  OAI22_X1 U24034 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput80), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(keyinput72), .ZN(n21117) );
  AOI221_X1 U24035 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput80), .C1(
        keyinput72), .C2(P3_M_IO_N_REG_SCAN_IN), .A(n21117), .ZN(n21122) );
  OAI22_X1 U24036 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(keyinput104), 
        .B1(keyinput67), .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n21118) );
  AOI221_X1 U24037 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput104), 
        .C1(P2_DATAO_REG_10__SCAN_IN), .C2(keyinput67), .A(n21118), .ZN(n21121) );
  OAI22_X1 U24038 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(keyinput87), 
        .B1(keyinput101), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n21119) );
  AOI221_X1 U24039 ( .B1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B2(keyinput87), 
        .C1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .C2(keyinput101), .A(n21119), 
        .ZN(n21120) );
  NAND4_X1 U24040 ( .A1(n21123), .A2(n21122), .A3(n21121), .A4(n21120), .ZN(
        n21146) );
  XOR2_X1 U24041 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B(keyinput64), .Z(
        n21128) );
  XNOR2_X1 U24042 ( .A(n21219), .B(keyinput108), .ZN(n21127) );
  INV_X1 U24043 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n21124) );
  XNOR2_X1 U24044 ( .A(n21124), .B(keyinput92), .ZN(n21126) );
  XOR2_X1 U24045 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B(keyinput83), .Z(
        n21125) );
  NOR4_X1 U24046 ( .A1(n21128), .A2(n21127), .A3(n21126), .A4(n21125), .ZN(
        n21134) );
  INV_X1 U24047 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n21130) );
  OAI22_X1 U24048 ( .A1(n21130), .A2(keyinput109), .B1(n21233), .B2(
        keyinput122), .ZN(n21129) );
  AOI221_X1 U24049 ( .B1(n21130), .B2(keyinput109), .C1(keyinput122), .C2(
        n21233), .A(n21129), .ZN(n21133) );
  OAI22_X1 U24050 ( .A1(n21234), .A2(keyinput110), .B1(n21188), .B2(keyinput82), .ZN(n21131) );
  AOI221_X1 U24051 ( .B1(n21234), .B2(keyinput110), .C1(keyinput82), .C2(
        n21188), .A(n21131), .ZN(n21132) );
  NAND3_X1 U24052 ( .A1(n21134), .A2(n21133), .A3(n21132), .ZN(n21145) );
  OAI22_X1 U24053 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(keyinput76), .B1(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput74), .ZN(n21135) );
  AOI221_X1 U24054 ( .B1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B2(keyinput76), 
        .C1(keyinput74), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(n21135), 
        .ZN(n21143) );
  OAI22_X1 U24055 ( .A1(READY12_REG_SCAN_IN), .A2(keyinput68), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput100), .ZN(n21136) );
  AOI221_X1 U24056 ( .B1(READY12_REG_SCAN_IN), .B2(keyinput68), .C1(
        keyinput100), .C2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(n21136), .ZN(
        n21142) );
  OAI22_X1 U24057 ( .A1(n21205), .A2(keyinput66), .B1(keyinput86), .B2(
        P3_EAX_REG_9__SCAN_IN), .ZN(n21137) );
  AOI221_X1 U24058 ( .B1(n21205), .B2(keyinput66), .C1(P3_EAX_REG_9__SCAN_IN), 
        .C2(keyinput86), .A(n21137), .ZN(n21141) );
  INV_X1 U24059 ( .A(DATAI_1_), .ZN(n21139) );
  OAI22_X1 U24060 ( .A1(n21139), .A2(keyinput125), .B1(keyinput69), .B2(READY2), .ZN(n21138) );
  AOI221_X1 U24061 ( .B1(n21139), .B2(keyinput125), .C1(READY2), .C2(
        keyinput69), .A(n21138), .ZN(n21140) );
  NAND4_X1 U24062 ( .A1(n21143), .A2(n21142), .A3(n21141), .A4(n21140), .ZN(
        n21144) );
  NOR4_X1 U24063 ( .A1(n21147), .A2(n21146), .A3(n21145), .A4(n21144), .ZN(
        n21253) );
  AOI22_X1 U24064 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput16), .B1(
        P1_EAX_REG_8__SCAN_IN), .B2(keyinput47), .ZN(n21148) );
  OAI221_X1 U24065 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput16), .C1(
        P1_EAX_REG_8__SCAN_IN), .C2(keyinput47), .A(n21148), .ZN(n21155) );
  AOI22_X1 U24066 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(keyinput30), .B1(READY2), 
        .B2(keyinput5), .ZN(n21149) );
  OAI221_X1 U24067 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(keyinput30), .C1(READY2), .C2(keyinput5), .A(n21149), .ZN(n21154) );
  AOI22_X1 U24068 ( .A1(DATAI_1_), .A2(keyinput61), .B1(
        P1_INSTQUEUE_REG_8__7__SCAN_IN), .B2(keyinput39), .ZN(n21150) );
  OAI221_X1 U24069 ( .B1(DATAI_1_), .B2(keyinput61), .C1(
        P1_INSTQUEUE_REG_8__7__SCAN_IN), .C2(keyinput39), .A(n21150), .ZN(
        n21153) );
  AOI22_X1 U24070 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(keyinput43), .B1(
        P2_INSTQUEUE_REG_10__1__SCAN_IN), .B2(keyinput23), .ZN(n21151) );
  OAI221_X1 U24071 ( .B1(P1_ADDRESS_REG_0__SCAN_IN), .B2(keyinput43), .C1(
        P2_INSTQUEUE_REG_10__1__SCAN_IN), .C2(keyinput23), .A(n21151), .ZN(
        n21152) );
  NOR4_X1 U24072 ( .A1(n21155), .A2(n21154), .A3(n21153), .A4(n21152), .ZN(
        n21185) );
  AOI22_X1 U24073 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput53), .B1(
        BUF1_REG_2__SCAN_IN), .B2(keyinput63), .ZN(n21156) );
  OAI221_X1 U24074 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput53), .C1(
        BUF1_REG_2__SCAN_IN), .C2(keyinput63), .A(n21156), .ZN(n21163) );
  AOI22_X1 U24075 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(keyinput45), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(keyinput54), .ZN(n21157) );
  OAI221_X1 U24076 ( .B1(P1_ADDRESS_REG_27__SCAN_IN), .B2(keyinput45), .C1(
        P2_EBX_REG_11__SCAN_IN), .C2(keyinput54), .A(n21157), .ZN(n21162) );
  AOI22_X1 U24077 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(keyinput21), 
        .B1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B2(keyinput31), .ZN(n21158) );
  OAI221_X1 U24078 ( .B1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B2(keyinput21), 
        .C1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .C2(keyinput31), .A(n21158), .ZN(
        n21161) );
  AOI22_X1 U24079 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(keyinput60), .B1(
        P1_INSTQUEUE_REG_2__3__SCAN_IN), .B2(keyinput12), .ZN(n21159) );
  OAI221_X1 U24080 ( .B1(P2_LWORD_REG_13__SCAN_IN), .B2(keyinput60), .C1(
        P1_INSTQUEUE_REG_2__3__SCAN_IN), .C2(keyinput12), .A(n21159), .ZN(
        n21160) );
  NOR4_X1 U24081 ( .A1(n21163), .A2(n21162), .A3(n21161), .A4(n21160), .ZN(
        n21184) );
  AOI22_X1 U24082 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(keyinput52), .B1(
        DATAI_13_), .B2(keyinput6), .ZN(n21164) );
  OAI221_X1 U24083 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(keyinput52), .C1(
        DATAI_13_), .C2(keyinput6), .A(n21164), .ZN(n21171) );
  AOI22_X1 U24084 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(keyinput41), .B1(
        P2_INSTQUEUE_REG_14__2__SCAN_IN), .B2(keyinput26), .ZN(n21165) );
  OAI221_X1 U24085 ( .B1(P3_DATAWIDTH_REG_16__SCAN_IN), .B2(keyinput41), .C1(
        P2_INSTQUEUE_REG_14__2__SCAN_IN), .C2(keyinput26), .A(n21165), .ZN(
        n21170) );
  AOI22_X1 U24086 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(keyinput28), 
        .B1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(keyinput49), .ZN(n21166) );
  OAI221_X1 U24087 ( .B1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B2(keyinput28), 
        .C1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .C2(keyinput49), .A(n21166), .ZN(
        n21169) );
  AOI22_X1 U24088 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(keyinput40), 
        .B1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(keyinput15), .ZN(n21167) );
  OAI221_X1 U24089 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput40), 
        .C1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .C2(keyinput15), .A(n21167), .ZN(
        n21168) );
  NOR4_X1 U24090 ( .A1(n21171), .A2(n21170), .A3(n21169), .A4(n21168), .ZN(
        n21183) );
  AOI22_X1 U24091 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput3), .B1(
        P3_STATE2_REG_0__SCAN_IN), .B2(keyinput38), .ZN(n21172) );
  OAI221_X1 U24092 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput3), .C1(
        P3_STATE2_REG_0__SCAN_IN), .C2(keyinput38), .A(n21172), .ZN(n21181) );
  AOI22_X1 U24093 ( .A1(BUF1_REG_28__SCAN_IN), .A2(keyinput42), .B1(
        P1_INSTQUEUE_REG_7__3__SCAN_IN), .B2(keyinput50), .ZN(n21173) );
  OAI221_X1 U24094 ( .B1(BUF1_REG_28__SCAN_IN), .B2(keyinput42), .C1(
        P1_INSTQUEUE_REG_7__3__SCAN_IN), .C2(keyinput50), .A(n21173), .ZN(
        n21180) );
  AOI22_X1 U24095 ( .A1(READY12_REG_SCAN_IN), .A2(keyinput4), .B1(
        P2_INSTQUEUE_REG_10__3__SCAN_IN), .B2(keyinput19), .ZN(n21174) );
  OAI221_X1 U24096 ( .B1(READY12_REG_SCAN_IN), .B2(keyinput4), .C1(
        P2_INSTQUEUE_REG_10__3__SCAN_IN), .C2(keyinput19), .A(n21174), .ZN(
        n21179) );
  AOI22_X1 U24097 ( .A1(n21177), .A2(keyinput17), .B1(keyinput13), .B2(n21176), 
        .ZN(n21175) );
  OAI221_X1 U24098 ( .B1(n21177), .B2(keyinput17), .C1(n21176), .C2(keyinput13), .A(n21175), .ZN(n21178) );
  NOR4_X1 U24099 ( .A1(n21181), .A2(n21180), .A3(n21179), .A4(n21178), .ZN(
        n21182) );
  NAND4_X1 U24100 ( .A1(n21185), .A2(n21184), .A3(n21183), .A4(n21182), .ZN(
        n21252) );
  INV_X1 U24101 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n21187) );
  AOI22_X1 U24102 ( .A1(n21188), .A2(keyinput18), .B1(n21187), .B2(keyinput35), 
        .ZN(n21186) );
  OAI221_X1 U24103 ( .B1(n21188), .B2(keyinput18), .C1(n21187), .C2(keyinput35), .A(n21186), .ZN(n21192) );
  XOR2_X1 U24104 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B(keyinput0), .Z(
        n21191) );
  XNOR2_X1 U24105 ( .A(n21189), .B(keyinput57), .ZN(n21190) );
  OR3_X1 U24106 ( .A1(n21192), .A2(n21191), .A3(n21190), .ZN(n21201) );
  AOI22_X1 U24107 ( .A1(n21195), .A2(keyinput56), .B1(keyinput27), .B2(n21194), 
        .ZN(n21193) );
  OAI221_X1 U24108 ( .B1(n21195), .B2(keyinput56), .C1(n21194), .C2(keyinput27), .A(n21193), .ZN(n21200) );
  AOI22_X1 U24109 ( .A1(n21198), .A2(keyinput34), .B1(n21197), .B2(keyinput33), 
        .ZN(n21196) );
  OAI221_X1 U24110 ( .B1(n21198), .B2(keyinput34), .C1(n21197), .C2(keyinput33), .A(n21196), .ZN(n21199) );
  NOR3_X1 U24111 ( .A1(n21201), .A2(n21200), .A3(n21199), .ZN(n21250) );
  AOI22_X1 U24112 ( .A1(n21203), .A2(keyinput1), .B1(n14353), .B2(keyinput62), 
        .ZN(n21202) );
  OAI221_X1 U24113 ( .B1(n21203), .B2(keyinput1), .C1(n14353), .C2(keyinput62), 
        .A(n21202), .ZN(n21216) );
  AOI22_X1 U24114 ( .A1(n21206), .A2(keyinput8), .B1(n21205), .B2(keyinput2), 
        .ZN(n21204) );
  OAI221_X1 U24115 ( .B1(n21206), .B2(keyinput8), .C1(n21205), .C2(keyinput2), 
        .A(n21204), .ZN(n21215) );
  AOI22_X1 U24116 ( .A1(n21209), .A2(keyinput10), .B1(n21208), .B2(keyinput11), 
        .ZN(n21207) );
  OAI221_X1 U24117 ( .B1(n21209), .B2(keyinput10), .C1(n21208), .C2(keyinput11), .A(n21207), .ZN(n21214) );
  AOI22_X1 U24118 ( .A1(n21212), .A2(keyinput59), .B1(keyinput24), .B2(n21211), 
        .ZN(n21210) );
  OAI221_X1 U24119 ( .B1(n21212), .B2(keyinput59), .C1(n21211), .C2(keyinput24), .A(n21210), .ZN(n21213) );
  NOR4_X1 U24120 ( .A1(n21216), .A2(n21215), .A3(n21214), .A4(n21213), .ZN(
        n21249) );
  AOI22_X1 U24121 ( .A1(n21219), .A2(keyinput44), .B1(n21218), .B2(keyinput9), 
        .ZN(n21217) );
  OAI221_X1 U24122 ( .B1(n21219), .B2(keyinput44), .C1(n21218), .C2(keyinput9), 
        .A(n21217), .ZN(n21231) );
  AOI22_X1 U24123 ( .A1(n21222), .A2(keyinput55), .B1(n21221), .B2(keyinput51), 
        .ZN(n21220) );
  OAI221_X1 U24124 ( .B1(n21222), .B2(keyinput55), .C1(n21221), .C2(keyinput51), .A(n21220), .ZN(n21230) );
  INV_X1 U24125 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n21225) );
  AOI22_X1 U24126 ( .A1(n21225), .A2(keyinput7), .B1(keyinput22), .B2(n21224), 
        .ZN(n21223) );
  OAI221_X1 U24127 ( .B1(n21225), .B2(keyinput7), .C1(n21224), .C2(keyinput22), 
        .A(n21223), .ZN(n21229) );
  AOI22_X1 U24128 ( .A1(n14390), .A2(keyinput25), .B1(keyinput36), .B2(n21227), 
        .ZN(n21226) );
  OAI221_X1 U24129 ( .B1(n14390), .B2(keyinput25), .C1(n21227), .C2(keyinput36), .A(n21226), .ZN(n21228) );
  NOR4_X1 U24130 ( .A1(n21231), .A2(n21230), .A3(n21229), .A4(n21228), .ZN(
        n21248) );
  AOI22_X1 U24131 ( .A1(n21234), .A2(keyinput46), .B1(n21233), .B2(keyinput58), 
        .ZN(n21232) );
  OAI221_X1 U24132 ( .B1(n21234), .B2(keyinput46), .C1(n21233), .C2(keyinput58), .A(n21232), .ZN(n21246) );
  AOI22_X1 U24133 ( .A1(n21237), .A2(keyinput20), .B1(n21236), .B2(keyinput32), 
        .ZN(n21235) );
  OAI221_X1 U24134 ( .B1(n21237), .B2(keyinput20), .C1(n21236), .C2(keyinput32), .A(n21235), .ZN(n21245) );
  AOI22_X1 U24135 ( .A1(n21240), .A2(keyinput29), .B1(n21239), .B2(keyinput48), 
        .ZN(n21238) );
  OAI221_X1 U24136 ( .B1(n21240), .B2(keyinput29), .C1(n21239), .C2(keyinput48), .A(n21238), .ZN(n21244) );
  XOR2_X1 U24137 ( .A(n13523), .B(keyinput14), .Z(n21242) );
  XNOR2_X1 U24138 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B(keyinput37), .ZN(
        n21241) );
  NAND2_X1 U24139 ( .A1(n21242), .A2(n21241), .ZN(n21243) );
  NOR4_X1 U24140 ( .A1(n21246), .A2(n21245), .A3(n21244), .A4(n21243), .ZN(
        n21247) );
  NAND4_X1 U24141 ( .A1(n21250), .A2(n21249), .A3(n21248), .A4(n21247), .ZN(
        n21251) );
  AOI211_X1 U24142 ( .C1(n21254), .C2(n21253), .A(n21252), .B(n21251), .ZN(
        n21257) );
  AOI22_X1 U24143 ( .A1(n21255), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(U215), .ZN(n21256) );
  XNOR2_X1 U24144 ( .A(n21257), .B(n21256), .ZN(U282) );
  AND2_X1 U11125 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13574) );
  AND2_X1 U12449 ( .A1(n10407), .A2(n10406), .ZN(n10559) );
  AND2_X1 U13243 ( .A1(n10408), .A2(n10406), .ZN(n10562) );
  INV_X2 U11203 ( .A(n9675), .ZN(n10452) );
  CLKBUF_X1 U11118 ( .A(n9694), .Z(n11934) );
  CLKBUF_X1 U11130 ( .A(n11148), .Z(n11891) );
  CLKBUF_X1 U11131 ( .A(n11078), .Z(n9694) );
  INV_X1 U11147 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10261) );
  CLKBUF_X1 U11148 ( .A(n10635), .Z(n13953) );
  CLKBUF_X1 U11151 ( .A(n9661), .Z(n12530) );
  CLKBUF_X1 U11156 ( .A(n18935), .Z(n9660) );
  CLKBUF_X1 U11161 ( .A(n11164), .Z(n13248) );
  NAND2_X1 U11181 ( .A1(n14093), .A2(n14092), .ZN(n15011) );
  CLKBUF_X1 U11199 ( .A(n11169), .Z(n15412) );
  CLKBUF_X1 U11258 ( .A(n10345), .Z(n10346) );
  CLKBUF_X1 U11466 ( .A(n10373), .Z(n10393) );
  CLKBUF_X1 U11673 ( .A(n15751), .Z(n15752) );
  CLKBUF_X1 U12485 ( .A(n13202), .Z(n9656) );
  CLKBUF_X1 U12726 ( .A(n15117), .Z(n15142) );
  CLKBUF_X1 U12750 ( .A(n13937), .Z(n9697) );
  CLKBUF_X1 U12938 ( .A(n15720), .Z(n15721) );
  AND3_X1 U13143 ( .A1(n10272), .A2(n10271), .A3(n10270), .ZN(n21259) );
endmodule

