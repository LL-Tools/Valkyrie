

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636;

  AOI211_X1 U4904 ( .C1(n6491), .C2(n6490), .A(n10407), .B(n9883), .ZN(n8623)
         );
  INV_X4 U4905 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X2 U4906 ( .A(n8999), .ZN(n8991) );
  INV_X2 U4907 ( .A(n6538), .ZN(n6732) );
  INV_X1 U4908 ( .A(n6143), .ZN(n6870) );
  CLKBUF_X2 U4909 ( .A(n5423), .Z(n7138) );
  INV_X1 U4910 ( .A(n6384), .ZN(n6337) );
  OAI211_X1 U4911 ( .C1(n7324), .C2(n7396), .A(n6152), .B(n6151), .ZN(n6539)
         );
  BUF_X1 U4912 ( .A(n6140), .Z(n6481) );
  NAND2_X1 U4913 ( .A1(n4449), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6378) );
  AND2_X1 U4914 ( .A1(n4947), .A2(n4946), .ZN(n5313) );
  CLKBUF_X1 U4915 ( .A(n9389), .Z(n4398) );
  NOR2_X1 U4916 ( .A1(n7979), .A2(n10531), .ZN(n9389) );
  AND2_X1 U4917 ( .A1(n9453), .A2(n9024), .ZN(n9009) );
  OAI21_X1 U4918 ( .B1(n8430), .B2(n5043), .A(n5041), .ZN(n5048) );
  INV_X1 U4919 ( .A(n8868), .ZN(n4730) );
  BUF_X1 U4920 ( .A(n5366), .Z(n5374) );
  OR2_X1 U4921 ( .A1(n9182), .A2(n9183), .ZN(n9196) );
  NAND2_X1 U4922 ( .A1(n4655), .A2(n7084), .ZN(n9354) );
  INV_X1 U4923 ( .A(n6732), .ZN(n6748) );
  INV_X1 U4924 ( .A(n4593), .ZN(n9656) );
  OAI21_X1 U4925 ( .B1(n9934), .B2(n4986), .A(n4984), .ZN(n9906) );
  XNOR2_X1 U4926 ( .A(n9291), .B(n9304), .ZN(n9290) );
  OR2_X1 U4927 ( .A1(n9507), .A2(n9358), .ZN(n9326) );
  INV_X1 U4928 ( .A(n4641), .ZN(n7896) );
  NAND2_X1 U4929 ( .A1(n6513), .A2(n7023), .ZN(n6515) );
  INV_X2 U4930 ( .A(n6485), .ZN(n6869) );
  AOI21_X1 U4931 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(n9907) );
  INV_X1 U4932 ( .A(n8332), .ZN(n10464) );
  CLKBUF_X3 U4933 ( .A(n9181), .Z(n4402) );
  OAI21_X1 U4934 ( .B1(n5220), .B2(n5218), .A(n5213), .ZN(n7088) );
  INV_X1 U4935 ( .A(n8837), .ZN(n9456) );
  NAND2_X1 U4936 ( .A1(n4752), .A2(n6138), .ZN(n6526) );
  AOI21_X1 U4937 ( .B1(n9931), .B2(n6337), .A(n6336), .ZN(n9702) );
  XNOR2_X1 U4938 ( .A(n6045), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6048) );
  NAND4_X2 U4939 ( .A1(n5465), .A2(n5464), .A3(n5463), .A4(n5462), .ZN(n9034)
         );
  MUX2_X1 U4940 ( .A(n9189), .B(n9188), .S(n9187), .Z(n9190) );
  MUX2_X1 U4941 ( .A(n9395), .B(n9454), .S(n10578), .Z(n9397) );
  MUX2_X1 U4942 ( .A(n9455), .B(n9454), .S(n10571), .Z(n9458) );
  AOI21_X1 U4943 ( .B1(n9966), .B2(n6337), .A(n6320), .ZN(n9663) );
  INV_X1 U4944 ( .A(n6513), .ZN(n8270) );
  OAI21_X4 U4945 ( .B1(n5845), .B2(n5844), .A(n5856), .ZN(n8455) );
  NAND2_X2 U4946 ( .A1(n4642), .A2(n7081), .ZN(n8430) );
  NAND2_X2 U4947 ( .A1(n4850), .A2(n4849), .ZN(n8275) );
  NAND2_X2 U4948 ( .A1(n8163), .A2(n8859), .ZN(n4850) );
  AND2_X2 U4949 ( .A1(n5314), .A2(n4513), .ZN(n5138) );
  NAND4_X2 U4950 ( .A1(n6022), .A2(n6021), .A3(n6020), .A4(n6019), .ZN(n6234)
         );
  AND3_X2 U4951 ( .A1(n6220), .A2(n4685), .A3(n4684), .ZN(n6022) );
  NAND2_X4 U4952 ( .A1(n5588), .A2(n5587), .ZN(n8485) );
  XNOR2_X2 U4953 ( .A(n4681), .B(n5753), .ZN(n8150) );
  XNOR2_X2 U4954 ( .A(n5792), .B(n5791), .ZN(n8426) );
  NAND3_X2 U4955 ( .A1(n4846), .A2(n4845), .A3(n8885), .ZN(n8064) );
  INV_X2 U4956 ( .A(n6885), .ZN(n10333) );
  NAND2_X2 U4957 ( .A1(n6563), .A2(n6562), .ZN(n8154) );
  NAND2_X2 U4958 ( .A1(n8676), .A2(n5805), .ZN(n8757) );
  NOR2_X2 U4959 ( .A1(n6208), .A2(n6207), .ZN(n6210) );
  NAND2_X2 U4960 ( .A1(n6274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6275) );
  NAND2_X2 U4961 ( .A1(n5295), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5297) );
  XNOR2_X2 U4962 ( .A(n6033), .B(n7745), .ZN(n6123) );
  NAND2_X2 U4963 ( .A1(n4606), .A2(n6295), .ZN(n10113) );
  NAND2_X2 U4964 ( .A1(n6115), .A2(n6123), .ZN(n7324) );
  NAND2_X2 U4965 ( .A1(n8192), .A2(n8901), .ZN(n8163) );
  OAI21_X2 U4966 ( .B1(n5310), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5325) );
  NAND2_X4 U4967 ( .A1(n5967), .A2(n9020), .ZN(n8999) );
  NAND2_X1 U4968 ( .A1(n5967), .A2(n8992), .ZN(n7104) );
  XNOR2_X2 U4969 ( .A(n5301), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5967) );
  INV_X1 U4970 ( .A(n5378), .ZN(n9199) );
  NAND2_X2 U4971 ( .A1(n5822), .A2(n5821), .ZN(n9291) );
  NAND2_X1 U4972 ( .A1(n7126), .A2(n7125), .ZN(n9278) );
  INV_X1 U4973 ( .A(n10079), .ZN(n7014) );
  NAND2_X1 U4974 ( .A1(n8259), .A2(n8260), .ZN(n5545) );
  NAND2_X1 U4975 ( .A1(n7258), .A2(n8010), .ZN(n8117) );
  NAND2_X1 U4976 ( .A1(n7249), .A2(n7865), .ZN(n7933) );
  INV_X4 U4977 ( .A(n6746), .ZN(n6726) );
  INV_X1 U4978 ( .A(n9030), .ZN(n8535) );
  INV_X1 U4979 ( .A(n5536), .ZN(n4399) );
  INV_X2 U4980 ( .A(n7022), .ZN(n7010) );
  AND3_X1 U4981 ( .A1(n5100), .A2(n5099), .A3(n7982), .ZN(n8867) );
  INV_X1 U4982 ( .A(n7060), .ZN(n10555) );
  INV_X1 U4983 ( .A(n5987), .ZN(n4407) );
  INV_X1 U4984 ( .A(n5624), .ZN(n5218) );
  NAND2_X4 U4985 ( .A1(n5971), .A2(n5743), .ZN(n7161) );
  CLKBUF_X1 U4986 ( .A(n6150), .Z(n4400) );
  BUF_X1 U4987 ( .A(n7176), .Z(n4746) );
  INV_X4 U4988 ( .A(n9198), .ZN(n5743) );
  INV_X2 U4989 ( .A(n8628), .ZN(n4966) );
  OAI21_X1 U4990 ( .B1(n7290), .B2(n4829), .A(n4828), .ZN(n4827) );
  NAND2_X1 U4991 ( .A1(n4791), .A2(n4720), .ZN(n5484) );
  NOR2_X1 U4992 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5308) );
  NOR2_X1 U4993 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5307) );
  AND2_X1 U4994 ( .A1(n4871), .A2(n7145), .ZN(n4425) );
  OAI21_X1 U4995 ( .B1(n8775), .B2(n4631), .A(n4629), .ZN(n6788) );
  OR2_X1 U4996 ( .A1(n8634), .A2(n6755), .ZN(n6781) );
  AND2_X1 U4997 ( .A1(n5025), .A2(n4598), .ZN(n8634) );
  AND2_X1 U4998 ( .A1(n5025), .A2(n5023), .ZN(n9700) );
  AND2_X1 U4999 ( .A1(n5028), .A2(n5026), .ZN(n9699) );
  AOI21_X1 U5000 ( .B1(n5071), .B2(n10541), .A(n4780), .ZN(n9454) );
  CLKBUF_X1 U5001 ( .A(n9656), .Z(n4751) );
  AOI21_X1 U5002 ( .B1(n4813), .B2(n10541), .A(n4811), .ZN(n9461) );
  AOI21_X1 U5003 ( .B1(n9247), .B2(n7097), .A(n7096), .ZN(n9236) );
  XNOR2_X1 U5004 ( .A(n9247), .B(n4958), .ZN(n4813) );
  XNOR2_X1 U5005 ( .A(n9899), .B(n9904), .ZN(n10163) );
  OAI21_X1 U5006 ( .B1(n9247), .B2(n5228), .A(n5225), .ZN(n7099) );
  OR2_X1 U5007 ( .A1(n9915), .A2(n9898), .ZN(n9899) );
  NAND2_X1 U5008 ( .A1(n4592), .A2(n4590), .ZN(n4595) );
  AOI21_X1 U5009 ( .B1(n4963), .B2(n4964), .A(n4479), .ZN(n4607) );
  OR2_X1 U5010 ( .A1(n10161), .A2(n10509), .ZN(n4756) );
  NAND2_X1 U5011 ( .A1(n4711), .A2(n4462), .ZN(n9914) );
  AND2_X1 U5012 ( .A1(n8616), .A2(n6492), .ZN(n6506) );
  AND2_X1 U5013 ( .A1(n4548), .A2(n4547), .ZN(n9942) );
  OR2_X1 U5014 ( .A1(n10093), .A2(n10402), .ZN(n4548) );
  AOI21_X1 U5015 ( .B1(n6489), .B2(n10399), .A(n6488), .ZN(n8616) );
  AND2_X1 U5016 ( .A1(n4550), .A2(n4549), .ZN(n10093) );
  NAND2_X1 U5017 ( .A1(n6391), .A2(n10399), .ZN(n4824) );
  AOI21_X1 U5018 ( .B1(n5005), .B2(n10528), .A(n5004), .ZN(n5003) );
  OAI21_X1 U5019 ( .B1(n4894), .B2(n10048), .A(n9926), .ZN(n10086) );
  NAND2_X1 U5020 ( .A1(n6868), .A2(n6867), .ZN(n7013) );
  AND2_X1 U5021 ( .A1(n6397), .A2(n4823), .ZN(n4822) );
  OR2_X1 U5022 ( .A1(n9907), .A2(n4578), .ZN(n5007) );
  AOI21_X1 U5023 ( .B1(n7014), .B2(n6874), .A(n7006), .ZN(n7035) );
  NAND2_X1 U5024 ( .A1(n8805), .A2(n8804), .ZN(n8840) );
  AOI21_X1 U5025 ( .B1(n10017), .B2(n6443), .A(n4704), .ZN(n10002) );
  NOR2_X1 U5026 ( .A1(n4456), .A2(n5010), .ZN(n5009) );
  OR2_X1 U5027 ( .A1(n4877), .A2(n7102), .ZN(n4876) );
  AND2_X1 U5028 ( .A1(n9887), .A2(n6396), .ZN(n6397) );
  AOI21_X1 U5029 ( .B1(n5123), .B2(n5122), .A(n5121), .ZN(n5120) );
  NAND2_X1 U5030 ( .A1(n9993), .A2(n4992), .ZN(n4989) );
  NAND2_X1 U5031 ( .A1(n6859), .A2(n6862), .ZN(n9533) );
  NOR2_X1 U5032 ( .A1(n7005), .A2(n7006), .ZN(n7008) );
  AOI21_X1 U5033 ( .B1(n4987), .B2(n4567), .A(n4566), .ZN(n4565) );
  NAND2_X1 U5034 ( .A1(n4703), .A2(n4701), .ZN(n10030) );
  AND2_X1 U5035 ( .A1(n4816), .A2(n6338), .ZN(n4820) );
  OR2_X1 U5036 ( .A1(n6858), .A2(n6857), .ZN(n6862) );
  INV_X1 U5037 ( .A(n8618), .ZN(n6491) );
  NAND2_X1 U5038 ( .A1(n7101), .A2(n7100), .ZN(n8646) );
  NAND2_X1 U5039 ( .A1(n10005), .A2(n10004), .ZN(n10003) );
  NOR2_X1 U5040 ( .A1(n8847), .A2(n5115), .ZN(n5114) );
  AOI21_X1 U5041 ( .B1(n5253), .B2(n9961), .A(n4475), .ZN(n5252) );
  NAND2_X1 U5042 ( .A1(n7129), .A2(n7128), .ZN(n9234) );
  OR2_X1 U5043 ( .A1(n5053), .A2(n5050), .ZN(n5049) );
  AND2_X1 U5044 ( .A1(n5940), .A2(n5939), .ZN(n8837) );
  AND2_X1 U5045 ( .A1(n6353), .A2(n6365), .ZN(n9891) );
  NAND2_X1 U5046 ( .A1(n9964), .A2(n9955), .ZN(n9949) );
  XNOR2_X1 U5047 ( .A(n6843), .B(SI_29_), .ZN(n9536) );
  OR2_X1 U5048 ( .A1(n9249), .A2(n9398), .ZN(n7129) );
  OR2_X1 U5049 ( .A1(n9469), .A2(n9026), .ZN(n8975) );
  NAND2_X1 U5050 ( .A1(n5927), .A2(n5926), .ZN(n9398) );
  OR2_X1 U5051 ( .A1(n9481), .A2(n9288), .ZN(n8845) );
  NOR2_X1 U5052 ( .A1(n9290), .A2(n5058), .ZN(n5057) );
  NAND2_X1 U5053 ( .A1(n5545), .A2(n4470), .ZN(n8340) );
  NAND3_X1 U5054 ( .A1(n6476), .A2(n6475), .A3(n6474), .ZN(n6843) );
  XNOR2_X1 U5055 ( .A(n6846), .B(n6845), .ZN(n8639) );
  AOI21_X1 U5056 ( .B1(n4854), .B2(n4857), .A(n4487), .ZN(n4851) );
  NAND2_X1 U5057 ( .A1(n5892), .A2(n5891), .ZN(n9469) );
  OR2_X1 U5058 ( .A1(n10087), .A2(n9603), .ZN(n6987) );
  OR2_X1 U5059 ( .A1(n9475), .A2(n8974), .ZN(n8971) );
  INV_X1 U5060 ( .A(n10102), .ZN(n9968) );
  OR2_X1 U5061 ( .A1(n6465), .A2(n6462), .ZN(n6476) );
  NAND2_X1 U5062 ( .A1(n6331), .A2(n6330), .ZN(n10091) );
  AND2_X1 U5063 ( .A1(n4855), .A2(n7122), .ZN(n4854) );
  INV_X2 U5064 ( .A(n7093), .ZN(n9481) );
  AOI21_X1 U5065 ( .B1(n5056), .B2(n4420), .A(n4472), .ZN(n5055) );
  INV_X1 U5066 ( .A(n7095), .ZN(n9463) );
  NAND2_X1 U5067 ( .A1(n5937), .A2(n5936), .ZN(n6465) );
  XNOR2_X1 U5068 ( .A(n5937), .B(n5936), .ZN(n8626) );
  INV_X1 U5069 ( .A(n9729), .ZN(n4609) );
  AND2_X1 U5070 ( .A1(n5847), .A2(n5846), .ZN(n7093) );
  OR2_X1 U5071 ( .A1(n10097), .A2(n9604), .ZN(n6825) );
  AND2_X1 U5072 ( .A1(n8955), .A2(n4860), .ZN(n4859) );
  OAI21_X1 U5073 ( .B1(n10046), .B2(n5107), .A(n10031), .ZN(n5106) );
  OR2_X1 U5074 ( .A1(n9491), .A2(n9317), .ZN(n8964) );
  NAND2_X1 U5075 ( .A1(n5921), .A2(n5920), .ZN(n5937) );
  NOR2_X1 U5076 ( .A1(n10118), .A2(n5077), .ZN(n5076) );
  OR2_X1 U5077 ( .A1(n10313), .A2(n6942), .ZN(n4571) );
  NAND2_X1 U5078 ( .A1(n7076), .A2(n7075), .ZN(n8308) );
  NAND2_X1 U5079 ( .A1(n6305), .A2(n6304), .ZN(n10108) );
  NAND2_X1 U5080 ( .A1(n4575), .A2(n4573), .ZN(n10313) );
  AND2_X1 U5081 ( .A1(n8849), .A2(n9326), .ZN(n8955) );
  NAND2_X1 U5082 ( .A1(n5794), .A2(n5793), .ZN(n9491) );
  AND2_X1 U5083 ( .A1(n6955), .A2(n6952), .ZN(n10031) );
  NAND2_X1 U5084 ( .A1(n9569), .A2(n6552), .ZN(n7996) );
  OAI21_X1 U5085 ( .B1(n5263), .B2(n4481), .A(n4417), .ZN(n4707) );
  AOI21_X1 U5086 ( .B1(n5014), .B2(n5019), .A(n5013), .ZN(n5012) );
  AND2_X1 U5087 ( .A1(n6817), .A2(n6818), .ZN(n10046) );
  OR2_X1 U5088 ( .A1(n9329), .A2(n9318), .ZN(n8849) );
  NAND2_X1 U5089 ( .A1(n9298), .A2(n8960), .ZN(n8810) );
  NAND2_X1 U5090 ( .A1(n8946), .A2(n8949), .ZN(n9355) );
  OR2_X1 U5091 ( .A1(n10325), .A2(n4576), .ZN(n4575) );
  NOR2_X1 U5092 ( .A1(n10128), .A2(n10123), .ZN(n5078) );
  OAI21_X1 U5093 ( .B1(n5264), .B2(n5266), .A(n4490), .ZN(n5263) );
  OAI21_X1 U5094 ( .B1(n5883), .B2(n4911), .A(n4908), .ZN(n5905) );
  INV_X1 U5095 ( .A(n5193), .ZN(n5192) );
  XNOR2_X1 U5096 ( .A(n5820), .B(n5831), .ZN(n8437) );
  NAND2_X1 U5097 ( .A1(n10326), .A2(n10333), .ZN(n10325) );
  AND2_X1 U5098 ( .A1(n8522), .A2(n5268), .ZN(n5265) );
  NAND2_X1 U5099 ( .A1(n5745), .A2(n5744), .ZN(n9329) );
  INV_X1 U5100 ( .A(n5091), .ZN(n5090) );
  INV_X1 U5101 ( .A(n4574), .ZN(n4573) );
  NAND2_X1 U5102 ( .A1(n7088), .A2(n9333), .ZN(n8960) );
  NAND2_X1 U5103 ( .A1(n4924), .A2(n4928), .ZN(n5856) );
  NAND2_X1 U5104 ( .A1(n5759), .A2(n5758), .ZN(n9507) );
  NAND2_X1 U5105 ( .A1(n6279), .A2(n6278), .ZN(n10123) );
  AND2_X1 U5106 ( .A1(n6940), .A2(n6813), .ZN(n10063) );
  NAND2_X1 U5107 ( .A1(n6266), .A2(n6265), .ZN(n10128) );
  AOI211_X1 U5108 ( .C1(n8332), .C2(n9693), .A(n8331), .B(n8330), .ZN(n8333)
         );
  NOR2_X1 U5109 ( .A1(n5082), .A2(n10143), .ZN(n5081) );
  NAND2_X1 U5110 ( .A1(n5843), .A2(n5840), .ZN(n5820) );
  AND2_X1 U5111 ( .A1(n5843), .A2(n5840), .ZN(n5832) );
  NAND2_X1 U5112 ( .A1(n4745), .A2(n4744), .ZN(n7868) );
  INV_X1 U5113 ( .A(n10133), .ZN(n10054) );
  NAND2_X1 U5114 ( .A1(n6254), .A2(n6253), .ZN(n10133) );
  AND2_X1 U5115 ( .A1(n5724), .A2(n5723), .ZN(n9363) );
  NAND2_X1 U5116 ( .A1(n5703), .A2(n5702), .ZN(n9514) );
  OR2_X1 U5117 ( .A1(n5806), .A2(n4930), .ZN(n5843) );
  OR2_X1 U5118 ( .A1(n6324), .A2(n6332), .ZN(n9640) );
  OR2_X1 U5119 ( .A1(n9521), .A2(n8708), .ZN(n8942) );
  AND2_X1 U5120 ( .A1(n8518), .A2(n6924), .ZN(n10318) );
  AND2_X1 U5121 ( .A1(n4577), .A2(n6804), .ZN(n10326) );
  NAND2_X1 U5122 ( .A1(n5769), .A2(n5768), .ZN(n5806) );
  AOI21_X1 U5123 ( .B1(n7985), .B2(n5036), .A(n6245), .ZN(n6250) );
  OR2_X1 U5124 ( .A1(n10317), .A2(n8417), .ZN(n8518) );
  AND2_X1 U5125 ( .A1(n8508), .A2(n10504), .ZN(n5083) );
  NAND2_X1 U5126 ( .A1(n6238), .A2(n6237), .ZN(n10143) );
  NAND2_X1 U5127 ( .A1(n5679), .A2(n5678), .ZN(n9521) );
  INV_X1 U5128 ( .A(n6926), .ZN(n6921) );
  OAI21_X1 U5129 ( .B1(n6884), .B2(n6188), .A(n6887), .ZN(n6804) );
  OAI21_X1 U5130 ( .B1(n8027), .B2(n7066), .A(n7065), .ZN(n8065) );
  OAI21_X1 U5131 ( .B1(n4559), .B2(n5132), .A(n4557), .ZN(n8179) );
  NAND2_X1 U5132 ( .A1(n5628), .A2(n5627), .ZN(n8921) );
  NAND2_X1 U5133 ( .A1(n4917), .A2(n4916), .ZN(n5769) );
  OAI211_X1 U5134 ( .C1(n5697), .C2(n4901), .A(n4897), .B(n4895), .ZN(n8127)
         );
  OR2_X1 U5135 ( .A1(n8485), .A2(n8535), .ZN(n8914) );
  OR2_X1 U5136 ( .A1(n5697), .A2(n4920), .ZN(n4915) );
  INV_X1 U5137 ( .A(n8590), .ZN(n10504) );
  AND2_X1 U5138 ( .A1(n5641), .A2(n5640), .ZN(n8926) );
  NAND2_X1 U5139 ( .A1(n6226), .A2(n6225), .ZN(n10147) );
  AND2_X1 U5140 ( .A1(n6912), .A2(n10341), .ZN(n8288) );
  AND2_X1 U5141 ( .A1(n4433), .A2(n10464), .ZN(n4779) );
  OAI21_X1 U5142 ( .B1(n4434), .B2(n6915), .A(n6927), .ZN(n6187) );
  NAND2_X1 U5143 ( .A1(n5659), .A2(n5658), .ZN(n8934) );
  AOI21_X1 U5144 ( .B1(n4560), .B2(n4558), .A(n6905), .ZN(n4557) );
  AND2_X1 U5145 ( .A1(n8895), .A2(n8897), .ZN(n8814) );
  NAND2_X1 U5146 ( .A1(n6908), .A2(n6903), .ZN(n8178) );
  OR2_X1 U5147 ( .A1(n10489), .A2(n8496), .ZN(n10310) );
  OR2_X1 U5148 ( .A1(n7321), .A2(n5218), .ZN(n5588) );
  OR2_X1 U5149 ( .A1(n7527), .A2(n5636), .ZN(n5641) );
  NAND2_X2 U5150 ( .A1(n4602), .A2(n5673), .ZN(n5697) );
  OR2_X1 U5151 ( .A1(n6101), .A2(n8553), .ZN(n6919) );
  NAND2_X1 U5152 ( .A1(n6904), .A2(n5281), .ZN(n8093) );
  NAND2_X1 U5153 ( .A1(n6206), .A2(n6205), .ZN(n10489) );
  OR2_X1 U5154 ( .A1(n7416), .A2(n7417), .ZN(n7429) );
  NAND2_X1 U5155 ( .A1(n5598), .A2(n5597), .ZN(n8530) );
  NAND2_X1 U5156 ( .A1(n5585), .A2(n5593), .ZN(n7321) );
  NAND2_X1 U5157 ( .A1(n5671), .A2(n5670), .ZN(n4602) );
  OR2_X1 U5158 ( .A1(n7111), .A2(n8059), .ZN(n8895) );
  NAND2_X2 U5159 ( .A1(n7979), .A2(n10533), .ZN(n9385) );
  NAND2_X1 U5160 ( .A1(n10391), .A2(n10446), .ZN(n10389) );
  NAND2_X1 U5161 ( .A1(n6383), .A2(n6382), .ZN(n10399) );
  AND2_X1 U5162 ( .A1(n5535), .A2(n5534), .ZN(n7070) );
  OAI211_X1 U5163 ( .C1(n7324), .C2(n7400), .A(n6176), .B(n6175), .ZN(n8094)
         );
  OR2_X1 U5164 ( .A1(n5616), .A2(n5615), .ZN(n5243) );
  NAND2_X1 U5165 ( .A1(n4996), .A2(n6083), .ZN(n8468) );
  AND2_X1 U5166 ( .A1(n5494), .A2(n5493), .ZN(n8059) );
  OAI21_X1 U5167 ( .B1(n5579), .B2(n4886), .A(n4883), .ZN(n5616) );
  INV_X1 U5168 ( .A(n5400), .ZN(n5760) );
  XNOR2_X1 U5169 ( .A(n5551), .B(n5550), .ZN(n7308) );
  NAND2_X1 U5170 ( .A1(n7185), .A2(n7296), .ZN(n7468) );
  INV_X2 U5171 ( .A(n4407), .ZN(n4408) );
  NAND3_X1 U5172 ( .A1(n4450), .A2(n6131), .A3(n6128), .ZN(n7335) );
  NAND2_X1 U5173 ( .A1(n7225), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7504) );
  NAND2_X1 U5174 ( .A1(n5209), .A2(n5207), .ZN(n5551) );
  BUF_X1 U5175 ( .A(n7054), .Z(n4404) );
  NAND4_X2 U5176 ( .A1(n5429), .A2(n5428), .A3(n5427), .A4(n5426), .ZN(n9035)
         );
  AOI22_X1 U5177 ( .A1(n4405), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6276), .B2(
        n9821), .ZN(n6083) );
  AND4_X1 U5178 ( .A1(n6158), .A2(n6157), .A3(n6156), .A4(n6155), .ZN(n7999)
         );
  OR2_X1 U5179 ( .A1(n7161), .A2(n5967), .ZN(n5328) );
  CLKBUF_X1 U5180 ( .A(n5421), .Z(n8403) );
  NAND2_X1 U5182 ( .A1(n4966), .A2(n7023), .ZN(n6509) );
  NAND2_X1 U5183 ( .A1(n6412), .A2(n6376), .ZN(n8438) );
  INV_X1 U5184 ( .A(n5660), .ZN(n5646) );
  OR2_X1 U5185 ( .A1(n5720), .A2(n7294), .ZN(n5390) );
  BUF_X1 U5186 ( .A(n9181), .Z(n4401) );
  AOI21_X1 U5187 ( .B1(n5515), .B2(n5208), .A(n5210), .ZN(n5207) );
  AND2_X1 U5188 ( .A1(n9534), .A2(n5374), .ZN(n5660) );
  XNOR2_X1 U5189 ( .A(n6406), .B(n6405), .ZN(n8489) );
  MUX2_X1 U5190 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10228), .S(n7324), .Z(n7953)
         );
  NAND2_X1 U5191 ( .A1(n5300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5301) );
  NAND2_X2 U5192 ( .A1(n6048), .A2(n6046), .ZN(n6384) );
  NAND2_X2 U5193 ( .A1(n10219), .A2(n6049), .ZN(n6143) );
  XNOR2_X1 U5194 ( .A(n5299), .B(n5298), .ZN(n5971) );
  NOR2_X1 U5195 ( .A1(n6049), .A2(n6048), .ZN(n6140) );
  NAND2_X1 U5196 ( .A1(n4449), .A2(n6381), .ZN(n7023) );
  XNOR2_X1 U5197 ( .A(n6409), .B(n6408), .ZN(n10227) );
  NOR2_X1 U5198 ( .A1(n4661), .A2(n4660), .ZN(n5507) );
  NAND2_X1 U5199 ( .A1(n5446), .A2(n5466), .ZN(n7431) );
  INV_X1 U5200 ( .A(n6048), .ZN(n10219) );
  INV_X1 U5201 ( .A(n4880), .ZN(n5515) );
  OAI21_X1 U5202 ( .B1(n6404), .B2(n6403), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6406) );
  XNOR2_X1 U5203 ( .A(n6400), .B(n6399), .ZN(n8580) );
  OAI21_X1 U5204 ( .B1(n4827), .B2(SI_7_), .A(n5531), .ZN(n4880) );
  INV_X1 U5205 ( .A(n5531), .ZN(n5210) );
  NAND2_X1 U5206 ( .A1(n4747), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U5207 ( .A1(n10212), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6045) );
  OAI21_X2 U5208 ( .B1(n5340), .B2(n5140), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5344) );
  NAND2_X1 U5209 ( .A1(n4536), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4535) );
  NAND2_X1 U5210 ( .A1(n4827), .A2(SI_7_), .ZN(n5531) );
  INV_X1 U5211 ( .A(n5657), .ZN(n5294) );
  AND2_X2 U5212 ( .A1(n5203), .A2(n4627), .ZN(n5637) );
  NOR2_X1 U5213 ( .A1(n5302), .A2(n5309), .ZN(n5968) );
  XNOR2_X1 U5214 ( .A(n5546), .B(SI_8_), .ZN(n5550) );
  NAND2_X1 U5215 ( .A1(n4616), .A2(n4614), .ZN(n7520) );
  NAND2_X2 U5216 ( .A1(n7290), .A2(P1_U3086), .ZN(n10224) );
  INV_X1 U5217 ( .A(n5484), .ZN(n4627) );
  AND3_X1 U5218 ( .A1(n4454), .A2(n4553), .A3(n4552), .ZN(n4554) );
  NOR2_X1 U5219 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  NAND2_X1 U5220 ( .A1(n4435), .A2(n7745), .ZN(n5137) );
  NAND2_X1 U5221 ( .A1(n7598), .A2(n5315), .ZN(n5140) );
  NAND2_X1 U5222 ( .A1(n6120), .A2(n6023), .ZN(n6135) );
  AND2_X1 U5223 ( .A1(n5293), .A2(n5292), .ZN(n4791) );
  NAND4_X1 U5224 ( .A1(n5308), .A2(n5307), .A3(n5291), .A4(n5290), .ZN(n5285)
         );
  NAND2_X2 U5225 ( .A1(n8370), .A2(n5329), .ZN(n5331) );
  INV_X1 U5226 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7626) );
  INV_X1 U5227 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5324) );
  INV_X1 U5228 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6408) );
  INV_X1 U5229 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6370) );
  INV_X1 U5230 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5291) );
  INV_X1 U5231 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5290) );
  NOR2_X1 U5232 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6024) );
  NOR2_X1 U5233 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6021) );
  NOR2_X1 U5234 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6020) );
  NOR2_X1 U5235 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6019) );
  INV_X1 U5236 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6220) );
  NOR2_X1 U5237 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5292) );
  NOR2_X1 U5238 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5293) );
  NOR2_X1 U5239 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6034) );
  INV_X1 U5240 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6402) );
  INV_X1 U5241 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4947) );
  INV_X1 U5242 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5675) );
  INV_X1 U5243 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6368) );
  INV_X4 U5244 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5245 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7562) );
  AND2_X1 U5246 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8369) );
  NOR2_X1 U5247 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4944) );
  NOR2_X1 U5248 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4942) );
  NOR2_X1 U5249 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4941) );
  NOR2_X1 U5250 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n4943) );
  AND2_X2 U5251 ( .A1(n4586), .A2(n4584), .ZN(n9570) );
  XNOR2_X1 U5252 ( .A(n8723), .B(n8722), .ZN(n8724) );
  OAI22_X1 U5253 ( .A1(n8724), .A2(n9269), .B1(n8723), .B2(n8722), .ZN(n8727)
         );
  INV_X4 U5254 ( .A(n5487), .ZN(n7290) );
  NAND2_X2 U5255 ( .A1(n9570), .A2(n9571), .ZN(n9569) );
  NAND2_X1 U5256 ( .A1(n7290), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n4828) );
  NAND2_X2 U5257 ( .A1(n9278), .A2(n8845), .ZN(n7127) );
  NOR2_X2 U5258 ( .A1(n9918), .A2(n10083), .ZN(n9900) );
  NOR2_X2 U5259 ( .A1(n6268), .A2(n6267), .ZN(n6288) );
  OAI21_X2 U5260 ( .B1(n9656), .B2(n9660), .A(n9559), .ZN(n9634) );
  NAND2_X2 U5261 ( .A1(n7556), .A2(n7557), .ZN(n7555) );
  INV_X2 U5262 ( .A(n9199), .ZN(n9181) );
  NAND2_X4 U5263 ( .A1(n5331), .A2(n5330), .ZN(n4414) );
  NAND2_X4 U5264 ( .A1(n8369), .A2(n7562), .ZN(n5330) );
  INV_X2 U5265 ( .A(n10535), .ZN(n4635) );
  NAND2_X2 U5266 ( .A1(n7108), .A2(n8874), .ZN(n10535) );
  OR2_X1 U5267 ( .A1(n6517), .A2(n6516), .ZN(n5272) );
  NAND2_X1 U5268 ( .A1(n6514), .A2(n7455), .ZN(n4403) );
  NAND3_X2 U5269 ( .A1(n4633), .A2(n4632), .A3(n7061), .ZN(n8027) );
  OAI22_X2 U5270 ( .A1(n10334), .A2(n10333), .B1(n9744), .B2(n10335), .ZN(
        n8412) );
  OR2_X1 U5271 ( .A1(n10102), .A2(n9663), .ZN(n6978) );
  NOR2_X2 U5272 ( .A1(n9949), .A2(n10091), .ZN(n5085) );
  INV_X1 U5273 ( .A(n4412), .ZN(n4405) );
  INV_X1 U5274 ( .A(n4412), .ZN(n4406) );
  OAI21_X2 U5275 ( .B1(n8248), .B2(n5015), .A(n5012), .ZN(n8550) );
  NAND3_X2 U5276 ( .A1(n6564), .A2(n8154), .A3(n6575), .ZN(n8248) );
  INV_X1 U5277 ( .A(n6364), .ZN(n4409) );
  INV_X1 U5278 ( .A(n6364), .ZN(n4410) );
  NAND2_X1 U5279 ( .A1(n7324), .A2(n5487), .ZN(n6364) );
  NAND2_X1 U5280 ( .A1(n4814), .A2(n7972), .ZN(n4411) );
  INV_X2 U5281 ( .A(n5760), .ZN(n5536) );
  NAND2_X1 U5282 ( .A1(n7324), .A2(n7290), .ZN(n6150) );
  NAND2_X1 U5283 ( .A1(n5331), .A2(n5330), .ZN(n4413) );
  XNOR2_X2 U5284 ( .A(n4700), .B(n6042), .ZN(n6115) );
  AOI21_X1 U5285 ( .B1(n5250), .B2(n5252), .A(n5249), .ZN(n5248) );
  INV_X1 U5286 ( .A(n5253), .ZN(n5250) );
  NAND2_X1 U5287 ( .A1(n4532), .A2(n6908), .ZN(n6909) );
  NAND2_X1 U5288 ( .A1(n6907), .A2(n6906), .ZN(n4532) );
  OR2_X1 U5289 ( .A1(n8646), .A2(n9025), .ZN(n9007) );
  OR2_X1 U5290 ( .A1(n5287), .A2(n7132), .ZN(n4877) );
  NAND2_X1 U5291 ( .A1(n9231), .A2(n4419), .ZN(n4878) );
  NOR2_X1 U5292 ( .A1(n5116), .A2(n5112), .ZN(n5111) );
  INV_X1 U5293 ( .A(n8971), .ZN(n5112) );
  AND2_X1 U5294 ( .A1(n5055), .A2(n4512), .ZN(n5053) );
  AND2_X1 U5295 ( .A1(n9475), .A2(n8974), .ZN(n8847) );
  OR2_X1 U5296 ( .A1(n9514), .A2(n9359), .ZN(n8948) );
  NAND2_X1 U5297 ( .A1(n4735), .A2(n4734), .ZN(n6530) );
  XNOR2_X1 U5298 ( .A(n6511), .B(n4750), .ZN(n4555) );
  NAND2_X1 U5299 ( .A1(n4906), .A2(n4469), .ZN(n5242) );
  NAND2_X1 U5300 ( .A1(n8995), .A2(n8994), .ZN(n8996) );
  INV_X1 U5301 ( .A(n10565), .ZN(n9443) );
  NAND2_X1 U5302 ( .A1(n8863), .A2(n8869), .ZN(n10565) );
  XNOR2_X1 U5303 ( .A(n4763), .B(n4403), .ZN(n6517) );
  AOI21_X1 U5304 ( .B1(n5248), .B2(n5251), .A(n4492), .ZN(n5246) );
  INV_X1 U5305 ( .A(n5252), .ZN(n5251) );
  NAND2_X1 U5306 ( .A1(n9960), .A2(n5248), .ZN(n4710) );
  AND2_X1 U5307 ( .A1(n8950), .A2(n9311), .ZN(n4955) );
  INV_X1 U5308 ( .A(n8965), .ZN(n4667) );
  NAND2_X1 U5309 ( .A1(n6171), .A2(n4463), .ZN(n6907) );
  NAND2_X1 U5310 ( .A1(n7440), .A2(n7184), .ZN(n7185) );
  NOR2_X1 U5311 ( .A1(n8004), .A2(n9750), .ZN(n6433) );
  INV_X1 U5312 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5735) );
  NOR2_X1 U5313 ( .A1(n5734), .A2(n4478), .ZN(n5237) );
  INV_X1 U5314 ( .A(n5512), .ZN(n4660) );
  NAND2_X1 U5315 ( .A1(n5190), .A2(n5653), .ZN(n5189) );
  NAND2_X1 U5316 ( .A1(n5192), .A2(n5194), .ZN(n5190) );
  NAND2_X1 U5317 ( .A1(n9058), .A2(n9059), .ZN(n9083) );
  INV_X1 U5318 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4946) );
  AOI21_X1 U5319 ( .B1(n9151), .B2(n9150), .A(n9149), .ZN(n9167) );
  NAND2_X1 U5320 ( .A1(n8641), .A2(n5986), .ZN(n8409) );
  NAND2_X1 U5321 ( .A1(n5929), .A2(n5928), .ZN(n5941) );
  INV_X1 U5322 ( .A(n9313), .ZN(n7092) );
  NAND2_X1 U5323 ( .A1(n5020), .A2(n4445), .ZN(n4592) );
  INV_X1 U5324 ( .A(n6818), .ZN(n5107) );
  AND2_X1 U5325 ( .A1(n5090), .A2(n4569), .ZN(n4568) );
  NAND2_X1 U5326 ( .A1(n4570), .A2(n6937), .ZN(n4569) );
  INV_X1 U5327 ( .A(n6219), .ZN(n4570) );
  AOI21_X1 U5328 ( .B1(n8178), .B2(n5255), .A(n4480), .ZN(n5254) );
  INV_X1 U5329 ( .A(n6437), .ZN(n5255) );
  INV_X1 U5330 ( .A(n6434), .ZN(n4561) );
  NOR2_X1 U5331 ( .A1(n6433), .A2(n5131), .ZN(n5130) );
  INV_X1 U5332 ( .A(n4712), .ZN(n5131) );
  OAI211_X1 U5333 ( .C1(n5036), .C2(n6363), .A(n4609), .B(n6366), .ZN(n6830)
         );
  OR2_X1 U5334 ( .A1(n10118), .A2(n9593), .ZN(n6965) );
  NAND2_X1 U5335 ( .A1(n6465), .A2(n6464), .ZN(n6475) );
  AND2_X1 U5336 ( .A1(n4904), .A2(n5734), .ZN(n4896) );
  NAND2_X1 U5337 ( .A1(n5617), .A2(SI_12_), .ZN(n4605) );
  OR2_X1 U5338 ( .A1(n6235), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U5339 ( .A1(n4639), .A2(n5002), .ZN(n5000) );
  OAI21_X1 U5340 ( .B1(n5487), .B2(n4580), .A(n4579), .ZN(n5469) );
  NAND2_X1 U5341 ( .A1(n4414), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4579) );
  OAI211_X1 U5342 ( .C1(n5331), .C2(n4640), .A(n4638), .B(n4637), .ZN(n5335)
         );
  NAND2_X1 U5343 ( .A1(n4639), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4638) );
  XNOR2_X1 U5344 ( .A(n8837), .B(n5948), .ZN(n6013) );
  NAND2_X1 U5345 ( .A1(n7819), .A2(n4648), .ZN(n4646) );
  INV_X1 U5346 ( .A(n9034), .ZN(n7947) );
  AND2_X1 U5347 ( .A1(n5199), .A2(n8698), .ZN(n5198) );
  NAND2_X1 U5348 ( .A1(n4453), .A2(n5881), .ZN(n5199) );
  AND2_X1 U5349 ( .A1(n9009), .A2(n9010), .ZN(n5108) );
  NOR2_X1 U5350 ( .A1(n9005), .A2(n9006), .ZN(n5109) );
  NAND2_X1 U5351 ( .A1(n4671), .A2(n8985), .ZN(n8987) );
  INV_X2 U5352 ( .A(n5421), .ZN(n7135) );
  INV_X1 U5354 ( .A(n8401), .ZN(n5987) );
  NAND2_X2 U5355 ( .A1(n5373), .A2(n9540), .ZN(n8401) );
  INV_X1 U5356 ( .A(n5101), .ZN(n5100) );
  OAI22_X1 U5357 ( .A1(n8401), .A2(n5371), .B1(n5423), .B2(n7223), .ZN(n5101)
         );
  NAND2_X1 U5358 ( .A1(n5180), .A2(n5181), .ZN(n5179) );
  INV_X1 U5359 ( .A(n7468), .ZN(n5180) );
  NOR2_X1 U5360 ( .A1(n9161), .A2(n9193), .ZN(n5154) );
  AOI21_X1 U5361 ( .B1(n4866), .B2(n4867), .A(n8808), .ZN(n4865) );
  AND2_X1 U5362 ( .A1(n4870), .A2(n8980), .ZN(n4866) );
  INV_X1 U5363 ( .A(n5062), .ZN(n5061) );
  NAND2_X1 U5364 ( .A1(n7078), .A2(n7077), .ZN(n5063) );
  NAND2_X1 U5365 ( .A1(n8308), .A2(n5064), .ZN(n5060) );
  NOR2_X1 U5366 ( .A1(n7080), .A2(n5065), .ZN(n5064) );
  INV_X1 U5367 ( .A(n7077), .ZN(n5065) );
  AND2_X1 U5368 ( .A1(n7290), .A2(n7176), .ZN(n5656) );
  NAND2_X1 U5369 ( .A1(n7176), .A2(n4414), .ZN(n5720) );
  AND2_X1 U5370 ( .A1(n9249), .A2(n9382), .ZN(n5070) );
  AND2_X2 U5371 ( .A1(n4644), .A2(n4466), .ZN(n9247) );
  INV_X1 U5372 ( .A(n8843), .ZN(n5115) );
  INV_X1 U5373 ( .A(n9302), .ZN(n5058) );
  INV_X1 U5374 ( .A(n9290), .ZN(n5056) );
  OR2_X1 U5375 ( .A1(n7088), .A2(n9333), .ZN(n9298) );
  NAND2_X1 U5376 ( .A1(n7119), .A2(n8948), .ZN(n9351) );
  NAND2_X1 U5377 ( .A1(n4859), .A2(n4856), .ZN(n4855) );
  AND2_X1 U5378 ( .A1(n6005), .A2(n7314), .ZN(n7151) );
  AOI22_X1 U5379 ( .A1(n6703), .A2(n6511), .B1(n4750), .B2(n6543), .ZN(n6516)
         );
  NAND2_X1 U5380 ( .A1(n8270), .A2(n8628), .ZN(n4807) );
  NAND2_X1 U5381 ( .A1(n7291), .A2(n4414), .ZN(n4914) );
  NAND2_X1 U5382 ( .A1(n4448), .A2(n5024), .ZN(n5023) );
  INV_X1 U5383 ( .A(n5026), .ZN(n5024) );
  AND2_X1 U5384 ( .A1(n7024), .A2(n4966), .ZN(n7322) );
  OR2_X1 U5385 ( .A1(n6763), .A2(n7326), .ZN(n6757) );
  INV_X1 U5386 ( .A(n8438), .ZN(n7024) );
  AOI21_X1 U5387 ( .B1(n7009), .B2(n7008), .A(n7007), .ZN(n7012) );
  NAND2_X1 U5388 ( .A1(n4541), .A2(n7004), .ZN(n7009) );
  OR2_X1 U5389 ( .A1(n7003), .A2(n7010), .ZN(n7004) );
  NAND2_X2 U5390 ( .A1(n8270), .A2(n7023), .ZN(n7044) );
  NAND3_X1 U5391 ( .A1(n7171), .A2(P1_STATE_REG_SCAN_IN), .A3(n7323), .ZN(
        n7326) );
  OR2_X1 U5392 ( .A1(n6485), .A2(n7394), .ZN(n6145) );
  NOR2_X2 U5393 ( .A1(n6490), .A2(n6491), .ZN(n9883) );
  INV_X1 U5394 ( .A(n6772), .ZN(n4823) );
  NAND2_X1 U5395 ( .A1(n6332), .A2(n4525), .ZN(n6354) );
  NAND2_X1 U5396 ( .A1(n8179), .A2(n6806), .ZN(n4577) );
  INV_X1 U5397 ( .A(n4412), .ZN(n6277) );
  INV_X1 U5398 ( .A(n7324), .ZN(n6276) );
  OR2_X1 U5399 ( .A1(n8468), .A2(n8566), .ZN(n10344) );
  NAND2_X1 U5400 ( .A1(n5132), .A2(n5130), .ZN(n6171) );
  NAND2_X1 U5401 ( .A1(n7961), .A2(n6133), .ZN(n10397) );
  OR2_X1 U5402 ( .A1(n6364), .A2(n7293), .ZN(n6138) );
  NAND2_X1 U5403 ( .A1(n6795), .A2(n6830), .ZN(n6897) );
  NAND2_X1 U5404 ( .A1(n4710), .A2(n4708), .ZN(n4711) );
  NOR2_X1 U5405 ( .A1(n6450), .A2(n4709), .ZN(n4708) );
  AND2_X2 U5406 ( .A1(n6027), .A2(n6026), .ZN(n6374) );
  AOI21_X1 U5407 ( .B1(n4416), .B2(n4920), .A(n4491), .ZN(n4916) );
  AOI21_X1 U5408 ( .B1(n5241), .B2(n5242), .A(n5634), .ZN(n5240) );
  NAND2_X1 U5409 ( .A1(n5474), .A2(n5434), .ZN(n5033) );
  NAND2_X1 U5410 ( .A1(n4649), .A2(n5201), .ZN(n8259) );
  NAND2_X1 U5411 ( .A1(n8054), .A2(n5202), .ZN(n4649) );
  NAND2_X1 U5412 ( .A1(n5984), .A2(n10533), .ZN(n8784) );
  XNOR2_X1 U5413 ( .A(n9198), .B(n9197), .ZN(n9206) );
  INV_X1 U5414 ( .A(n5009), .ZN(n5005) );
  NAND2_X1 U5415 ( .A1(n6909), .A2(n8288), .ZN(n4531) );
  INV_X1 U5416 ( .A(n6974), .ZN(n4979) );
  NAND2_X1 U5417 ( .A1(n4978), .A2(n4975), .ZN(n4974) );
  AOI21_X1 U5418 ( .B1(n4538), .B2(n4976), .A(n6951), .ZN(n4975) );
  AND2_X1 U5419 ( .A1(n6976), .A2(n9980), .ZN(n4981) );
  INV_X1 U5420 ( .A(n4666), .ZN(n4665) );
  NAND2_X1 U5421 ( .A1(n5075), .A2(n9664), .ZN(n6966) );
  INV_X1 U5422 ( .A(n7129), .ZN(n8984) );
  INV_X1 U5423 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U5424 ( .A1(n6999), .A2(n4604), .ZN(n4603) );
  NAND2_X1 U5425 ( .A1(n6996), .A2(n7022), .ZN(n4604) );
  INV_X1 U5426 ( .A(n6991), .ZN(n6999) );
  OAI211_X1 U5427 ( .C1(n6990), .C2(n6996), .A(n6795), .B(n6989), .ZN(n6991)
         );
  OR2_X1 U5428 ( .A1(n6975), .A2(n6328), .ZN(n6824) );
  AND2_X1 U5429 ( .A1(n6250), .A2(n9737), .ZN(n6949) );
  INV_X1 U5430 ( .A(n4929), .ZN(n4927) );
  AND3_X1 U5431 ( .A1(n5237), .A2(n4451), .A3(n4922), .ZN(n4921) );
  NAND2_X1 U5432 ( .A1(n5696), .A2(n5695), .ZN(n4922) );
  NOR2_X1 U5433 ( .A1(n4443), .A2(n4919), .ZN(n4904) );
  OAI21_X1 U5434 ( .B1(n5196), .B2(n5194), .A(n8744), .ZN(n5193) );
  INV_X1 U5435 ( .A(n5607), .ZN(n4653) );
  NAND2_X1 U5436 ( .A1(n7512), .A2(n7181), .ZN(n4613) );
  NAND2_X1 U5437 ( .A1(n7515), .A2(n7201), .ZN(n7202) );
  INV_X1 U5438 ( .A(n7203), .ZN(n4714) );
  AND2_X1 U5439 ( .A1(n4625), .A2(n7468), .ZN(n7363) );
  INV_X1 U5440 ( .A(n7923), .ZN(n4729) );
  AND2_X1 U5441 ( .A1(n4762), .A2(n4761), .ZN(n7189) );
  NAND2_X1 U5442 ( .A1(n8111), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4761) );
  INV_X1 U5443 ( .A(n5172), .ZN(n5171) );
  NAND2_X1 U5444 ( .A1(n5168), .A2(n4526), .ZN(n4622) );
  OAI21_X1 U5445 ( .B1(n9085), .B2(n4726), .A(n4724), .ZN(n9128) );
  INV_X1 U5446 ( .A(n4725), .ZN(n4724) );
  OAI21_X1 U5447 ( .B1(n9086), .B2(n4726), .A(n9104), .ZN(n4725) );
  INV_X1 U5448 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5311) );
  INV_X1 U5449 ( .A(n7131), .ZN(n4879) );
  NOR2_X1 U5450 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n4831) );
  INV_X1 U5451 ( .A(n4444), .ZN(n5867) );
  NOR2_X1 U5452 ( .A1(n5772), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n4844) );
  INV_X1 U5453 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5680) );
  INV_X1 U5454 ( .A(n5682), .ZN(n5681) );
  INV_X1 U5455 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7595) );
  NOR2_X1 U5456 ( .A1(n5599), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U5457 ( .A1(n8611), .A2(n8309), .ZN(n8855) );
  INV_X1 U5458 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5521) );
  INV_X1 U5459 ( .A(n5523), .ZN(n5522) );
  AND2_X1 U5460 ( .A1(n4834), .A2(n4833), .ZN(n5458) );
  INV_X1 U5461 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n4834) );
  NAND2_X1 U5462 ( .A1(n7109), .A2(n7060), .ZN(n8890) );
  NAND2_X1 U5463 ( .A1(n4730), .A2(n10538), .ZN(n7107) );
  NAND2_X1 U5464 ( .A1(n7107), .A2(n5072), .ZN(n4641) );
  NAND2_X1 U5465 ( .A1(n8868), .A2(n4404), .ZN(n5072) );
  NOR2_X1 U5466 ( .A1(n8984), .A2(n5230), .ZN(n5229) );
  INV_X1 U5467 ( .A(n7097), .ZN(n5230) );
  NAND2_X1 U5468 ( .A1(n9481), .A2(n9269), .ZN(n5059) );
  AND2_X1 U5469 ( .A1(n5057), .A2(n5059), .ZN(n5052) );
  NAND2_X1 U5470 ( .A1(n9355), .A2(n8949), .ZN(n4860) );
  INV_X1 U5471 ( .A(n7117), .ZN(n5097) );
  NOR2_X1 U5472 ( .A1(n8938), .A2(n5094), .ZN(n5093) );
  INV_X1 U5473 ( .A(n7116), .ZN(n5094) );
  AND2_X1 U5474 ( .A1(n8165), .A2(n8168), .ZN(n8170) );
  NOR2_X1 U5475 ( .A1(n5186), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n5184) );
  AND2_X1 U5476 ( .A1(n5553), .A2(n5552), .ZN(n5556) );
  INV_X1 U5477 ( .A(n8325), .ZN(n5016) );
  NOR2_X1 U5478 ( .A1(n7016), .A2(n7015), .ZN(n7019) );
  NOR2_X1 U5479 ( .A1(n7014), .A2(n7022), .ZN(n7015) );
  NAND2_X1 U5480 ( .A1(n4494), .A2(n4430), .ZN(n4973) );
  NAND2_X1 U5481 ( .A1(n9872), .A2(n8438), .ZN(n7022) );
  NOR2_X1 U5482 ( .A1(n5124), .A2(n9925), .ZN(n5118) );
  NAND2_X1 U5483 ( .A1(n4988), .A2(n6329), .ZN(n4816) );
  NAND2_X1 U5484 ( .A1(n4610), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6315) );
  INV_X1 U5485 ( .A(n6306), .ZN(n4610) );
  NAND2_X1 U5486 ( .A1(n10504), .A2(n9741), .ZN(n6943) );
  INV_X1 U5487 ( .A(n10310), .ZN(n4576) );
  INV_X1 U5488 ( .A(n5130), .ZN(n4558) );
  NAND2_X1 U5489 ( .A1(n9904), .A2(n6829), .ZN(n5125) );
  NOR2_X1 U5490 ( .A1(n4461), .A2(n5259), .ZN(n5258) );
  INV_X1 U5491 ( .A(n6441), .ZN(n5259) );
  INV_X1 U5492 ( .A(n6949), .ZN(n6940) );
  OR2_X1 U5493 ( .A1(n10143), .A2(n9739), .ZN(n6439) );
  OR2_X1 U5494 ( .A1(n9726), .A2(n8512), .ZN(n5277) );
  NAND2_X1 U5495 ( .A1(n6465), .A2(n6466), .ZN(n6846) );
  AOI21_X1 U5496 ( .B1(n5888), .B2(n4910), .A(n4909), .ZN(n4908) );
  INV_X1 U5497 ( .A(n5888), .ZN(n4911) );
  INV_X1 U5498 ( .A(n5882), .ZN(n4910) );
  AND2_X1 U5499 ( .A1(n5920), .A2(n5904), .ZN(n5919) );
  INV_X1 U5500 ( .A(n5768), .ZN(n5222) );
  NAND2_X1 U5501 ( .A1(n5733), .A2(n5719), .ZN(n5734) );
  NAND2_X1 U5502 ( .A1(n4903), .A2(n4899), .ZN(n4898) );
  NAND2_X1 U5503 ( .A1(n4900), .A2(n4902), .ZN(n4899) );
  INV_X1 U5504 ( .A(n4904), .ZN(n4900) );
  AOI21_X1 U5505 ( .B1(n4904), .B2(n5696), .A(n4478), .ZN(n4903) );
  INV_X1 U5506 ( .A(n5734), .ZN(n4902) );
  AOI21_X1 U5507 ( .B1(n4887), .B2(n4885), .A(n4884), .ZN(n4883) );
  INV_X1 U5508 ( .A(n5592), .ZN(n4884) );
  INV_X1 U5509 ( .A(n5578), .ZN(n4885) );
  NAND2_X1 U5510 ( .A1(n5620), .A2(n4605), .ZN(n5621) );
  AOI21_X1 U5511 ( .B1(n5513), .B2(n5512), .A(n5511), .ZN(n5514) );
  NAND2_X1 U5512 ( .A1(n5746), .A2(n8671), .ZN(n5772) );
  INV_X1 U5513 ( .A(n5763), .ZN(n5746) );
  XNOR2_X1 U5514 ( .A(n10560), .B(n5536), .ZN(n5454) );
  XNOR2_X1 U5515 ( .A(n4730), .B(n4411), .ZN(n5380) );
  AND2_X1 U5516 ( .A1(n5975), .A2(n7969), .ZN(n6005) );
  NAND2_X1 U5517 ( .A1(n4422), .A2(n4455), .ZN(n5309) );
  AND2_X1 U5518 ( .A1(n8409), .A2(n5992), .ZN(n9025) );
  AND4_X1 U5519 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .ZN(n8708)
         );
  INV_X1 U5520 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5142) );
  XNOR2_X1 U5521 ( .A(n7520), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n7514) );
  OR2_X1 U5522 ( .A1(n4613), .A2(n7418), .ZN(n7182) );
  XNOR2_X1 U5523 ( .A(n7202), .B(n7234), .ZN(n7421) );
  NAND2_X1 U5524 ( .A1(n4717), .A2(n4716), .ZN(n7435) );
  OR2_X1 U5525 ( .A1(n7431), .A2(n7205), .ZN(n4717) );
  NAND2_X1 U5526 ( .A1(n4624), .A2(n4625), .ZN(n5176) );
  AND2_X1 U5527 ( .A1(n4436), .A2(n7468), .ZN(n4624) );
  NAND2_X1 U5528 ( .A1(n7363), .A2(n4421), .ZN(n5178) );
  OAI21_X1 U5529 ( .B1(n7208), .B2(n4723), .A(n4721), .ZN(n7210) );
  INV_X1 U5530 ( .A(n4722), .ZN(n4721) );
  OAI21_X1 U5531 ( .B1(n7207), .B2(n4723), .A(n7209), .ZN(n4722) );
  NOR2_X1 U5532 ( .A1(n7189), .A2(n7264), .ZN(n7194) );
  NAND2_X1 U5533 ( .A1(n5169), .A2(n5174), .ZN(n5168) );
  INV_X1 U5534 ( .A(n9067), .ZN(n5169) );
  XNOR2_X1 U5535 ( .A(n9128), .B(n9115), .ZN(n9127) );
  AND2_X1 U5536 ( .A1(n5947), .A2(n5946), .ZN(n8836) );
  INV_X1 U5537 ( .A(n10544), .ZN(n4872) );
  INV_X1 U5538 ( .A(n9234), .ZN(n9235) );
  NAND2_X1 U5539 ( .A1(n9237), .A2(n9380), .ZN(n9239) );
  INV_X1 U5540 ( .A(n9345), .ZN(n9318) );
  OR2_X1 U5541 ( .A1(n5761), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5763) );
  CLKBUF_X1 U5542 ( .A(n9351), .Z(n9352) );
  OR2_X1 U5543 ( .A1(n5661), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5682) );
  AND4_X1 U5544 ( .A1(n5650), .A2(n5649), .A3(n5648), .A4(n5647), .ZN(n8925)
         );
  AND2_X1 U5545 ( .A1(n7113), .A2(n8854), .ZN(n4849) );
  NAND2_X1 U5546 ( .A1(n5522), .A2(n5521), .ZN(n5537) );
  NAND2_X1 U5547 ( .A1(n5458), .A2(n5457), .ZN(n5495) );
  NAND2_X1 U5548 ( .A1(n8803), .A2(n8802), .ZN(n9010) );
  NAND2_X1 U5549 ( .A1(n4643), .A2(n5227), .ZN(n9226) );
  NAND2_X1 U5550 ( .A1(n9247), .A2(n5229), .ZN(n4643) );
  XNOR2_X1 U5551 ( .A(n8837), .B(n8836), .ZN(n9225) );
  INV_X1 U5552 ( .A(n8970), .ZN(n4868) );
  INV_X1 U5553 ( .A(n5114), .ZN(n4869) );
  NAND2_X1 U5554 ( .A1(n9273), .A2(n8974), .ZN(n4645) );
  AND2_X1 U5555 ( .A1(n8809), .A2(n8971), .ZN(n9267) );
  INV_X1 U5556 ( .A(n4859), .ZN(n4857) );
  INV_X1 U5557 ( .A(n9027), .ZN(n9358) );
  INV_X1 U5558 ( .A(n9380), .ZN(n10539) );
  AOI21_X1 U5559 ( .B1(n5045), .B2(n8928), .A(n4459), .ZN(n5044) );
  AND2_X1 U5560 ( .A1(n8751), .A2(n8691), .ZN(n8928) );
  NAND2_X1 U5561 ( .A1(n5060), .A2(n4432), .ZN(n4642) );
  OR2_X1 U5562 ( .A1(n5605), .A2(n7080), .ZN(n8823) );
  AND2_X1 U5563 ( .A1(n8991), .A2(n7142), .ZN(n9380) );
  OR2_X1 U5564 ( .A1(n8999), .A2(n5993), .ZN(n7974) );
  NAND2_X1 U5565 ( .A1(n4414), .A2(n5332), .ZN(n4782) );
  NAND2_X2 U5566 ( .A1(n7104), .A2(n7105), .ZN(n10541) );
  OR2_X1 U5567 ( .A1(n5325), .A2(n4757), .ZN(n5323) );
  INV_X1 U5568 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5315) );
  NOR2_X1 U5569 ( .A1(n5285), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5203) );
  INV_X1 U5570 ( .A(n7335), .ZN(n7552) );
  INV_X1 U5571 ( .A(n6556), .ZN(n5022) );
  NAND2_X1 U5572 ( .A1(n6638), .A2(n4431), .ZN(n4596) );
  NOR2_X1 U5573 ( .A1(n4787), .A2(n4786), .ZN(n4785) );
  INV_X1 U5574 ( .A(n9615), .ZN(n4787) );
  INV_X1 U5575 ( .A(n6655), .ZN(n4786) );
  XNOR2_X1 U5576 ( .A(n6551), .B(n6549), .ZN(n9571) );
  NOR2_X1 U5577 ( .A1(n4591), .A2(n6706), .ZN(n4590) );
  INV_X1 U5578 ( .A(n6699), .ZN(n4591) );
  NAND2_X1 U5579 ( .A1(n7012), .A2(n4963), .ZN(n4608) );
  AND4_X1 U5580 ( .A1(n6054), .A2(n6053), .A3(n6052), .A4(n6051), .ZN(n8511)
         );
  AND4_X1 U5581 ( .A1(n6216), .A2(n6215), .A3(n6214), .A4(n6213), .ZN(n8496)
         );
  AND4_X1 U5582 ( .A1(n6100), .A2(n6099), .A3(n6098), .A4(n6097), .ZN(n8464)
         );
  AND4_X1 U5583 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n8293)
         );
  NAND2_X1 U5584 ( .A1(n10219), .A2(n4426), .ZN(n5245) );
  NAND2_X1 U5585 ( .A1(n6114), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4533) );
  NAND2_X1 U5586 ( .A1(n4796), .A2(n4795), .ZN(n9755) );
  NAND2_X1 U5587 ( .A1(n7392), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4795) );
  OR2_X1 U5588 ( .A1(n7392), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4796) );
  OR2_X1 U5589 ( .A1(n7489), .A2(n7490), .ZN(n7878) );
  OR2_X1 U5590 ( .A1(n8042), .A2(n8043), .ZN(n9845) );
  AND2_X1 U5591 ( .A1(n10267), .A2(n9861), .ZN(n10279) );
  NAND2_X1 U5592 ( .A1(n9900), .A2(n9891), .ZN(n6490) );
  AOI21_X1 U5593 ( .B1(n9536), .B2(n5036), .A(n6477), .ZN(n8618) );
  NAND2_X1 U5594 ( .A1(n4819), .A2(n4820), .ZN(n9938) );
  OR2_X1 U5595 ( .A1(n4989), .A2(n4566), .ZN(n4819) );
  INV_X1 U5596 ( .A(n4992), .ZN(n4567) );
  INV_X1 U5597 ( .A(n6831), .ZN(n4993) );
  INV_X1 U5598 ( .A(n6962), .ZN(n4994) );
  INV_X1 U5599 ( .A(n4995), .ZN(n4991) );
  NAND2_X1 U5600 ( .A1(n4989), .A2(n4987), .ZN(n9969) );
  INV_X1 U5601 ( .A(n6952), .ZN(n5103) );
  NAND2_X1 U5602 ( .A1(n10133), .A2(n6661), .ZN(n6818) );
  NAND2_X1 U5603 ( .A1(n10045), .A2(n10046), .ZN(n5104) );
  AOI21_X1 U5604 ( .B1(n5090), .B2(n6797), .A(n5088), .ZN(n5087) );
  NAND2_X1 U5605 ( .A1(n4571), .A2(n4568), .ZN(n4572) );
  INV_X1 U5606 ( .A(n6796), .ZN(n5088) );
  NAND2_X1 U5607 ( .A1(n10061), .A2(n10063), .ZN(n10062) );
  NAND2_X1 U5608 ( .A1(n10313), .A2(n6219), .ZN(n8519) );
  NOR2_X1 U5609 ( .A1(n10318), .A2(n8411), .ZN(n5268) );
  INV_X1 U5610 ( .A(n5267), .ZN(n5266) );
  OAI21_X1 U5611 ( .B1(n10318), .B2(n5271), .A(n5270), .ZN(n5267) );
  NAND2_X1 U5612 ( .A1(n10499), .A2(n8417), .ZN(n5270) );
  NAND2_X1 U5613 ( .A1(n6943), .A2(n6937), .ZN(n8522) );
  NAND2_X1 U5614 ( .A1(n4698), .A2(n4696), .ZN(n10355) );
  NAND2_X1 U5615 ( .A1(n4697), .A2(n8566), .ZN(n4696) );
  INV_X1 U5616 ( .A(n10370), .ZN(n4686) );
  OR2_X1 U5617 ( .A1(n6364), .A2(n7297), .ZN(n6175) );
  NAND2_X1 U5618 ( .A1(n10397), .A2(n6800), .ZN(n4529) );
  AND2_X1 U5619 ( .A1(n5129), .A2(n6430), .ZN(n5133) );
  NAND2_X1 U5620 ( .A1(n4556), .A2(n4555), .ZN(n7961) );
  INV_X1 U5621 ( .A(n7958), .ZN(n4556) );
  OR2_X1 U5622 ( .A1(n6515), .A2(n7455), .ZN(n6759) );
  NOR2_X1 U5623 ( .A1(n9914), .A2(n9897), .ZN(n9915) );
  AND2_X1 U5624 ( .A1(n6448), .A2(n6447), .ZN(n5253) );
  NAND2_X1 U5625 ( .A1(n10113), .A2(n9664), .ZN(n4781) );
  AND2_X2 U5626 ( .A1(n4705), .A2(n4464), .ZN(n10017) );
  NAND2_X1 U5627 ( .A1(n10030), .A2(n6442), .ZN(n4705) );
  NAND2_X1 U5628 ( .A1(n6440), .A2(n6439), .ZN(n10059) );
  NAND2_X1 U5629 ( .A1(n8297), .A2(n10492), .ZN(n10507) );
  INV_X1 U5630 ( .A(n7326), .ZN(n10209) );
  INV_X1 U5631 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U5632 ( .A1(n5889), .A2(n5888), .ZN(n5901) );
  NAND2_X1 U5633 ( .A1(n4601), .A2(n4599), .ZN(n6404) );
  AND2_X1 U5634 ( .A1(n6377), .A2(n4600), .ZN(n4599) );
  INV_X1 U5635 ( .A(n6379), .ZN(n4601) );
  INV_X1 U5636 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6405) );
  INV_X1 U5637 ( .A(n5806), .ZN(n4932) );
  NOR2_X1 U5638 ( .A1(n5276), .A2(n4930), .ZN(n4929) );
  AND2_X1 U5639 ( .A1(n5855), .A2(n5837), .ZN(n5844) );
  NAND2_X1 U5640 ( .A1(n6375), .A2(n6402), .ZN(n6412) );
  INV_X2 U5641 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6377) );
  INV_X1 U5642 ( .A(n7023), .ZN(n7042) );
  NAND2_X1 U5643 ( .A1(n4682), .A2(n5235), .ZN(n4681) );
  NAND2_X1 U5644 ( .A1(n4680), .A2(n4678), .ZN(n4682) );
  AOI21_X1 U5645 ( .B1(n5696), .B2(n5695), .A(n4679), .ZN(n4678) );
  OAI21_X1 U5646 ( .B1(n5697), .B2(n5696), .A(n5695), .ZN(n5715) );
  OR2_X1 U5647 ( .A1(n6203), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6223) );
  INV_X1 U5648 ( .A(n5242), .ZN(n5239) );
  INV_X1 U5649 ( .A(n4905), .ZN(n5241) );
  OAI21_X1 U5650 ( .B1(n5242), .B2(n5244), .A(n4605), .ZN(n4905) );
  NOR2_X1 U5651 ( .A1(n6068), .A2(n6036), .ZN(n6189) );
  INV_X1 U5652 ( .A(n5436), .ZN(n5437) );
  INV_X1 U5653 ( .A(SI_5_), .ZN(n4658) );
  INV_X1 U5654 ( .A(n5469), .ZN(n4659) );
  OR2_X1 U5655 ( .A1(n6149), .A2(n6044), .ZN(n6160) );
  INV_X1 U5656 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6023) );
  INV_X1 U5657 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5074) );
  INV_X1 U5658 ( .A(SI_0_), .ZN(n5073) );
  NAND2_X1 U5659 ( .A1(n5334), .A2(n5333), .ZN(n5401) );
  INV_X1 U5660 ( .A(n5335), .ZN(n5334) );
  NAND2_X1 U5661 ( .A1(n5335), .A2(SI_1_), .ZN(n5403) );
  NAND2_X1 U5662 ( .A1(n8056), .A2(n5202), .ZN(n8202) );
  INV_X1 U5663 ( .A(n7817), .ZN(n5430) );
  AND2_X1 U5664 ( .A1(n5778), .A2(n5777), .ZN(n9333) );
  AND2_X1 U5665 ( .A1(n6786), .A2(n4630), .ZN(n4629) );
  OR2_X1 U5666 ( .A1(n5917), .A2(n4631), .ZN(n4630) );
  INV_X1 U5667 ( .A(n5918), .ZN(n4631) );
  AND2_X1 U5668 ( .A1(n7814), .A2(n5400), .ZN(n5379) );
  AND3_X1 U5669 ( .A1(n5710), .A2(n5709), .A3(n5708), .ZN(n9359) );
  XNOR2_X1 U5670 ( .A(n5454), .B(n7110), .ZN(n7945) );
  OR2_X1 U5671 ( .A1(n6009), .A2(n5996), .ZN(n8795) );
  AND2_X1 U5672 ( .A1(n5854), .A2(n5853), .ZN(n9288) );
  NAND2_X1 U5673 ( .A1(n4647), .A2(n7987), .ZN(n5483) );
  INV_X1 U5674 ( .A(n8786), .ZN(n8790) );
  INV_X1 U5675 ( .A(n9025), .ZN(n9227) );
  INV_X1 U5676 ( .A(n8836), .ZN(n9237) );
  NAND2_X1 U5677 ( .A1(n9233), .A2(n5986), .ZN(n4843) );
  NAND2_X1 U5678 ( .A1(n5827), .A2(n5826), .ZN(n9304) );
  AND2_X1 U5679 ( .A1(n5802), .A2(n5801), .ZN(n9317) );
  INV_X1 U5680 ( .A(n8708), .ZN(n9370) );
  XNOR2_X1 U5681 ( .A(n7935), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7923) );
  OR2_X1 U5682 ( .A1(n9165), .A2(n5147), .ZN(n5146) );
  INV_X1 U5683 ( .A(n5150), .ZN(n5147) );
  NAND2_X1 U5684 ( .A1(n5152), .A2(n5150), .ZN(n5145) );
  NOR2_X1 U5685 ( .A1(n9217), .A2(n4528), .ZN(n5148) );
  INV_X1 U5686 ( .A(n5153), .ZN(n5149) );
  NAND2_X1 U5687 ( .A1(n9211), .A2(n9212), .ZN(n4806) );
  NOR2_X1 U5688 ( .A1(n9187), .A2(n9427), .ZN(n4808) );
  OR2_X1 U5689 ( .A1(n7505), .A2(n9199), .ZN(n9213) );
  NAND2_X1 U5690 ( .A1(n5770), .A2(n5624), .ZN(n5217) );
  AND2_X1 U5691 ( .A1(n8024), .A2(n7314), .ZN(n5983) );
  NAND2_X1 U5692 ( .A1(n5224), .A2(n4415), .ZN(n4862) );
  INV_X1 U5693 ( .A(n8926), .ZN(n8751) );
  NAND2_X1 U5694 ( .A1(n10578), .A2(n9443), .ZN(n9424) );
  AND2_X1 U5695 ( .A1(n7174), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7317) );
  INV_X1 U5696 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5296) );
  INV_X1 U5697 ( .A(n8631), .ZN(n4794) );
  INV_X1 U5698 ( .A(n8632), .ZN(n4793) );
  NAND2_X1 U5699 ( .A1(n10083), .A2(n9693), .ZN(n4789) );
  AND2_X1 U5700 ( .A1(n4458), .A2(n5023), .ZN(n4598) );
  NAND2_X1 U5701 ( .A1(n4914), .A2(n4912), .ZN(n6124) );
  NAND2_X1 U5702 ( .A1(n7831), .A2(n6118), .ZN(n5086) );
  NAND2_X1 U5703 ( .A1(n5471), .A2(n5032), .ZN(n6165) );
  AND2_X1 U5704 ( .A1(n4409), .A2(n5037), .ZN(n5032) );
  OAI21_X1 U5705 ( .B1(n7527), .B2(n6364), .A(n6039), .ZN(n8590) );
  NOR2_X1 U5706 ( .A1(n9699), .A2(n9698), .ZN(n4733) );
  INV_X1 U5707 ( .A(n9697), .ZN(n4732) );
  NAND2_X1 U5708 ( .A1(n10087), .A2(n9693), .ZN(n4767) );
  NAND2_X1 U5709 ( .A1(n6771), .A2(n6770), .ZN(n9719) );
  NOR2_X2 U5710 ( .A1(n6757), .A2(n6754), .ZN(n9716) );
  NAND2_X1 U5711 ( .A1(n6769), .A2(n8456), .ZN(n9721) );
  AND4_X1 U5712 ( .A1(n6170), .A2(n6169), .A3(n6168), .A4(n6167), .ZN(n9750)
         );
  OR2_X1 U5713 ( .A1(n7385), .A2(n7386), .ZN(n7487) );
  OR2_X1 U5714 ( .A1(n7881), .A2(n7882), .ZN(n8040) );
  AOI21_X1 U5715 ( .B1(n9867), .B2(n10293), .A(n4739), .ZN(n9874) );
  AND2_X1 U5716 ( .A1(n9869), .A2(n10284), .ZN(n4739) );
  CLKBUF_X1 U5717 ( .A(n6513), .Z(n9872) );
  OAI21_X1 U5718 ( .B1(n10308), .B2(n9876), .A(n9875), .ZN(n4772) );
  NAND2_X1 U5719 ( .A1(n6487), .A2(n6486), .ZN(n6488) );
  INV_X1 U5720 ( .A(n6341), .ZN(n6342) );
  INV_X1 U5721 ( .A(n10382), .ZN(n10401) );
  NAND2_X1 U5722 ( .A1(n8438), .A2(n8628), .ZN(n7455) );
  NAND2_X1 U5723 ( .A1(n4824), .A2(n4424), .ZN(n4821) );
  AND2_X1 U5724 ( .A1(n9904), .A2(n9905), .ZN(n4578) );
  XNOR2_X1 U5725 ( .A(n6454), .B(n6897), .ZN(n10158) );
  INV_X1 U5726 ( .A(n9908), .ZN(n5010) );
  NAND3_X1 U5727 ( .A1(n4962), .A2(n6918), .A3(n4961), .ZN(n6928) );
  NAND2_X1 U5728 ( .A1(n4531), .A2(n4530), .ZN(n4961) );
  NOR2_X1 U5729 ( .A1(n8917), .A2(n8999), .ZN(n4936) );
  NOR2_X1 U5730 ( .A1(n8502), .A2(n6942), .ZN(n4977) );
  NOR2_X1 U5731 ( .A1(n6949), .A2(n4427), .ZN(n4976) );
  OAI21_X1 U5732 ( .B1(n4677), .B2(n4956), .A(n8959), .ZN(n4676) );
  NOR2_X1 U5733 ( .A1(n4981), .A2(n6328), .ZN(n4980) );
  OR2_X1 U5734 ( .A1(n6959), .A2(n4983), .ZN(n4982) );
  INV_X1 U5735 ( .A(n5713), .ZN(n5714) );
  INV_X1 U5736 ( .A(n5195), .ZN(n5194) );
  AOI21_X1 U5737 ( .B1(n4669), .B2(n4668), .A(n9280), .ZN(n8968) );
  INV_X1 U5738 ( .A(n9087), .ZN(n4726) );
  AND2_X1 U5739 ( .A1(n6351), .A2(n6987), .ZN(n6839) );
  INV_X1 U5740 ( .A(n6996), .ZN(n7001) );
  INV_X1 U5741 ( .A(n6187), .ZN(n6887) );
  INV_X1 U5742 ( .A(n5078), .ZN(n5077) );
  INV_X1 U5743 ( .A(n5083), .ZN(n5082) );
  INV_X1 U5744 ( .A(n5900), .ZN(n4909) );
  OAI21_X1 U5745 ( .B1(n5487), .B2(P1_DATAO_REG_17__SCAN_IN), .A(n4784), .ZN(
        n5717) );
  NAND2_X1 U5746 ( .A1(n5487), .A2(n8129), .ZN(n4784) );
  OAI21_X1 U5747 ( .B1(n5487), .B2(P1_DATAO_REG_9__SCAN_IN), .A(n4792), .ZN(
        n5575) );
  NAND2_X1 U5748 ( .A1(n5487), .A2(n7787), .ZN(n4792) );
  OAI21_X1 U5749 ( .B1(n5487), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n5038), .ZN(
        n5385) );
  NAND2_X1 U5750 ( .A1(n4414), .A2(n5039), .ZN(n5038) );
  INV_X1 U5751 ( .A(n7972), .ZN(n5974) );
  NAND2_X1 U5752 ( .A1(n4755), .A2(n4753), .ZN(n4671) );
  NAND2_X1 U5753 ( .A1(n7363), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7362) );
  NAND2_X1 U5754 ( .A1(n4626), .A2(n4800), .ZN(n4625) );
  INV_X1 U5755 ( .A(n7185), .ZN(n4626) );
  INV_X1 U5756 ( .A(n7467), .ZN(n4723) );
  NOR2_X1 U5757 ( .A1(n7924), .A2(n4623), .ZN(n7188) );
  NOR2_X1 U5758 ( .A1(n7935), .A2(n8212), .ZN(n4623) );
  NAND2_X1 U5759 ( .A1(n5174), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5172) );
  OR2_X1 U5760 ( .A1(n5941), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5985) );
  AND2_X1 U5761 ( .A1(n4867), .A2(n8980), .ZN(n4863) );
  INV_X1 U5762 ( .A(n8819), .ZN(n7113) );
  NAND2_X1 U5763 ( .A1(n4635), .A2(n7058), .ZN(n4634) );
  INV_X1 U5764 ( .A(n7058), .ZN(n4636) );
  INV_X1 U5765 ( .A(n7057), .ZN(n7056) );
  NAND2_X1 U5766 ( .A1(n10536), .A2(n10535), .ZN(n10534) );
  OR2_X1 U5767 ( .A1(n8999), .A2(n6000), .ZN(n7159) );
  INV_X1 U5768 ( .A(n8949), .ZN(n4856) );
  AND2_X1 U5769 ( .A1(n8994), .A2(n9198), .ZN(n6000) );
  NAND2_X1 U5770 ( .A1(n4429), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4757) );
  INV_X1 U5771 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U5772 ( .A1(n5204), .A2(n4627), .ZN(n5657) );
  NOR2_X1 U5773 ( .A1(n5285), .A2(n5205), .ZN(n5204) );
  NAND2_X1 U5774 ( .A1(n5206), .A2(n7626), .ZN(n5205) );
  INV_X1 U5775 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5187) );
  AND2_X1 U5776 ( .A1(n5556), .A2(n5555), .ZN(n5595) );
  NOR2_X1 U5777 ( .A1(n6058), .A2(n6040), .ZN(n4799) );
  AND2_X1 U5778 ( .A1(n6534), .A2(n7912), .ZN(n4582) );
  NOR2_X1 U5779 ( .A1(n6723), .A2(n5031), .ZN(n5030) );
  INV_X1 U5780 ( .A(n9633), .ZN(n5031) );
  INV_X1 U5781 ( .A(SI_15_), .ZN(n7672) );
  INV_X1 U5782 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8671) );
  INV_X1 U5783 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4685) );
  NOR2_X1 U5784 ( .A1(n4993), .A2(n4994), .ZN(n4992) );
  OAI21_X1 U5785 ( .B1(n8509), .B2(n6797), .A(n8598), .ZN(n5091) );
  AND2_X1 U5786 ( .A1(n6239), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6246) );
  NOR2_X1 U5787 ( .A1(n6187), .A2(n8289), .ZN(n6806) );
  NAND2_X1 U5788 ( .A1(n5126), .A2(n9925), .ZN(n5119) );
  INV_X1 U5789 ( .A(n5246), .ZN(n4709) );
  NAND2_X1 U5790 ( .A1(n10036), .A2(n5076), .ZN(n10008) );
  NAND2_X1 U5791 ( .A1(n8524), .A2(n5081), .ZN(n10068) );
  NAND2_X1 U5792 ( .A1(n7552), .A2(n7953), .ZN(n7958) );
  AND2_X1 U5793 ( .A1(n6466), .A2(n5925), .ZN(n5936) );
  AND2_X1 U5794 ( .A1(n5900), .A2(n5887), .ZN(n5888) );
  AOI21_X1 U5795 ( .B1(n4927), .B2(n4928), .A(n4926), .ZN(n4925) );
  INV_X1 U5796 ( .A(n5855), .ZN(n4926) );
  NAND2_X1 U5797 ( .A1(n6374), .A2(n6373), .ZN(n6379) );
  NOR2_X1 U5798 ( .A1(n6372), .A2(n6371), .ZN(n6373) );
  INV_X1 U5799 ( .A(SI_21_), .ZN(n7675) );
  INV_X1 U5800 ( .A(n4921), .ZN(n4920) );
  NAND2_X1 U5801 ( .A1(n5234), .A2(n4451), .ZN(n5233) );
  NAND2_X1 U5802 ( .A1(n4921), .A2(n4919), .ZN(n4918) );
  NAND2_X1 U5803 ( .A1(n5235), .A2(n5753), .ZN(n5234) );
  AOI21_X1 U5804 ( .B1(n5237), .B2(n4443), .A(n5236), .ZN(n5235) );
  INV_X1 U5805 ( .A(n5733), .ZN(n5236) );
  INV_X1 U5806 ( .A(n5237), .ZN(n4679) );
  NAND2_X1 U5807 ( .A1(n5697), .A2(n5695), .ZN(n4680) );
  INV_X1 U5808 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U5809 ( .A1(n4656), .A2(n5654), .ZN(n5671) );
  OAI21_X1 U5810 ( .B1(n4414), .B2(n4810), .A(n4809), .ZN(n5580) );
  NAND2_X1 U5811 ( .A1(n5487), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n4809) );
  INV_X1 U5812 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5329) );
  OR2_X1 U5813 ( .A1(n5189), .A2(n5192), .ZN(n4651) );
  NOR2_X1 U5814 ( .A1(n5189), .A2(n4653), .ZN(n4652) );
  NAND2_X1 U5815 ( .A1(n8686), .A2(n9028), .ZN(n5195) );
  XNOR2_X1 U5816 ( .A(n5400), .B(n4774), .ZN(n5397) );
  AND2_X1 U5817 ( .A1(n4836), .A2(n4673), .ZN(n4672) );
  AND2_X1 U5818 ( .A1(n8409), .A2(n8408), .ZN(n9219) );
  OR2_X1 U5819 ( .A1(n7349), .A2(n7179), .ZN(n7350) );
  NAND2_X1 U5820 ( .A1(n4615), .A2(n4467), .ZN(n7197) );
  NAND2_X1 U5821 ( .A1(n7183), .A2(n7436), .ZN(n7440) );
  OAI21_X1 U5822 ( .B1(n7204), .B2(n4715), .A(n4713), .ZN(n7206) );
  AOI21_X1 U5823 ( .B1(n7435), .B2(n4714), .A(n4473), .ZN(n4713) );
  INV_X1 U5824 ( .A(n7435), .ZN(n4715) );
  NAND2_X1 U5825 ( .A1(n5178), .A2(n5179), .ZN(n7471) );
  INV_X1 U5826 ( .A(n7463), .ZN(n4744) );
  AOI21_X1 U5827 ( .B1(n7927), .B2(n7925), .A(n7926), .ZN(n7924) );
  OAI21_X1 U5828 ( .B1(n7212), .B2(n4729), .A(n4727), .ZN(n7214) );
  INV_X1 U5829 ( .A(n4728), .ZN(n4727) );
  OAI21_X1 U5830 ( .B1(n7211), .B2(n4729), .A(n7213), .ZN(n4728) );
  AOI21_X1 U5831 ( .B1(n7218), .B2(n4719), .A(n4718), .ZN(n7220) );
  OR2_X1 U5832 ( .A1(n7264), .A2(n8380), .ZN(n4719) );
  AND2_X1 U5833 ( .A1(n7264), .A2(n8380), .ZN(n4718) );
  NAND2_X1 U5834 ( .A1(n7220), .A2(n7219), .ZN(n9058) );
  OAI21_X1 U5835 ( .B1(n5161), .B2(n5164), .A(n5160), .ZN(n9040) );
  NAND2_X1 U5836 ( .A1(n5157), .A2(n7193), .ZN(n5161) );
  NAND2_X1 U5837 ( .A1(n9040), .A2(n9084), .ZN(n9067) );
  OR2_X1 U5838 ( .A1(n9042), .A2(n5172), .ZN(n5170) );
  NAND2_X1 U5839 ( .A1(n4622), .A2(n5173), .ZN(n4620) );
  NAND2_X1 U5840 ( .A1(n4619), .A2(n4524), .ZN(n4618) );
  NAND2_X1 U5841 ( .A1(n9130), .A2(n9129), .ZN(n9151) );
  NOR2_X1 U5842 ( .A1(n9161), .A2(n5165), .ZN(n9145) );
  XNOR2_X1 U5843 ( .A(n9167), .B(n9176), .ZN(n9169) );
  AND2_X1 U5844 ( .A1(n5153), .A2(n5151), .ZN(n5150) );
  NAND2_X1 U5845 ( .A1(n9163), .A2(n9192), .ZN(n5153) );
  AND2_X1 U5846 ( .A1(n8409), .A2(n7141), .ZN(n8839) );
  AND2_X1 U5847 ( .A1(n4877), .A2(n7102), .ZN(n4875) );
  NAND2_X1 U5848 ( .A1(n9231), .A2(n4428), .ZN(n4873) );
  INV_X1 U5849 ( .A(n5985), .ZN(n8641) );
  AOI21_X1 U5850 ( .B1(n5227), .B2(n5226), .A(n4482), .ZN(n5225) );
  INV_X1 U5851 ( .A(n5229), .ZN(n5226) );
  INV_X1 U5852 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U5853 ( .A1(n4844), .A2(n5795), .ZN(n5848) );
  INV_X1 U5854 ( .A(n4844), .ZN(n5796) );
  INV_X1 U5855 ( .A(n5216), .ZN(n5215) );
  AND2_X1 U5856 ( .A1(n4439), .A2(n4840), .ZN(n4839) );
  INV_X1 U5857 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n4840) );
  NAND2_X1 U5858 ( .A1(n5681), .A2(n4439), .ZN(n5725) );
  NAND2_X1 U5859 ( .A1(n5681), .A2(n5680), .ZN(n5704) );
  NAND2_X1 U5860 ( .A1(n5643), .A2(n5642), .ZN(n5661) );
  INV_X1 U5861 ( .A(n5644), .ZN(n5643) );
  NAND2_X1 U5862 ( .A1(n4842), .A2(n7595), .ZN(n5644) );
  INV_X1 U5863 ( .A(n4842), .ZN(n5608) );
  AND2_X1 U5864 ( .A1(n4423), .A2(n7763), .ZN(n4837) );
  OR2_X1 U5865 ( .A1(n5569), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U5866 ( .A1(n5522), .A2(n4423), .ZN(n5560) );
  AND2_X1 U5867 ( .A1(n4835), .A2(n5457), .ZN(n4832) );
  INV_X1 U5868 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4835) );
  OAI211_X1 U5869 ( .C1(n5636), .C2(n7298), .A(n5447), .B(n4489), .ZN(n8138)
         );
  NAND2_X1 U5870 ( .A1(n10534), .A2(n7058), .ZN(n8075) );
  NAND2_X1 U5871 ( .A1(n7134), .A2(n7974), .ZN(n10544) );
  NAND2_X1 U5872 ( .A1(n4641), .A2(n7053), .ZN(n7899) );
  NAND2_X1 U5873 ( .A1(n7896), .A2(n8867), .ZN(n7897) );
  AOI21_X1 U5874 ( .B1(n8593), .B2(n5624), .A(n4518), .ZN(n7095) );
  INV_X1 U5875 ( .A(n5111), .ZN(n4870) );
  INV_X1 U5876 ( .A(n5059), .ZN(n5050) );
  OR2_X1 U5877 ( .A1(n9313), .A2(n9330), .ZN(n9332) );
  AND2_X1 U5878 ( .A1(n8849), .A2(n9311), .ZN(n9330) );
  NAND2_X1 U5879 ( .A1(n4654), .A2(n7085), .ZN(n9344) );
  OR2_X1 U5880 ( .A1(n9352), .A2(n9355), .ZN(n4858) );
  INV_X1 U5881 ( .A(n9363), .ZN(n9431) );
  AND2_X1 U5882 ( .A1(n5096), .A2(n8936), .ZN(n5095) );
  NAND2_X1 U5883 ( .A1(n8827), .A2(n5097), .ZN(n5096) );
  NOR2_X1 U5884 ( .A1(n8911), .A2(n5136), .ZN(n5135) );
  INV_X1 U5885 ( .A(n8912), .ZN(n5136) );
  INV_X1 U5886 ( .A(n10562), .ZN(n10567) );
  INV_X1 U5887 ( .A(n8138), .ZN(n10560) );
  NAND2_X1 U5888 ( .A1(n4414), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U5889 ( .A1(n5310), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5966) );
  INV_X1 U5890 ( .A(n5140), .ZN(n5139) );
  INV_X1 U5891 ( .A(n5186), .ZN(n5185) );
  AND2_X1 U5892 ( .A1(n5441), .A2(n5440), .ZN(n5445) );
  OAI21_X1 U5893 ( .B1(n4720), .B2(n9528), .A(P2_IR_REG_2__SCAN_IN), .ZN(n4616) );
  AND2_X1 U5894 ( .A1(n4799), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6239) );
  INV_X1 U5895 ( .A(n4799), .ZN(n6228) );
  NAND2_X1 U5896 ( .A1(n6638), .A2(n6637), .ZN(n9550) );
  NOR2_X1 U5897 ( .A1(n6123), .A2(n4913), .ZN(n4912) );
  NOR2_X1 U5898 ( .A1(n5487), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4913) );
  NOR2_X1 U5899 ( .A1(n5027), .A2(n9602), .ZN(n5026) );
  INV_X1 U5900 ( .A(n5029), .ZN(n5027) );
  NAND2_X1 U5901 ( .A1(n9632), .A2(n6722), .ZN(n5029) );
  NAND2_X1 U5902 ( .A1(n9634), .A2(n5030), .ZN(n5028) );
  OR2_X1 U5903 ( .A1(n6315), .A2(n9564), .ZN(n6323) );
  NAND2_X1 U5904 ( .A1(n8248), .A2(n5018), .ZN(n5017) );
  INV_X1 U5905 ( .A(n9657), .ZN(n4594) );
  INV_X1 U5906 ( .A(n6600), .ZN(n5013) );
  NAND2_X1 U5907 ( .A1(n4589), .A2(n4588), .ZN(n4587) );
  INV_X1 U5908 ( .A(n6532), .ZN(n4588) );
  INV_X1 U5909 ( .A(n9703), .ZN(n9649) );
  AND2_X1 U5910 ( .A1(n7044), .A2(n7322), .ZN(n6765) );
  INV_X1 U5911 ( .A(n7019), .ZN(n4972) );
  AOI21_X1 U5912 ( .B1(n7019), .B2(n10079), .A(n7018), .ZN(n4970) );
  AND4_X1 U5913 ( .A1(n6350), .A2(n6349), .A3(n6348), .A4(n6347), .ZN(n9704)
         );
  AND4_X1 U5914 ( .A1(n6346), .A2(n6345), .A3(n6344), .A4(n6343), .ZN(n9603)
         );
  AND2_X1 U5915 ( .A1(n6312), .A2(n6311), .ZN(n9594) );
  AND4_X1 U5916 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6078), .ZN(n8553)
         );
  AND4_X1 U5917 ( .A1(n6185), .A2(n6184), .A3(n6183), .A4(n6182), .ZN(n8181)
         );
  NAND2_X1 U5918 ( .A1(n9755), .A2(n9754), .ZN(n9753) );
  NAND2_X1 U5919 ( .A1(n4741), .A2(n4740), .ZN(n7493) );
  INV_X1 U5920 ( .A(n7407), .ZN(n4740) );
  OR2_X1 U5921 ( .A1(n7495), .A2(n7496), .ZN(n7886) );
  NAND2_X1 U5922 ( .A1(n4743), .A2(n4742), .ZN(n8046) );
  INV_X1 U5923 ( .A(n7889), .ZN(n4742) );
  NAND2_X1 U5924 ( .A1(n4737), .A2(n4736), .ZN(n9855) );
  INV_X1 U5925 ( .A(n8049), .ZN(n4736) );
  INV_X1 U5926 ( .A(n8048), .ZN(n4737) );
  AND2_X1 U5927 ( .A1(n10240), .A2(n10239), .ZN(n10242) );
  AOI21_X1 U5928 ( .B1(n10243), .B2(P1_REG1_REG_14__SCAN_IN), .A(n10247), .ZN(
        n9847) );
  OR2_X1 U5929 ( .A1(n10271), .A2(n10270), .ZN(n10267) );
  AND2_X1 U5930 ( .A1(n10278), .A2(n9863), .ZN(n10296) );
  INV_X1 U5931 ( .A(n6830), .ZN(n5121) );
  NAND2_X1 U5932 ( .A1(n6332), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6341) );
  NAND2_X1 U5933 ( .A1(n5085), .A2(n5084), .ZN(n9918) );
  AND2_X1 U5934 ( .A1(n6288), .A2(n6287), .ZN(n6296) );
  NAND2_X1 U5935 ( .A1(n6296), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U5936 ( .A1(n5102), .A2(n6961), .ZN(n4562) );
  AOI21_X1 U5937 ( .B1(n5102), .B2(n5106), .A(n10018), .ZN(n4564) );
  NAND2_X1 U5938 ( .A1(n6246), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6256) );
  OR2_X1 U5939 ( .A1(n6256), .A2(n6255), .ZN(n6268) );
  NAND2_X1 U5940 ( .A1(n8510), .A2(n8509), .ZN(n5089) );
  NAND2_X1 U5941 ( .A1(n8519), .A2(n6937), .ZN(n8510) );
  OR2_X1 U5942 ( .A1(n7455), .A2(n7042), .ZN(n10407) );
  INV_X1 U5943 ( .A(n8522), .ZN(n5264) );
  OAI21_X1 U5944 ( .B1(n6218), .B2(n4576), .A(n10318), .ZN(n4574) );
  INV_X1 U5945 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U5946 ( .A1(n10325), .A2(n6218), .ZN(n10311) );
  NAND2_X1 U5947 ( .A1(n4612), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6196) );
  INV_X1 U5948 ( .A(n6085), .ZN(n4612) );
  NAND2_X1 U5949 ( .A1(n4611), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6208) );
  INV_X1 U5950 ( .A(n6196), .ZN(n4611) );
  AND2_X1 U5951 ( .A1(n10344), .A2(n10343), .ZN(n10370) );
  NOR2_X1 U5952 ( .A1(n4695), .A2(n4693), .ZN(n4691) );
  NOR2_X1 U5953 ( .A1(n4695), .A2(n4441), .ZN(n4689) );
  NAND2_X1 U5954 ( .A1(n6177), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6106) );
  NOR2_X1 U5955 ( .A1(n6106), .A2(n6094), .ZN(n6095) );
  AND3_X1 U5956 ( .A1(n6392), .A2(n10464), .A3(n4440), .ZN(n10373) );
  INV_X1 U5957 ( .A(n4560), .ZN(n4559) );
  NOR2_X1 U5958 ( .A1(n8093), .A2(n4561), .ZN(n4560) );
  AND3_X1 U5959 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6177) );
  AND2_X1 U5960 ( .A1(n6753), .A2(n10210), .ZN(n7449) );
  NOR2_X1 U5961 ( .A1(n7326), .A2(n6765), .ZN(n7534) );
  INV_X1 U5962 ( .A(n4985), .ZN(n4984) );
  OAI21_X1 U5963 ( .B1(n6338), .B2(n4986), .A(n9897), .ZN(n4985) );
  NAND2_X1 U5964 ( .A1(n9914), .A2(n6451), .ZN(n6503) );
  NAND2_X1 U5965 ( .A1(n6322), .A2(n6321), .ZN(n10097) );
  NOR2_X1 U5966 ( .A1(n9978), .A2(n6973), .ZN(n9977) );
  NAND2_X1 U5967 ( .A1(n8426), .A2(n5036), .ZN(n4606) );
  AND2_X1 U5968 ( .A1(n6965), .A2(n6832), .ZN(n10004) );
  NAND2_X1 U5969 ( .A1(n5257), .A2(n4702), .ZN(n4701) );
  NAND2_X1 U5970 ( .A1(n6440), .A2(n4474), .ZN(n4703) );
  INV_X1 U5971 ( .A(n5258), .ZN(n4702) );
  INV_X1 U5972 ( .A(n10063), .ZN(n5260) );
  INV_X1 U5973 ( .A(n10059), .ZN(n5261) );
  INV_X1 U5974 ( .A(n10507), .ZN(n10153) );
  AND2_X1 U5975 ( .A1(n6031), .A2(n4454), .ZN(n4537) );
  XNOR2_X1 U5976 ( .A(n5905), .B(n5919), .ZN(n8593) );
  NAND2_X1 U5977 ( .A1(n4903), .A2(n4902), .ZN(n4901) );
  OAI21_X1 U5978 ( .B1(n5734), .B2(n4903), .A(n4898), .ZN(n4897) );
  NAND2_X1 U5979 ( .A1(n5243), .A2(n5239), .ZN(n5629) );
  NAND2_X1 U5980 ( .A1(n5243), .A2(n4469), .ZN(n5622) );
  NAND2_X1 U5981 ( .A1(n5579), .A2(n5578), .ZN(n4889) );
  XNOR2_X1 U5982 ( .A(n5579), .B(n5578), .ZN(n7328) );
  INV_X1 U5983 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U5984 ( .A1(n5516), .A2(n5515), .ZN(n5532) );
  NAND2_X1 U5985 ( .A1(n4581), .A2(n5514), .ZN(n5516) );
  INV_X1 U5986 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U5987 ( .A1(n5474), .A2(n5034), .ZN(n5037) );
  NOR2_X1 U5988 ( .A1(n5438), .A2(n5035), .ZN(n5034) );
  INV_X1 U5989 ( .A(n5434), .ZN(n5035) );
  NAND2_X1 U5990 ( .A1(n4628), .A2(n5918), .ZN(n6787) );
  NAND2_X1 U5991 ( .A1(n8775), .A2(n5917), .ZN(n4628) );
  NAND2_X1 U5992 ( .A1(n8531), .A2(n5607), .ZN(n4765) );
  NAND2_X1 U5993 ( .A1(n5197), .A2(n5712), .ZN(n8715) );
  AND2_X1 U5994 ( .A1(n7819), .A2(n5433), .ZN(n7944) );
  NAND2_X1 U5995 ( .A1(n5545), .A2(n5544), .ZN(n8339) );
  NAND2_X1 U5996 ( .A1(n5191), .A2(n5195), .ZN(n8745) );
  NAND2_X1 U5997 ( .A1(n4765), .A2(n5196), .ZN(n5191) );
  OR2_X1 U5998 ( .A1(n5380), .A2(n4404), .ZN(n5381) );
  INV_X1 U5999 ( .A(n8782), .ZN(n8793) );
  NAND2_X1 U6000 ( .A1(n5502), .A2(n5501), .ZN(n8056) );
  INV_X1 U6001 ( .A(n8054), .ZN(n5502) );
  OR2_X1 U6002 ( .A1(n6009), .A2(n7142), .ZN(n8782) );
  AND2_X1 U6003 ( .A1(n5979), .A2(n5978), .ZN(n8786) );
  NAND2_X1 U6004 ( .A1(n6008), .A2(n6007), .ZN(n8797) );
  INV_X1 U6005 ( .A(n9288), .ZN(n9269) );
  NAND2_X1 U6006 ( .A1(n5752), .A2(n5751), .ZN(n9345) );
  OAI211_X1 U6007 ( .C1(n7138), .C2(n9427), .A(n5765), .B(n5764), .ZN(n9027)
         );
  INV_X1 U6008 ( .A(n8309), .ZN(n9031) );
  NAND4_X1 U6009 ( .A1(n5528), .A2(n5527), .A3(n5526), .A4(n5525), .ZN(n9033)
         );
  OR2_X1 U6010 ( .A1(n5423), .A2(n5461), .ZN(n5462) );
  OR2_X1 U6011 ( .A1(n5423), .A2(n7205), .ZN(n5450) );
  OR2_X1 U6012 ( .A1(n5421), .A2(n5422), .ZN(n5429) );
  OR2_X1 U6013 ( .A1(n5646), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5428) );
  INV_X1 U6014 ( .A(P2_U3893), .ZN(n9036) );
  XNOR2_X1 U6015 ( .A(n7226), .B(n7222), .ZN(n7346) );
  NAND2_X1 U6016 ( .A1(n7420), .A2(n5182), .ZN(n7423) );
  NAND2_X1 U6017 ( .A1(n7434), .A2(n7435), .ZN(n7433) );
  NAND2_X1 U6018 ( .A1(n7204), .A2(n7203), .ZN(n7434) );
  XNOR2_X1 U6019 ( .A(n7206), .B(n4800), .ZN(n7361) );
  NAND2_X1 U6020 ( .A1(n7208), .A2(n7207), .ZN(n7466) );
  NAND2_X1 U6021 ( .A1(n7466), .A2(n7467), .ZN(n7465) );
  AND3_X1 U6022 ( .A1(n5178), .A2(n4497), .A3(n5179), .ZN(n7186) );
  NAND2_X1 U6023 ( .A1(n7861), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7927) );
  XNOR2_X1 U6024 ( .A(n7214), .B(n8016), .ZN(n8007) );
  NAND2_X1 U6025 ( .A1(n5157), .A2(n5163), .ZN(n8229) );
  XNOR2_X1 U6026 ( .A(n7218), .B(n7264), .ZN(n8239) );
  NAND2_X1 U6027 ( .A1(n5159), .A2(n5158), .ZN(n9039) );
  AOI21_X1 U6028 ( .B1(n5156), .B2(n5163), .A(n5162), .ZN(n5158) );
  NAND2_X1 U6029 ( .A1(n5155), .A2(n5163), .ZN(n5159) );
  NAND2_X1 U6030 ( .A1(n5170), .A2(n5168), .ZN(n9093) );
  NAND2_X1 U6031 ( .A1(n9088), .A2(n9087), .ZN(n9103) );
  NAND2_X1 U6032 ( .A1(n9085), .A2(n9086), .ZN(n9088) );
  AND2_X1 U6033 ( .A1(n4465), .A2(n4617), .ZN(n9095) );
  OR2_X1 U6034 ( .A1(P2_U3150), .A2(n7281), .ZN(n9171) );
  NAND2_X1 U6035 ( .A1(n9239), .A2(n9238), .ZN(n9240) );
  AOI21_X1 U6036 ( .B1(n9303), .B2(n9302), .A(n4420), .ZN(n9286) );
  NAND2_X1 U6037 ( .A1(n5060), .A2(n5061), .ZN(n8391) );
  NAND2_X1 U6038 ( .A1(n4850), .A2(n8854), .ZN(n8276) );
  CLKBUF_X1 U6039 ( .A(n8138), .Z(n4764) );
  OR2_X1 U6040 ( .A1(n10565), .A2(n8024), .ZN(n10531) );
  INV_X1 U6041 ( .A(n9424), .ZN(n9438) );
  NAND2_X1 U6042 ( .A1(n9231), .A2(n7131), .ZN(n9224) );
  INV_X1 U6043 ( .A(n5069), .ZN(n4780) );
  AOI21_X1 U6044 ( .B1(n9227), .B2(n9380), .A(n5070), .ZN(n5069) );
  OAI21_X1 U6045 ( .B1(n9026), .B2(n10537), .A(n4812), .ZN(n4811) );
  NAND2_X1 U6046 ( .A1(n9249), .A2(n9380), .ZN(n4812) );
  NAND2_X1 U6047 ( .A1(n5113), .A2(n8971), .ZN(n9254) );
  NAND2_X1 U6048 ( .A1(n7127), .A2(n5114), .ZN(n5113) );
  NAND2_X1 U6049 ( .A1(n7127), .A2(n8843), .ZN(n9265) );
  NAND2_X1 U6050 ( .A1(n9303), .A2(n5057), .ZN(n5054) );
  NAND2_X1 U6051 ( .A1(n4853), .A2(n4854), .ZN(n9299) );
  OR2_X1 U6052 ( .A1(n9351), .A2(n4857), .ZN(n4853) );
  NAND2_X1 U6053 ( .A1(n8150), .A2(n5624), .ZN(n5759) );
  NAND2_X1 U6054 ( .A1(n5040), .A2(n5044), .ZN(n9379) );
  NAND2_X1 U6055 ( .A1(n8430), .A2(n5045), .ZN(n5040) );
  NAND2_X1 U6056 ( .A1(n8927), .A2(n5047), .ZN(n8543) );
  OR2_X1 U6057 ( .A1(n8430), .A2(n8928), .ZN(n5047) );
  NAND2_X1 U6058 ( .A1(n8428), .A2(n7116), .ZN(n5098) );
  OAI21_X1 U6059 ( .B1(n8308), .B2(n7078), .A(n7077), .ZN(n8319) );
  NAND2_X1 U6060 ( .A1(n7114), .A2(n8912), .ZN(n8318) );
  NAND2_X1 U6061 ( .A1(n7314), .A2(n7313), .ZN(n7319) );
  NAND2_X1 U6062 ( .A1(n5340), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5316) );
  INV_X1 U6063 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8579) );
  OR2_X1 U6064 ( .A1(n5325), .A2(n5324), .ZN(n5326) );
  INV_X1 U6065 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8493) );
  INV_X1 U6066 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8454) );
  INV_X1 U6067 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8441) );
  INV_X1 U6068 ( .A(n9020), .ZN(n8869) );
  INV_X1 U6069 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8336) );
  INV_X1 U6070 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8274) );
  INV_X1 U6071 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n8211) );
  INV_X1 U6072 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n8037) );
  INV_X1 U6073 ( .A(n7234), .ZN(n7418) );
  INV_X1 U6074 ( .A(n6768), .ZN(n7323) );
  NAND2_X1 U6075 ( .A1(n7308), .A2(n5036), .ZN(n4996) );
  NAND2_X1 U6076 ( .A1(n5020), .A2(n6691), .ZN(n9591) );
  NAND2_X1 U6077 ( .A1(n5028), .A2(n5029), .ZN(n9601) );
  NAND2_X1 U6078 ( .A1(n4597), .A2(n6659), .ZN(n9627) );
  NAND2_X1 U6079 ( .A1(n4596), .A2(n4785), .ZN(n4597) );
  AOI21_X1 U6080 ( .B1(n9634), .B2(n9633), .A(n9632), .ZN(n9636) );
  INV_X1 U6081 ( .A(n9716), .ZN(n9695) );
  NAND2_X1 U6082 ( .A1(n6564), .A2(n8154), .ZN(n8250) );
  NAND2_X1 U6083 ( .A1(n7041), .A2(n7040), .ZN(n7043) );
  NAND2_X1 U6084 ( .A1(n4545), .A2(n7027), .ZN(n4544) );
  INV_X1 U6085 ( .A(n7026), .ZN(n7027) );
  NAND2_X1 U6086 ( .A1(n4608), .A2(n4607), .ZN(n4545) );
  AOI21_X1 U6087 ( .B1(n9952), .B2(n6337), .A(n6327), .ZN(n9604) );
  INV_X1 U6088 ( .A(n9594), .ZN(n9733) );
  AND2_X1 U6089 ( .A1(n6294), .A2(n6293), .ZN(n9593) );
  NAND2_X1 U6090 ( .A1(n6869), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4534) );
  OR2_X1 U6091 ( .A1(n6485), .A2(n7829), .ZN(n6131) );
  NAND2_X1 U6092 ( .A1(n9813), .A2(n9814), .ZN(n9812) );
  NAND2_X1 U6093 ( .A1(n7487), .A2(n7486), .ZN(n7489) );
  NAND2_X1 U6094 ( .A1(n8040), .A2(n8039), .ZN(n8042) );
  AND2_X1 U6095 ( .A1(n10238), .A2(n10237), .ZN(n10247) );
  INV_X1 U6096 ( .A(n7013), .ZN(n10076) );
  INV_X1 U6097 ( .A(n6354), .ZN(n6356) );
  NAND2_X1 U6098 ( .A1(n4824), .A2(n4823), .ZN(n9894) );
  XNOR2_X1 U6099 ( .A(n9924), .B(n9925), .ZN(n4894) );
  NAND2_X1 U6100 ( .A1(n4551), .A2(n10399), .ZN(n4550) );
  NAND2_X1 U6101 ( .A1(n9939), .A2(n9938), .ZN(n4551) );
  NAND2_X1 U6102 ( .A1(n4710), .A2(n5246), .ZN(n9929) );
  INV_X1 U6103 ( .A(n9640), .ZN(n9952) );
  AOI21_X1 U6104 ( .B1(n4995), .B2(n4994), .A(n4993), .ZN(n4990) );
  NAND2_X1 U6105 ( .A1(n4563), .A2(n5102), .ZN(n10019) );
  NAND2_X1 U6106 ( .A1(n10045), .A2(n5105), .ZN(n4563) );
  NAND2_X1 U6107 ( .A1(n5104), .A2(n6818), .ZN(n10032) );
  INV_X1 U6108 ( .A(n6244), .ZN(n6245) );
  NAND2_X1 U6109 ( .A1(n5262), .A2(n5266), .ZN(n8517) );
  NAND2_X1 U6110 ( .A1(n8412), .A2(n5268), .ZN(n5262) );
  AOI21_X1 U6111 ( .B1(n8412), .B2(n8414), .A(n5269), .ZN(n10319) );
  OR2_X1 U6112 ( .A1(n10402), .A2(n9872), .ZN(n10411) );
  NAND2_X1 U6113 ( .A1(n5256), .A2(n6437), .ZN(n8177) );
  NAND2_X1 U6114 ( .A1(n6171), .A2(n6434), .ZN(n8088) );
  OAI21_X1 U6115 ( .B1(n10397), .B2(n6148), .A(n6800), .ZN(n8099) );
  INV_X1 U6116 ( .A(n10412), .ZN(n10394) );
  NAND2_X1 U6117 ( .A1(n10209), .A2(n6760), .ZN(n10382) );
  NAND2_X1 U6118 ( .A1(n7458), .A2(n10382), .ZN(n10324) );
  INV_X1 U6119 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n4826) );
  NAND2_X1 U6120 ( .A1(n10075), .A2(n4777), .ZN(n10151) );
  INV_X1 U6121 ( .A(n4778), .ZN(n4777) );
  OAI21_X1 U6122 ( .B1(n10076), .B2(n10503), .A(n10077), .ZN(n4778) );
  NAND2_X1 U6123 ( .A1(n4804), .A2(n6506), .ZN(n4683) );
  NAND2_X1 U6124 ( .A1(n4824), .A2(n4822), .ZN(n10154) );
  NOR2_X1 U6125 ( .A1(n10086), .A2(n4891), .ZN(n10164) );
  NAND2_X1 U6126 ( .A1(n4893), .A2(n4892), .ZN(n4891) );
  NAND2_X1 U6127 ( .A1(n10087), .A2(n10490), .ZN(n4892) );
  INV_X1 U6128 ( .A(n10085), .ZN(n4893) );
  OAI21_X1 U6129 ( .B1(n9917), .B2(n9925), .A(n9916), .ZN(n10167) );
  NAND2_X1 U6130 ( .A1(n5247), .A2(n5252), .ZN(n9943) );
  NAND2_X1 U6131 ( .A1(n9960), .A2(n5253), .ZN(n5247) );
  AND2_X1 U6132 ( .A1(n10209), .A2(n10208), .ZN(n10423) );
  INV_X1 U6133 ( .A(n6030), .ZN(n4552) );
  NOR2_X1 U6134 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(n6029), .ZN(n4553) );
  NAND2_X1 U6135 ( .A1(n6862), .A2(n6861), .ZN(n6866) );
  INV_X1 U6136 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10225) );
  INV_X1 U6137 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8582) );
  INV_X1 U6138 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8490) );
  INV_X1 U6139 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8458) );
  NAND2_X1 U6140 ( .A1(n4932), .A2(n4929), .ZN(n4924) );
  INV_X1 U6141 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8439) );
  OR2_X1 U6142 ( .A1(n6375), .A2(n6402), .ZN(n6376) );
  NAND2_X1 U6143 ( .A1(n5220), .A2(n5211), .ZN(n8335) );
  INV_X1 U6144 ( .A(n5212), .ZN(n5211) );
  INV_X1 U6145 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U6146 ( .A1(n5238), .A2(n4471), .ZN(n5635) );
  NAND2_X1 U6147 ( .A1(n5616), .A2(n5239), .ZN(n5238) );
  XNOR2_X1 U6148 ( .A(n6038), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9853) );
  AND2_X1 U6149 ( .A1(n6192), .A2(n6203), .ZN(n7884) );
  INV_X1 U6150 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U6151 ( .A1(n4657), .A2(n5509), .ZN(n5476) );
  NAND2_X1 U6152 ( .A1(n5471), .A2(n5037), .ZN(n7298) );
  XNOR2_X1 U6153 ( .A(n6163), .B(n6162), .ZN(n7856) );
  NAND2_X1 U6154 ( .A1(n6136), .A2(n6135), .ZN(n7839) );
  OAI22_X1 U6155 ( .A1(n6120), .A2(n4738), .B1(P1_IR_REG_2__SCAN_IN), .B2(
        P1_IR_REG_31__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U6156 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4738) );
  NAND2_X1 U6157 ( .A1(n6122), .A2(n6121), .ZN(n7392) );
  NAND2_X1 U6158 ( .A1(n5401), .A2(n5403), .ZN(n5337) );
  NAND2_X1 U6159 ( .A1(n5487), .A2(SI_0_), .ZN(n6132) );
  NAND2_X1 U6160 ( .A1(n6788), .A2(n5286), .ZN(n6017) );
  NAND2_X1 U6161 ( .A1(n7212), .A2(n7211), .ZN(n7922) );
  AOI21_X1 U6162 ( .B1(n9216), .B2(n9215), .A(n4806), .ZN(n4805) );
  OAI21_X1 U6163 ( .B1(n9454), .B2(n10550), .A(n5066), .ZN(P2_U3205) );
  INV_X1 U6164 ( .A(n5067), .ZN(n5066) );
  OAI21_X1 U6165 ( .B1(n9459), .B2(n9366), .A(n5068), .ZN(n5067) );
  AND2_X1 U6166 ( .A1(n9230), .A2(n4515), .ZN(n5068) );
  OR2_X1 U6167 ( .A1(n7170), .A2(n9424), .ZN(n5278) );
  NAND2_X1 U6168 ( .A1(n4862), .A2(n7169), .ZN(n4861) );
  OR2_X1 U6169 ( .A1(n7170), .A2(n9500), .ZN(n5275) );
  AND2_X1 U6170 ( .A1(n8638), .A2(n4789), .ZN(n4788) );
  AND2_X1 U6171 ( .A1(n9712), .A2(n4767), .ZN(n4766) );
  INV_X1 U6172 ( .A(n4772), .ZN(n4771) );
  OR2_X1 U6173 ( .A1(n9873), .A2(n8270), .ZN(n4773) );
  NAND2_X1 U6174 ( .A1(n4776), .A2(n4775), .ZN(P1_U3553) );
  NAND2_X1 U6175 ( .A1(n10526), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n4775) );
  NAND2_X1 U6176 ( .A1(n10151), .A2(n10528), .ZN(n4776) );
  NAND2_X1 U6177 ( .A1(n10526), .A2(n4826), .ZN(n4825) );
  NOR2_X1 U6178 ( .A1(n10528), .A2(n10084), .ZN(n5004) );
  NAND2_X1 U6179 ( .A1(n4760), .A2(n4758), .ZN(P1_U3545) );
  OR2_X1 U6180 ( .A1(n10528), .A2(n4759), .ZN(n4758) );
  INV_X1 U6181 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n4759) );
  AND2_X2 U6182 ( .A1(n7171), .A2(n6510), .ZN(n6543) );
  AND3_X1 U6183 ( .A1(n7147), .A2(n4425), .A3(n10578), .ZN(n4415) );
  CLKBUF_X3 U6184 ( .A(n5656), .Z(n5624) );
  AND2_X1 U6185 ( .A1(n5233), .A2(n4918), .ZN(n4416) );
  INV_X1 U6186 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U6187 ( .A1(n10147), .A2(n9740), .ZN(n4417) );
  OR2_X1 U6189 ( .A1(n7188), .A2(n8016), .ZN(n4418) );
  INV_X1 U6190 ( .A(n5695), .ZN(n4919) );
  INV_X1 U6191 ( .A(n6329), .ZN(n4566) );
  NOR2_X1 U6192 ( .A1(n5287), .A2(n4879), .ZN(n4419) );
  OAI21_X1 U6193 ( .B1(n9084), .B2(n9040), .A(n9067), .ZN(n9042) );
  INV_X1 U6194 ( .A(n9042), .ZN(n4619) );
  AND2_X1 U6195 ( .A1(n8685), .A2(n9317), .ZN(n4420) );
  AND2_X1 U6196 ( .A1(n5181), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4421) );
  INV_X1 U6197 ( .A(n5809), .ZN(n4930) );
  NAND2_X1 U6198 ( .A1(n4619), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9066) );
  AND4_X1 U6199 ( .A1(n5307), .A2(n5313), .A3(n5308), .A4(n5306), .ZN(n4422)
         );
  INV_X1 U6200 ( .A(n9273), .ZN(n9475) );
  AND2_X1 U6201 ( .A1(n5865), .A2(n5864), .ZN(n9273) );
  NAND2_X1 U6202 ( .A1(n5100), .A2(n5099), .ZN(n7529) );
  INV_X1 U6203 ( .A(n8411), .ZN(n8414) );
  AND2_X1 U6204 ( .A1(n10310), .A2(n6923), .ZN(n8411) );
  AND2_X1 U6205 ( .A1(n5521), .A2(n4838), .ZN(n4423) );
  AND2_X1 U6206 ( .A1(n4822), .A2(n10528), .ZN(n4424) );
  AND2_X1 U6207 ( .A1(n6049), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U6208 ( .A1(n6987), .A2(n9905), .ZN(n9925) );
  NAND2_X1 U6209 ( .A1(n6057), .A2(n6056), .ZN(n10317) );
  AOI21_X1 U6210 ( .B1(n10063), .B2(n5258), .A(n4484), .ZN(n5257) );
  AOI21_X2 U6211 ( .B1(n9533), .B2(n4410), .A(n4522), .ZN(n10079) );
  OR3_X1 U6212 ( .A1(n6946), .A2(n6945), .A3(n7010), .ZN(n4427) );
  NOR2_X1 U6213 ( .A1(n6352), .A2(n5127), .ZN(n5126) );
  INV_X1 U6214 ( .A(n5126), .ZN(n5122) );
  INV_X1 U6215 ( .A(n8468), .ZN(n4697) );
  INV_X1 U6216 ( .A(n5106), .ZN(n5105) );
  AND2_X1 U6217 ( .A1(n8988), .A2(n4419), .ZN(n4428) );
  INV_X1 U6218 ( .A(n8194), .ZN(n8901) );
  XOR2_X1 U6219 ( .A(n5317), .B(P2_IR_REG_24__SCAN_IN), .Z(n4429) );
  AND2_X1 U6220 ( .A1(n5283), .A2(n7011), .ZN(n4430) );
  AND2_X1 U6221 ( .A1(n4493), .A2(n6637), .ZN(n4431) );
  AND2_X1 U6222 ( .A1(n5061), .A2(n4483), .ZN(n4432) );
  NAND2_X1 U6223 ( .A1(n7095), .A2(n4907), .ZN(n8981) );
  AND3_X1 U6224 ( .A1(n5079), .A2(n4697), .A3(n10453), .ZN(n4433) );
  AND2_X1 U6225 ( .A1(n10343), .A2(n10341), .ZN(n4434) );
  AND2_X1 U6226 ( .A1(n6399), .A2(n6408), .ZN(n4435) );
  AND2_X1 U6227 ( .A1(n4421), .A2(n5177), .ZN(n4436) );
  INV_X1 U6228 ( .A(n4720), .ZN(n4615) );
  INV_X1 U6229 ( .A(n10113), .ZN(n5075) );
  NAND2_X1 U6230 ( .A1(n8524), .A2(n10504), .ZN(n4437) );
  AND2_X1 U6231 ( .A1(n6392), .A2(n10453), .ZN(n4438) );
  AOI21_X1 U6232 ( .B1(n8626), .B2(n5036), .A(n4514), .ZN(n9902) );
  INV_X1 U6233 ( .A(n9902), .ZN(n10083) );
  AND2_X1 U6234 ( .A1(n5680), .A2(n4841), .ZN(n4439) );
  AND2_X1 U6235 ( .A1(n5079), .A2(n10453), .ZN(n4440) );
  INV_X1 U6236 ( .A(n9026), .ZN(n9268) );
  AND2_X1 U6237 ( .A1(n5899), .A2(n5898), .ZN(n9026) );
  INV_X1 U6238 ( .A(n7193), .ZN(n5162) );
  INV_X1 U6239 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6044) );
  INV_X1 U6240 ( .A(n7296), .ZN(n4800) );
  NOR2_X1 U6241 ( .A1(n5046), .A2(n7082), .ZN(n5045) );
  AND2_X1 U6242 ( .A1(n8093), .A2(n8178), .ZN(n4441) );
  INV_X1 U6243 ( .A(n6529), .ZN(n6703) );
  INV_X1 U6244 ( .A(n6529), .ZN(n4734) );
  XNOR2_X1 U6245 ( .A(n6866), .B(n6865), .ZN(n9527) );
  AND4_X1 U6246 ( .A1(n5500), .A2(n5499), .A3(n5498), .A4(n5497), .ZN(n7990)
         );
  NAND2_X1 U6247 ( .A1(n5469), .A2(SI_5_), .ZN(n5509) );
  INV_X1 U6248 ( .A(n5720), .ZN(n5906) );
  AND2_X1 U6249 ( .A1(n4858), .A2(n8949), .ZN(n4442) );
  NOR2_X1 U6250 ( .A1(n5714), .A2(SI_16_), .ZN(n4443) );
  OR3_X1 U6251 ( .A1(n5848), .A2(P2_REG3_REG_22__SCAN_IN), .A3(
        P2_REG3_REG_23__SCAN_IN), .ZN(n4444) );
  AOI21_X1 U6252 ( .B1(n5111), .B2(n4869), .A(n4868), .ZN(n4867) );
  AND2_X1 U6253 ( .A1(n6696), .A2(n6691), .ZN(n4445) );
  AND2_X1 U6254 ( .A1(n5167), .A2(n5166), .ZN(n9161) );
  AND3_X1 U6255 ( .A1(n6987), .A2(n7022), .A3(n6992), .ZN(n4446) );
  OAI21_X1 U6256 ( .B1(n7321), .B2(n6364), .A(n6193), .ZN(n10335) );
  INV_X1 U6257 ( .A(n10335), .ZN(n10484) );
  NOR2_X1 U6258 ( .A1(n5155), .A2(n5156), .ZN(n7192) );
  AND3_X1 U6259 ( .A1(n8958), .A2(n8960), .A3(n8957), .ZN(n4447) );
  NOR2_X1 U6260 ( .A1(n9697), .A2(n9698), .ZN(n4448) );
  OR2_X1 U6261 ( .A1(n6379), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U6262 ( .A1(n10062), .A2(n6813), .ZN(n10045) );
  AND2_X1 U6263 ( .A1(n6129), .A2(n6130), .ZN(n4450) );
  INV_X1 U6264 ( .A(n6994), .ZN(n4986) );
  NAND2_X1 U6265 ( .A1(n5737), .A2(SI_18_), .ZN(n4451) );
  NAND2_X1 U6266 ( .A1(n5055), .A2(n5054), .ZN(n9279) );
  NAND2_X1 U6267 ( .A1(n5089), .A2(n6233), .ZN(n8597) );
  AND2_X1 U6268 ( .A1(n10083), .A2(n10490), .ZN(n4452) );
  NAND2_X1 U6269 ( .A1(n5877), .A2(n5876), .ZN(n4453) );
  AND4_X1 U6270 ( .A1(n7745), .A2(n6399), .A3(n6408), .A4(n6042), .ZN(n4454)
         );
  AND4_X1 U6271 ( .A1(n5305), .A2(n5304), .A3(n5303), .A4(n5675), .ZN(n4455)
         );
  INV_X1 U6272 ( .A(n8988), .ZN(n7102) );
  NAND2_X1 U6273 ( .A1(n10087), .A2(n9603), .ZN(n9905) );
  INV_X1 U6274 ( .A(n9905), .ZN(n5127) );
  OR2_X1 U6275 ( .A1(n10082), .A2(n4452), .ZN(n4456) );
  NAND2_X1 U6276 ( .A1(n6351), .A2(n6829), .ZN(n9904) );
  INV_X1 U6277 ( .A(n9904), .ZN(n5128) );
  AND2_X1 U6278 ( .A1(n5873), .A2(n5872), .ZN(n8974) );
  NAND2_X1 U6279 ( .A1(n6374), .A2(n6031), .ZN(n6398) );
  NAND2_X1 U6280 ( .A1(n10036), .A2(n5078), .ZN(n4457) );
  INV_X1 U6281 ( .A(n7017), .ZN(n7018) );
  NOR2_X1 U6282 ( .A1(n8632), .A2(n8631), .ZN(n4458) );
  AND2_X1 U6283 ( .A1(n8934), .A2(n9383), .ZN(n4459) );
  INV_X1 U6284 ( .A(n9249), .ZN(n7130) );
  NAND2_X1 U6285 ( .A1(n4843), .A2(n5935), .ZN(n9249) );
  INV_X1 U6286 ( .A(n6250), .ZN(n10138) );
  NAND2_X1 U6287 ( .A1(n6286), .A2(n6285), .ZN(n10118) );
  AND3_X1 U6288 ( .A1(n4949), .A2(n4950), .A3(n4948), .ZN(n4460) );
  INV_X1 U6289 ( .A(n5276), .ZN(n4931) );
  AND2_X1 U6290 ( .A1(n10133), .A2(n9736), .ZN(n4461) );
  OR2_X1 U6291 ( .A1(n9732), .A2(n10091), .ZN(n4462) );
  NAND2_X1 U6292 ( .A1(n5369), .A2(n5368), .ZN(n7054) );
  AND2_X1 U6293 ( .A1(n5281), .A2(n6434), .ZN(n4463) );
  NAND2_X1 U6294 ( .A1(n10128), .A2(n9735), .ZN(n4464) );
  XNOR2_X1 U6295 ( .A(n5736), .B(SI_18_), .ZN(n5753) );
  NAND2_X1 U6296 ( .A1(n4572), .A2(n5087), .ZN(n10061) );
  XNOR2_X1 U6297 ( .A(n5316), .B(n5315), .ZN(n8595) );
  AND2_X1 U6298 ( .A1(n5913), .A2(n5912), .ZN(n8701) );
  INV_X1 U6299 ( .A(n8701), .ZN(n4907) );
  NAND2_X1 U6300 ( .A1(n4595), .A2(n4594), .ZN(n4593) );
  AND2_X1 U6301 ( .A1(n9891), .A2(n9729), .ZN(n7000) );
  INV_X1 U6302 ( .A(n7000), .ZN(n6795) );
  AND2_X1 U6303 ( .A1(n4620), .A2(n4618), .ZN(n4465) );
  NAND2_X1 U6304 ( .A1(n9260), .A2(n9026), .ZN(n4466) );
  AND4_X1 U6305 ( .A1(n6089), .A2(n6088), .A3(n6087), .A4(n6086), .ZN(n8566)
         );
  NAND2_X1 U6306 ( .A1(n10083), .A2(n9704), .ZN(n6829) );
  AND2_X1 U6307 ( .A1(n5142), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4467) );
  AND2_X1 U6308 ( .A1(n6113), .A2(n5245), .ZN(n4468) );
  INV_X1 U6309 ( .A(n5019), .ZN(n5018) );
  NAND2_X1 U6310 ( .A1(n6576), .A2(n8324), .ZN(n5019) );
  OR2_X1 U6311 ( .A1(n5614), .A2(SI_11_), .ZN(n4469) );
  AND2_X1 U6312 ( .A1(n5566), .A2(n5544), .ZN(n4470) );
  INV_X1 U6313 ( .A(n5085), .ZN(n9930) );
  NAND2_X1 U6314 ( .A1(n6825), .A2(n6983), .ZN(n9944) );
  INV_X1 U6315 ( .A(n9944), .ZN(n5249) );
  AND2_X1 U6316 ( .A1(n5241), .A2(n5634), .ZN(n4471) );
  NOR2_X1 U6317 ( .A1(n9291), .A2(n9304), .ZN(n4472) );
  AND2_X1 U6318 ( .A1(n7431), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4473) );
  OR2_X1 U6319 ( .A1(n8094), .A2(n8181), .ZN(n6904) );
  AND2_X1 U6320 ( .A1(n5257), .A2(n6439), .ZN(n4474) );
  AND2_X1 U6321 ( .A1(n10102), .A2(n6449), .ZN(n4475) );
  AND2_X1 U6322 ( .A1(n4533), .A2(n4468), .ZN(n4476) );
  INV_X1 U6323 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7745) );
  INV_X1 U6324 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5343) );
  AND2_X1 U6325 ( .A1(n4416), .A2(n4915), .ZN(n4477) );
  NAND2_X1 U6326 ( .A1(n5583), .A2(n5592), .ZN(n4888) );
  AND2_X1 U6327 ( .A1(n5504), .A2(n8203), .ZN(n5202) );
  INV_X1 U6328 ( .A(n4699), .ZN(n4693) );
  NAND2_X1 U6329 ( .A1(n10464), .A2(n8464), .ZN(n4699) );
  INV_X1 U6330 ( .A(n5330), .ZN(n4639) );
  AND2_X1 U6331 ( .A1(n5714), .A2(SI_16_), .ZN(n4478) );
  NOR2_X1 U6332 ( .A1(n7017), .A2(n7022), .ZN(n4479) );
  NOR2_X1 U6333 ( .A1(n8256), .A2(n9748), .ZN(n4480) );
  AND2_X1 U6334 ( .A1(n8508), .A2(n6810), .ZN(n4481) );
  AND2_X1 U6335 ( .A1(n8837), .A2(n8836), .ZN(n4482) );
  OR2_X1 U6336 ( .A1(n8921), .A2(n9028), .ZN(n4483) );
  AND4_X1 U6337 ( .A1(n6145), .A2(n6146), .A3(n6144), .A4(n6147), .ZN(n8100)
         );
  INV_X1 U6338 ( .A(n8100), .ZN(n4735) );
  INV_X1 U6339 ( .A(n5124), .ZN(n5123) );
  NAND2_X1 U6340 ( .A1(n5125), .A2(n6795), .ZN(n5124) );
  INV_X1 U6341 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7389) );
  INV_X1 U6342 ( .A(n5228), .ZN(n5227) );
  OAI21_X1 U6343 ( .B1(n5231), .B2(n8984), .A(n7128), .ZN(n5228) );
  INV_X1 U6344 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5950) );
  INV_X1 U6345 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6043) );
  AOI21_X1 U6346 ( .B1(n5105), .B2(n5107), .A(n5103), .ZN(n5102) );
  AND2_X1 U6347 ( .A1(n10054), .A2(n6661), .ZN(n4484) );
  OR3_X1 U6348 ( .A1(n9009), .A2(n8992), .A3(n8991), .ZN(n4485) );
  OR2_X1 U6349 ( .A1(n6398), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4486) );
  NAND2_X1 U6350 ( .A1(n8964), .A2(n9298), .ZN(n4487) );
  AND2_X1 U6351 ( .A1(n5530), .A2(n8058), .ZN(n4488) );
  AND3_X1 U6352 ( .A1(n5086), .A2(n6124), .A3(n6125), .ZN(n10429) );
  INV_X1 U6353 ( .A(n10429), .ZN(n4750) );
  OR2_X1 U6354 ( .A1(n4746), .A2(n7431), .ZN(n4489) );
  INV_X1 U6355 ( .A(n5271), .ZN(n5269) );
  NAND2_X1 U6356 ( .A1(n6395), .A2(n8496), .ZN(n5271) );
  NAND2_X1 U6357 ( .A1(n10504), .A2(n8511), .ZN(n4490) );
  INV_X1 U6358 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n8131) );
  INV_X1 U6359 ( .A(n5015), .ZN(n5014) );
  OR2_X1 U6360 ( .A1(n6601), .A2(n5016), .ZN(n5015) );
  NAND2_X1 U6361 ( .A1(n5768), .A2(n5741), .ZN(n4491) );
  AND2_X1 U6362 ( .A1(n9326), .A2(n8946), .ZN(n4956) );
  NOR2_X1 U6363 ( .A1(n9955), .A2(n9604), .ZN(n4492) );
  NAND2_X1 U6364 ( .A1(n9610), .A2(n6644), .ZN(n4493) );
  AND2_X1 U6365 ( .A1(n6491), .A2(n6478), .ZN(n7006) );
  INV_X1 U6366 ( .A(n7096), .ZN(n5231) );
  NAND2_X1 U6367 ( .A1(n10076), .A2(n9878), .ZN(n4494) );
  NOR3_X1 U6368 ( .A1(n9248), .A2(n9255), .A3(n8834), .ZN(n4495) );
  NAND2_X1 U6369 ( .A1(n9007), .A2(n8806), .ZN(n8988) );
  NAND2_X1 U6370 ( .A1(n5840), .A2(n5839), .ZN(n4496) );
  INV_X1 U6371 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6399) );
  OR2_X1 U6372 ( .A1(n7472), .A2(n8067), .ZN(n4497) );
  INV_X1 U6373 ( .A(n8986), .ZN(n4836) );
  OAI21_X1 U6374 ( .B1(n7127), .B2(n4870), .A(n4867), .ZN(n9246) );
  OR2_X1 U6375 ( .A1(n5127), .A2(n6995), .ZN(n4498) );
  AND2_X1 U6376 ( .A1(n10103), .A2(n10104), .ZN(n4499) );
  OR2_X1 U6377 ( .A1(n8808), .A2(n8979), .ZN(n9248) );
  INV_X1 U6378 ( .A(n9248), .ZN(n4958) );
  AND3_X1 U6379 ( .A1(n5565), .A2(n5563), .A3(n5564), .ZN(n4500) );
  INV_X1 U6380 ( .A(n6942), .ZN(n6937) );
  AND2_X1 U6381 ( .A1(n8590), .A2(n8511), .ZN(n6942) );
  AND2_X1 U6382 ( .A1(n6393), .A2(n8553), .ZN(n4501) );
  AND2_X1 U6383 ( .A1(n5081), .A2(n6250), .ZN(n4502) );
  AND2_X1 U6384 ( .A1(n9463), .A2(n8701), .ZN(n8979) );
  AND2_X1 U6385 ( .A1(n6914), .A2(n7022), .ZN(n4503) );
  AND2_X1 U6386 ( .A1(n6914), .A2(n7010), .ZN(n4504) );
  OR2_X1 U6387 ( .A1(n7324), .A2(n7839), .ZN(n4505) );
  AND2_X1 U6388 ( .A1(n4448), .A2(n5030), .ZN(n4506) );
  AND2_X1 U6389 ( .A1(n8976), .A2(n8977), .ZN(n4507) );
  AND2_X1 U6390 ( .A1(n5732), .A2(n5712), .ZN(n4508) );
  AND2_X1 U6391 ( .A1(n5125), .A2(n5119), .ZN(n4509) );
  AND2_X1 U6392 ( .A1(n5265), .A2(n4417), .ZN(n4510) );
  NAND2_X1 U6393 ( .A1(n4496), .A2(n4931), .ZN(n4928) );
  AND2_X1 U6394 ( .A1(n4876), .A2(n4872), .ZN(n4511) );
  NOR2_X1 U6395 ( .A1(n4888), .A2(n5577), .ZN(n4887) );
  NAND2_X1 U6396 ( .A1(n7093), .A2(n9288), .ZN(n4512) );
  NAND2_X1 U6397 ( .A1(n4954), .A2(n4955), .ZN(n4677) );
  AND2_X1 U6398 ( .A1(n6738), .A2(n6737), .ZN(n8631) );
  INV_X1 U6399 ( .A(n5577), .ZN(n4890) );
  INV_X1 U6400 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5206) );
  INV_X1 U6401 ( .A(n4754), .ZN(n4753) );
  NAND2_X1 U6402 ( .A1(n8982), .A2(n9234), .ZN(n4754) );
  INV_X1 U6403 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4600) );
  INV_X1 U6404 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9528) );
  AND2_X1 U6405 ( .A1(n5139), .A2(n5343), .ZN(n4513) );
  INV_X2 U6406 ( .A(n10324), .ZN(n10402) );
  OR2_X1 U6407 ( .A1(n6783), .A2(n7448), .ZN(n10526) );
  NAND2_X1 U6408 ( .A1(n6340), .A2(n6339), .ZN(n10087) );
  INV_X1 U6409 ( .A(n10087), .ZN(n5084) );
  NAND2_X1 U6410 ( .A1(n5017), .A2(n8325), .ZN(n8459) );
  NAND2_X1 U6411 ( .A1(n8009), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8008) );
  AND2_X1 U6412 ( .A1(n5279), .A2(n10499), .ZN(n8524) );
  INV_X1 U6413 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4580) );
  NOR2_X1 U6414 ( .A1(n4412), .A2(n8627), .ZN(n4514) );
  AND3_X1 U6415 ( .A1(n5323), .A2(n5322), .A3(n5321), .ZN(n7312) );
  INV_X1 U6416 ( .A(n9940), .ZN(n4549) );
  INV_X1 U6417 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5002) );
  INV_X1 U6418 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5039) );
  INV_X1 U6419 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n4829) );
  AND2_X1 U6420 ( .A1(n8248), .A2(n6576), .ZN(n8326) );
  OR3_X2 U6421 ( .A1(n8489), .A2(n10227), .A3(n8580), .ZN(n7171) );
  NAND2_X1 U6422 ( .A1(n5098), .A2(n7117), .ZN(n8542) );
  NAND2_X1 U6423 ( .A1(n4694), .A2(n5254), .ZN(n8287) );
  OR2_X1 U6424 ( .A1(n9385), .A2(n9228), .ZN(n4515) );
  AND2_X1 U6425 ( .A1(n10057), .A2(n6441), .ZN(n4516) );
  OR2_X1 U6426 ( .A1(n10510), .A2(n10162), .ZN(n4517) );
  NAND2_X1 U6427 ( .A1(n10036), .A2(n10042), .ZN(n10022) );
  NAND2_X1 U6428 ( .A1(n8524), .A2(n5083), .ZN(n8504) );
  INV_X1 U6429 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4684) );
  AOI21_X1 U6430 ( .B1(n8008), .B2(n4418), .A(n8113), .ZN(n8112) );
  NAND2_X1 U6431 ( .A1(n5294), .A2(n5274), .ZN(n5754) );
  AND4_X1 U6432 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n8417)
         );
  NAND2_X1 U6433 ( .A1(n5261), .A2(n5260), .ZN(n10057) );
  NAND2_X1 U6434 ( .A1(n6392), .A2(n4440), .ZN(n5080) );
  AND2_X1 U6435 ( .A1(n5906), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n4518) );
  INV_X1 U6436 ( .A(n5157), .ZN(n5156) );
  OR2_X1 U6437 ( .A1(n7191), .A2(n8230), .ZN(n5157) );
  INV_X2 U6438 ( .A(n10573), .ZN(n10571) );
  NOR2_X1 U6439 ( .A1(n9038), .A2(n9037), .ZN(n4519) );
  AND2_X1 U6440 ( .A1(n4831), .A2(n4830), .ZN(n4520) );
  AND2_X1 U6441 ( .A1(n8056), .A2(n5504), .ZN(n4521) );
  INV_X1 U6442 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6227) );
  INV_X1 U6443 ( .A(n9385), .ZN(n10550) );
  OAI211_X1 U6444 ( .C1(n7324), .C2(n9790), .A(n6105), .B(n6104), .ZN(n8256)
         );
  INV_X1 U6445 ( .A(n8256), .ZN(n5079) );
  INV_X1 U6446 ( .A(n9725), .ZN(n9693) );
  INV_X1 U6447 ( .A(n10537), .ZN(n9382) );
  OR2_X1 U6448 ( .A1(n8999), .A2(n7142), .ZN(n10537) );
  INV_X1 U6449 ( .A(n9115), .ZN(n5173) );
  INV_X1 U6450 ( .A(n9217), .ZN(n9146) );
  NOR2_X1 U6451 ( .A1(n4412), .A2(n10221), .ZN(n4522) );
  OR2_X1 U6452 ( .A1(n10571), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4523) );
  AND2_X1 U6453 ( .A1(n5171), .A2(n5173), .ZN(n4524) );
  AND2_X1 U6454 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P1_REG3_REG_26__SCAN_IN), 
        .ZN(n4525) );
  INV_X1 U6455 ( .A(n9068), .ZN(n5174) );
  OR2_X1 U6456 ( .A1(n9102), .A2(n9071), .ZN(n4526) );
  AND2_X1 U6457 ( .A1(n4583), .A2(n7914), .ZN(n4527) );
  AND3_X2 U6458 ( .A1(n7971), .A2(n7166), .A3(n7165), .ZN(n10578) );
  INV_X1 U6459 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4833) );
  INV_X1 U6460 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n4841) );
  INV_X1 U6461 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6102) );
  XNOR2_X1 U6462 ( .A(n5722), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9176) );
  INV_X1 U6463 ( .A(n9176), .ZN(n5166) );
  INV_X1 U6464 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4838) );
  AND2_X1 U6465 ( .A1(n5149), .A2(n9200), .ZN(n4528) );
  INV_X1 U6466 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5001) );
  INV_X1 U6467 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4881) );
  INV_X1 U6468 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n4810) );
  INV_X1 U6469 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4640) );
  AOI21_X1 U6470 ( .B1(n10090), .B2(n10393), .A(n9941), .ZN(n4547) );
  XNOR2_X1 U6471 ( .A(n7210), .B(n7862), .ZN(n7860) );
  AOI21_X1 U6472 ( .B1(n7186), .B2(n7862), .A(n7187), .ZN(n7861) );
  OAI211_X1 U6473 ( .C1(n5179), .C2(n7862), .A(n5176), .B(n5175), .ZN(n7187)
         );
  OR2_X1 U6474 ( .A1(n4497), .A2(n7862), .ZN(n5175) );
  INV_X1 U6475 ( .A(n7862), .ZN(n5177) );
  NAND2_X1 U6476 ( .A1(n5133), .A2(n4529), .ZN(n5132) );
  AND2_X1 U6477 ( .A1(n4503), .A2(n4434), .ZN(n4530) );
  INV_X2 U6478 ( .A(n4555), .ZN(n7959) );
  NAND2_X2 U6479 ( .A1(n4534), .A2(n4476), .ZN(n6511) );
  XNOR2_X2 U6480 ( .A(n4535), .B(n6043), .ZN(n6049) );
  NAND2_X1 U6481 ( .A1(n6374), .A2(n4537), .ZN(n4536) );
  NAND2_X1 U6482 ( .A1(n4539), .A2(n4977), .ZN(n4538) );
  NAND2_X1 U6483 ( .A1(n6944), .A2(n6943), .ZN(n4539) );
  NAND2_X1 U6484 ( .A1(n6936), .A2(n4540), .ZN(n6944) );
  AND2_X1 U6485 ( .A1(n6935), .A2(n6934), .ZN(n4540) );
  NAND2_X1 U6486 ( .A1(n6998), .A2(n4542), .ZN(n4541) );
  AOI21_X1 U6487 ( .B1(n4543), .B2(n4446), .A(n4603), .ZN(n4542) );
  NAND2_X1 U6488 ( .A1(n6993), .A2(n6994), .ZN(n4543) );
  NAND4_X1 U6489 ( .A1(n4546), .A2(n7052), .A3(n7051), .A4(n4544), .ZN(
        P1_U3242) );
  NAND4_X1 U6490 ( .A1(n4965), .A2(n5282), .A3(n9872), .A4(n7021), .ZN(n4546)
         );
  INV_X1 U6491 ( .A(n6374), .ZN(n6243) );
  NAND2_X1 U6492 ( .A1(n4554), .A2(n6374), .ZN(n10212) );
  OAI22_X2 U6493 ( .A1(n10045), .A2(n4562), .B1(n4564), .B2(n6284), .ZN(n10005) );
  OAI21_X2 U6494 ( .B1(n9993), .B2(n4988), .A(n4565), .ZN(n9934) );
  INV_X1 U6495 ( .A(n9934), .ZN(n9937) );
  NAND2_X4 U6496 ( .A1(n5331), .A2(n5330), .ZN(n5487) );
  OR2_X1 U6497 ( .A1(n6186), .A2(n6915), .ZN(n6884) );
  OR2_X1 U6498 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  NAND2_X1 U6499 ( .A1(n5507), .A2(n5508), .ZN(n4581) );
  NAND2_X1 U6500 ( .A1(n5474), .A2(n5473), .ZN(n5508) );
  NAND2_X1 U6501 ( .A1(n7555), .A2(n4582), .ZN(n4586) );
  AND2_X1 U6502 ( .A1(n4587), .A2(n6534), .ZN(n7914) );
  NAND2_X1 U6503 ( .A1(n7555), .A2(n7912), .ZN(n4583) );
  NAND2_X1 U6504 ( .A1(n4585), .A2(n6534), .ZN(n4584) );
  INV_X1 U6505 ( .A(n4587), .ZN(n4585) );
  INV_X1 U6506 ( .A(n6533), .ZN(n4589) );
  NAND2_X1 U6507 ( .A1(n4592), .A2(n6699), .ZN(n6707) );
  INV_X1 U6508 ( .A(n4595), .ZN(n9658) );
  NAND2_X1 U6509 ( .A1(n9627), .A2(n9625), .ZN(n6666) );
  NAND2_X1 U6510 ( .A1(n4882), .A2(n5240), .ZN(n4656) );
  NAND2_X1 U6511 ( .A1(n6830), .A2(n6829), .ZN(n6996) );
  NAND2_X1 U6512 ( .A1(n4613), .A2(n7418), .ZN(n7437) );
  NAND3_X1 U6513 ( .A1(n4615), .A2(n5417), .A3(P2_IR_REG_31__SCAN_IN), .ZN(
        n4614) );
  AND2_X4 U6514 ( .A1(n5142), .A2(n5141), .ZN(n4720) );
  NAND3_X1 U6515 ( .A1(n4465), .A2(P2_REG2_REG_15__SCAN_IN), .A3(n4617), .ZN(
        n9122) );
  NAND3_X1 U6516 ( .A1(n5170), .A2(n4621), .A3(n9115), .ZN(n4617) );
  INV_X1 U6517 ( .A(n4622), .ZN(n4621) );
  XNOR2_X2 U6518 ( .A(n7188), .B(n7330), .ZN(n8009) );
  NAND3_X1 U6519 ( .A1(n4791), .A2(n4720), .A3(n5206), .ZN(n5302) );
  NAND3_X1 U6520 ( .A1(n4634), .A2(n7059), .A3(n4636), .ZN(n4632) );
  NAND3_X1 U6521 ( .A1(n4634), .A2(n7059), .A3(n10536), .ZN(n4633) );
  NAND3_X1 U6522 ( .A1(n5331), .A2(n5330), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n4637) );
  AND2_X1 U6523 ( .A1(n7896), .A2(n8992), .ZN(n8813) );
  NAND2_X1 U6524 ( .A1(n9256), .A2(n9255), .ZN(n4644) );
  NAND2_X1 U6525 ( .A1(n7094), .A2(n4645), .ZN(n9256) );
  NAND2_X1 U6526 ( .A1(n4646), .A2(n5456), .ZN(n4647) );
  AND2_X1 U6527 ( .A1(n7945), .A2(n5433), .ZN(n4648) );
  NAND2_X2 U6528 ( .A1(n5431), .A2(n5430), .ZN(n7819) );
  NAND2_X1 U6529 ( .A1(n7943), .A2(n5456), .ZN(n7988) );
  NAND2_X1 U6530 ( .A1(n4648), .A2(n7819), .ZN(n7943) );
  NAND2_X1 U6531 ( .A1(n8531), .A2(n4652), .ZN(n4650) );
  NAND2_X1 U6532 ( .A1(n4650), .A2(n4651), .ZN(n5188) );
  NAND2_X1 U6533 ( .A1(n9354), .A2(n9355), .ZN(n4654) );
  NAND2_X1 U6534 ( .A1(n9368), .A2(n8811), .ZN(n4655) );
  NAND3_X1 U6535 ( .A1(n5401), .A2(n5403), .A3(n5402), .ZN(n5383) );
  NAND2_X2 U6536 ( .A1(n5339), .A2(n5383), .ZN(n7291) );
  NAND2_X1 U6537 ( .A1(n5635), .A2(n4656), .ZN(n7527) );
  NAND3_X1 U6538 ( .A1(n5509), .A2(n4657), .A3(n5475), .ZN(n4661) );
  NAND2_X1 U6539 ( .A1(n4659), .A2(n4658), .ZN(n4657) );
  INV_X1 U6540 ( .A(n4661), .ZN(n5506) );
  OAI211_X1 U6541 ( .C1(n4665), .C2(n4460), .A(n8966), .B(n4662), .ZN(n4669)
         );
  NAND2_X1 U6542 ( .A1(n4663), .A2(n4666), .ZN(n4662) );
  INV_X1 U6543 ( .A(n4952), .ZN(n4663) );
  NAND2_X1 U6544 ( .A1(n4664), .A2(n8965), .ZN(n4670) );
  NAND2_X1 U6545 ( .A1(n4460), .A2(n4952), .ZN(n4664) );
  NOR2_X1 U6546 ( .A1(n4667), .A2(n8967), .ZN(n4666) );
  NAND2_X1 U6547 ( .A1(n4670), .A2(n4472), .ZN(n4668) );
  OAI21_X1 U6548 ( .B1(n4755), .B2(n4674), .A(n4672), .ZN(n4675) );
  NAND2_X1 U6549 ( .A1(n4754), .A2(n8985), .ZN(n4673) );
  INV_X1 U6550 ( .A(n8985), .ZN(n4674) );
  NAND2_X1 U6551 ( .A1(n4675), .A2(n7102), .ZN(n9003) );
  INV_X1 U6552 ( .A(n4676), .ZN(n4953) );
  OAI21_X4 U6553 ( .B1(n5551), .B2(n5550), .A(n5549), .ZN(n5579) );
  NAND2_X1 U6554 ( .A1(n4683), .A2(n10528), .ZN(n6508) );
  NAND2_X1 U6555 ( .A1(n4683), .A2(n10510), .ZN(n6785) );
  INV_X1 U6556 ( .A(n8092), .ZN(n4692) );
  NAND3_X1 U6557 ( .A1(n4688), .A2(n4690), .A3(n4687), .ZN(n10371) );
  NAND4_X1 U6558 ( .A1(n4688), .A2(n4687), .A3(n4690), .A4(n4686), .ZN(n4698)
         );
  NAND2_X1 U6559 ( .A1(n4692), .A2(n4691), .ZN(n4687) );
  NAND2_X1 U6560 ( .A1(n4689), .A2(n4699), .ZN(n4688) );
  OR2_X1 U6561 ( .A1(n6438), .A2(n4693), .ZN(n4690) );
  NAND2_X1 U6562 ( .A1(n8092), .A2(n4441), .ZN(n4694) );
  INV_X1 U6563 ( .A(n5254), .ZN(n4695) );
  OAI21_X2 U6564 ( .B1(n6398), .B2(n5137), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4700) );
  AND2_X1 U6565 ( .A1(n10027), .A2(n9686), .ZN(n4704) );
  AOI21_X1 U6566 ( .B1(n8412), .B2(n5265), .A(n5263), .ZN(n8503) );
  NAND2_X1 U6567 ( .A1(n4707), .A2(n4706), .ZN(n8596) );
  NAND2_X1 U6568 ( .A1(n8412), .A2(n4510), .ZN(n4706) );
  OR2_X1 U6569 ( .A1(n6539), .A2(n7999), .ZN(n4712) );
  NAND2_X1 U6570 ( .A1(n4712), .A2(n6430), .ZN(n8103) );
  NAND2_X1 U6571 ( .A1(n6798), .A2(n4712), .ZN(n6802) );
  NAND2_X1 U6572 ( .A1(n5132), .A2(n4712), .ZN(n10377) );
  NAND2_X1 U6573 ( .A1(n7431), .A2(n7205), .ZN(n4716) );
  NAND2_X1 U6574 ( .A1(n4720), .A2(n5417), .ZN(n5439) );
  NAND2_X1 U6575 ( .A1(n4720), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7180) );
  NAND2_X1 U6576 ( .A1(n4720), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7199) );
  XNOR2_X1 U6577 ( .A(n5380), .B(n10538), .ZN(n7545) );
  NAND2_X1 U6578 ( .A1(n5197), .A2(n4508), .ZN(n8713) );
  NAND2_X1 U6579 ( .A1(n5589), .A2(n8535), .ZN(n8477) );
  XNOR2_X2 U6580 ( .A(n5370), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9534) );
  NAND3_X1 U6581 ( .A1(n5138), .A2(n5351), .A3(n5637), .ZN(n9529) );
  NAND2_X1 U6582 ( .A1(n8789), .A2(n5692), .ZN(n8706) );
  OR2_X1 U6583 ( .A1(n6902), .A2(n6812), .ZN(n6815) );
  NAND2_X1 U6584 ( .A1(n4974), .A2(n10046), .ZN(n6957) );
  NAND3_X2 U6585 ( .A1(n5349), .A2(n4769), .A3(n5350), .ZN(n8868) );
  NAND2_X1 U6586 ( .A1(n6947), .A2(n7010), .ZN(n4978) );
  AOI21_X1 U6587 ( .B1(n6993), .B2(n6992), .A(n4498), .ZN(n6997) );
  OAI21_X1 U6588 ( .B1(n4982), .B2(n6960), .A(n4980), .ZN(n6982) );
  AND2_X1 U6589 ( .A1(n4731), .A2(n6524), .ZN(n7557) );
  NAND2_X1 U6590 ( .A1(n7532), .A2(n7533), .ZN(n4731) );
  AOI21_X2 U6591 ( .B1(n10002), .B2(n6445), .A(n6444), .ZN(n9991) );
  NAND2_X1 U6592 ( .A1(n6436), .A2(n6435), .ZN(n8092) );
  INV_X1 U6593 ( .A(n9909), .ZN(n5008) );
  OAI211_X1 U6594 ( .C1(n4733), .C2(n4732), .A(n9700), .B(n9716), .ZN(n4768)
         );
  AOI21_X1 U6595 ( .B1(n9700), .B2(n4794), .A(n4793), .ZN(n8633) );
  NAND2_X1 U6596 ( .A1(n9648), .A2(n6688), .ZN(n5020) );
  NAND2_X1 U6597 ( .A1(n6512), .A2(n4749), .ZN(n4763) );
  AND2_X2 U6598 ( .A1(n5272), .A2(n7912), .ZN(n7556) );
  NAND2_X2 U6599 ( .A1(n4814), .A2(n7972), .ZN(n5400) );
  AND2_X2 U6600 ( .A1(n5327), .A2(n7315), .ZN(n7972) );
  MUX2_X1 U6601 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9549), .S(n7176), .Z(n7982) );
  NAND2_X2 U6602 ( .A1(n5378), .A2(n7278), .ZN(n7176) );
  XNOR2_X1 U6603 ( .A(n9866), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9871) );
  AOI21_X1 U6604 ( .B1(n10243), .B2(P1_REG2_REG_14__SCAN_IN), .A(n10242), .ZN(
        n9859) );
  MUX2_X1 U6605 ( .A(n7394), .B(P1_REG2_REG_2__SCAN_IN), .S(n7839), .Z(n7838)
         );
  INV_X1 U6606 ( .A(n7408), .ZN(n4741) );
  INV_X1 U6607 ( .A(n7890), .ZN(n4743) );
  NOR2_X1 U6608 ( .A1(n9860), .A2(n10255), .ZN(n10271) );
  NAND2_X1 U6609 ( .A1(n7886), .A2(n7885), .ZN(n9836) );
  NAND2_X1 U6610 ( .A1(n9118), .A2(n9117), .ZN(n9139) );
  AOI21_X2 U6611 ( .B1(n9180), .B2(n9179), .A(n9178), .ZN(n9182) );
  NAND2_X1 U6612 ( .A1(n9097), .A2(n9096), .ZN(n9099) );
  INV_X1 U6613 ( .A(n7464), .ZN(n4745) );
  NOR2_X2 U6614 ( .A1(n9184), .A2(n9195), .ZN(n9186) );
  NAND2_X1 U6615 ( .A1(n9075), .A2(n9076), .ZN(n9097) );
  NAND2_X1 U6616 ( .A1(n7253), .A2(n7930), .ZN(n8013) );
  NAND2_X1 U6617 ( .A1(n7263), .A2(n8119), .ZN(n8234) );
  NAND2_X1 U6618 ( .A1(n7272), .A2(n7273), .ZN(n9053) );
  NAND2_X1 U6619 ( .A1(n9049), .A2(n9050), .ZN(n9079) );
  NAND2_X1 U6620 ( .A1(n7268), .A2(n8231), .ZN(n8236) );
  NAND2_X1 U6621 ( .A1(n8677), .A2(n8678), .ZN(n8676) );
  AOI21_X2 U6622 ( .B1(n8757), .B2(n5830), .A(n5829), .ZN(n8723) );
  NAND2_X1 U6623 ( .A1(n8533), .A2(n8532), .ZN(n8531) );
  NAND2_X1 U6624 ( .A1(n5184), .A2(n5294), .ZN(n4747) );
  NAND2_X1 U6625 ( .A1(n5274), .A2(n5187), .ZN(n5186) );
  NAND2_X1 U6626 ( .A1(n4861), .A2(n5278), .ZN(P2_U3488) );
  NAND2_X2 U6627 ( .A1(n4748), .A2(n7056), .ZN(n7108) );
  INV_X1 U6628 ( .A(n4774), .ZN(n4748) );
  AND3_X4 U6629 ( .A1(n5390), .A2(n5391), .A3(n5389), .ZN(n4774) );
  NAND2_X1 U6630 ( .A1(n5787), .A2(n5786), .ZN(n8735) );
  NAND2_X1 U6631 ( .A1(n8735), .A2(n5788), .ZN(n8677) );
  NAND2_X1 U6632 ( .A1(n8275), .A2(n8858), .ZN(n7114) );
  NAND2_X1 U6633 ( .A1(n9008), .A2(n9007), .ZN(n5110) );
  NAND2_X2 U6634 ( .A1(n9232), .A2(n9234), .ZN(n9231) );
  INV_X1 U6635 ( .A(n6525), .ZN(n6542) );
  NAND2_X1 U6636 ( .A1(n4750), .A2(n6525), .ZN(n4749) );
  AND2_X4 U6637 ( .A1(n7171), .A2(n6509), .ZN(n6525) );
  NAND2_X1 U6638 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  AND2_X1 U6639 ( .A1(n6139), .A2(n4505), .ZN(n4752) );
  NAND2_X1 U6640 ( .A1(n4959), .A2(n4958), .ZN(n4755) );
  OAI211_X1 U6641 ( .C1(n10163), .C2(n10205), .A(n4517), .B(n4756), .ZN(
        P1_U3517) );
  NAND2_X1 U6642 ( .A1(n5591), .A2(n8476), .ZN(n8533) );
  NAND2_X1 U6643 ( .A1(n8706), .A2(n8705), .ZN(n5197) );
  XNOR2_X1 U6644 ( .A(n5388), .B(n5387), .ZN(n6137) );
  NAND2_X1 U6645 ( .A1(n10173), .A2(n10528), .ZN(n4760) );
  OAI21_X1 U6646 ( .B1(n10105), .B2(n10153), .A(n4499), .ZN(n10173) );
  NAND2_X1 U6647 ( .A1(n9991), .A2(n4781), .ZN(n9960) );
  NAND3_X1 U6648 ( .A1(n5401), .A2(n5402), .A3(n5404), .ZN(n5408) );
  AOI21_X1 U6649 ( .B1(n10355), .B2(n10354), .A(n4501), .ZN(n10334) );
  NAND2_X1 U6650 ( .A1(n6523), .A2(n5273), .ZN(n7533) );
  AND2_X1 U6651 ( .A1(n6978), .A2(n6823), .ZN(n6975) );
  NAND2_X1 U6652 ( .A1(n10296), .A2(n10295), .ZN(n10294) );
  AOI21_X1 U6653 ( .B1(n9186), .B2(P2_U3893), .A(n9209), .ZN(n9188) );
  NAND2_X1 U6654 ( .A1(n7493), .A2(n7492), .ZN(n7495) );
  NAND2_X1 U6655 ( .A1(n8046), .A2(n8045), .ZN(n8048) );
  OR2_X1 U6656 ( .A1(n9874), .A2(n9872), .ZN(n4770) );
  NAND2_X1 U6657 ( .A1(n9810), .A2(n9811), .ZN(n9809) );
  NAND2_X1 U6658 ( .A1(n7190), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5164) );
  NOR2_X1 U6659 ( .A1(n5167), .A2(n5166), .ZN(n5165) );
  INV_X1 U6660 ( .A(n8112), .ZN(n4762) );
  NAND2_X1 U6661 ( .A1(n5188), .A2(n5667), .ZN(n8650) );
  OAI21_X1 U6662 ( .B1(n4798), .B2(n4797), .A(n9353), .ZN(n8953) );
  NAND2_X1 U6663 ( .A1(n4937), .A2(n4936), .ZN(n4935) );
  NAND2_X1 U6664 ( .A1(n4768), .A2(n4766), .ZN(P1_U3240) );
  AND2_X1 U6665 ( .A1(n6521), .A2(n6520), .ZN(n6523) );
  NAND2_X1 U6666 ( .A1(n5342), .A2(n9199), .ZN(n4769) );
  NAND3_X1 U6667 ( .A1(n8026), .A2(n4847), .A3(n8891), .ZN(n4845) );
  NAND2_X1 U6668 ( .A1(n10529), .A2(n7108), .ZN(n8026) );
  AOI21_X2 U6669 ( .B1(n8064), .B2(n8814), .A(n7112), .ZN(n8192) );
  NAND2_X1 U6670 ( .A1(n4852), .A2(n4851), .ZN(n7123) );
  NAND2_X1 U6671 ( .A1(n7897), .A2(n7107), .ZN(n10530) );
  AOI21_X1 U6672 ( .B1(n5110), .B2(n5109), .A(n5108), .ZN(n9012) );
  NAND3_X1 U6673 ( .A1(n4773), .A2(n4771), .A3(n4770), .ZN(P1_U3262) );
  NOR2_X1 U6674 ( .A1(n10252), .A2(n9848), .ZN(n10264) );
  NOR2_X2 U6675 ( .A1(n10409), .A2(n6539), .ZN(n10391) );
  NOR2_X2 U6676 ( .A1(n10372), .A2(n6394), .ZN(n8421) );
  NAND2_X1 U6678 ( .A1(n7456), .A2(n10429), .ZN(n10408) );
  AND3_X2 U6679 ( .A1(n10036), .A2(n5075), .A3(n5076), .ZN(n9996) );
  NAND2_X1 U6680 ( .A1(n5049), .A2(n5051), .ZN(n9266) );
  OAI21_X1 U6681 ( .B1(n5043), .B2(n5045), .A(n8932), .ZN(n5042) );
  NAND2_X1 U6682 ( .A1(n6788), .A2(n8790), .ZN(n4803) );
  NOR2_X1 U6683 ( .A1(n6787), .A2(n6786), .ZN(n4802) );
  NAND2_X1 U6684 ( .A1(n4783), .A2(n4782), .ZN(n5342) );
  NAND2_X1 U6685 ( .A1(n7291), .A2(n7290), .ZN(n4783) );
  NAND2_X1 U6686 ( .A1(n4790), .A2(n4788), .ZN(P1_U3214) );
  OAI21_X1 U6687 ( .B1(n8633), .B2(n8634), .A(n9716), .ZN(n4790) );
  NAND2_X1 U6688 ( .A1(n9144), .A2(n9143), .ZN(n5167) );
  AOI21_X1 U6689 ( .B1(n4820), .B2(n4566), .A(n4986), .ZN(n4817) );
  OAI211_X1 U6690 ( .C1(n9214), .C2(n9213), .A(n5143), .B(n4805), .ZN(P2_U3201) );
  NAND2_X2 U6691 ( .A1(n10003), .A2(n6965), .ZN(n9993) );
  NAND2_X1 U6692 ( .A1(n4956), .A2(n8947), .ZN(n4954) );
  NAND2_X1 U6693 ( .A1(n4953), .A2(n4677), .ZN(n4949) );
  OAI211_X1 U6694 ( .C1(n4886), .C2(n5579), .A(n5241), .B(n4883), .ZN(n4882)
         );
  AOI21_X1 U6695 ( .B1(n8990), .B2(n8999), .A(n8989), .ZN(n9002) );
  NAND2_X1 U6696 ( .A1(n8943), .A2(n8948), .ZN(n4797) );
  INV_X1 U6697 ( .A(n8944), .ZN(n4798) );
  NAND2_X1 U6698 ( .A1(n4939), .A2(n8999), .ZN(n4938) );
  NAND2_X1 U6699 ( .A1(n4934), .A2(n8924), .ZN(n4933) );
  OAI21_X1 U6700 ( .B1(n9002), .B2(n4485), .A(n8996), .ZN(n8997) );
  NAND2_X1 U6701 ( .A1(n10154), .A2(n10510), .ZN(n10156) );
  NAND2_X1 U6702 ( .A1(n4818), .A2(n4817), .ZN(n9924) );
  NAND3_X1 U6703 ( .A1(n4801), .A2(n9191), .A3(n9190), .ZN(P2_U3200) );
  OAI21_X1 U6704 ( .B1(n9166), .B2(n9194), .A(n9146), .ZN(n4801) );
  NAND2_X1 U6705 ( .A1(n9124), .A2(n9123), .ZN(n9144) );
  NAND2_X2 U6706 ( .A1(n5637), .A2(n5314), .ZN(n5340) );
  OAI21_X1 U6707 ( .B1(n4803), .B2(n4802), .A(n6794), .ZN(P2_U3154) );
  AND2_X1 U6708 ( .A1(n5011), .A2(n5009), .ZN(n10161) );
  NAND2_X1 U6709 ( .A1(n5011), .A2(n9908), .ZN(n10081) );
  NAND2_X1 U6710 ( .A1(n8617), .A2(n10507), .ZN(n4804) );
  NAND2_X1 U6711 ( .A1(n7520), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4815) );
  OAI21_X1 U6712 ( .B1(n7042), .B2(n8628), .A(n4807), .ZN(n6514) );
  XNOR2_X1 U6713 ( .A(n9083), .B(n9060), .ZN(n9061) );
  OAI21_X1 U6714 ( .B1(n7520), .B2(P2_REG1_REG_2__SCAN_IN), .A(n4815), .ZN(
        n7517) );
  INV_X1 U6715 ( .A(n5621), .ZN(n4906) );
  OAI21_X1 U6716 ( .B1(n8968), .B2(n8969), .A(n4960), .ZN(n4959) );
  AOI21_X1 U6717 ( .B1(n9205), .B2(n9204), .A(n4808), .ZN(n9207) );
  INV_X1 U6718 ( .A(n4887), .ZN(n4886) );
  INV_X1 U6719 ( .A(n5044), .ZN(n5043) );
  NAND2_X1 U6720 ( .A1(n5048), .A2(n7083), .ZN(n9368) );
  INV_X1 U6721 ( .A(n5042), .ZN(n5041) );
  AND2_X1 U6722 ( .A1(n8914), .A2(n8306), .ZN(n8858) );
  NAND2_X1 U6723 ( .A1(n4889), .A2(n4890), .ZN(n5584) );
  NAND2_X1 U6724 ( .A1(n8913), .A2(n8916), .ZN(n4939) );
  NAND2_X1 U6725 ( .A1(n8918), .A2(n7115), .ZN(n4937) );
  AOI21_X1 U6726 ( .B1(n4933), .B2(n8931), .A(n8930), .ZN(n8939) );
  OAI21_X1 U6727 ( .B1(n4953), .B2(n4957), .A(n8953), .ZN(n4952) );
  AND2_X2 U6728 ( .A1(n5328), .A2(n7104), .ZN(n4814) );
  OR2_X1 U6729 ( .A1(n8867), .A2(n5379), .ZN(n7546) );
  NAND2_X1 U6730 ( .A1(n4989), .A2(n4820), .ZN(n4818) );
  NAND2_X1 U6731 ( .A1(n4821), .A2(n4825), .ZN(n6458) );
  NAND2_X1 U6732 ( .A1(n5867), .A2(n4831), .ZN(n5907) );
  NAND2_X1 U6733 ( .A1(n5867), .A2(n4520), .ZN(n5930) );
  NAND2_X1 U6734 ( .A1(n5867), .A2(n5866), .ZN(n5893) );
  NAND2_X1 U6735 ( .A1(n5458), .A2(n4832), .ZN(n5523) );
  NAND2_X1 U6736 ( .A1(n5522), .A2(n4837), .ZN(n5569) );
  NAND2_X1 U6737 ( .A1(n5681), .A2(n4839), .ZN(n5761) );
  NAND3_X1 U6738 ( .A1(n4847), .A2(n4848), .A3(n8891), .ZN(n4846) );
  NAND2_X1 U6739 ( .A1(n8886), .A2(n8889), .ZN(n4847) );
  NAND2_X1 U6740 ( .A1(n8886), .A2(n8890), .ZN(n4848) );
  INV_X2 U6741 ( .A(n7176), .ZN(n5756) );
  NAND2_X1 U6742 ( .A1(n9351), .A2(n4854), .ZN(n4852) );
  OAI21_X2 U6743 ( .B1(n5340), .B2(P2_IR_REG_26__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6744 ( .A1(n7127), .A2(n4863), .ZN(n4864) );
  NAND2_X1 U6745 ( .A1(n4864), .A2(n4865), .ZN(n9232) );
  NAND2_X1 U6746 ( .A1(n4878), .A2(n4875), .ZN(n4874) );
  NAND3_X1 U6747 ( .A1(n4874), .A2(n4873), .A3(n4511), .ZN(n4871) );
  NAND2_X1 U6748 ( .A1(n4878), .A2(n4877), .ZN(n9008) );
  NAND3_X1 U6749 ( .A1(n4874), .A2(n4873), .A3(n4876), .ZN(n7146) );
  NAND2_X1 U6750 ( .A1(n4889), .A2(n4887), .ZN(n5593) );
  NAND2_X1 U6751 ( .A1(n5697), .A2(n4896), .ZN(n4895) );
  NAND2_X1 U6752 ( .A1(n5883), .A2(n5882), .ZN(n5889) );
  MUX2_X1 U6753 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4414), .Z(n5617) );
  MUX2_X1 U6754 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5487), .Z(n5614) );
  MUX2_X1 U6755 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5487), .Z(n5630) );
  MUX2_X1 U6756 ( .A(n8037), .B(n5698), .S(n4414), .Z(n5713) );
  MUX2_X1 U6757 ( .A(n8211), .B(n5735), .S(n4414), .Z(n5736) );
  MUX2_X1 U6758 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4413), .Z(n5672) );
  MUX2_X1 U6759 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4413), .Z(n5693) );
  MUX2_X1 U6760 ( .A(n8274), .B(n8272), .S(n5487), .Z(n5739) );
  MUX2_X1 U6761 ( .A(n8441), .B(n8439), .S(n5487), .Z(n5817) );
  MUX2_X1 U6762 ( .A(n8336), .B(n8317), .S(n5487), .Z(n5810) );
  MUX2_X1 U6763 ( .A(n8454), .B(n8458), .S(n4414), .Z(n5835) );
  MUX2_X1 U6764 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4413), .Z(n5814) );
  MUX2_X1 U6765 ( .A(n8493), .B(n8490), .S(n5487), .Z(n5858) );
  MUX2_X1 U6766 ( .A(n8579), .B(n8582), .S(n4414), .Z(n5885) );
  MUX2_X1 U6767 ( .A(n8594), .B(n10225), .S(n4413), .Z(n5902) );
  MUX2_X1 U6768 ( .A(n7736), .B(n8627), .S(n5487), .Z(n5923) );
  MUX2_X1 U6769 ( .A(n5938), .B(n8640), .S(n4414), .Z(n6467) );
  MUX2_X1 U6770 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4413), .Z(n6848) );
  NAND2_X1 U6771 ( .A1(n5697), .A2(n4416), .ZN(n4917) );
  NAND2_X1 U6772 ( .A1(n5806), .A2(n4928), .ZN(n4923) );
  NAND2_X1 U6773 ( .A1(n4923), .A2(n4925), .ZN(n5862) );
  NAND3_X1 U6774 ( .A1(n4938), .A2(n4935), .A3(n8919), .ZN(n4934) );
  NOR2_X2 U6775 ( .A1(n4945), .A2(n4940), .ZN(n5314) );
  NAND4_X1 U6776 ( .A1(n4944), .A2(n4943), .A3(n4942), .A4(n4941), .ZN(n4940)
         );
  NAND4_X1 U6777 ( .A1(n5313), .A2(n5311), .A3(n5324), .A4(n5312), .ZN(n4945)
         );
  AND2_X1 U6778 ( .A1(n5637), .A2(n5138), .ZN(n5357) );
  NAND2_X2 U6779 ( .A1(n9529), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6780 ( .A1(n4487), .A2(n8991), .ZN(n4948) );
  AND2_X1 U6781 ( .A1(n8962), .A2(n4951), .ZN(n4950) );
  AOI21_X1 U6782 ( .B1(n4957), .B2(n8954), .A(n4447), .ZN(n4951) );
  AND2_X1 U6783 ( .A1(n8952), .A2(n8960), .ZN(n4957) );
  AND2_X1 U6784 ( .A1(n8978), .A2(n4507), .ZN(n4960) );
  NAND2_X2 U6785 ( .A1(n8306), .A2(n8855), .ZN(n8819) );
  OR2_X2 U6786 ( .A1(n8611), .A2(n8309), .ZN(n8306) );
  AND2_X2 U6787 ( .A1(n4500), .A2(n5562), .ZN(n8309) );
  NAND2_X1 U6788 ( .A1(n6928), .A2(n6919), .ZN(n6920) );
  NAND2_X1 U6789 ( .A1(n6911), .A2(n4504), .ZN(n4962) );
  INV_X1 U6790 ( .A(n4969), .ZN(n4963) );
  INV_X1 U6791 ( .A(n4971), .ZN(n4964) );
  OAI211_X1 U6792 ( .C1(n7012), .C2(n4968), .A(n4967), .B(n4966), .ZN(n4965)
         );
  NAND2_X1 U6793 ( .A1(n4969), .A2(n7024), .ZN(n4967) );
  NAND2_X1 U6794 ( .A1(n4971), .A2(n7024), .ZN(n4968) );
  OAI21_X2 U6795 ( .B1(n4973), .B2(n10079), .A(n4970), .ZN(n4969) );
  NAND2_X1 U6796 ( .A1(n4973), .A2(n4972), .ZN(n4971) );
  NAND2_X1 U6797 ( .A1(n4979), .A2(n6976), .ZN(n4983) );
  INV_X1 U6798 ( .A(n4988), .ZN(n4987) );
  OAI21_X1 U6799 ( .B1(n4995), .B2(n4993), .A(n9971), .ZN(n4988) );
  OAI21_X1 U6800 ( .B1(n9993), .B2(n4991), .A(n4990), .ZN(n9970) );
  OAI21_X1 U6801 ( .B1(n9993), .B2(n6303), .A(n6962), .ZN(n9981) );
  AOI21_X1 U6802 ( .B1(n6962), .B2(n6303), .A(n9980), .ZN(n4995) );
  NAND3_X1 U6803 ( .A1(n5000), .A2(n4998), .A3(n4997), .ZN(n5436) );
  NAND3_X1 U6804 ( .A1(n5331), .A2(n5330), .A3(n5001), .ZN(n4997) );
  NAND2_X1 U6805 ( .A1(n4999), .A2(n5002), .ZN(n4998) );
  INV_X1 U6806 ( .A(n5331), .ZN(n4999) );
  OAI211_X1 U6807 ( .C1(n10163), .C2(n10145), .A(n5006), .B(n5003), .ZN(
        P1_U3549) );
  NAND3_X1 U6808 ( .A1(n5008), .A2(n5007), .A3(n10528), .ZN(n5006) );
  NAND2_X1 U6809 ( .A1(n5007), .A2(n5008), .ZN(n5011) );
  NAND2_X1 U6810 ( .A1(n7996), .A2(n6556), .ZN(n6563) );
  NAND2_X1 U6811 ( .A1(n7996), .A2(n5021), .ZN(n8153) );
  NOR2_X1 U6812 ( .A1(n5022), .A2(n6562), .ZN(n5021) );
  NAND2_X1 U6813 ( .A1(n9634), .A2(n4506), .ZN(n5025) );
  NAND2_X1 U6814 ( .A1(n5033), .A2(n5438), .ZN(n5471) );
  INV_X2 U6815 ( .A(n6364), .ZN(n5036) );
  INV_X1 U6816 ( .A(n8927), .ZN(n5046) );
  NAND2_X1 U6817 ( .A1(n9301), .A2(n5052), .ZN(n5051) );
  OAI21_X2 U6818 ( .B1(n9344), .B2(n7086), .A(n7087), .ZN(n9313) );
  OAI21_X1 U6819 ( .B1(n7080), .B2(n5063), .A(n7079), .ZN(n5062) );
  XNOR2_X1 U6820 ( .A(n9226), .B(n9225), .ZN(n5071) );
  AOI21_X1 U6821 ( .B1(n4413), .B2(n5074), .A(n5073), .ZN(n5336) );
  OAI21_X2 U6822 ( .B1(n9578), .B2(n6683), .A(n6682), .ZN(n9648) );
  INV_X2 U6823 ( .A(n6140), .ZN(n6126) );
  OAI211_X2 U6824 ( .C1(n7044), .C2(n7024), .A(n8090), .B(n7171), .ZN(n6529)
         );
  OAI211_X1 U6825 ( .C1(n7552), .C2(n6529), .A(n6519), .B(n6518), .ZN(n7532)
         );
  NAND2_X1 U6826 ( .A1(n6666), .A2(n9624), .ZN(n9578) );
  INV_X1 U6827 ( .A(n5080), .ZN(n8300) );
  AND2_X2 U6828 ( .A1(n4502), .A2(n8524), .ZN(n10067) );
  NAND4_X1 U6829 ( .A1(n6027), .A2(n6031), .A3(n4435), .A4(n6026), .ZN(n6032)
         );
  NAND2_X1 U6830 ( .A1(n8428), .A2(n5093), .ZN(n5092) );
  NAND2_X1 U6831 ( .A1(n5092), .A2(n5095), .ZN(n9377) );
  AND2_X1 U6832 ( .A1(n5375), .A2(n5376), .ZN(n5099) );
  INV_X1 U6833 ( .A(n8975), .ZN(n5116) );
  NAND2_X1 U6834 ( .A1(n9924), .A2(n5118), .ZN(n5117) );
  NAND2_X1 U6835 ( .A1(n5117), .A2(n5120), .ZN(n6479) );
  OAI21_X1 U6836 ( .B1(n9924), .B2(n5122), .A(n4509), .ZN(n6459) );
  NAND2_X1 U6837 ( .A1(n6148), .A2(n6800), .ZN(n5129) );
  NAND2_X1 U6838 ( .A1(n7114), .A2(n5135), .ZN(n5134) );
  NAND2_X1 U6839 ( .A1(n5134), .A2(n8916), .ZN(n8390) );
  INV_X2 U6840 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5141) );
  NAND4_X1 U6841 ( .A1(n5146), .A2(n5145), .A3(n5148), .A4(n5144), .ZN(n5143)
         );
  NAND3_X1 U6842 ( .A1(n5154), .A2(n9165), .A3(n9200), .ZN(n5144) );
  AOI21_X1 U6843 ( .B1(n9165), .B2(n9164), .A(n9163), .ZN(n9194) );
  INV_X1 U6844 ( .A(n9200), .ZN(n5151) );
  INV_X1 U6845 ( .A(n5154), .ZN(n5152) );
  INV_X1 U6846 ( .A(n7194), .ZN(n5163) );
  AOI21_X1 U6847 ( .B1(n7194), .B2(n7193), .A(n4519), .ZN(n5160) );
  CLKBUF_X1 U6848 ( .A(n5164), .Z(n5155) );
  INV_X1 U6849 ( .A(n7469), .ZN(n5181) );
  NAND3_X1 U6850 ( .A1(n7182), .A2(n7437), .A3(P2_REG2_REG_3__SCAN_IN), .ZN(
        n7420) );
  NAND2_X1 U6851 ( .A1(n7182), .A2(n7437), .ZN(n5183) );
  NAND2_X1 U6852 ( .A1(n5183), .A2(n5422), .ZN(n5182) );
  NAND2_X1 U6853 ( .A1(n5294), .A2(n5185), .ZN(n5295) );
  INV_X1 U6854 ( .A(n5188), .ZN(n8649) );
  OR2_X1 U6855 ( .A1(n8686), .A2(n9028), .ZN(n5196) );
  OAI21_X1 U6856 ( .B1(n8723), .B2(n4453), .A(n5881), .ZN(n8697) );
  NAND2_X1 U6857 ( .A1(n5200), .A2(n5198), .ZN(n8775) );
  NAND2_X1 U6858 ( .A1(n8723), .A2(n5881), .ZN(n5200) );
  AND2_X2 U6859 ( .A1(n8340), .A2(n5568), .ZN(n5589) );
  AOI21_X1 U6860 ( .B1(n5202), .B2(n8055), .A(n4488), .ZN(n5201) );
  INV_X1 U6861 ( .A(n5514), .ZN(n5208) );
  NAND3_X1 U6862 ( .A1(n5508), .A2(n5507), .A3(n5515), .ZN(n5209) );
  OAI21_X1 U6863 ( .B1(n5769), .B2(n5223), .A(n5219), .ZN(n5212) );
  INV_X1 U6864 ( .A(n5214), .ZN(n5213) );
  OAI21_X1 U6865 ( .B1(n5769), .B2(n5217), .A(n5215), .ZN(n5214) );
  OAI21_X1 U6866 ( .B1(n5219), .B2(n5218), .A(n5771), .ZN(n5216) );
  NAND2_X1 U6867 ( .A1(n5770), .A2(n5222), .ZN(n5219) );
  NAND2_X1 U6868 ( .A1(n5769), .A2(n5221), .ZN(n5220) );
  NOR2_X1 U6869 ( .A1(n5770), .A2(n5222), .ZN(n5221) );
  INV_X1 U6870 ( .A(n5770), .ZN(n5223) );
  NAND2_X1 U6871 ( .A1(n7106), .A2(n10541), .ZN(n5224) );
  NAND4_X1 U6872 ( .A1(n5224), .A2(n4425), .A3(n10571), .A4(n7147), .ZN(n7155)
         );
  AND2_X1 U6873 ( .A1(n5224), .A2(n4425), .ZN(n8648) );
  NAND2_X1 U6874 ( .A1(n5411), .A2(SI_3_), .ZN(n5434) );
  OAI21_X1 U6875 ( .B1(n5487), .B2(n5410), .A(n5232), .ZN(n5411) );
  NAND2_X1 U6876 ( .A1(n4414), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5232) );
  INV_X1 U6877 ( .A(n5615), .ZN(n5244) );
  NAND2_X1 U6878 ( .A1(n8092), .A2(n8093), .ZN(n5256) );
  INV_X1 U6879 ( .A(n8840), .ZN(n9453) );
  INV_X1 U6880 ( .A(n9010), .ZN(n9450) );
  OAI21_X1 U6881 ( .B1(n4494), .B2(n8270), .A(n7025), .ZN(n7026) );
  NAND2_X1 U6882 ( .A1(n10158), .A2(n10080), .ZN(n6457) );
  XNOR2_X1 U6883 ( .A(n5358), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5366) );
  NOR2_X1 U6884 ( .A1(n7088), .A2(n9305), .ZN(n7089) );
  CLKBUF_X1 U6885 ( .A(n9301), .Z(n9303) );
  INV_X1 U6886 ( .A(n5366), .ZN(n5372) );
  OR2_X1 U6887 ( .A1(n5357), .A2(n9528), .ZN(n5358) );
  AND2_X1 U6888 ( .A1(P2_U3893), .A2(n7278), .ZN(n9215) );
  NOR2_X1 U6889 ( .A1(n8998), .A2(n8997), .ZN(n9015) );
  INV_X1 U6890 ( .A(n9534), .ZN(n5373) );
  OAI21_X2 U6891 ( .B1(n7092), .B2(n7091), .A(n7090), .ZN(n9301) );
  INV_X1 U6892 ( .A(n5967), .ZN(n8863) );
  NAND2_X1 U6893 ( .A1(n6243), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6251) );
  OR2_X1 U6894 ( .A1(n6143), .A2(n6127), .ZN(n6129) );
  NAND2_X1 U6895 ( .A1(n9527), .A2(n5036), .ZN(n6868) );
  CLKBUF_X1 U6896 ( .A(n5971), .Z(n8994) );
  INV_X1 U6897 ( .A(n5971), .ZN(n8992) );
  INV_X1 U6898 ( .A(n8895), .ZN(n7112) );
  OR2_X1 U6899 ( .A1(n7171), .A2(n6522), .ZN(n5273) );
  NOR2_X1 U6900 ( .A1(n10402), .A2(n7952), .ZN(n10332) );
  AND3_X1 U6901 ( .A1(n5313), .A2(n5675), .A3(n5311), .ZN(n5274) );
  NOR2_X1 U6902 ( .A1(n5842), .A2(n5841), .ZN(n5276) );
  AND2_X2 U6903 ( .A1(n8421), .A2(n6395), .ZN(n5279) );
  NAND2_X1 U6904 ( .A1(n9385), .A2(n8025), .ZN(n9366) );
  AND2_X1 U6905 ( .A1(n6848), .A2(n6466), .ZN(n5280) );
  INV_X1 U6906 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8317) );
  INV_X1 U6907 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5410) );
  INV_X1 U6908 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5468) );
  INV_X1 U6909 ( .A(n6049), .ZN(n6046) );
  AND2_X1 U6910 ( .A1(n7044), .A2(n7483), .ZN(n10490) );
  NAND2_X1 U6911 ( .A1(n8094), .A2(n8181), .ZN(n5281) );
  INV_X1 U6912 ( .A(n10489), .ZN(n6395) );
  AND2_X1 U6913 ( .A1(n7049), .A2(n7047), .ZN(n5282) );
  OR2_X1 U6914 ( .A1(n10079), .A2(n7010), .ZN(n5283) );
  AND2_X1 U6915 ( .A1(n9330), .A2(n9314), .ZN(n5284) );
  AND3_X1 U6916 ( .A1(n5982), .A2(n6013), .A3(n8790), .ZN(n5286) );
  AND2_X1 U6917 ( .A1(n8837), .A2(n9237), .ZN(n5287) );
  NOR2_X1 U6918 ( .A1(n6501), .A2(n6500), .ZN(n5288) );
  INV_X1 U6919 ( .A(n8725), .ZN(n5875) );
  BUF_X1 U6920 ( .A(n6115), .Z(n6116) );
  NAND2_X1 U6921 ( .A1(n6977), .A2(n7022), .ZN(n5289) );
  INV_X1 U6922 ( .A(n6904), .ZN(n6905) );
  NOR2_X1 U6923 ( .A1(n6188), .A2(n6905), .ZN(n6906) );
  INV_X1 U6924 ( .A(n9980), .ZN(n6973) );
  OR2_X1 U6925 ( .A1(n6975), .A2(n7022), .ZN(n6976) );
  NAND2_X1 U6926 ( .A1(n6979), .A2(n7022), .ZN(n6980) );
  NAND2_X1 U6927 ( .A1(n5249), .A2(n6980), .ZN(n6981) );
  NAND2_X1 U6928 ( .A1(n6994), .A2(n7010), .ZN(n6995) );
  INV_X1 U6929 ( .A(n7034), .ZN(n7011) );
  AOI22_X1 U6930 ( .A1(n7036), .A2(n7035), .B1(n10079), .B2(n7034), .ZN(n7037)
         );
  INV_X1 U6931 ( .A(n6101), .ZN(n6393) );
  INV_X1 U6932 ( .A(n8974), .ZN(n5874) );
  AOI21_X1 U6933 ( .B1(n8810), .B2(n5284), .A(n7089), .ZN(n7090) );
  OAI21_X1 U6934 ( .B1(n6538), .B2(n8100), .A(n6527), .ZN(n6528) );
  OAI21_X1 U6935 ( .B1(n8776), .B2(n4907), .A(n8774), .ZN(n5916) );
  INV_X1 U6936 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7763) );
  NAND2_X1 U6937 ( .A1(n9142), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U6938 ( .A1(n9456), .A2(n9237), .ZN(n7098) );
  INV_X1 U6939 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5642) );
  AND2_X1 U6940 ( .A1(n9463), .A2(n4907), .ZN(n7096) );
  OR2_X1 U6941 ( .A1(n8167), .A2(n8901), .ZN(n8193) );
  NAND2_X1 U6942 ( .A1(n7335), .A2(n6543), .ZN(n6520) );
  NOR2_X1 U6943 ( .A1(n7018), .A2(n7039), .ZN(n7040) );
  INV_X1 U6944 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6040) );
  INV_X1 U6945 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U6946 ( .A1(n9902), .A2(n9730), .ZN(n6351) );
  AND2_X1 U6947 ( .A1(n6847), .A2(n5280), .ZN(n6464) );
  INV_X1 U6948 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5698) );
  INV_X1 U6949 ( .A(n8652), .ZN(n5667) );
  INV_X1 U6950 ( .A(n7138), .ZN(n5988) );
  INV_X1 U6951 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7598) );
  INV_X1 U6952 ( .A(n7144), .ZN(n7145) );
  NAND2_X1 U6953 ( .A1(n4907), .A2(n9382), .ZN(n9238) );
  INV_X1 U6954 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6094) );
  AND2_X1 U6955 ( .A1(n5882), .A2(n5860), .ZN(n5861) );
  NAND2_X1 U6956 ( .A1(n5739), .A2(n5738), .ZN(n5768) );
  INV_X1 U6957 ( .A(n5880), .ZN(n5881) );
  INV_X1 U6958 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5457) );
  OR2_X1 U6959 ( .A1(n5421), .A2(n7224), .ZN(n5376) );
  INV_X1 U6960 ( .A(n9209), .ZN(n9154) );
  NAND2_X1 U6961 ( .A1(n9443), .A2(n5983), .ZN(n10533) );
  AND2_X1 U6962 ( .A1(n8999), .A2(n7162), .ZN(n7973) );
  OR2_X1 U6963 ( .A1(n9219), .A2(n9218), .ZN(n9448) );
  AND2_X1 U6964 ( .A1(n8875), .A2(n8890), .ZN(n8816) );
  AND2_X1 U6965 ( .A1(n5997), .A2(n7314), .ZN(n7150) );
  INV_X1 U6966 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5965) );
  OR2_X1 U6967 ( .A1(n5595), .A2(n9528), .ZN(n5586) );
  AND2_X1 U6968 ( .A1(n7997), .A2(n7995), .ZN(n6552) );
  NAND2_X1 U6969 ( .A1(n6074), .A2(n6073), .ZN(n6101) );
  INV_X1 U6970 ( .A(n6757), .ZN(n6771) );
  AND2_X1 U6971 ( .A1(n6333), .A2(n6341), .ZN(n9931) );
  AND2_X1 U6972 ( .A1(n6302), .A2(n6301), .ZN(n6827) );
  INV_X1 U6973 ( .A(n9701), .ZN(n9687) );
  INV_X1 U6974 ( .A(n6759), .ZN(n6760) );
  OR2_X1 U6975 ( .A1(n10208), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U6976 ( .A1(n10138), .A2(n9737), .ZN(n6441) );
  INV_X1 U6977 ( .A(n10399), .ZN(n10048) );
  NAND2_X1 U6978 ( .A1(n6404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6375) );
  XNOR2_X1 U6979 ( .A(n5614), .B(SI_11_), .ZN(n5615) );
  INV_X1 U6980 ( .A(n6135), .ZN(n6149) );
  INV_X1 U6981 ( .A(n8795), .ZN(n8779) );
  INV_X1 U6982 ( .A(n9333), .ZN(n9305) );
  INV_X1 U6983 ( .A(n8925), .ZN(n8691) );
  INV_X1 U6984 ( .A(n9171), .ZN(n9210) );
  INV_X1 U6985 ( .A(n9144), .ZN(n9126) );
  INV_X1 U6986 ( .A(n9213), .ZN(n9173) );
  INV_X1 U6987 ( .A(n10533), .ZN(n9388) );
  AND2_X1 U6988 ( .A1(n7160), .A2(n7159), .ZN(n7971) );
  AND2_X1 U6989 ( .A1(n9326), .A2(n8950), .ZN(n9343) );
  INV_X1 U6990 ( .A(n9500), .ZN(n9520) );
  NAND2_X1 U6991 ( .A1(n10544), .A2(n8191), .ZN(n10562) );
  OR3_X1 U6992 ( .A1(n8578), .A2(n8595), .A3(n8491), .ZN(n7173) );
  XNOR2_X1 U6993 ( .A(n5970), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9020) );
  NOR2_X1 U6994 ( .A1(n5557), .A2(n5595), .ZN(n8016) );
  XNOR2_X1 U6995 ( .A(n6413), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U6996 ( .A1(n6095), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6085) );
  INV_X1 U6997 ( .A(n9719), .ZN(n9710) );
  INV_X1 U6998 ( .A(n6827), .ZN(n9664) );
  INV_X1 U6999 ( .A(n10269), .ZN(n10293) );
  INV_X1 U7000 ( .A(n10299), .ZN(n10284) );
  OR2_X1 U7001 ( .A1(n10235), .A2(n7409), .ZN(n10269) );
  INV_X1 U7002 ( .A(n9868), .ZN(n10305) );
  INV_X1 U7003 ( .A(n10407), .ZN(n10390) );
  INV_X1 U7004 ( .A(n6893), .ZN(n9971) );
  INV_X1 U7005 ( .A(n10411), .ZN(n10393) );
  NAND2_X1 U7006 ( .A1(n6425), .A2(n10211), .ZN(n7448) );
  INV_X1 U7007 ( .A(n10490), .ZN(n10503) );
  INV_X1 U7008 ( .A(n7448), .ZN(n6782) );
  NAND2_X1 U7009 ( .A1(n6411), .A2(n6410), .ZN(n10208) );
  NOR2_X1 U7010 ( .A1(n7173), .A2(n8452), .ZN(n7281) );
  INV_X1 U7011 ( .A(n8797), .ZN(n8748) );
  INV_X1 U7012 ( .A(n8784), .ZN(n8800) );
  INV_X1 U7013 ( .A(n9215), .ZN(n9159) );
  OR2_X1 U7014 ( .A1(n7505), .A2(n4402), .ZN(n9217) );
  NAND2_X1 U7015 ( .A1(n10578), .A2(n10562), .ZN(n9441) );
  INV_X1 U7016 ( .A(n8200), .ZN(n8247) );
  OR2_X1 U7017 ( .A1(n10573), .A2(n10565), .ZN(n9500) );
  OR2_X1 U7018 ( .A1(n10573), .A2(n10567), .ZN(n9524) );
  AND2_X1 U7019 ( .A1(n7154), .A2(n7153), .ZN(n10573) );
  AND2_X1 U7020 ( .A1(n7173), .A2(n7317), .ZN(n7314) );
  INV_X1 U7021 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7329) );
  AND2_X1 U7022 ( .A1(n7327), .A2(n7388), .ZN(n10233) );
  INV_X1 U7023 ( .A(n10097), .ZN(n9955) );
  INV_X1 U7024 ( .A(n9721), .ZN(n9708) );
  INV_X1 U7025 ( .A(n10108), .ZN(n9988) );
  AND2_X1 U7026 ( .A1(n6761), .A2(n10382), .ZN(n9725) );
  INV_X1 U7027 ( .A(P1_U3973), .ZN(n9738) );
  OR2_X1 U7028 ( .A1(n10235), .A2(n10230), .ZN(n10299) );
  INV_X1 U7029 ( .A(n10233), .ZN(n10308) );
  AND2_X1 U7030 ( .A1(n10315), .A2(n10314), .ZN(n10498) );
  OR2_X1 U7031 ( .A1(n10402), .A2(n8091), .ZN(n10412) );
  INV_X1 U7032 ( .A(n10080), .ZN(n10145) );
  INV_X2 U7033 ( .A(n10526), .ZN(n10528) );
  NAND2_X1 U7034 ( .A1(n10509), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6784) );
  INV_X1 U7035 ( .A(n10160), .ZN(n10205) );
  OR2_X1 U7036 ( .A1(n6783), .A2(n6782), .ZN(n10509) );
  INV_X2 U7037 ( .A(n10509), .ZN(n10510) );
  INV_X1 U7038 ( .A(n10423), .ZN(n10424) );
  INV_X1 U7039 ( .A(n7047), .ZN(n8456) );
  INV_X1 U7040 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n8129) );
  AND2_X2 U7041 ( .A1(n7281), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3893) );
  OR4_X1 U7042 ( .A1(n7289), .A2(n7288), .A3(n7287), .A4(n7286), .ZN(P2_U3194)
         );
  AND2_X2 U7043 ( .A1(n7172), .A2(n7323), .ZN(P1_U3973) );
  XNOR2_X2 U7044 ( .A(n5297), .B(n5296), .ZN(n9198) );
  NAND2_X1 U7045 ( .A1(n5299), .A2(n5298), .ZN(n5300) );
  NOR2_X1 U7046 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5305) );
  NOR2_X1 U7047 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5304) );
  NOR2_X1 U7048 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5303) );
  NOR2_X1 U7049 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5306) );
  NAND2_X1 U7050 ( .A1(n5968), .A2(n5312), .ZN(n5310) );
  INV_X1 U7051 ( .A(P2_B_REG_SCAN_IN), .ZN(n5317) );
  INV_X1 U7052 ( .A(n8595), .ZN(n5322) );
  NAND3_X1 U7053 ( .A1(n5950), .A2(n5324), .A3(P2_B_REG_SCAN_IN), .ZN(n5319)
         );
  NAND2_X1 U7054 ( .A1(n5317), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U7055 ( .A1(n5319), .A2(n5318), .ZN(n5320) );
  NAND2_X1 U7056 ( .A1(n5325), .A2(n5320), .ZN(n5321) );
  INV_X1 U7057 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7318) );
  NAND2_X1 U7058 ( .A1(n7312), .A2(n7318), .ZN(n5327) );
  NAND2_X1 U7059 ( .A1(n5325), .A2(n5324), .ZN(n5949) );
  NAND2_X1 U7060 ( .A1(n5949), .A2(n5326), .ZN(n8491) );
  NAND2_X1 U7061 ( .A1(n8491), .A2(n8595), .ZN(n7315) );
  NOR2_X4 U7062 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8370) );
  INV_X1 U7063 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5332) );
  INV_X1 U7064 ( .A(SI_1_), .ZN(n5333) );
  OAI21_X1 U7065 ( .B1(n5487), .B2(P1_DATAO_REG_0__SCAN_IN), .A(n5336), .ZN(
        n5338) );
  NAND2_X1 U7066 ( .A1(n5337), .A2(n5338), .ZN(n5339) );
  INV_X1 U7067 ( .A(n5338), .ZN(n5402) );
  XNOR2_X2 U7068 ( .A(n5341), .B(n7598), .ZN(n5378) );
  XNOR2_X2 U7069 ( .A(n5344), .B(n5343), .ZN(n7278) );
  NAND2_X1 U7070 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5345) );
  XNOR2_X2 U7071 ( .A(n5345), .B(n5141), .ZN(n7347) );
  NAND3_X1 U7072 ( .A1(n7278), .A2(n5378), .A3(n7347), .ZN(n5350) );
  INV_X1 U7073 ( .A(n7278), .ZN(n9017) );
  INV_X1 U7074 ( .A(n7291), .ZN(n5346) );
  NAND2_X1 U7075 ( .A1(n5346), .A2(n7290), .ZN(n5347) );
  NAND3_X1 U7076 ( .A1(n9017), .A2(n5348), .A3(n5347), .ZN(n5349) );
  INV_X1 U7077 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5351) );
  INV_X1 U7078 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5360) );
  AOI22_X1 U7079 ( .A1(n5360), .A2(P2_REG2_REG_1__SCAN_IN), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(P2_REG0_REG_1__SCAN_IN), .ZN(n5356) );
  INV_X1 U7080 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U7081 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG2_REG_1__SCAN_IN), 
        .ZN(n5352) );
  OAI21_X1 U7082 ( .B1(n5353), .B2(P2_IR_REG_30__SCAN_IN), .A(n5352), .ZN(
        n5354) );
  NAND2_X1 U7083 ( .A1(n5370), .A2(n5354), .ZN(n5355) );
  OAI21_X1 U7084 ( .B1(n5370), .B2(n5356), .A(n5355), .ZN(n5359) );
  NAND2_X1 U7086 ( .A1(n5359), .A2(n9540), .ZN(n5369) );
  AOI22_X1 U7087 ( .A1(n5360), .A2(P2_REG3_REG_1__SCAN_IN), .B1(
        P2_REG1_REG_1__SCAN_IN), .B2(P2_IR_REG_30__SCAN_IN), .ZN(n5365) );
  INV_X1 U7088 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U7089 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG3_REG_1__SCAN_IN), 
        .ZN(n5361) );
  OAI21_X1 U7090 ( .B1(n5362), .B2(P2_IR_REG_30__SCAN_IN), .A(n5361), .ZN(
        n5363) );
  NAND2_X1 U7091 ( .A1(n5370), .A2(n5363), .ZN(n5364) );
  OAI21_X1 U7092 ( .B1(n5370), .B2(n5365), .A(n5364), .ZN(n5367) );
  NAND2_X1 U7093 ( .A1(n5367), .A2(n5374), .ZN(n5368) );
  INV_X1 U7094 ( .A(n7054), .ZN(n10538) );
  INV_X1 U7095 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U7096 ( .A1(n9534), .A2(n5372), .ZN(n5421) );
  INV_X1 U7097 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7224) );
  NAND2_X2 U7098 ( .A1(n5373), .A2(n5374), .ZN(n5423) );
  INV_X1 U7099 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7223) );
  NAND2_X1 U7100 ( .A1(n5660), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U7101 ( .A1(n7290), .A2(SI_0_), .ZN(n5377) );
  XNOR2_X1 U7102 ( .A(n5377), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9549) );
  INV_X1 U7103 ( .A(n7982), .ZN(n7814) );
  NAND2_X1 U7104 ( .A1(n7545), .A2(n7546), .ZN(n5382) );
  NAND2_X1 U7105 ( .A1(n5382), .A2(n5381), .ZN(n7539) );
  NAND2_X1 U7106 ( .A1(n5383), .A2(n5403), .ZN(n5388) );
  INV_X1 U7107 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7294) );
  INV_X1 U7108 ( .A(SI_2_), .ZN(n5384) );
  NAND2_X1 U7109 ( .A1(n5385), .A2(n5384), .ZN(n5404) );
  INV_X1 U7110 ( .A(n5385), .ZN(n5386) );
  NAND2_X1 U7111 ( .A1(n5386), .A2(SI_2_), .ZN(n5406) );
  NAND2_X1 U7112 ( .A1(n5404), .A2(n5406), .ZN(n5387) );
  NAND2_X1 U7113 ( .A1(n5656), .A2(n6137), .ZN(n5391) );
  OR2_X1 U7114 ( .A1(n7176), .A2(n7292), .ZN(n5389) );
  INV_X1 U7115 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5392) );
  OR2_X2 U7116 ( .A1(n8401), .A2(n5392), .ZN(n5396) );
  INV_X1 U7117 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10549) );
  OR2_X1 U7118 ( .A1(n5421), .A2(n10549), .ZN(n5395) );
  NAND2_X1 U7119 ( .A1(n5660), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5394) );
  INV_X1 U7120 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7196) );
  OR2_X1 U7121 ( .A1(n5423), .A2(n7196), .ZN(n5393) );
  NAND4_X2 U7122 ( .A1(n5396), .A2(n5395), .A3(n5394), .A4(n5393), .ZN(n7057)
         );
  XNOR2_X1 U7123 ( .A(n5397), .B(n7057), .ZN(n7540) );
  NAND2_X1 U7124 ( .A1(n7539), .A2(n7540), .ZN(n5399) );
  INV_X1 U7125 ( .A(n7057), .ZN(n7901) );
  NAND2_X1 U7126 ( .A1(n5397), .A2(n7901), .ZN(n5398) );
  NAND2_X1 U7127 ( .A1(n5399), .A2(n5398), .ZN(n7818) );
  INV_X1 U7128 ( .A(n7818), .ZN(n5431) );
  INV_X1 U7129 ( .A(n5656), .ZN(n5636) );
  INV_X1 U7130 ( .A(n5403), .ZN(n5405) );
  NAND2_X1 U7131 ( .A1(n5405), .A2(n5404), .ZN(n5407) );
  NAND3_X1 U7132 ( .A1(n5408), .A2(n5407), .A3(n5406), .ZN(n5415) );
  INV_X1 U7133 ( .A(n5415), .ZN(n5412) );
  INV_X1 U7134 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5409) );
  OAI21_X1 U7135 ( .B1(n5411), .B2(SI_3_), .A(n5434), .ZN(n5413) );
  NAND2_X1 U7136 ( .A1(n5412), .A2(n5413), .ZN(n5416) );
  INV_X1 U7137 ( .A(n5413), .ZN(n5414) );
  NAND2_X1 U7138 ( .A1(n5415), .A2(n5414), .ZN(n5474) );
  NAND2_X1 U7139 ( .A1(n5416), .A2(n5474), .ZN(n7295) );
  NAND2_X1 U7140 ( .A1(n5906), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U7141 ( .A1(n5439), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5418) );
  XNOR2_X1 U7142 ( .A(n5418), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7234) );
  NAND2_X1 U7143 ( .A1(n5756), .A2(n7234), .ZN(n5419) );
  OAI211_X1 U7144 ( .C1(n5636), .C2(n7295), .A(n5420), .B(n5419), .ZN(n7060)
         );
  XNOR2_X1 U7145 ( .A(n5536), .B(n7060), .ZN(n5432) );
  INV_X1 U7146 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5422) );
  INV_X1 U7147 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5424) );
  OR2_X1 U7148 ( .A1(n5423), .A2(n5424), .ZN(n5427) );
  INV_X1 U7149 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5425) );
  OR2_X1 U7150 ( .A1(n8401), .A2(n5425), .ZN(n5426) );
  XNOR2_X1 U7151 ( .A(n5432), .B(n9035), .ZN(n7817) );
  NAND2_X1 U7152 ( .A1(n5432), .A2(n9035), .ZN(n5433) );
  INV_X1 U7153 ( .A(SI_4_), .ZN(n5435) );
  NAND2_X1 U7154 ( .A1(n5436), .A2(n5435), .ZN(n5475) );
  NAND2_X1 U7155 ( .A1(n5437), .A2(SI_4_), .ZN(n5472) );
  AND2_X1 U7156 ( .A1(n5475), .A2(n5472), .ZN(n5438) );
  NAND2_X1 U7157 ( .A1(n5906), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5447) );
  INV_X1 U7158 ( .A(n5439), .ZN(n5441) );
  INV_X1 U7159 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5440) );
  INV_X1 U7160 ( .A(n5445), .ZN(n5442) );
  NAND2_X1 U7161 ( .A1(n5442), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5443) );
  MUX2_X1 U7162 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5443), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5446) );
  INV_X1 U7163 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U7164 ( .A1(n5445), .A2(n5444), .ZN(n5466) );
  INV_X1 U7165 ( .A(n7431), .ZN(n7232) );
  NAND2_X1 U7166 ( .A1(n7135), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5453) );
  INV_X1 U7167 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5448) );
  OR2_X1 U7168 ( .A1(n8401), .A2(n5448), .ZN(n5452) );
  INV_X1 U7169 ( .A(n5458), .ZN(n5459) );
  NAND2_X1 U7170 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5449) );
  AND2_X1 U7171 ( .A1(n5459), .A2(n5449), .ZN(n8031) );
  OR2_X1 U7172 ( .A1(n5646), .A2(n8031), .ZN(n5451) );
  INV_X1 U7173 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7205) );
  NAND4_X2 U7174 ( .A1(n5453), .A2(n5452), .A3(n5451), .A4(n5450), .ZN(n7110)
         );
  INV_X1 U7175 ( .A(n5454), .ZN(n5455) );
  OR2_X1 U7176 ( .A1(n7110), .A2(n5455), .ZN(n5456) );
  NAND2_X1 U7177 ( .A1(n4408), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5465) );
  INV_X1 U7178 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n8144) );
  OR2_X1 U7179 ( .A1(n5421), .A2(n8144), .ZN(n5464) );
  NAND2_X1 U7180 ( .A1(n5459), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5460) );
  AND2_X1 U7181 ( .A1(n5495), .A2(n5460), .ZN(n8145) );
  OR2_X1 U7182 ( .A1(n5646), .A2(n8145), .ZN(n5463) );
  INV_X1 U7183 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U7184 ( .A1(n5466), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5467) );
  INV_X1 U7185 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7611) );
  XNOR2_X1 U7186 ( .A(n5467), .B(n7611), .ZN(n7296) );
  OAI22_X1 U7187 ( .A1(n5720), .A2(n4580), .B1(n4746), .B2(n7296), .ZN(n5479)
         );
  AND2_X1 U7188 ( .A1(n5476), .A2(n5472), .ZN(n5470) );
  NAND2_X1 U7189 ( .A1(n5471), .A2(n5470), .ZN(n5477) );
  AND2_X1 U7190 ( .A1(n5434), .A2(n5472), .ZN(n5473) );
  NAND2_X1 U7191 ( .A1(n5508), .A2(n5506), .ZN(n5486) );
  NAND2_X1 U7192 ( .A1(n5477), .A2(n5486), .ZN(n7297) );
  NOR2_X1 U7193 ( .A1(n7297), .A2(n5636), .ZN(n5478) );
  OR2_X2 U7194 ( .A1(n5479), .A2(n5478), .ZN(n8147) );
  XNOR2_X1 U7195 ( .A(n5536), .B(n8147), .ZN(n5480) );
  XNOR2_X1 U7196 ( .A(n7947), .B(n5480), .ZN(n7987) );
  INV_X1 U7197 ( .A(n5480), .ZN(n5481) );
  NAND2_X1 U7198 ( .A1(n5481), .A2(n7947), .ZN(n5482) );
  NAND2_X1 U7199 ( .A1(n5483), .A2(n5482), .ZN(n8054) );
  INV_X2 U7200 ( .A(n5720), .ZN(n5757) );
  NAND2_X1 U7201 ( .A1(n5484), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5485) );
  XNOR2_X1 U7202 ( .A(n5485), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7472) );
  AOI22_X1 U7203 ( .A1(n5757), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5756), .B2(
        n7472), .ZN(n5494) );
  NAND2_X1 U7204 ( .A1(n5486), .A2(n5509), .ZN(n5492) );
  INV_X1 U7205 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7304) );
  INV_X1 U7206 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7306) );
  MUX2_X1 U7207 ( .A(n7304), .B(n7306), .S(n4414), .Z(n5489) );
  INV_X1 U7208 ( .A(SI_6_), .ZN(n5488) );
  NAND2_X1 U7209 ( .A1(n5489), .A2(n5488), .ZN(n5512) );
  INV_X1 U7210 ( .A(n5489), .ZN(n5490) );
  NAND2_X1 U7211 ( .A1(n5490), .A2(SI_6_), .ZN(n5510) );
  NAND2_X1 U7212 ( .A1(n5512), .A2(n5510), .ZN(n5491) );
  XNOR2_X1 U7213 ( .A(n5492), .B(n5491), .ZN(n7302) );
  NAND2_X1 U7214 ( .A1(n7302), .A2(n5624), .ZN(n5493) );
  XNOR2_X1 U7215 ( .A(n8059), .B(n5536), .ZN(n5503) );
  NAND2_X1 U7216 ( .A1(n5987), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5500) );
  INV_X1 U7217 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n8067) );
  OR2_X1 U7218 ( .A1(n5421), .A2(n8067), .ZN(n5499) );
  NAND2_X1 U7219 ( .A1(n5495), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5496) );
  AND2_X1 U7220 ( .A1(n5523), .A2(n5496), .ZN(n8068) );
  OR2_X1 U7221 ( .A1(n5646), .A2(n8068), .ZN(n5498) );
  INV_X1 U7222 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7242) );
  OR2_X1 U7223 ( .A1(n5423), .A2(n7242), .ZN(n5497) );
  XNOR2_X1 U7224 ( .A(n5503), .B(n7990), .ZN(n8055) );
  INV_X1 U7225 ( .A(n8055), .ZN(n5501) );
  OR2_X1 U7226 ( .A1(n5503), .A2(n7990), .ZN(n5504) );
  INV_X1 U7227 ( .A(n4399), .ZN(n5520) );
  NAND2_X1 U7228 ( .A1(n5302), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5505) );
  XNOR2_X1 U7229 ( .A(n5505), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7862) );
  AOI22_X1 U7230 ( .A1(n5757), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5756), .B2(
        n7862), .ZN(n5519) );
  INV_X1 U7231 ( .A(n5509), .ZN(n5513) );
  INV_X1 U7232 ( .A(n5510), .ZN(n5511) );
  AND2_X1 U7233 ( .A1(n5532), .A2(n5517), .ZN(n7301) );
  NAND2_X1 U7234 ( .A1(n7301), .A2(n5624), .ZN(n5518) );
  NAND2_X1 U7235 ( .A1(n5519), .A2(n5518), .ZN(n8200) );
  XNOR2_X1 U7236 ( .A(n5536), .B(n8200), .ZN(n5529) );
  NAND2_X1 U7237 ( .A1(n7135), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5528) );
  INV_X1 U7238 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8245) );
  OR2_X1 U7239 ( .A1(n5423), .A2(n8245), .ZN(n5527) );
  NAND2_X1 U7240 ( .A1(n5523), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5524) );
  AND2_X1 U7241 ( .A1(n5537), .A2(n5524), .ZN(n8221) );
  OR2_X1 U7242 ( .A1(n5646), .A2(n8221), .ZN(n5526) );
  INV_X1 U7243 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7648) );
  OR2_X1 U7244 ( .A1(n8401), .A2(n7648), .ZN(n5525) );
  INV_X1 U7245 ( .A(n9033), .ZN(n8058) );
  XNOR2_X1 U7246 ( .A(n5529), .B(n8058), .ZN(n8203) );
  INV_X1 U7247 ( .A(n5529), .ZN(n5530) );
  MUX2_X1 U7248 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n4414), .Z(n5546) );
  NAND2_X1 U7249 ( .A1(n7308), .A2(n5624), .ZN(n5535) );
  NOR2_X1 U7250 ( .A1(n5302), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5553) );
  OR2_X1 U7251 ( .A1(n5553), .A2(n9528), .ZN(n5533) );
  XNOR2_X1 U7252 ( .A(n5533), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7935) );
  AOI22_X1 U7253 ( .A1(n5757), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5756), .B2(
        n7935), .ZN(n5534) );
  XNOR2_X1 U7254 ( .A(n7070), .B(n5536), .ZN(n5543) );
  NAND2_X1 U7255 ( .A1(n7135), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5542) );
  INV_X1 U7256 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8217) );
  OR2_X1 U7257 ( .A1(n5423), .A2(n8217), .ZN(n5541) );
  NAND2_X1 U7258 ( .A1(n5537), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5538) );
  AND2_X1 U7259 ( .A1(n5560), .A2(n5538), .ZN(n8263) );
  OR2_X1 U7260 ( .A1(n5646), .A2(n8263), .ZN(n5540) );
  INV_X1 U7261 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7693) );
  OR2_X1 U7262 ( .A1(n8401), .A2(n7693), .ZN(n5539) );
  NAND4_X1 U7263 ( .A1(n5542), .A2(n5541), .A3(n5540), .A4(n5539), .ZN(n9032)
         );
  XNOR2_X1 U7264 ( .A(n5543), .B(n9032), .ZN(n8260) );
  INV_X1 U7265 ( .A(n9032), .ZN(n8205) );
  NAND2_X1 U7266 ( .A1(n5543), .A2(n8205), .ZN(n5544) );
  INV_X1 U7267 ( .A(n5546), .ZN(n5548) );
  INV_X1 U7268 ( .A(SI_8_), .ZN(n5547) );
  NAND2_X1 U7269 ( .A1(n5548), .A2(n5547), .ZN(n5549) );
  XNOR2_X1 U7270 ( .A(n5575), .B(SI_9_), .ZN(n5578) );
  NAND2_X1 U7271 ( .A1(n7328), .A2(n5624), .ZN(n5559) );
  INV_X1 U7272 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5552) );
  NOR2_X1 U7273 ( .A1(n5556), .A2(n9528), .ZN(n5554) );
  MUX2_X1 U7274 ( .A(n9528), .B(n5554), .S(P2_IR_REG_9__SCAN_IN), .Z(n5557) );
  INV_X1 U7275 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5555) );
  AOI22_X1 U7276 ( .A1(n5757), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5756), .B2(
        n8016), .ZN(n5558) );
  NAND2_X2 U7277 ( .A1(n5559), .A2(n5558), .ZN(n8611) );
  XNOR2_X1 U7278 ( .A(n8611), .B(n5536), .ZN(n5567) );
  NAND2_X1 U7279 ( .A1(n4408), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5565) );
  INV_X1 U7280 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7254) );
  OR2_X1 U7281 ( .A1(n8403), .A2(n7254), .ZN(n5564) );
  NAND2_X1 U7282 ( .A1(n5560), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5561) );
  AND2_X1 U7283 ( .A1(n5569), .A2(n5561), .ZN(n8609) );
  OR2_X1 U7284 ( .A1(n5646), .A2(n8609), .ZN(n5563) );
  INV_X1 U7285 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8348) );
  OR2_X1 U7286 ( .A1(n7138), .A2(n8348), .ZN(n5562) );
  XNOR2_X1 U7287 ( .A(n5567), .B(n9031), .ZN(n8338) );
  INV_X1 U7288 ( .A(n8338), .ZN(n5566) );
  NAND2_X1 U7289 ( .A1(n5567), .A2(n9031), .ZN(n5568) );
  NAND2_X1 U7290 ( .A1(n4408), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5574) );
  INV_X1 U7291 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8375) );
  OR2_X1 U7292 ( .A1(n5421), .A2(n8375), .ZN(n5573) );
  NAND2_X1 U7293 ( .A1(n5569), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5570) );
  AND2_X1 U7294 ( .A1(n5599), .A2(n5570), .ZN(n8483) );
  OR2_X1 U7295 ( .A1(n5646), .A2(n8483), .ZN(n5572) );
  INV_X1 U7296 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8397) );
  OR2_X1 U7297 ( .A1(n7138), .A2(n8397), .ZN(n5571) );
  NAND4_X1 U7298 ( .A1(n5574), .A2(n5573), .A3(n5572), .A4(n5571), .ZN(n9030)
         );
  INV_X1 U7299 ( .A(n5575), .ZN(n5576) );
  NOR2_X1 U7300 ( .A1(n5576), .A2(SI_9_), .ZN(n5577) );
  NAND2_X1 U7301 ( .A1(n5580), .A2(SI_10_), .ZN(n5592) );
  INV_X1 U7302 ( .A(n5580), .ZN(n5582) );
  INV_X1 U7303 ( .A(SI_10_), .ZN(n5581) );
  NAND2_X1 U7304 ( .A1(n5582), .A2(n5581), .ZN(n5583) );
  NAND2_X1 U7305 ( .A1(n5584), .A2(n4888), .ZN(n5585) );
  XNOR2_X1 U7306 ( .A(n5586), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7259) );
  AOI22_X1 U7307 ( .A1(n5757), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5756), .B2(
        n7259), .ZN(n5587) );
  XNOR2_X1 U7308 ( .A(n8485), .B(n4411), .ZN(n8479) );
  NAND2_X1 U7309 ( .A1(n8477), .A2(n8479), .ZN(n5591) );
  INV_X1 U7310 ( .A(n5589), .ZN(n5590) );
  NAND2_X1 U7311 ( .A1(n5590), .A2(n9030), .ZN(n8476) );
  XNOR2_X1 U7312 ( .A(n5616), .B(n5615), .ZN(n7338) );
  NAND2_X1 U7313 ( .A1(n7338), .A2(n5624), .ZN(n5598) );
  INV_X1 U7314 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7315 ( .A1(n5595), .A2(n5594), .ZN(n5625) );
  NAND2_X1 U7316 ( .A1(n5625), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5596) );
  XNOR2_X1 U7317 ( .A(n5596), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7264) );
  AOI22_X1 U7318 ( .A1(n5757), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5756), .B2(
        n7264), .ZN(n5597) );
  NAND2_X1 U7319 ( .A1(n4408), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5604) );
  INV_X1 U7320 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8384) );
  OR2_X1 U7321 ( .A1(n8403), .A2(n8384), .ZN(n5603) );
  NAND2_X1 U7322 ( .A1(n5599), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5600) );
  AND2_X1 U7323 ( .A1(n5608), .A2(n5600), .ZN(n8536) );
  OR2_X1 U7324 ( .A1(n5646), .A2(n8536), .ZN(n5602) );
  INV_X1 U7325 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8380) );
  OR2_X1 U7326 ( .A1(n7138), .A2(n8380), .ZN(n5601) );
  NAND4_X1 U7327 ( .A1(n5604), .A2(n5603), .A3(n5602), .A4(n5601), .ZN(n9029)
         );
  OR2_X1 U7328 ( .A1(n8530), .A2(n9029), .ZN(n7079) );
  INV_X1 U7329 ( .A(n7079), .ZN(n5605) );
  AND2_X1 U7330 ( .A1(n8530), .A2(n9029), .ZN(n7080) );
  XNOR2_X1 U7331 ( .A(n8823), .B(n5760), .ZN(n8532) );
  INV_X1 U7332 ( .A(n8532), .ZN(n5606) );
  NAND2_X1 U7333 ( .A1(n5606), .A2(n9029), .ZN(n5607) );
  NAND2_X1 U7334 ( .A1(n4408), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5613) );
  INV_X1 U7335 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9037) );
  OR2_X1 U7336 ( .A1(n5421), .A2(n9037), .ZN(n5612) );
  NAND2_X1 U7337 ( .A1(n5608), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5609) );
  AND2_X1 U7338 ( .A1(n5644), .A2(n5609), .ZN(n8693) );
  OR2_X1 U7339 ( .A1(n5646), .A2(n8693), .ZN(n5611) );
  INV_X1 U7340 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8443) );
  OR2_X1 U7341 ( .A1(n7138), .A2(n8443), .ZN(n5610) );
  NAND4_X1 U7342 ( .A1(n5613), .A2(n5612), .A3(n5611), .A4(n5610), .ZN(n9028)
         );
  INV_X1 U7343 ( .A(n5617), .ZN(n5619) );
  INV_X1 U7344 ( .A(SI_12_), .ZN(n5618) );
  NAND2_X1 U7345 ( .A1(n5619), .A2(n5618), .ZN(n5620) );
  NAND2_X1 U7346 ( .A1(n5622), .A2(n5621), .ZN(n5623) );
  AND2_X1 U7347 ( .A1(n5623), .A2(n5629), .ZN(n7342) );
  NAND2_X1 U7348 ( .A1(n7342), .A2(n5624), .ZN(n5628) );
  OAI21_X1 U7349 ( .B1(n5625), .B2(P2_IR_REG_11__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5626) );
  XNOR2_X1 U7350 ( .A(n5626), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9038) );
  AOI22_X1 U7351 ( .A1(n5757), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9038), .B2(
        n5756), .ZN(n5627) );
  XNOR2_X1 U7352 ( .A(n8921), .B(n5536), .ZN(n8686) );
  NAND2_X1 U7353 ( .A1(n5630), .A2(SI_13_), .ZN(n5654) );
  INV_X1 U7354 ( .A(n5630), .ZN(n5632) );
  INV_X1 U7355 ( .A(SI_13_), .ZN(n5631) );
  NAND2_X1 U7356 ( .A1(n5632), .A2(n5631), .ZN(n5633) );
  NAND2_X1 U7357 ( .A1(n5654), .A2(n5633), .ZN(n5634) );
  INV_X1 U7358 ( .A(n5637), .ZN(n5638) );
  NAND2_X1 U7359 ( .A1(n5638), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5639) );
  XNOR2_X1 U7360 ( .A(n5639), .B(n7626), .ZN(n9084) );
  INV_X1 U7361 ( .A(n9084), .ZN(n9060) );
  AOI22_X1 U7362 ( .A1(n5757), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5756), .B2(
        n9060), .ZN(n5640) );
  XNOR2_X1 U7363 ( .A(n8926), .B(n5400), .ZN(n5651) );
  NAND2_X1 U7364 ( .A1(n4408), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5650) );
  INV_X1 U7365 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9045) );
  OR2_X1 U7366 ( .A1(n8403), .A2(n9045), .ZN(n5649) );
  NAND2_X1 U7367 ( .A1(n5644), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5645) );
  AND2_X1 U7368 ( .A1(n5661), .A2(n5645), .ZN(n8749) );
  OR2_X1 U7369 ( .A1(n5646), .A2(n8749), .ZN(n5648) );
  INV_X1 U7370 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9044) );
  OR2_X1 U7371 ( .A1(n7138), .A2(n9044), .ZN(n5647) );
  XNOR2_X1 U7372 ( .A(n5651), .B(n8691), .ZN(n8744) );
  INV_X1 U7373 ( .A(n5651), .ZN(n5652) );
  NAND2_X1 U7374 ( .A1(n5652), .A2(n8691), .ZN(n5653) );
  XNOR2_X1 U7375 ( .A(n5672), .B(SI_14_), .ZN(n5655) );
  XNOR2_X1 U7376 ( .A(n5671), .B(n5655), .ZN(n7825) );
  NAND2_X1 U7377 ( .A1(n7825), .A2(n5624), .ZN(n5659) );
  NAND2_X1 U7378 ( .A1(n5657), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5701) );
  XNOR2_X1 U7379 ( .A(n5701), .B(P2_IR_REG_14__SCAN_IN), .ZN(n9102) );
  AOI22_X1 U7380 ( .A1(n5757), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5756), .B2(
        n9102), .ZN(n5658) );
  XNOR2_X1 U7381 ( .A(n8934), .B(n5520), .ZN(n5688) );
  NAND2_X1 U7382 ( .A1(n5661), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7383 ( .A1(n5682), .A2(n5662), .ZN(n8655) );
  NAND2_X1 U7384 ( .A1(n5986), .A2(n8655), .ZN(n5666) );
  INV_X1 U7385 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9071) );
  OR2_X1 U7386 ( .A1(n5421), .A2(n9071), .ZN(n5665) );
  INV_X1 U7387 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9101) );
  OR2_X1 U7388 ( .A1(n7138), .A2(n9101), .ZN(n5664) );
  INV_X1 U7389 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8547) );
  OR2_X1 U7390 ( .A1(n8401), .A2(n8547), .ZN(n5663) );
  NAND4_X1 U7391 ( .A1(n5666), .A2(n5665), .A3(n5664), .A4(n5663), .ZN(n9383)
         );
  XNOR2_X1 U7392 ( .A(n5688), .B(n9383), .ZN(n8652) );
  INV_X1 U7393 ( .A(n5672), .ZN(n5669) );
  INV_X1 U7394 ( .A(SI_14_), .ZN(n5668) );
  NAND2_X1 U7395 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  NAND2_X1 U7396 ( .A1(n5672), .A2(SI_14_), .ZN(n5673) );
  XNOR2_X1 U7397 ( .A(n5693), .B(SI_15_), .ZN(n5674) );
  XNOR2_X1 U7398 ( .A(n5697), .B(n5674), .ZN(n7908) );
  NAND2_X1 U7399 ( .A1(n7908), .A2(n5624), .ZN(n5679) );
  NAND2_X1 U7400 ( .A1(n5701), .A2(n5675), .ZN(n5676) );
  NAND2_X1 U7401 ( .A1(n5676), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5677) );
  XNOR2_X1 U7402 ( .A(n5677), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9115) );
  AOI22_X1 U7403 ( .A1(n5757), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5756), .B2(
        n9115), .ZN(n5678) );
  XNOR2_X1 U7404 ( .A(n9521), .B(n5520), .ZN(n5691) );
  NAND2_X1 U7405 ( .A1(n5682), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7406 ( .A1(n5704), .A2(n5683), .ZN(n9387) );
  NAND2_X1 U7407 ( .A1(n9387), .A2(n5986), .ZN(n5687) );
  NAND2_X1 U7408 ( .A1(n4408), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7409 ( .A1(n7135), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5685) );
  INV_X1 U7410 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9437) );
  OR2_X1 U7411 ( .A1(n7138), .A2(n9437), .ZN(n5684) );
  XNOR2_X1 U7412 ( .A(n5691), .B(n8708), .ZN(n8791) );
  INV_X1 U7413 ( .A(n5688), .ZN(n5689) );
  INV_X1 U7414 ( .A(n9383), .ZN(n8933) );
  NAND2_X1 U7415 ( .A1(n5689), .A2(n8933), .ZN(n8788) );
  AND2_X1 U7416 ( .A1(n8791), .A2(n8788), .ZN(n5690) );
  NAND2_X1 U7417 ( .A1(n8650), .A2(n5690), .ZN(n8789) );
  NAND2_X1 U7418 ( .A1(n5691), .A2(n9370), .ZN(n5692) );
  AND2_X1 U7419 ( .A1(n5693), .A2(SI_15_), .ZN(n5696) );
  INV_X1 U7420 ( .A(n5693), .ZN(n5694) );
  NAND2_X1 U7421 ( .A1(n5694), .A2(n7672), .ZN(n5695) );
  XNOR2_X1 U7422 ( .A(n5713), .B(SI_16_), .ZN(n5699) );
  XNOR2_X1 U7423 ( .A(n5715), .B(n5699), .ZN(n7985) );
  NAND2_X1 U7424 ( .A1(n7985), .A2(n5624), .ZN(n5703) );
  OAI21_X1 U7425 ( .B1(P2_IR_REG_14__SCAN_IN), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7426 ( .A1(n5701), .A2(n5700), .ZN(n5721) );
  XNOR2_X1 U7427 ( .A(n5721), .B(n4947), .ZN(n9148) );
  AOI22_X1 U7428 ( .A1(n5757), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5756), .B2(
        n9148), .ZN(n5702) );
  XNOR2_X1 U7429 ( .A(n9514), .B(n5520), .ZN(n5711) );
  NAND2_X1 U7430 ( .A1(n5704), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U7431 ( .A1(n5725), .A2(n5705), .ZN(n9374) );
  NAND2_X1 U7432 ( .A1(n9374), .A2(n5986), .ZN(n5710) );
  INV_X1 U7433 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9513) );
  OR2_X1 U7434 ( .A1(n8401), .A2(n9513), .ZN(n5707) );
  INV_X1 U7435 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9373) );
  OR2_X1 U7436 ( .A1(n8403), .A2(n9373), .ZN(n5706) );
  AND2_X1 U7437 ( .A1(n5707), .A2(n5706), .ZN(n5709) );
  NAND2_X1 U7438 ( .A1(n5988), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5708) );
  XNOR2_X1 U7439 ( .A(n5711), .B(n9359), .ZN(n8705) );
  INV_X1 U7440 ( .A(n9359), .ZN(n9381) );
  NAND2_X1 U7441 ( .A1(n5711), .A2(n9381), .ZN(n5712) );
  INV_X1 U7442 ( .A(SI_17_), .ZN(n5716) );
  NAND2_X1 U7443 ( .A1(n5717), .A2(n5716), .ZN(n5733) );
  INV_X1 U7444 ( .A(n5717), .ZN(n5718) );
  NAND2_X1 U7445 ( .A1(n5718), .A2(SI_17_), .ZN(n5719) );
  NAND2_X1 U7446 ( .A1(n8127), .A2(n5624), .ZN(n5724) );
  OAI21_X1 U7447 ( .B1(n5721), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5722) );
  AOI22_X1 U7448 ( .A1(n5757), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5756), .B2(
        n9176), .ZN(n5723) );
  XNOR2_X1 U7449 ( .A(n9363), .B(n5520), .ZN(n5729) );
  INV_X1 U7450 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U7451 ( .A1(n5725), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U7452 ( .A1(n5761), .A2(n5726), .ZN(n9360) );
  NAND2_X1 U7453 ( .A1(n9360), .A2(n5986), .ZN(n5728) );
  AOI22_X1 U7454 ( .A1(n4408), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n7135), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n5727) );
  OAI211_X1 U7455 ( .C1(n7138), .C2(n9168), .A(n5728), .B(n5727), .ZN(n9371)
         );
  INV_X1 U7456 ( .A(n9371), .ZN(n8769) );
  NAND2_X1 U7457 ( .A1(n5729), .A2(n8769), .ZN(n8665) );
  INV_X1 U7458 ( .A(n5729), .ZN(n5730) );
  NAND2_X1 U7459 ( .A1(n5730), .A2(n9371), .ZN(n5731) );
  NAND2_X1 U7460 ( .A1(n8665), .A2(n5731), .ZN(n8716) );
  INV_X1 U7461 ( .A(n8716), .ZN(n5732) );
  INV_X1 U7462 ( .A(n5736), .ZN(n5737) );
  INV_X1 U7463 ( .A(SI_19_), .ZN(n5738) );
  INV_X1 U7464 ( .A(n5739), .ZN(n5740) );
  NAND2_X1 U7465 ( .A1(n5740), .A2(SI_19_), .ZN(n5741) );
  NAND2_X1 U7466 ( .A1(n4477), .A2(n4491), .ZN(n5742) );
  NAND2_X1 U7467 ( .A1(n5769), .A2(n5742), .ZN(n8269) );
  NAND2_X1 U7468 ( .A1(n8269), .A2(n5624), .ZN(n5745) );
  AOI22_X1 U7469 ( .A1(n5757), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5743), .B2(
        n5756), .ZN(n5744) );
  XNOR2_X1 U7470 ( .A(n9329), .B(n5520), .ZN(n8667) );
  NAND2_X1 U7471 ( .A1(n5763), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5747) );
  NAND2_X1 U7472 ( .A1(n5772), .A2(n5747), .ZN(n9337) );
  NAND2_X1 U7473 ( .A1(n9337), .A2(n5986), .ZN(n5752) );
  INV_X1 U7474 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9197) );
  NAND2_X1 U7475 ( .A1(n4408), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U7476 ( .A1(n7135), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5748) );
  OAI211_X1 U7477 ( .C1(n9197), .C2(n7138), .A(n5749), .B(n5748), .ZN(n5750)
         );
  INV_X1 U7478 ( .A(n5750), .ZN(n5751) );
  NAND2_X1 U7479 ( .A1(n5754), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5755) );
  XNOR2_X1 U7480 ( .A(n5755), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9187) );
  AOI22_X1 U7481 ( .A1(n5757), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5756), .B2(
        n9187), .ZN(n5758) );
  XNOR2_X1 U7482 ( .A(n9507), .B(n4399), .ZN(n8666) );
  INV_X1 U7483 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9427) );
  NAND2_X1 U7484 ( .A1(n5761), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7485 ( .A1(n5763), .A2(n5762), .ZN(n9348) );
  NAND2_X1 U7486 ( .A1(n9348), .A2(n5986), .ZN(n5765) );
  AOI22_X1 U7487 ( .A1(n4408), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n7135), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U7488 ( .A1(n8666), .A2(n9358), .ZN(n8668) );
  OAI211_X1 U7489 ( .C1(n8667), .C2(n9345), .A(n8665), .B(n8668), .ZN(n5766)
         );
  INV_X1 U7490 ( .A(n5766), .ZN(n5767) );
  NAND2_X1 U7491 ( .A1(n8713), .A2(n5767), .ZN(n5787) );
  XNOR2_X1 U7492 ( .A(n5810), .B(SI_20_), .ZN(n5770) );
  NAND2_X1 U7493 ( .A1(n5757), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5771) );
  XNOR2_X1 U7494 ( .A(n7088), .B(n4399), .ZN(n5779) );
  NAND2_X1 U7495 ( .A1(n5772), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U7496 ( .A1(n5796), .A2(n5773), .ZN(n9319) );
  NAND2_X1 U7497 ( .A1(n9319), .A2(n5986), .ZN(n5778) );
  INV_X1 U7498 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U7499 ( .A1(n7135), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U7500 ( .A1(n4408), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5774) );
  OAI211_X1 U7501 ( .C1(n7138), .C2(n9422), .A(n5775), .B(n5774), .ZN(n5776)
         );
  INV_X1 U7502 ( .A(n5776), .ZN(n5777) );
  NAND2_X1 U7503 ( .A1(n5779), .A2(n9333), .ZN(n5788) );
  INV_X1 U7504 ( .A(n5779), .ZN(n5780) );
  NAND2_X1 U7505 ( .A1(n5780), .A2(n9305), .ZN(n5781) );
  NAND2_X1 U7506 ( .A1(n5788), .A2(n5781), .ZN(n8737) );
  INV_X1 U7507 ( .A(n8667), .ZN(n8734) );
  INV_X1 U7508 ( .A(n8666), .ZN(n5782) );
  AOI21_X1 U7509 ( .B1(n5782), .B2(n9027), .A(n9345), .ZN(n5784) );
  NAND3_X1 U7510 ( .A1(n5782), .A2(n9027), .A3(n9345), .ZN(n5783) );
  OAI21_X1 U7511 ( .B1(n8734), .B2(n5784), .A(n5783), .ZN(n5785) );
  NOR2_X1 U7512 ( .A1(n8737), .A2(n5785), .ZN(n5786) );
  INV_X1 U7513 ( .A(SI_20_), .ZN(n5808) );
  OAI21_X1 U7514 ( .B1(n5806), .B2(n5808), .A(n5810), .ZN(n5790) );
  NAND2_X1 U7515 ( .A1(n5806), .A2(n5808), .ZN(n5789) );
  NAND2_X1 U7516 ( .A1(n5790), .A2(n5789), .ZN(n5792) );
  XNOR2_X1 U7517 ( .A(n5814), .B(n7675), .ZN(n5791) );
  NAND2_X1 U7518 ( .A1(n8426), .A2(n5624), .ZN(n5794) );
  NAND2_X1 U7519 ( .A1(n5757), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5793) );
  XNOR2_X1 U7520 ( .A(n9491), .B(n5520), .ZN(n5803) );
  INV_X1 U7521 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7522 ( .A1(n5796), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U7523 ( .A1(n5848), .A2(n5797), .ZN(n9308) );
  NAND2_X1 U7524 ( .A1(n9308), .A2(n5986), .ZN(n5802) );
  INV_X1 U7525 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U7526 ( .A1(n4408), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7527 ( .A1(n5988), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5798) );
  OAI211_X1 U7528 ( .C1(n8403), .C2(n9307), .A(n5799), .B(n5798), .ZN(n5800)
         );
  INV_X1 U7529 ( .A(n5800), .ZN(n5801) );
  XNOR2_X1 U7530 ( .A(n5803), .B(n9317), .ZN(n8678) );
  INV_X1 U7531 ( .A(n5803), .ZN(n5804) );
  NAND2_X1 U7532 ( .A1(n5804), .A2(n9317), .ZN(n5805) );
  INV_X1 U7533 ( .A(n5814), .ZN(n5807) );
  AOI22_X1 U7534 ( .A1(n5808), .A2(n5810), .B1(n5807), .B2(n7675), .ZN(n5809)
         );
  INV_X1 U7535 ( .A(n5810), .ZN(n5813) );
  NAND2_X1 U7536 ( .A1(n5813), .A2(SI_20_), .ZN(n5811) );
  NAND2_X1 U7537 ( .A1(n5811), .A2(n7675), .ZN(n5815) );
  AND2_X1 U7538 ( .A1(SI_20_), .A2(SI_21_), .ZN(n5812) );
  AOI22_X1 U7539 ( .A1(n5815), .A2(n5814), .B1(n5813), .B2(n5812), .ZN(n5840)
         );
  INV_X1 U7540 ( .A(SI_22_), .ZN(n5816) );
  NAND2_X1 U7541 ( .A1(n5817), .A2(n5816), .ZN(n5841) );
  INV_X1 U7542 ( .A(n5817), .ZN(n5818) );
  NAND2_X1 U7543 ( .A1(n5818), .A2(SI_22_), .ZN(n5819) );
  NAND2_X1 U7544 ( .A1(n5841), .A2(n5819), .ZN(n5831) );
  NAND2_X1 U7545 ( .A1(n8437), .A2(n5624), .ZN(n5822) );
  NAND2_X1 U7546 ( .A1(n5757), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5821) );
  XNOR2_X1 U7547 ( .A(n9291), .B(n4399), .ZN(n8755) );
  INV_X1 U7548 ( .A(n8755), .ZN(n5828) );
  XNOR2_X1 U7549 ( .A(n5848), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U7550 ( .A1(n9292), .A2(n5986), .ZN(n5827) );
  INV_X1 U7551 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9416) );
  NAND2_X1 U7552 ( .A1(n7135), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7553 ( .A1(n4408), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5823) );
  OAI211_X1 U7554 ( .C1(n7138), .C2(n9416), .A(n5824), .B(n5823), .ZN(n5825)
         );
  INV_X1 U7555 ( .A(n5825), .ZN(n5826) );
  NAND2_X1 U7556 ( .A1(n5828), .A2(n9304), .ZN(n5830) );
  INV_X1 U7557 ( .A(n9304), .ZN(n8754) );
  AND2_X1 U7558 ( .A1(n8755), .A2(n8754), .ZN(n5829) );
  INV_X1 U7559 ( .A(n5831), .ZN(n5838) );
  NAND2_X1 U7560 ( .A1(n5832), .A2(n5838), .ZN(n5833) );
  NAND2_X1 U7561 ( .A1(n5833), .A2(n5841), .ZN(n5845) );
  INV_X1 U7562 ( .A(SI_23_), .ZN(n5834) );
  NAND2_X1 U7563 ( .A1(n5835), .A2(n5834), .ZN(n5855) );
  INV_X1 U7564 ( .A(n5835), .ZN(n5836) );
  NAND2_X1 U7565 ( .A1(n5836), .A2(SI_23_), .ZN(n5837) );
  AND2_X1 U7566 ( .A1(n5838), .A2(n5844), .ZN(n5839) );
  INV_X1 U7567 ( .A(n5844), .ZN(n5842) );
  NAND2_X1 U7568 ( .A1(n8455), .A2(n5624), .ZN(n5847) );
  NAND2_X1 U7569 ( .A1(n5906), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5846) );
  XNOR2_X1 U7570 ( .A(n7093), .B(n5520), .ZN(n8659) );
  INV_X1 U7571 ( .A(n8659), .ZN(n8722) );
  OAI21_X1 U7572 ( .B1(n5848), .B2(P2_REG3_REG_22__SCAN_IN), .A(
        P2_REG3_REG_23__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7573 ( .A1(n5849), .A2(n4444), .ZN(n9283) );
  NAND2_X1 U7574 ( .A1(n9283), .A2(n5986), .ZN(n5854) );
  INV_X1 U7575 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9411) );
  NAND2_X1 U7576 ( .A1(n4408), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U7577 ( .A1(n7135), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5850) );
  OAI211_X1 U7578 ( .C1(n9411), .C2(n7138), .A(n5851), .B(n5850), .ZN(n5852)
         );
  INV_X1 U7579 ( .A(n5852), .ZN(n5853) );
  NAND2_X1 U7580 ( .A1(n8722), .A2(n9269), .ZN(n5877) );
  INV_X1 U7581 ( .A(SI_24_), .ZN(n5857) );
  NAND2_X1 U7582 ( .A1(n5858), .A2(n5857), .ZN(n5882) );
  INV_X1 U7583 ( .A(n5858), .ZN(n5859) );
  NAND2_X1 U7584 ( .A1(n5859), .A2(SI_24_), .ZN(n5860) );
  NAND2_X1 U7585 ( .A1(n5862), .A2(n5861), .ZN(n5883) );
  OR2_X1 U7586 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  NAND2_X1 U7587 ( .A1(n5883), .A2(n5863), .ZN(n8488) );
  NAND2_X1 U7588 ( .A1(n8488), .A2(n5624), .ZN(n5865) );
  NAND2_X1 U7589 ( .A1(n5757), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5864) );
  XNOR2_X1 U7590 ( .A(n9273), .B(n5520), .ZN(n8725) );
  INV_X1 U7591 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7592 ( .A1(n4444), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7593 ( .A1(n5893), .A2(n5868), .ZN(n9271) );
  NAND2_X1 U7594 ( .A1(n9271), .A2(n5986), .ZN(n5873) );
  INV_X1 U7595 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U7596 ( .A1(n5988), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U7597 ( .A1(n7135), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5869) );
  OAI211_X1 U7598 ( .C1(n8401), .C2(n9474), .A(n5870), .B(n5869), .ZN(n5871)
         );
  INV_X1 U7599 ( .A(n5871), .ZN(n5872) );
  NAND2_X1 U7600 ( .A1(n5875), .A2(n5874), .ZN(n5876) );
  AOI21_X1 U7601 ( .B1(n8659), .B2(n9288), .A(n8974), .ZN(n5879) );
  NAND3_X1 U7602 ( .A1(n8659), .A2(n9288), .A3(n8974), .ZN(n5878) );
  OAI21_X1 U7603 ( .B1(n5879), .B2(n5875), .A(n5878), .ZN(n5880) );
  INV_X1 U7604 ( .A(SI_25_), .ZN(n5884) );
  NAND2_X1 U7605 ( .A1(n5885), .A2(n5884), .ZN(n5900) );
  INV_X1 U7606 ( .A(n5885), .ZN(n5886) );
  NAND2_X1 U7607 ( .A1(n5886), .A2(SI_25_), .ZN(n5887) );
  OR2_X1 U7608 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  NAND2_X1 U7609 ( .A1(n5901), .A2(n5890), .ZN(n8577) );
  NAND2_X1 U7610 ( .A1(n8577), .A2(n5624), .ZN(n5892) );
  NAND2_X1 U7611 ( .A1(n5757), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5891) );
  XNOR2_X1 U7612 ( .A(n9469), .B(n5520), .ZN(n5914) );
  NAND2_X1 U7613 ( .A1(n5893), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7614 ( .A1(n5907), .A2(n5894), .ZN(n9258) );
  NAND2_X1 U7615 ( .A1(n9258), .A2(n5986), .ZN(n5899) );
  INV_X1 U7616 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9405) );
  NAND2_X1 U7617 ( .A1(n4408), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7618 ( .A1(n7135), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5895) );
  OAI211_X1 U7619 ( .C1(n9405), .C2(n7138), .A(n5896), .B(n5895), .ZN(n5897)
         );
  INV_X1 U7620 ( .A(n5897), .ZN(n5898) );
  XNOR2_X1 U7621 ( .A(n5914), .B(n9026), .ZN(n8698) );
  INV_X1 U7622 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8594) );
  INV_X1 U7623 ( .A(SI_26_), .ZN(n7673) );
  NAND2_X1 U7624 ( .A1(n5902), .A2(n7673), .ZN(n5920) );
  INV_X1 U7625 ( .A(n5902), .ZN(n5903) );
  NAND2_X1 U7626 ( .A1(n5903), .A2(SI_26_), .ZN(n5904) );
  XNOR2_X1 U7627 ( .A(n7095), .B(n4399), .ZN(n8776) );
  NAND2_X1 U7628 ( .A1(n5907), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7629 ( .A1(n5930), .A2(n5908), .ZN(n9251) );
  NAND2_X1 U7630 ( .A1(n9251), .A2(n5986), .ZN(n5913) );
  INV_X1 U7631 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9462) );
  NAND2_X1 U7632 ( .A1(n5988), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7633 ( .A1(n7135), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5909) );
  OAI211_X1 U7634 ( .C1(n8401), .C2(n9462), .A(n5910), .B(n5909), .ZN(n5911)
         );
  INV_X1 U7635 ( .A(n5911), .ZN(n5912) );
  INV_X1 U7636 ( .A(n5914), .ZN(n5915) );
  NAND2_X1 U7637 ( .A1(n5915), .A2(n9026), .ZN(n8774) );
  INV_X1 U7638 ( .A(n5916), .ZN(n5917) );
  NAND2_X1 U7639 ( .A1(n8776), .A2(n4907), .ZN(n5918) );
  NAND2_X1 U7640 ( .A1(n5905), .A2(n5919), .ZN(n5921) );
  INV_X1 U7641 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7736) );
  INV_X1 U7642 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8627) );
  INV_X1 U7643 ( .A(SI_27_), .ZN(n5922) );
  NAND2_X1 U7644 ( .A1(n5923), .A2(n5922), .ZN(n6466) );
  INV_X1 U7645 ( .A(n5923), .ZN(n5924) );
  NAND2_X1 U7646 ( .A1(n5924), .A2(SI_27_), .ZN(n5925) );
  NAND2_X1 U7647 ( .A1(n8626), .A2(n5624), .ZN(n5927) );
  NAND2_X1 U7648 ( .A1(n5757), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5926) );
  XNOR2_X1 U7649 ( .A(n9398), .B(n4399), .ZN(n6012) );
  INV_X1 U7650 ( .A(n5930), .ZN(n5929) );
  INV_X1 U7651 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7652 ( .A1(n5930), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7653 ( .A1(n5941), .A2(n5931), .ZN(n9233) );
  INV_X1 U7654 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7721) );
  NAND2_X1 U7655 ( .A1(n4408), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7656 ( .A1(n7135), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5932) );
  OAI211_X1 U7657 ( .C1(n7721), .C2(n7138), .A(n5933), .B(n5932), .ZN(n5934)
         );
  INV_X1 U7658 ( .A(n5934), .ZN(n5935) );
  NOR2_X1 U7659 ( .A1(n6012), .A2(n7130), .ZN(n5981) );
  AOI21_X1 U7660 ( .B1(n6012), .B2(n7130), .A(n5981), .ZN(n6786) );
  INV_X1 U7661 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5938) );
  INV_X1 U7662 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8640) );
  XNOR2_X1 U7663 ( .A(n6467), .B(SI_28_), .ZN(n6845) );
  NAND2_X1 U7664 ( .A1(n8639), .A2(n5624), .ZN(n5940) );
  NAND2_X1 U7665 ( .A1(n5757), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7666 ( .A1(n5941), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U7667 ( .A1(n5985), .A2(n5942), .ZN(n9229) );
  NAND2_X1 U7668 ( .A1(n9229), .A2(n5986), .ZN(n5947) );
  INV_X1 U7669 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9395) );
  NAND2_X1 U7670 ( .A1(n4408), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7671 ( .A1(n7135), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5943) );
  OAI211_X1 U7672 ( .C1(n9395), .C2(n7138), .A(n5944), .B(n5943), .ZN(n5945)
         );
  INV_X1 U7673 ( .A(n5945), .ZN(n5946) );
  XNOR2_X1 U7674 ( .A(n8836), .B(n4399), .ZN(n5948) );
  INV_X1 U7675 ( .A(n6013), .ZN(n5980) );
  NAND2_X1 U7676 ( .A1(n5949), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5951) );
  XNOR2_X1 U7677 ( .A(n5951), .B(n5950), .ZN(n8578) );
  NAND2_X1 U7678 ( .A1(n8578), .A2(n8595), .ZN(n5954) );
  INV_X1 U7679 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n5952) );
  NAND2_X1 U7680 ( .A1(n7312), .A2(n5952), .ZN(n5953) );
  NAND2_X1 U7681 ( .A1(n5954), .A2(n5953), .ZN(n7969) );
  OR2_X1 U7682 ( .A1(n7969), .A2(n5974), .ZN(n7158) );
  NOR2_X1 U7683 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .ZN(
        n7574) );
  NOR4_X1 U7684 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5957) );
  NOR4_X1 U7685 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5956) );
  NOR4_X1 U7686 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5955) );
  NAND4_X1 U7687 ( .A1(n7574), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(n5963)
         );
  NOR4_X1 U7688 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5961) );
  NOR4_X1 U7689 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5960) );
  NOR4_X1 U7690 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n5959) );
  NOR4_X1 U7691 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5958) );
  NAND4_X1 U7692 ( .A1(n5961), .A2(n5960), .A3(n5959), .A4(n5958), .ZN(n5962)
         );
  OAI21_X1 U7693 ( .B1(n5963), .B2(n5962), .A(n7312), .ZN(n7157) );
  INV_X1 U7694 ( .A(n7157), .ZN(n5964) );
  NOR2_X1 U7695 ( .A1(n7158), .A2(n5964), .ZN(n5997) );
  XNOR2_X1 U7696 ( .A(n5966), .B(n5965), .ZN(n7174) );
  INV_X1 U7697 ( .A(n5968), .ZN(n5969) );
  NAND2_X1 U7698 ( .A1(n5969), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7699 ( .A1(n5743), .A2(n9020), .ZN(n7105) );
  NOR2_X1 U7700 ( .A1(n8994), .A2(n7105), .ZN(n5976) );
  INV_X1 U7701 ( .A(n5976), .ZN(n5972) );
  NAND3_X1 U7702 ( .A1(n10565), .A2(n8999), .A3(n5972), .ZN(n5998) );
  INV_X1 U7703 ( .A(n5998), .ZN(n5973) );
  NAND2_X1 U7704 ( .A1(n7150), .A2(n5973), .ZN(n5979) );
  AND2_X1 U7705 ( .A1(n5974), .A2(n7157), .ZN(n5975) );
  NAND2_X1 U7706 ( .A1(n8863), .A2(n5976), .ZN(n7148) );
  INV_X1 U7707 ( .A(n7148), .ZN(n5977) );
  NAND2_X1 U7708 ( .A1(n7151), .A2(n5977), .ZN(n5978) );
  NAND2_X1 U7709 ( .A1(n5980), .A2(n8790), .ZN(n6018) );
  INV_X1 U7710 ( .A(n5981), .ZN(n5982) );
  NAND2_X1 U7711 ( .A1(n7150), .A2(n9443), .ZN(n5984) );
  INV_X1 U7712 ( .A(n7161), .ZN(n8024) );
  INV_X1 U7713 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U7714 ( .A1(n4408), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7715 ( .A1(n5988), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5989) );
  OAI211_X1 U7716 ( .C1(n8403), .C2(n8642), .A(n5990), .B(n5989), .ZN(n5991)
         );
  INV_X1 U7717 ( .A(n5991), .ZN(n5992) );
  INV_X1 U7718 ( .A(n6000), .ZN(n5993) );
  INV_X1 U7719 ( .A(n7974), .ZN(n5994) );
  NAND2_X1 U7720 ( .A1(n5994), .A2(n7151), .ZN(n6009) );
  NAND2_X1 U7721 ( .A1(n9017), .A2(n9199), .ZN(n5995) );
  NAND2_X1 U7722 ( .A1(n4746), .A2(n5995), .ZN(n7142) );
  INV_X1 U7723 ( .A(n7142), .ZN(n5996) );
  INV_X1 U7724 ( .A(n5997), .ZN(n5999) );
  NAND2_X1 U7725 ( .A1(n5998), .A2(n10531), .ZN(n7152) );
  NAND2_X1 U7726 ( .A1(n5999), .A2(n7152), .ZN(n6002) );
  AND3_X1 U7727 ( .A1(n7159), .A2(n7173), .A3(n7174), .ZN(n6001) );
  OAI211_X1 U7728 ( .C1(n6005), .C2(n7148), .A(n6002), .B(n6001), .ZN(n6003)
         );
  NAND2_X1 U7729 ( .A1(n6003), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6008) );
  INV_X1 U7730 ( .A(n7314), .ZN(n6004) );
  NOR2_X1 U7731 ( .A1(n7974), .A2(n6004), .ZN(n9018) );
  INV_X1 U7732 ( .A(n6005), .ZN(n6006) );
  NAND2_X1 U7733 ( .A1(n9018), .A2(n6006), .ZN(n6007) );
  AOI22_X1 U7734 ( .A1(n9229), .A2(n8797), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n6011) );
  NAND2_X1 U7735 ( .A1(n9249), .A2(n8793), .ZN(n6010) );
  OAI211_X1 U7736 ( .C1(n9025), .C2(n8795), .A(n6011), .B(n6010), .ZN(n6015)
         );
  NOR4_X1 U7737 ( .A1(n6013), .A2(n8786), .A3(n7130), .A4(n6012), .ZN(n6014)
         );
  AOI211_X1 U7738 ( .C1(n8784), .C2(n9456), .A(n6015), .B(n6014), .ZN(n6016)
         );
  OAI211_X1 U7739 ( .C1(n6788), .C2(n6018), .A(n6017), .B(n6016), .ZN(P2_U3160) );
  INV_X1 U7740 ( .A(n6234), .ZN(n6027) );
  NOR2_X4 U7741 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6120) );
  NAND2_X1 U7742 ( .A1(n6034), .A2(n6024), .ZN(n6025) );
  NOR2_X2 U7743 ( .A1(n6135), .A2(n6025), .ZN(n6026) );
  NOR2_X1 U7744 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6028) );
  NAND4_X1 U7745 ( .A1(n6028), .A2(n6377), .A3(n6402), .A4(n6405), .ZN(n6030)
         );
  INV_X2 U7746 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6367) );
  NAND4_X1 U7747 ( .A1(n6368), .A2(n6367), .A3(n6370), .A4(n4600), .ZN(n6029)
         );
  NAND2_X1 U7748 ( .A1(n6032), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6033) );
  AND2_X1 U7749 ( .A1(n6149), .A2(n6034), .ZN(n6172) );
  NAND2_X1 U7750 ( .A1(n6172), .A2(n6173), .ZN(n6235) );
  INV_X1 U7751 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6070) );
  INV_X1 U7752 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6035) );
  NAND3_X1 U7753 ( .A1(n6070), .A2(n6090), .A3(n6035), .ZN(n6036) );
  NAND2_X1 U7754 ( .A1(n6189), .A2(n4684), .ZN(n6203) );
  NAND2_X1 U7755 ( .A1(n6223), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6055) );
  INV_X1 U7756 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7757 ( .A1(n6055), .A2(n6221), .ZN(n6037) );
  NAND2_X1 U7758 ( .A1(n6037), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6038) );
  AOI22_X1 U7759 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n6277), .B1(n9853), .B2(
        n6276), .ZN(n6039) );
  NAND2_X1 U7760 ( .A1(n6210), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7761 ( .A1(n6058), .A2(n6040), .ZN(n6041) );
  AND2_X1 U7762 ( .A1(n6228), .A2(n6041), .ZN(n8585) );
  NAND2_X1 U7763 ( .A1(n8585), .A2(n6337), .ZN(n6054) );
  INV_X1 U7764 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8038) );
  OR2_X1 U7765 ( .A1(n6126), .A2(n8038), .ZN(n6053) );
  NAND2_X2 U7766 ( .A1(n6048), .A2(n6049), .ZN(n6485) );
  INV_X1 U7767 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6047) );
  OR2_X1 U7768 ( .A1(n6485), .A2(n6047), .ZN(n6052) );
  INV_X1 U7769 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n6050) );
  OR2_X1 U7770 ( .A1(n6143), .A2(n6050), .ZN(n6051) );
  INV_X1 U7771 ( .A(n8511), .ZN(n9741) );
  NAND2_X1 U7772 ( .A1(n7342), .A2(n5036), .ZN(n6057) );
  XNOR2_X1 U7773 ( .A(n6055), .B(P1_IR_REG_12__SCAN_IN), .ZN(n8044) );
  AOI22_X1 U7774 ( .A1(n6277), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6276), .B2(
        n8044), .ZN(n6056) );
  OR2_X1 U7775 ( .A1(n6210), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6059) );
  AND2_X1 U7776 ( .A1(n6059), .A2(n6058), .ZN(n10316) );
  NAND2_X1 U7777 ( .A1(n6337), .A2(n10316), .ZN(n6066) );
  INV_X1 U7778 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6060) );
  OR2_X1 U7779 ( .A1(n6126), .A2(n6060), .ZN(n6065) );
  INV_X1 U7780 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6061) );
  OR2_X1 U7781 ( .A1(n6143), .A2(n6061), .ZN(n6064) );
  INV_X1 U7782 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6062) );
  OR2_X1 U7783 ( .A1(n6485), .A2(n6062), .ZN(n6063) );
  INV_X1 U7784 ( .A(n8518), .ZN(n6067) );
  NOR2_X1 U7785 ( .A1(n8522), .A2(n6067), .ZN(n6219) );
  NAND2_X1 U7786 ( .A1(n7328), .A2(n5036), .ZN(n6074) );
  NAND2_X1 U7787 ( .A1(n6068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7788 ( .A1(n6091), .A2(n6090), .ZN(n6069) );
  NAND2_X1 U7789 ( .A1(n6069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U7790 ( .A1(n6082), .A2(n6070), .ZN(n6071) );
  NAND2_X1 U7791 ( .A1(n6071), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6072) );
  XNOR2_X1 U7792 ( .A(n6072), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7491) );
  AOI22_X1 U7793 ( .A1(n4406), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6276), .B2(
        n7491), .ZN(n6073) );
  NAND2_X1 U7794 ( .A1(n6870), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6081) );
  INV_X1 U7795 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6075) );
  OR2_X1 U7796 ( .A1(n6126), .A2(n6075), .ZN(n6080) );
  NAND2_X1 U7797 ( .A1(n6085), .A2(n7389), .ZN(n6076) );
  NAND2_X1 U7798 ( .A1(n6196), .A2(n6076), .ZN(n10350) );
  OR2_X1 U7799 ( .A1(n6384), .A2(n10350), .ZN(n6079) );
  INV_X1 U7800 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6077) );
  OR2_X1 U7801 ( .A1(n6485), .A2(n6077), .ZN(n6078) );
  XNOR2_X1 U7802 ( .A(n6082), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9821) );
  NAND2_X1 U7803 ( .A1(n6870), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6089) );
  INV_X1 U7804 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7382) );
  OR2_X1 U7805 ( .A1(n6126), .A2(n7382), .ZN(n6088) );
  OR2_X1 U7806 ( .A1(n6095), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7807 ( .A1(n6085), .A2(n6084), .ZN(n10366) );
  OR2_X1 U7808 ( .A1(n6384), .A2(n10366), .ZN(n6087) );
  INV_X1 U7809 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7563) );
  OR2_X1 U7810 ( .A1(n6485), .A2(n7563), .ZN(n6086) );
  NAND2_X1 U7811 ( .A1(n6919), .A2(n10344), .ZN(n6915) );
  NAND2_X1 U7812 ( .A1(n8468), .A2(n8566), .ZN(n10343) );
  XNOR2_X1 U7813 ( .A(n6091), .B(n6090), .ZN(n9804) );
  NAND2_X1 U7814 ( .A1(n7301), .A2(n5036), .ZN(n6093) );
  OR2_X1 U7815 ( .A1(n4412), .A2(n4829), .ZN(n6092) );
  OAI211_X1 U7816 ( .C1(n7324), .C2(n9804), .A(n6093), .B(n6092), .ZN(n8332)
         );
  NAND2_X1 U7817 ( .A1(n6870), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6100) );
  INV_X1 U7818 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7380) );
  OR2_X1 U7819 ( .A1(n6126), .A2(n7380), .ZN(n6099) );
  AND2_X1 U7820 ( .A1(n6106), .A2(n6094), .ZN(n6096) );
  OR2_X1 U7821 ( .A1(n6096), .A2(n6095), .ZN(n8329) );
  OR2_X1 U7822 ( .A1(n6384), .A2(n8329), .ZN(n6098) );
  INV_X1 U7823 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7404) );
  OR2_X1 U7824 ( .A1(n6485), .A2(n7404), .ZN(n6097) );
  NAND2_X1 U7825 ( .A1(n8332), .A2(n8464), .ZN(n10341) );
  NAND2_X1 U7826 ( .A1(n6101), .A2(n8553), .ZN(n6927) );
  NAND2_X1 U7827 ( .A1(n6235), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6103) );
  XNOR2_X1 U7828 ( .A(n6103), .B(n6102), .ZN(n9790) );
  NAND2_X1 U7829 ( .A1(n7302), .A2(n4410), .ZN(n6105) );
  OR2_X1 U7830 ( .A1(n4400), .A2(n7306), .ZN(n6104) );
  NAND2_X1 U7831 ( .A1(n6481), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6111) );
  INV_X1 U7832 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7402) );
  OR2_X1 U7833 ( .A1(n6485), .A2(n7402), .ZN(n6110) );
  OAI21_X1 U7834 ( .B1(n6177), .B2(P1_REG3_REG_6__SCAN_IN), .A(n6106), .ZN(
        n8253) );
  OR2_X1 U7835 ( .A1(n6384), .A2(n8253), .ZN(n6109) );
  INV_X1 U7836 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6107) );
  OR2_X1 U7837 ( .A1(n6143), .A2(n6107), .ZN(n6108) );
  NAND2_X1 U7838 ( .A1(n8256), .A2(n8293), .ZN(n6908) );
  INV_X1 U7839 ( .A(n6908), .ZN(n8289) );
  NAND2_X1 U7840 ( .A1(n6140), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6113) );
  INV_X1 U7841 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6112) );
  INV_X1 U7842 ( .A(n6384), .ZN(n6114) );
  INV_X1 U7843 ( .A(n6116), .ZN(n7831) );
  NAND2_X1 U7844 ( .A1(n7290), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6117) );
  OAI21_X1 U7845 ( .B1(n7291), .B2(n7290), .A(n6117), .ZN(n6118) );
  NAND2_X1 U7846 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6119) );
  MUX2_X1 U7847 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6119), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n6122) );
  INV_X1 U7848 ( .A(n6120), .ZN(n6121) );
  INV_X1 U7849 ( .A(n7392), .ZN(n9759) );
  NAND3_X1 U7850 ( .A1(n6116), .A2(n9759), .A3(n6123), .ZN(n6125) );
  INV_X1 U7851 ( .A(n6123), .ZN(n10230) );
  INV_X1 U7852 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7829) );
  INV_X1 U7853 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6522) );
  OR2_X1 U7854 ( .A1(n6126), .A2(n6522), .ZN(n6130) );
  INV_X1 U7855 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6127) );
  INV_X1 U7856 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7454) );
  OR2_X1 U7857 ( .A1(n6384), .A2(n7454), .ZN(n6128) );
  XNOR2_X1 U7858 ( .A(n6132), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10228) );
  OR2_X1 U7859 ( .A1(n6511), .A2(n10429), .ZN(n6133) );
  INV_X1 U7860 ( .A(n6134), .ZN(n6136) );
  OR2_X1 U7861 ( .A1(n6150), .A2(n5039), .ZN(n6139) );
  INV_X1 U7862 ( .A(n6137), .ZN(n7293) );
  NAND2_X1 U7863 ( .A1(n6140), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6147) );
  INV_X1 U7864 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6141) );
  OR2_X1 U7865 ( .A1(n6384), .A2(n6141), .ZN(n6146) );
  INV_X1 U7866 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7394) );
  INV_X1 U7867 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6142) );
  OR2_X1 U7868 ( .A1(n6143), .A2(n6142), .ZN(n6144) );
  AND2_X1 U7869 ( .A1(n6526), .A2(n8100), .ZN(n6148) );
  OR2_X1 U7870 ( .A1(n6526), .A2(n8100), .ZN(n6800) );
  INV_X1 U7871 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6159) );
  XNOR2_X1 U7872 ( .A(n6160), .B(n6159), .ZN(n7396) );
  OR2_X1 U7873 ( .A1(n4400), .A2(n5409), .ZN(n6152) );
  OR2_X1 U7874 ( .A1(n6364), .A2(n7295), .ZN(n6151) );
  NAND2_X1 U7875 ( .A1(n6481), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6158) );
  INV_X1 U7876 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6153) );
  OR2_X1 U7877 ( .A1(n6485), .A2(n6153), .ZN(n6157) );
  INV_X1 U7878 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6154) );
  OR2_X1 U7879 ( .A1(n6143), .A2(n6154), .ZN(n6156) );
  OR2_X1 U7880 ( .A1(n6384), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7881 ( .A1(n6539), .A2(n7999), .ZN(n6430) );
  NAND2_X1 U7882 ( .A1(n6160), .A2(n6159), .ZN(n6161) );
  NAND2_X1 U7883 ( .A1(n6161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6163) );
  INV_X1 U7884 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6162) );
  OR2_X1 U7885 ( .A1(n4400), .A2(n5002), .ZN(n6164) );
  OAI211_X1 U7886 ( .C1(n7324), .C2(n7856), .A(n6165), .B(n6164), .ZN(n8004)
         );
  NAND2_X1 U7887 ( .A1(n6481), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6170) );
  INV_X1 U7888 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7398) );
  OR2_X1 U7889 ( .A1(n6485), .A2(n7398), .ZN(n6169) );
  XNOR2_X1 U7890 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10381) );
  OR2_X1 U7891 ( .A1(n6384), .A2(n10381), .ZN(n6168) );
  INV_X1 U7892 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6166) );
  OR2_X1 U7893 ( .A1(n6143), .A2(n6166), .ZN(n6167) );
  NAND2_X1 U7894 ( .A1(n8004), .A2(n9750), .ZN(n6434) );
  OR2_X1 U7895 ( .A1(n6172), .A2(n6044), .ZN(n6174) );
  XNOR2_X1 U7896 ( .A(n6174), .B(n6173), .ZN(n7400) );
  OR2_X1 U7897 ( .A1(n4400), .A2(n5468), .ZN(n6176) );
  AOI21_X1 U7898 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6178) );
  NOR2_X1 U7899 ( .A1(n6178), .A2(n6177), .ZN(n8160) );
  NAND2_X1 U7900 ( .A1(n6337), .A2(n8160), .ZN(n6185) );
  INV_X1 U7901 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6179) );
  OR2_X1 U7902 ( .A1(n6126), .A2(n6179), .ZN(n6184) );
  INV_X1 U7903 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6180) );
  OR2_X1 U7904 ( .A1(n6485), .A2(n6180), .ZN(n6183) );
  INV_X1 U7905 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6181) );
  OR2_X1 U7906 ( .A1(n6143), .A2(n6181), .ZN(n6182) );
  OR2_X1 U7907 ( .A1(n8256), .A2(n8293), .ZN(n6903) );
  INV_X1 U7908 ( .A(n6903), .ZN(n6188) );
  INV_X1 U7909 ( .A(n8464), .ZN(n9747) );
  NAND2_X1 U7910 ( .A1(n10464), .A2(n9747), .ZN(n6912) );
  INV_X1 U7911 ( .A(n6912), .ZN(n6186) );
  INV_X1 U7912 ( .A(n6189), .ZN(n6190) );
  NAND2_X1 U7913 ( .A1(n6190), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6191) );
  MUX2_X1 U7914 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6191), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n6192) );
  AOI22_X1 U7915 ( .A1(n6277), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6276), .B2(
        n7884), .ZN(n6193) );
  NAND2_X1 U7916 ( .A1(n6481), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6202) );
  INV_X1 U7917 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6194) );
  OR2_X1 U7918 ( .A1(n6143), .A2(n6194), .ZN(n6201) );
  NAND2_X1 U7919 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  NAND2_X1 U7920 ( .A1(n6208), .A2(n6197), .ZN(n10330) );
  OR2_X1 U7921 ( .A1(n6384), .A2(n10330), .ZN(n6200) );
  INV_X1 U7922 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6198) );
  OR2_X1 U7923 ( .A1(n6485), .A2(n6198), .ZN(n6199) );
  NAND4_X1 U7924 ( .A1(n6202), .A2(n6201), .A3(n6200), .A4(n6199), .ZN(n9744)
         );
  AND2_X1 U7925 ( .A1(n10484), .A2(n9744), .ZN(n6926) );
  INV_X1 U7926 ( .A(n9744), .ZN(n6607) );
  NAND2_X1 U7927 ( .A1(n10335), .A2(n6607), .ZN(n8413) );
  NAND2_X1 U7928 ( .A1(n6921), .A2(n8413), .ZN(n6885) );
  NAND2_X1 U7929 ( .A1(n7338), .A2(n5036), .ZN(n6206) );
  NAND2_X1 U7930 ( .A1(n6203), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6204) );
  XNOR2_X1 U7931 ( .A(n6204), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U7932 ( .A1(n4406), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6276), .B2(
        n9840), .ZN(n6205) );
  AND2_X1 U7933 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  NOR2_X1 U7934 ( .A1(n6210), .A2(n6209), .ZN(n9677) );
  NAND2_X1 U7935 ( .A1(n6337), .A2(n9677), .ZN(n6216) );
  INV_X1 U7936 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6211) );
  OR2_X1 U7937 ( .A1(n6126), .A2(n6211), .ZN(n6215) );
  INV_X1 U7938 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7887) );
  OR2_X1 U7939 ( .A1(n6485), .A2(n7887), .ZN(n6214) );
  INV_X1 U7940 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6212) );
  OR2_X1 U7941 ( .A1(n6143), .A2(n6212), .ZN(n6213) );
  NAND2_X1 U7942 ( .A1(n10489), .A2(n8496), .ZN(n6923) );
  INV_X1 U7943 ( .A(n8413), .ZN(n6217) );
  NOR2_X1 U7944 ( .A1(n8414), .A2(n6217), .ZN(n6218) );
  NAND2_X1 U7945 ( .A1(n10317), .A2(n8417), .ZN(n6924) );
  NAND2_X1 U7946 ( .A1(n7825), .A2(n5036), .ZN(n6226) );
  NAND2_X1 U7947 ( .A1(n6221), .A2(n6220), .ZN(n6222) );
  OAI21_X1 U7948 ( .B1(n6223), .B2(n6222), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6224) );
  XNOR2_X1 U7949 ( .A(n6224), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U7950 ( .A1(n6277), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n10243), 
        .B2(n6276), .ZN(n6225) );
  AND2_X1 U7951 ( .A1(n6228), .A2(n6227), .ZN(n6229) );
  OR2_X1 U7952 ( .A1(n6229), .A2(n6239), .ZN(n9555) );
  AOI22_X1 U7953 ( .A1(n6481), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n6870), .B2(
        P1_REG0_REG_14__SCAN_IN), .ZN(n6232) );
  INV_X1 U7954 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6230) );
  OR2_X1 U7955 ( .A1(n6485), .A2(n6230), .ZN(n6231) );
  OAI211_X1 U7956 ( .C1(n9555), .C2(n6384), .A(n6232), .B(n6231), .ZN(n9740)
         );
  INV_X1 U7957 ( .A(n9740), .ZN(n6810) );
  XNOR2_X1 U7958 ( .A(n10147), .B(n6810), .ZN(n8502) );
  INV_X1 U7959 ( .A(n8502), .ZN(n8509) );
  AND2_X1 U7960 ( .A1(n10147), .A2(n6810), .ZN(n6797) );
  INV_X1 U7961 ( .A(n6797), .ZN(n6233) );
  NAND2_X1 U7962 ( .A1(n7908), .A2(n5036), .ZN(n6238) );
  OAI21_X1 U7963 ( .B1(n6235), .B2(n6234), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6236) );
  XNOR2_X1 U7964 ( .A(n6236), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U7965 ( .A1(n4406), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6276), .B2(
        n10260), .ZN(n6237) );
  NOR2_X1 U7966 ( .A1(n6239), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6240) );
  OR2_X1 U7967 ( .A1(n6246), .A2(n6240), .ZN(n8603) );
  AOI22_X1 U7968 ( .A1(n6481), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n6870), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U7969 ( .A1(n6869), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6241) );
  OAI211_X1 U7970 ( .C1(n8603), .C2(n6384), .A(n6242), .B(n6241), .ZN(n9739)
         );
  XNOR2_X1 U7971 ( .A(n10143), .B(n9739), .ZN(n8598) );
  INV_X1 U7972 ( .A(n9739), .ZN(n8512) );
  NAND2_X1 U7973 ( .A1(n10143), .A2(n8512), .ZN(n6796) );
  XNOR2_X1 U7974 ( .A(n6251), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10274) );
  AOI22_X1 U7975 ( .A1(n6277), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6276), .B2(
        n10274), .ZN(n6244) );
  OR2_X1 U7976 ( .A1(n6246), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7977 ( .A1(n6256), .A2(n6247), .ZN(n10069) );
  AOI22_X1 U7978 ( .A1(n6481), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n6869), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n6249) );
  INV_X1 U7979 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10199) );
  OR2_X1 U7980 ( .A1(n6143), .A2(n10199), .ZN(n6248) );
  OAI211_X1 U7981 ( .C1(n10069), .C2(n6384), .A(n6249), .B(n6248), .ZN(n9737)
         );
  INV_X1 U7982 ( .A(n9737), .ZN(n6651) );
  NAND2_X1 U7983 ( .A1(n10138), .A2(n6651), .ZN(n6813) );
  NAND2_X1 U7984 ( .A1(n8127), .A2(n5036), .ZN(n6254) );
  NAND2_X1 U7985 ( .A1(n6251), .A2(n6369), .ZN(n6252) );
  NAND2_X1 U7986 ( .A1(n6252), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6263) );
  XNOR2_X1 U7987 ( .A(n6263), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10286) );
  AOI22_X1 U7988 ( .A1(n4406), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6276), .B2(
        n10286), .ZN(n6253) );
  INV_X1 U7989 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7990 ( .A1(n6256), .A2(n6255), .ZN(n6257) );
  AND2_X1 U7991 ( .A1(n6268), .A2(n6257), .ZN(n10051) );
  NAND2_X1 U7992 ( .A1(n10051), .A2(n6337), .ZN(n6262) );
  INV_X1 U7993 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10134) );
  NAND2_X1 U7994 ( .A1(n6869), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7995 ( .A1(n6870), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6258) );
  OAI211_X1 U7996 ( .C1(n6126), .C2(n10134), .A(n6259), .B(n6258), .ZN(n6260)
         );
  INV_X1 U7997 ( .A(n6260), .ZN(n6261) );
  NAND2_X1 U7998 ( .A1(n6262), .A2(n6261), .ZN(n9736) );
  NAND2_X1 U7999 ( .A1(n10054), .A2(n9736), .ZN(n6817) );
  INV_X1 U8000 ( .A(n9736), .ZN(n6661) );
  NAND2_X1 U8001 ( .A1(n8150), .A2(n5036), .ZN(n6266) );
  NAND2_X1 U8002 ( .A1(n6263), .A2(n6370), .ZN(n6264) );
  NAND2_X1 U8003 ( .A1(n6264), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6273) );
  XNOR2_X1 U8004 ( .A(n6273), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U8005 ( .A1(n6277), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6276), .B2(
        n10304), .ZN(n6265) );
  INV_X1 U8006 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6267) );
  AND2_X1 U8007 ( .A1(n6268), .A2(n6267), .ZN(n6269) );
  OR2_X1 U8008 ( .A1(n6269), .A2(n6288), .ZN(n9691) );
  INV_X1 U8009 ( .A(n9691), .ZN(n10039) );
  INV_X1 U8010 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10129) );
  NAND2_X1 U8011 ( .A1(n6870), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U8012 ( .A1(n6869), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6270) );
  OAI211_X1 U8013 ( .C1(n6126), .C2(n10129), .A(n6271), .B(n6270), .ZN(n6272)
         );
  AOI21_X1 U8014 ( .B1(n10039), .B2(n6337), .A(n6272), .ZN(n9584) );
  OR2_X1 U8015 ( .A1(n10128), .A2(n9584), .ZN(n6955) );
  NAND2_X1 U8016 ( .A1(n10128), .A2(n9584), .ZN(n6952) );
  NAND2_X1 U8017 ( .A1(n8269), .A2(n5036), .ZN(n6279) );
  NAND2_X1 U8018 ( .A1(n6273), .A2(n6367), .ZN(n6274) );
  XNOR2_X2 U8019 ( .A(n6275), .B(P1_IR_REG_19__SCAN_IN), .ZN(n6513) );
  AOI22_X1 U8020 ( .A1(n4406), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9872), .B2(
        n6276), .ZN(n6278) );
  INV_X1 U8021 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6280) );
  XNOR2_X1 U8022 ( .A(n6288), .B(n6280), .ZN(n10024) );
  INV_X1 U8023 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10124) );
  NAND2_X1 U8024 ( .A1(n6870), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U8025 ( .A1(n6869), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6281) );
  OAI211_X1 U8026 ( .C1(n6126), .C2(n10124), .A(n6282), .B(n6281), .ZN(n6283)
         );
  AOI21_X1 U8027 ( .B1(n10024), .B2(n6337), .A(n6283), .ZN(n9686) );
  OR2_X1 U8028 ( .A1(n10123), .A2(n9686), .ZN(n6964) );
  NAND2_X1 U8029 ( .A1(n10123), .A2(n9686), .ZN(n6961) );
  NAND2_X1 U8030 ( .A1(n6964), .A2(n6961), .ZN(n10018) );
  INV_X1 U8031 ( .A(n10018), .ZN(n10016) );
  INV_X1 U8032 ( .A(n6961), .ZN(n6284) );
  NAND2_X1 U8033 ( .A1(n8335), .A2(n5036), .ZN(n6286) );
  OR2_X1 U8034 ( .A1(n4412), .A2(n8317), .ZN(n6285) );
  AND2_X1 U8035 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n6287) );
  AOI21_X1 U8036 ( .B1(n6288), .B2(P1_REG3_REG_19__SCAN_IN), .A(
        P1_REG3_REG_20__SCAN_IN), .ZN(n6289) );
  OR2_X1 U8037 ( .A1(n6296), .A2(n6289), .ZN(n9652) );
  INV_X1 U8038 ( .A(n9652), .ZN(n10010) );
  NAND2_X1 U8039 ( .A1(n10010), .A2(n6337), .ZN(n6294) );
  INV_X1 U8040 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10183) );
  NAND2_X1 U8041 ( .A1(n6869), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U8042 ( .A1(n6481), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6290) );
  OAI211_X1 U8043 ( .C1(n6143), .C2(n10183), .A(n6291), .B(n6290), .ZN(n6292)
         );
  INV_X1 U8044 ( .A(n6292), .ZN(n6293) );
  NAND2_X1 U8045 ( .A1(n10118), .A2(n9593), .ZN(n6832) );
  INV_X1 U8046 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8630) );
  OR2_X1 U8047 ( .A1(n4412), .A2(n8630), .ZN(n6295) );
  OR2_X1 U8048 ( .A1(n6296), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6297) );
  AND2_X1 U8049 ( .A1(n6306), .A2(n6297), .ZN(n9997) );
  NAND2_X1 U8050 ( .A1(n9997), .A2(n6337), .ZN(n6302) );
  INV_X1 U8051 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10179) );
  NAND2_X1 U8052 ( .A1(n6481), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U8053 ( .A1(n6869), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6298) );
  OAI211_X1 U8054 ( .C1(n6143), .C2(n10179), .A(n6299), .B(n6298), .ZN(n6300)
         );
  INV_X1 U8055 ( .A(n6300), .ZN(n6301) );
  XNOR2_X1 U8056 ( .A(n10113), .B(n9664), .ZN(n9992) );
  INV_X1 U8057 ( .A(n9992), .ZN(n6303) );
  NAND2_X1 U8058 ( .A1(n10113), .A2(n6827), .ZN(n6962) );
  NAND2_X1 U8059 ( .A1(n8437), .A2(n5036), .ZN(n6305) );
  OR2_X1 U8060 ( .A1(n4412), .A2(n8439), .ZN(n6304) );
  INV_X1 U8061 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9667) );
  NAND2_X1 U8062 ( .A1(n6306), .A2(n9667), .ZN(n6307) );
  NAND2_X1 U8063 ( .A1(n6315), .A2(n6307), .ZN(n9662) );
  OR2_X1 U8064 ( .A1(n9662), .A2(n6384), .ZN(n6312) );
  INV_X1 U8065 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U8066 ( .A1(n6870), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U8067 ( .A1(n6869), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6308) );
  OAI211_X1 U8068 ( .C1(n6126), .C2(n10109), .A(n6309), .B(n6308), .ZN(n6310)
         );
  INV_X1 U8069 ( .A(n6310), .ZN(n6311) );
  XNOR2_X1 U8070 ( .A(n10108), .B(n9594), .ZN(n9980) );
  NAND2_X1 U8071 ( .A1(n10108), .A2(n9594), .ZN(n6831) );
  NAND2_X1 U8072 ( .A1(n8455), .A2(n5036), .ZN(n6314) );
  OR2_X1 U8073 ( .A1(n4412), .A2(n8458), .ZN(n6313) );
  NAND2_X2 U8074 ( .A1(n6314), .A2(n6313), .ZN(n10102) );
  INV_X1 U8075 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9564) );
  NAND2_X1 U8076 ( .A1(n6315), .A2(n9564), .ZN(n6316) );
  AND2_X1 U8077 ( .A1(n6323), .A2(n6316), .ZN(n9966) );
  INV_X1 U8078 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U8079 ( .A1(n6870), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U8080 ( .A1(n6481), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6317) );
  OAI211_X1 U8081 ( .C1(n6319), .C2(n6485), .A(n6318), .B(n6317), .ZN(n6320)
         );
  NAND2_X1 U8082 ( .A1(n10102), .A2(n9663), .ZN(n9945) );
  NAND2_X1 U8083 ( .A1(n6978), .A2(n9945), .ZN(n6893) );
  NAND2_X1 U8084 ( .A1(n8488), .A2(n5036), .ZN(n6322) );
  OR2_X1 U8085 ( .A1(n4412), .A2(n8490), .ZN(n6321) );
  INV_X1 U8086 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9639) );
  AND2_X1 U8087 ( .A1(n6323), .A2(n9639), .ZN(n6324) );
  NOR2_X2 U8088 ( .A1(n6323), .A2(n9639), .ZN(n6332) );
  INV_X1 U8089 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10098) );
  NAND2_X1 U8090 ( .A1(n6869), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U8091 ( .A1(n6870), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6325) );
  OAI211_X1 U8092 ( .C1(n6126), .C2(n10098), .A(n6326), .B(n6325), .ZN(n6327)
         );
  NAND2_X1 U8093 ( .A1(n10097), .A2(n9604), .ZN(n6983) );
  INV_X1 U8094 ( .A(n9945), .ZN(n6328) );
  NOR2_X1 U8095 ( .A1(n9944), .A2(n6328), .ZN(n6329) );
  NAND2_X1 U8096 ( .A1(n8577), .A2(n5036), .ZN(n6331) );
  OR2_X1 U8097 ( .A1(n4412), .A2(n8582), .ZN(n6330) );
  OR2_X1 U8098 ( .A1(n6332), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6333) );
  INV_X1 U8099 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7684) );
  NAND2_X1 U8100 ( .A1(n6869), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U8101 ( .A1(n6870), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6334) );
  OAI211_X1 U8102 ( .C1(n6126), .C2(n7684), .A(n6335), .B(n6334), .ZN(n6336)
         );
  OR2_X1 U8103 ( .A1(n10091), .A2(n9702), .ZN(n6992) );
  NAND2_X1 U8104 ( .A1(n10091), .A2(n9702), .ZN(n6994) );
  NAND2_X1 U8105 ( .A1(n6992), .A2(n6994), .ZN(n9935) );
  INV_X1 U8106 ( .A(n6825), .ZN(n9936) );
  NOR2_X1 U8107 ( .A1(n9935), .A2(n9936), .ZN(n6338) );
  NAND2_X1 U8108 ( .A1(n8593), .A2(n5036), .ZN(n6340) );
  OR2_X1 U8109 ( .A1(n4412), .A2(n10225), .ZN(n6339) );
  NAND2_X1 U8110 ( .A1(n6481), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6346) );
  INV_X1 U8111 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10165) );
  OR2_X1 U8112 ( .A1(n6143), .A2(n10165), .ZN(n6345) );
  OAI21_X1 U8113 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n6342), .A(n6354), .ZN(
        n9920) );
  OR2_X1 U8114 ( .A1(n6384), .A2(n9920), .ZN(n6344) );
  INV_X1 U8115 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9921) );
  OR2_X1 U8116 ( .A1(n6485), .A2(n9921), .ZN(n6343) );
  INV_X1 U8117 ( .A(n9925), .ZN(n9897) );
  NAND2_X1 U8118 ( .A1(n6481), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6350) );
  INV_X1 U8119 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10162) );
  OR2_X1 U8120 ( .A1(n6143), .A2(n10162), .ZN(n6349) );
  INV_X1 U8121 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8635) );
  XNOR2_X1 U8122 ( .A(n6354), .B(n8635), .ZN(n9910) );
  OR2_X1 U8123 ( .A1(n6384), .A2(n9910), .ZN(n6348) );
  INV_X1 U8124 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9901) );
  OR2_X1 U8125 ( .A1(n6485), .A2(n9901), .ZN(n6347) );
  INV_X1 U8126 ( .A(n9704), .ZN(n9730) );
  INV_X1 U8127 ( .A(n6351), .ZN(n7002) );
  INV_X1 U8128 ( .A(n6829), .ZN(n6352) );
  NAND2_X1 U8129 ( .A1(n8639), .A2(n5036), .ZN(n6353) );
  NOR2_X1 U8130 ( .A1(n4412), .A2(n8640), .ZN(n6363) );
  INV_X1 U8131 ( .A(n6363), .ZN(n6365) );
  NAND2_X1 U8132 ( .A1(n6481), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6362) );
  INV_X1 U8133 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7670) );
  OR2_X1 U8134 ( .A1(n6143), .A2(n7670), .ZN(n6361) );
  INV_X1 U8135 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7714) );
  OAI21_X1 U8136 ( .B1(n6354), .B2(n8635), .A(n7714), .ZN(n6357) );
  AND2_X1 U8137 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6355) );
  NAND2_X1 U8138 ( .A1(n6356), .A2(n6355), .ZN(n8619) );
  NAND2_X1 U8139 ( .A1(n6357), .A2(n8619), .ZN(n9888) );
  OR2_X1 U8140 ( .A1(n6384), .A2(n9888), .ZN(n6360) );
  INV_X1 U8141 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6358) );
  OR2_X1 U8142 ( .A1(n6485), .A2(n6358), .ZN(n6359) );
  NAND4_X1 U8143 ( .A1(n6362), .A2(n6361), .A3(n6360), .A4(n6359), .ZN(n9729)
         );
  OR2_X1 U8144 ( .A1(n8639), .A2(n6363), .ZN(n6366) );
  XNOR2_X1 U8145 ( .A(n6459), .B(n6897), .ZN(n6391) );
  NAND2_X1 U8146 ( .A1(n6368), .A2(n6367), .ZN(n6372) );
  NAND2_X1 U8147 ( .A1(n6370), .A2(n6369), .ZN(n6371) );
  NAND2_X1 U8148 ( .A1(n9872), .A2(n7024), .ZN(n6383) );
  XNOR2_X2 U8149 ( .A(n6378), .B(n6377), .ZN(n8628) );
  NAND2_X1 U8150 ( .A1(n6379), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6380) );
  MUX2_X1 U8151 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6380), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n6381) );
  NAND2_X1 U8152 ( .A1(n4966), .A2(n7042), .ZN(n6382) );
  NAND2_X1 U8153 ( .A1(n7322), .A2(n7831), .ZN(n9701) );
  OR2_X1 U8154 ( .A1(n9704), .A2(n9701), .ZN(n6390) );
  NAND2_X1 U8155 ( .A1(n6870), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U8156 ( .A1(n6481), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6387) );
  OR2_X1 U8157 ( .A1(n6384), .A2(n8619), .ZN(n6386) );
  INV_X1 U8158 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8620) );
  OR2_X1 U8159 ( .A1(n6485), .A2(n8620), .ZN(n6385) );
  NAND4_X1 U8160 ( .A1(n6388), .A2(n6387), .A3(n6386), .A4(n6385), .ZN(n9728)
         );
  NAND2_X1 U8161 ( .A1(n7322), .A2(n6115), .ZN(n9703) );
  NAND2_X1 U8162 ( .A1(n9728), .A2(n9649), .ZN(n6389) );
  NAND2_X1 U8163 ( .A1(n6390), .A2(n6389), .ZN(n6772) );
  OR2_X1 U8164 ( .A1(n10408), .A2(n6526), .ZN(n10409) );
  INV_X1 U8165 ( .A(n8004), .ZN(n10446) );
  INV_X2 U8166 ( .A(n10389), .ZN(n6392) );
  NAND2_X1 U8167 ( .A1(n10484), .A2(n6393), .ZN(n6394) );
  INV_X1 U8168 ( .A(n10317), .ZN(n10499) );
  INV_X1 U8169 ( .A(n10147), .ZN(n8508) );
  AND2_X2 U8170 ( .A1(n10067), .A2(n10054), .ZN(n10036) );
  INV_X1 U8171 ( .A(n10128), .ZN(n10042) );
  AND2_X2 U8172 ( .A1(n9996), .A2(n9988), .ZN(n9963) );
  AND2_X2 U8173 ( .A1(n9963), .A2(n9968), .ZN(n9964) );
  OAI211_X1 U8174 ( .C1(n9891), .C2(n9900), .A(n10390), .B(n6490), .ZN(n9887)
         );
  INV_X1 U8175 ( .A(n7455), .ZN(n7483) );
  NAND2_X1 U8176 ( .A1(n6778), .A2(n10490), .ZN(n6396) );
  NAND2_X1 U8177 ( .A1(n6398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U8178 ( .A1(n8580), .A2(P1_B_REG_SCAN_IN), .ZN(n6407) );
  INV_X1 U8179 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U8180 ( .A1(n6402), .A2(n6401), .ZN(n6403) );
  MUX2_X1 U8181 ( .A(P1_B_REG_SCAN_IN), .B(n6407), .S(n8489), .Z(n6411) );
  NAND2_X1 U8182 ( .A1(n4486), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6409) );
  INV_X1 U8183 ( .A(n10227), .ZN(n6410) );
  NAND2_X1 U8184 ( .A1(n10227), .A2(n8580), .ZN(n10210) );
  OAI21_X1 U8185 ( .B1(n10208), .B2(P1_D_REG_1__SCAN_IN), .A(n10210), .ZN(
        n6424) );
  NAND2_X1 U8186 ( .A1(n6412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6413) );
  NOR4_X1 U8187 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6417) );
  NOR4_X1 U8188 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6416) );
  NOR4_X1 U8189 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6415) );
  NOR4_X1 U8190 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6414) );
  NAND4_X1 U8191 ( .A1(n6417), .A2(n6416), .A3(n6415), .A4(n6414), .ZN(n6422)
         );
  NOR2_X1 U8192 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .ZN(
        n7573) );
  NOR4_X1 U8193 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6420) );
  NOR4_X1 U8194 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6419) );
  NOR4_X1 U8195 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6418) );
  NAND4_X1 U8196 ( .A1(n7573), .A2(n6420), .A3(n6419), .A4(n6418), .ZN(n6421)
         );
  NOR2_X1 U8197 ( .A1(n6422), .A2(n6421), .ZN(n6751) );
  OR2_X1 U8198 ( .A1(n10208), .A2(n6751), .ZN(n6423) );
  NAND4_X1 U8199 ( .A1(n6424), .A2(n7534), .A3(n6423), .A4(n6759), .ZN(n6783)
         );
  NAND2_X1 U8200 ( .A1(n8489), .A2(n10227), .ZN(n10211) );
  NAND2_X1 U8201 ( .A1(n7335), .A2(n7953), .ZN(n7957) );
  NAND2_X1 U8202 ( .A1(n7959), .A2(n7957), .ZN(n6427) );
  INV_X1 U8203 ( .A(n6511), .ZN(n7451) );
  NAND2_X1 U8204 ( .A1(n7451), .A2(n10429), .ZN(n6426) );
  NAND2_X1 U8205 ( .A1(n6427), .A2(n6426), .ZN(n10405) );
  XNOR2_X1 U8206 ( .A(n6526), .B(n8100), .ZN(n10406) );
  NAND2_X1 U8207 ( .A1(n10405), .A2(n10406), .ZN(n6429) );
  OR2_X1 U8208 ( .A1(n4735), .A2(n6526), .ZN(n6428) );
  NAND2_X1 U8209 ( .A1(n6429), .A2(n6428), .ZN(n8102) );
  NAND2_X1 U8210 ( .A1(n8102), .A2(n8103), .ZN(n6432) );
  INV_X1 U8211 ( .A(n7999), .ZN(n9752) );
  OR2_X1 U8212 ( .A1(n9752), .A2(n6539), .ZN(n6431) );
  NAND2_X1 U8213 ( .A1(n6432), .A2(n6431), .ZN(n10387) );
  INV_X1 U8214 ( .A(n6433), .ZN(n6798) );
  NAND2_X1 U8215 ( .A1(n6798), .A2(n6434), .ZN(n10388) );
  NAND2_X1 U8216 ( .A1(n10387), .A2(n10388), .ZN(n6436) );
  NAND2_X1 U8217 ( .A1(n10446), .A2(n9750), .ZN(n6435) );
  INV_X1 U8218 ( .A(n8181), .ZN(n9749) );
  OR2_X1 U8219 ( .A1(n8094), .A2(n9749), .ZN(n6437) );
  INV_X1 U8220 ( .A(n8293), .ZN(n9748) );
  INV_X1 U8221 ( .A(n8288), .ZN(n6438) );
  INV_X1 U8222 ( .A(n8566), .ZN(n9746) );
  NAND2_X1 U8223 ( .A1(n6919), .A2(n6927), .ZN(n10354) );
  INV_X1 U8224 ( .A(n8417), .ZN(n9742) );
  INV_X1 U8225 ( .A(n10143), .ZN(n9726) );
  NAND2_X1 U8226 ( .A1(n8596), .A2(n5277), .ZN(n6440) );
  NAND2_X1 U8227 ( .A1(n10042), .A2(n9584), .ZN(n6442) );
  INV_X1 U8228 ( .A(n9584), .ZN(n9735) );
  INV_X1 U8229 ( .A(n9686), .ZN(n9734) );
  NAND2_X1 U8230 ( .A1(n10123), .A2(n9734), .ZN(n6443) );
  INV_X1 U8231 ( .A(n10123), .ZN(n10027) );
  INV_X1 U8232 ( .A(n10118), .ZN(n10013) );
  NAND2_X1 U8233 ( .A1(n10013), .A2(n9593), .ZN(n6445) );
  NOR2_X1 U8234 ( .A1(n10013), .A2(n9593), .ZN(n6444) );
  NAND2_X1 U8235 ( .A1(n10108), .A2(n9733), .ZN(n6446) );
  INV_X1 U8236 ( .A(n6446), .ZN(n9961) );
  AOI22_X1 U8237 ( .A1(n9968), .A2(n9663), .B1(n9594), .B2(n9988), .ZN(n6448)
         );
  NOR2_X1 U8238 ( .A1(n10113), .A2(n9664), .ZN(n9958) );
  NAND2_X1 U8239 ( .A1(n9958), .A2(n6446), .ZN(n6447) );
  INV_X1 U8240 ( .A(n9663), .ZN(n6449) );
  INV_X1 U8241 ( .A(n10091), .ZN(n9933) );
  NOR2_X1 U8242 ( .A1(n9933), .A2(n9702), .ZN(n6450) );
  INV_X1 U8243 ( .A(n9702), .ZN(n9732) );
  INV_X1 U8244 ( .A(n9603), .ZN(n9731) );
  AND2_X1 U8245 ( .A1(n10087), .A2(n9731), .ZN(n9898) );
  NOR2_X1 U8246 ( .A1(n5128), .A2(n9898), .ZN(n6451) );
  NOR2_X1 U8247 ( .A1(n9925), .A2(n9898), .ZN(n6453) );
  NOR2_X1 U8248 ( .A1(n10083), .A2(n9730), .ZN(n6452) );
  AOI21_X1 U8249 ( .B1(n9904), .B2(n6453), .A(n6452), .ZN(n6495) );
  NAND2_X1 U8250 ( .A1(n6503), .A2(n6495), .ZN(n6454) );
  INV_X1 U8251 ( .A(n7044), .ZN(n6770) );
  NAND2_X1 U8252 ( .A1(n6770), .A2(n7322), .ZN(n7450) );
  OR2_X1 U8253 ( .A1(n9872), .A2(n8438), .ZN(n6455) );
  AOI21_X1 U8254 ( .B1(n7044), .B2(n6455), .A(n7483), .ZN(n6456) );
  NAND2_X1 U8255 ( .A1(n7450), .A2(n6456), .ZN(n8297) );
  OR2_X1 U8256 ( .A1(n6515), .A2(n7024), .ZN(n10492) );
  NOR2_X1 U8257 ( .A1(n10526), .A2(n10153), .ZN(n10080) );
  NAND2_X1 U8258 ( .A1(n6458), .A2(n6457), .ZN(P1_U3550) );
  INV_X1 U8259 ( .A(n6467), .ZN(n6468) );
  NAND2_X1 U8260 ( .A1(n6468), .A2(SI_28_), .ZN(n6461) );
  INV_X1 U8261 ( .A(n6848), .ZN(n6460) );
  AND2_X1 U8262 ( .A1(n6461), .A2(n6460), .ZN(n6473) );
  INV_X1 U8263 ( .A(n6473), .ZN(n6462) );
  INV_X1 U8264 ( .A(SI_28_), .ZN(n6463) );
  NAND2_X1 U8265 ( .A1(n6467), .A2(n6463), .ZN(n6847) );
  INV_X1 U8266 ( .A(n6466), .ZN(n6472) );
  OAI21_X1 U8267 ( .B1(n6848), .B2(SI_28_), .A(n6467), .ZN(n6471) );
  NAND2_X1 U8268 ( .A1(n6848), .A2(SI_28_), .ZN(n6469) );
  NAND2_X1 U8269 ( .A1(n6469), .A2(n6468), .ZN(n6470) );
  AOI22_X1 U8270 ( .A1(n6473), .A2(n6472), .B1(n6471), .B2(n6470), .ZN(n6474)
         );
  INV_X1 U8271 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10223) );
  NOR2_X1 U8272 ( .A1(n4412), .A2(n10223), .ZN(n6477) );
  AND2_X1 U8273 ( .A1(n8618), .A2(n9728), .ZN(n7005) );
  INV_X1 U8274 ( .A(n9728), .ZN(n6478) );
  XNOR2_X1 U8275 ( .A(n6479), .B(n7008), .ZN(n6489) );
  NAND2_X1 U8276 ( .A1(n9729), .A2(n9687), .ZN(n6487) );
  INV_X1 U8277 ( .A(P1_B_REG_SCAN_IN), .ZN(n7046) );
  NOR2_X1 U8278 ( .A1(n6123), .A2(n7046), .ZN(n6480) );
  NOR2_X1 U8279 ( .A1(n9703), .A2(n6480), .ZN(n9879) );
  INV_X1 U8280 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n6484) );
  NAND2_X1 U8281 ( .A1(n6481), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U8282 ( .A1(n6870), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6482) );
  OAI211_X1 U8283 ( .C1(n6485), .C2(n6484), .A(n6483), .B(n6482), .ZN(n9727)
         );
  NAND2_X1 U8284 ( .A1(n9879), .A2(n9727), .ZN(n6486) );
  AOI21_X1 U8285 ( .B1(n10490), .B2(n6491), .A(n8623), .ZN(n6492) );
  INV_X1 U8286 ( .A(n6503), .ZN(n6494) );
  INV_X1 U8287 ( .A(n7008), .ZN(n6493) );
  NOR2_X1 U8288 ( .A1(n9891), .A2(n4609), .ZN(n6499) );
  NAND3_X1 U8289 ( .A1(n6494), .A2(n6493), .A3(n6497), .ZN(n6505) );
  AND2_X1 U8290 ( .A1(n6495), .A2(n6897), .ZN(n6496) );
  AND2_X1 U8291 ( .A1(n6496), .A2(n7008), .ZN(n6502) );
  INV_X1 U8292 ( .A(n6496), .ZN(n6498) );
  INV_X1 U8293 ( .A(n6499), .ZN(n6497) );
  AOI21_X1 U8294 ( .B1(n6498), .B2(n6497), .A(n7008), .ZN(n6501) );
  NOR2_X1 U8295 ( .A1(n6493), .A2(n6499), .ZN(n6500) );
  AOI21_X1 U8296 ( .B1(n6503), .B2(n6502), .A(n5288), .ZN(n6504) );
  NAND2_X1 U8297 ( .A1(n6505), .A2(n6504), .ZN(n8617) );
  NAND2_X1 U8298 ( .A1(n10526), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U8299 ( .A1(n6508), .A2(n6507), .ZN(P1_U3551) );
  INV_X1 U8300 ( .A(n6509), .ZN(n6510) );
  NAND2_X1 U8301 ( .A1(n6511), .A2(n6543), .ZN(n6512) );
  NAND2_X4 U8302 ( .A1(n6514), .A2(n7455), .ZN(n6746) );
  OR2_X2 U8303 ( .A1(n6515), .A2(n8628), .ZN(n8090) );
  NAND2_X1 U8304 ( .A1(n6517), .A2(n6516), .ZN(n7912) );
  NAND2_X1 U8305 ( .A1(n7953), .A2(n6543), .ZN(n6519) );
  INV_X1 U8306 ( .A(n7171), .ZN(n6764) );
  NAND2_X1 U8307 ( .A1(n6764), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U8308 ( .A1(n7953), .A2(n6525), .ZN(n6521) );
  NAND2_X1 U8309 ( .A1(n6523), .A2(n6746), .ZN(n6524) );
  XNOR2_X1 U8310 ( .A(n6528), .B(n6746), .ZN(n6533) );
  NAND2_X1 U8311 ( .A1(n6526), .A2(n6543), .ZN(n6531) );
  AND2_X1 U8312 ( .A1(n6530), .A2(n6531), .ZN(n6532) );
  NAND2_X1 U8313 ( .A1(n6533), .A2(n6532), .ZN(n6534) );
  NAND2_X1 U8314 ( .A1(n6539), .A2(n6525), .ZN(n6536) );
  OR2_X1 U8315 ( .A1(n7999), .A2(n6538), .ZN(n6535) );
  NAND2_X1 U8316 ( .A1(n6536), .A2(n6535), .ZN(n6537) );
  XNOR2_X1 U8317 ( .A(n6537), .B(n6746), .ZN(n6551) );
  NAND2_X1 U8318 ( .A1(n6539), .A2(n6732), .ZN(n6541) );
  INV_X4 U8319 ( .A(n6703), .ZN(n6745) );
  OR2_X1 U8320 ( .A1(n6745), .A2(n7999), .ZN(n6540) );
  NAND2_X1 U8321 ( .A1(n6541), .A2(n6540), .ZN(n6549) );
  NAND2_X1 U8322 ( .A1(n8004), .A2(n6525), .ZN(n6545) );
  OR2_X1 U8323 ( .A1(n9750), .A2(n6538), .ZN(n6544) );
  NAND2_X1 U8324 ( .A1(n6545), .A2(n6544), .ZN(n6546) );
  XNOR2_X1 U8325 ( .A(n6546), .B(n6746), .ZN(n6553) );
  NAND2_X1 U8326 ( .A1(n8004), .A2(n6732), .ZN(n6548) );
  OR2_X1 U8327 ( .A1(n6745), .A2(n9750), .ZN(n6547) );
  NAND2_X1 U8328 ( .A1(n6548), .A2(n6547), .ZN(n6554) );
  XNOR2_X1 U8329 ( .A(n6553), .B(n6554), .ZN(n7997) );
  INV_X1 U8330 ( .A(n6549), .ZN(n6550) );
  NAND2_X1 U8331 ( .A1(n6551), .A2(n6550), .ZN(n7995) );
  INV_X1 U8332 ( .A(n6553), .ZN(n6555) );
  NAND2_X1 U8333 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  NAND2_X1 U8334 ( .A1(n8094), .A2(n6525), .ZN(n6558) );
  OR2_X1 U8335 ( .A1(n8181), .A2(n6538), .ZN(n6557) );
  NAND2_X1 U8336 ( .A1(n6558), .A2(n6557), .ZN(n6559) );
  XNOR2_X1 U8337 ( .A(n6559), .B(n6726), .ZN(n6562) );
  NAND2_X1 U8338 ( .A1(n8094), .A2(n6732), .ZN(n6561) );
  OR2_X1 U8339 ( .A1(n6745), .A2(n8181), .ZN(n6560) );
  NAND2_X1 U8340 ( .A1(n6561), .A2(n6560), .ZN(n8156) );
  NAND2_X1 U8341 ( .A1(n8153), .A2(n8156), .ZN(n6564) );
  NAND2_X1 U8342 ( .A1(n8256), .A2(n6525), .ZN(n6566) );
  OR2_X1 U8343 ( .A1(n8293), .A2(n6538), .ZN(n6565) );
  NAND2_X1 U8344 ( .A1(n6566), .A2(n6565), .ZN(n6567) );
  XNOR2_X1 U8345 ( .A(n6567), .B(n6746), .ZN(n6570) );
  NAND2_X1 U8346 ( .A1(n8256), .A2(n6732), .ZN(n6569) );
  OR2_X1 U8347 ( .A1(n6745), .A2(n8293), .ZN(n6568) );
  AND2_X1 U8348 ( .A1(n6569), .A2(n6568), .ZN(n6571) );
  NAND2_X1 U8349 ( .A1(n6570), .A2(n6571), .ZN(n6576) );
  INV_X1 U8350 ( .A(n6570), .ZN(n6573) );
  INV_X1 U8351 ( .A(n6571), .ZN(n6572) );
  NAND2_X1 U8352 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  NAND2_X1 U8353 ( .A1(n6576), .A2(n6574), .ZN(n8251) );
  INV_X1 U8354 ( .A(n8251), .ZN(n6575) );
  NAND2_X1 U8355 ( .A1(n8332), .A2(n6525), .ZN(n6578) );
  OR2_X1 U8356 ( .A1(n8464), .A2(n6538), .ZN(n6577) );
  NAND2_X1 U8357 ( .A1(n6578), .A2(n6577), .ZN(n6579) );
  XNOR2_X1 U8358 ( .A(n6579), .B(n6746), .ZN(n6582) );
  NAND2_X1 U8359 ( .A1(n8332), .A2(n6732), .ZN(n6581) );
  OR2_X1 U8360 ( .A1(n6745), .A2(n8464), .ZN(n6580) );
  AND2_X1 U8361 ( .A1(n6581), .A2(n6580), .ZN(n6583) );
  NAND2_X1 U8362 ( .A1(n6582), .A2(n6583), .ZN(n8324) );
  INV_X1 U8363 ( .A(n6582), .ZN(n6585) );
  INV_X1 U8364 ( .A(n6583), .ZN(n6584) );
  NAND2_X1 U8365 ( .A1(n6585), .A2(n6584), .ZN(n8325) );
  NAND2_X1 U8366 ( .A1(n6101), .A2(n6525), .ZN(n6587) );
  OR2_X1 U8367 ( .A1(n8553), .A2(n6538), .ZN(n6586) );
  NAND2_X1 U8368 ( .A1(n6587), .A2(n6586), .ZN(n6588) );
  XNOR2_X1 U8369 ( .A(n6588), .B(n6746), .ZN(n8562) );
  NAND2_X1 U8370 ( .A1(n6101), .A2(n6732), .ZN(n6590) );
  OR2_X1 U8371 ( .A1(n6745), .A2(n8553), .ZN(n6589) );
  NAND2_X1 U8372 ( .A1(n6590), .A2(n6589), .ZN(n8561) );
  INV_X1 U8373 ( .A(n8561), .ZN(n6596) );
  NAND2_X1 U8374 ( .A1(n8468), .A2(n6732), .ZN(n6592) );
  OR2_X1 U8375 ( .A1(n6745), .A2(n8566), .ZN(n6591) );
  NAND2_X1 U8376 ( .A1(n6592), .A2(n6591), .ZN(n6597) );
  INV_X1 U8377 ( .A(n6597), .ZN(n8462) );
  NAND2_X1 U8378 ( .A1(n8468), .A2(n6525), .ZN(n6594) );
  OR2_X1 U8379 ( .A1(n8566), .A2(n6538), .ZN(n6593) );
  NAND2_X1 U8380 ( .A1(n6594), .A2(n6593), .ZN(n6595) );
  XNOR2_X1 U8381 ( .A(n6595), .B(n6726), .ZN(n8560) );
  INV_X1 U8382 ( .A(n8560), .ZN(n8460) );
  OAI22_X1 U8383 ( .A1(n8562), .A2(n6596), .B1(n8462), .B2(n8460), .ZN(n6601)
         );
  OAI21_X1 U8384 ( .B1(n8560), .B2(n6597), .A(n8561), .ZN(n6599) );
  NOR2_X1 U8385 ( .A1(n8561), .A2(n6597), .ZN(n6598) );
  AOI22_X1 U8386 ( .A1(n8562), .A2(n6599), .B1(n6598), .B2(n8460), .ZN(n6600)
         );
  NAND2_X1 U8387 ( .A1(n10489), .A2(n6525), .ZN(n6603) );
  OR2_X1 U8388 ( .A1(n8496), .A2(n6538), .ZN(n6602) );
  NAND2_X1 U8389 ( .A1(n6603), .A2(n6602), .ZN(n6604) );
  XNOR2_X1 U8390 ( .A(n6604), .B(n6726), .ZN(n9674) );
  NAND2_X1 U8391 ( .A1(n10489), .A2(n6732), .ZN(n6606) );
  OR2_X1 U8392 ( .A1(n6745), .A2(n8496), .ZN(n6605) );
  NAND2_X1 U8393 ( .A1(n6606), .A2(n6605), .ZN(n6615) );
  OAI22_X1 U8394 ( .A1(n10484), .A2(n6542), .B1(n6607), .B2(n6748), .ZN(n6608)
         );
  XNOR2_X1 U8395 ( .A(n6608), .B(n6726), .ZN(n6612) );
  OR2_X1 U8396 ( .A1(n10484), .A2(n6538), .ZN(n6610) );
  NAND2_X1 U8397 ( .A1(n4734), .A2(n9744), .ZN(n6609) );
  NAND2_X1 U8398 ( .A1(n6610), .A2(n6609), .ZN(n8552) );
  AOI22_X1 U8399 ( .A1(n9674), .A2(n6615), .B1(n6612), .B2(n8552), .ZN(n6611)
         );
  NAND2_X1 U8400 ( .A1(n8550), .A2(n6611), .ZN(n6620) );
  INV_X1 U8401 ( .A(n9674), .ZN(n6618) );
  INV_X1 U8402 ( .A(n6612), .ZN(n9672) );
  INV_X1 U8403 ( .A(n8552), .ZN(n6613) );
  NAND2_X1 U8404 ( .A1(n9672), .A2(n6613), .ZN(n6614) );
  NAND2_X1 U8405 ( .A1(n6614), .A2(n6615), .ZN(n6617) );
  INV_X1 U8406 ( .A(n6614), .ZN(n6616) );
  INV_X1 U8407 ( .A(n6615), .ZN(n9673) );
  AOI22_X1 U8408 ( .A1(n6618), .A2(n6617), .B1(n6616), .B2(n9673), .ZN(n6619)
         );
  NAND2_X1 U8409 ( .A1(n6620), .A2(n6619), .ZN(n8495) );
  NAND2_X1 U8410 ( .A1(n10317), .A2(n6525), .ZN(n6622) );
  OR2_X1 U8411 ( .A1(n8417), .A2(n6538), .ZN(n6621) );
  NAND2_X1 U8412 ( .A1(n6622), .A2(n6621), .ZN(n6623) );
  XNOR2_X1 U8413 ( .A(n6623), .B(n6726), .ZN(n6625) );
  NOR2_X1 U8414 ( .A1(n8417), .A2(n6745), .ZN(n6624) );
  AOI21_X1 U8415 ( .B1(n10317), .B2(n6732), .A(n6624), .ZN(n6626) );
  XNOR2_X1 U8416 ( .A(n6625), .B(n6626), .ZN(n8494) );
  NAND2_X1 U8417 ( .A1(n8495), .A2(n8494), .ZN(n6629) );
  INV_X1 U8418 ( .A(n6625), .ZN(n6627) );
  NAND2_X1 U8419 ( .A1(n6627), .A2(n6626), .ZN(n6628) );
  NAND2_X1 U8420 ( .A1(n6629), .A2(n6628), .ZN(n8584) );
  NAND2_X1 U8421 ( .A1(n8590), .A2(n6525), .ZN(n6631) );
  OR2_X1 U8422 ( .A1(n8511), .A2(n6748), .ZN(n6630) );
  NAND2_X1 U8423 ( .A1(n6631), .A2(n6630), .ZN(n6632) );
  XNOR2_X1 U8424 ( .A(n6632), .B(n6726), .ZN(n6634) );
  NOR2_X1 U8425 ( .A1(n8511), .A2(n6745), .ZN(n6633) );
  AOI21_X1 U8426 ( .B1(n8590), .B2(n6543), .A(n6633), .ZN(n6635) );
  XNOR2_X1 U8427 ( .A(n6634), .B(n6635), .ZN(n8583) );
  NAND2_X1 U8428 ( .A1(n8584), .A2(n8583), .ZN(n6638) );
  INV_X1 U8429 ( .A(n6634), .ZN(n6636) );
  NAND2_X1 U8430 ( .A1(n6636), .A2(n6635), .ZN(n6637) );
  NAND2_X1 U8431 ( .A1(n10147), .A2(n6525), .ZN(n6640) );
  NAND2_X1 U8432 ( .A1(n9740), .A2(n6732), .ZN(n6639) );
  NAND2_X1 U8433 ( .A1(n6640), .A2(n6639), .ZN(n6641) );
  XNOR2_X1 U8434 ( .A(n6641), .B(n6726), .ZN(n6650) );
  INV_X1 U8435 ( .A(n6650), .ZN(n9610) );
  NAND2_X1 U8436 ( .A1(n10147), .A2(n6732), .ZN(n6643) );
  NAND2_X1 U8437 ( .A1(n9740), .A2(n4734), .ZN(n6642) );
  NAND2_X1 U8438 ( .A1(n6643), .A2(n6642), .ZN(n9552) );
  INV_X1 U8439 ( .A(n9552), .ZN(n6644) );
  NAND2_X1 U8440 ( .A1(n10143), .A2(n6525), .ZN(n6646) );
  NAND2_X1 U8441 ( .A1(n9739), .A2(n6732), .ZN(n6645) );
  NAND2_X1 U8442 ( .A1(n6646), .A2(n6645), .ZN(n6647) );
  XNOR2_X1 U8443 ( .A(n6647), .B(n6726), .ZN(n9614) );
  NAND2_X1 U8444 ( .A1(n10143), .A2(n6732), .ZN(n6649) );
  NAND2_X1 U8445 ( .A1(n9739), .A2(n4734), .ZN(n6648) );
  NAND2_X1 U8446 ( .A1(n6649), .A2(n6648), .ZN(n9612) );
  AOI22_X1 U8447 ( .A1(n9614), .A2(n9612), .B1(n6650), .B2(n9552), .ZN(n6655)
         );
  OAI22_X1 U8448 ( .A1(n6250), .A2(n6542), .B1(n6651), .B2(n6748), .ZN(n6652)
         );
  XNOR2_X1 U8449 ( .A(n6652), .B(n6726), .ZN(n9617) );
  OR2_X1 U8450 ( .A1(n6250), .A2(n6748), .ZN(n6654) );
  NAND2_X1 U8451 ( .A1(n9737), .A2(n4734), .ZN(n6653) );
  NAND2_X1 U8452 ( .A1(n6654), .A2(n6653), .ZN(n9616) );
  NAND2_X1 U8453 ( .A1(n9617), .A2(n9616), .ZN(n9615) );
  INV_X1 U8454 ( .A(n9617), .ZN(n6658) );
  OAI21_X1 U8455 ( .B1(n9614), .B2(n9612), .A(n9616), .ZN(n6657) );
  NOR2_X1 U8456 ( .A1(n9616), .A2(n9612), .ZN(n6656) );
  INV_X1 U8457 ( .A(n9614), .ZN(n9611) );
  AOI22_X1 U8458 ( .A1(n6658), .A2(n6657), .B1(n6656), .B2(n9611), .ZN(n6659)
         );
  OAI22_X1 U8459 ( .A1(n10054), .A2(n6542), .B1(n6661), .B2(n6748), .ZN(n6660)
         );
  XNOR2_X1 U8460 ( .A(n6660), .B(n6726), .ZN(n6662) );
  OAI22_X1 U8461 ( .A1(n10054), .A2(n6748), .B1(n6661), .B2(n6745), .ZN(n6663)
         );
  NAND2_X1 U8462 ( .A1(n6662), .A2(n6663), .ZN(n9625) );
  INV_X1 U8463 ( .A(n6662), .ZN(n6665) );
  INV_X1 U8464 ( .A(n6663), .ZN(n6664) );
  NAND2_X1 U8465 ( .A1(n6665), .A2(n6664), .ZN(n9624) );
  NAND2_X1 U8466 ( .A1(n10123), .A2(n6525), .ZN(n6668) );
  OR2_X1 U8467 ( .A1(n9686), .A2(n6748), .ZN(n6667) );
  NAND2_X1 U8468 ( .A1(n6668), .A2(n6667), .ZN(n6669) );
  XNOR2_X1 U8469 ( .A(n6669), .B(n6726), .ZN(n9581) );
  NAND2_X1 U8470 ( .A1(n10123), .A2(n6732), .ZN(n6671) );
  OR2_X1 U8471 ( .A1(n9686), .A2(n6745), .ZN(n6670) );
  NAND2_X1 U8472 ( .A1(n6671), .A2(n6670), .ZN(n6678) );
  NAND2_X1 U8473 ( .A1(n10128), .A2(n6525), .ZN(n6673) );
  OR2_X1 U8474 ( .A1(n9584), .A2(n6748), .ZN(n6672) );
  NAND2_X1 U8475 ( .A1(n6673), .A2(n6672), .ZN(n6674) );
  XNOR2_X1 U8476 ( .A(n6674), .B(n6726), .ZN(n6680) );
  NAND2_X1 U8477 ( .A1(n10128), .A2(n6732), .ZN(n6676) );
  OR2_X1 U8478 ( .A1(n9584), .A2(n6745), .ZN(n6675) );
  NAND2_X1 U8479 ( .A1(n6676), .A2(n6675), .ZN(n9685) );
  OAI22_X1 U8480 ( .A1(n9581), .A2(n6678), .B1(n6680), .B2(n9685), .ZN(n6683)
         );
  INV_X1 U8481 ( .A(n6680), .ZN(n9579) );
  INV_X1 U8482 ( .A(n9685), .ZN(n6677) );
  INV_X1 U8483 ( .A(n6678), .ZN(n9580) );
  OAI21_X1 U8484 ( .B1(n9579), .B2(n6677), .A(n9580), .ZN(n6681) );
  AND2_X1 U8485 ( .A1(n6678), .A2(n9685), .ZN(n6679) );
  AOI22_X1 U8486 ( .A1(n6681), .A2(n9581), .B1(n6680), .B2(n6679), .ZN(n6682)
         );
  NAND2_X1 U8487 ( .A1(n10118), .A2(n6525), .ZN(n6685) );
  OR2_X1 U8488 ( .A1(n9593), .A2(n6748), .ZN(n6684) );
  NAND2_X1 U8489 ( .A1(n6685), .A2(n6684), .ZN(n6686) );
  XNOR2_X1 U8490 ( .A(n6686), .B(n6746), .ZN(n9646) );
  NOR2_X1 U8491 ( .A1(n9593), .A2(n6745), .ZN(n6687) );
  AOI21_X1 U8492 ( .B1(n10118), .B2(n6543), .A(n6687), .ZN(n6689) );
  NAND2_X1 U8493 ( .A1(n9646), .A2(n6689), .ZN(n6688) );
  INV_X1 U8494 ( .A(n9646), .ZN(n6690) );
  INV_X1 U8495 ( .A(n6689), .ZN(n9645) );
  NAND2_X1 U8496 ( .A1(n6690), .A2(n9645), .ZN(n6691) );
  NAND2_X1 U8497 ( .A1(n10113), .A2(n6525), .ZN(n6693) );
  NAND2_X1 U8498 ( .A1(n9664), .A2(n6732), .ZN(n6692) );
  NAND2_X1 U8499 ( .A1(n6693), .A2(n6692), .ZN(n6694) );
  XNOR2_X1 U8500 ( .A(n6694), .B(n6746), .ZN(n6698) );
  NOR2_X1 U8501 ( .A1(n6827), .A2(n6745), .ZN(n6695) );
  AOI21_X1 U8502 ( .B1(n10113), .B2(n6732), .A(n6695), .ZN(n6697) );
  XNOR2_X1 U8503 ( .A(n6698), .B(n6697), .ZN(n9592) );
  INV_X1 U8504 ( .A(n9592), .ZN(n6696) );
  NAND2_X1 U8505 ( .A1(n6698), .A2(n6697), .ZN(n6699) );
  NAND2_X1 U8506 ( .A1(n10108), .A2(n6525), .ZN(n6701) );
  NAND2_X1 U8507 ( .A1(n9733), .A2(n6732), .ZN(n6700) );
  NAND2_X1 U8508 ( .A1(n6701), .A2(n6700), .ZN(n6702) );
  XNOR2_X1 U8509 ( .A(n6702), .B(n6746), .ZN(n6706) );
  NAND2_X1 U8510 ( .A1(n10108), .A2(n6732), .ZN(n6705) );
  NAND2_X1 U8511 ( .A1(n9733), .A2(n4734), .ZN(n6704) );
  NAND2_X1 U8512 ( .A1(n6705), .A2(n6704), .ZN(n9657) );
  AND2_X2 U8513 ( .A1(n6707), .A2(n6706), .ZN(n9660) );
  NAND2_X1 U8514 ( .A1(n10102), .A2(n6525), .ZN(n6709) );
  OR2_X1 U8515 ( .A1(n9663), .A2(n6748), .ZN(n6708) );
  NAND2_X1 U8516 ( .A1(n6709), .A2(n6708), .ZN(n6710) );
  XNOR2_X1 U8517 ( .A(n6710), .B(n6746), .ZN(n6713) );
  NOR2_X1 U8518 ( .A1(n9663), .A2(n6745), .ZN(n6711) );
  AOI21_X1 U8519 ( .B1(n10102), .B2(n6543), .A(n6711), .ZN(n6712) );
  NAND2_X1 U8520 ( .A1(n6713), .A2(n6712), .ZN(n9633) );
  OR2_X1 U8521 ( .A1(n6713), .A2(n6712), .ZN(n6714) );
  AND2_X1 U8522 ( .A1(n9633), .A2(n6714), .ZN(n9559) );
  NAND2_X1 U8523 ( .A1(n10097), .A2(n6525), .ZN(n6716) );
  OR2_X1 U8524 ( .A1(n9604), .A2(n6748), .ZN(n6715) );
  NAND2_X1 U8525 ( .A1(n6716), .A2(n6715), .ZN(n6717) );
  XNOR2_X1 U8526 ( .A(n6717), .B(n6746), .ZN(n6720) );
  NOR2_X1 U8527 ( .A1(n9604), .A2(n6745), .ZN(n6718) );
  AOI21_X1 U8528 ( .B1(n10097), .B2(n6543), .A(n6718), .ZN(n6719) );
  NAND2_X1 U8529 ( .A1(n6720), .A2(n6719), .ZN(n6722) );
  OR2_X1 U8530 ( .A1(n6720), .A2(n6719), .ZN(n6721) );
  NAND2_X1 U8531 ( .A1(n6722), .A2(n6721), .ZN(n9632) );
  INV_X1 U8532 ( .A(n6722), .ZN(n6723) );
  NAND2_X1 U8533 ( .A1(n10091), .A2(n6525), .ZN(n6725) );
  OR2_X1 U8534 ( .A1(n9702), .A2(n6748), .ZN(n6724) );
  NAND2_X1 U8535 ( .A1(n6725), .A2(n6724), .ZN(n6727) );
  XNOR2_X1 U8536 ( .A(n6727), .B(n6726), .ZN(n6734) );
  OAI22_X1 U8537 ( .A1(n9933), .A2(n6748), .B1(n9702), .B2(n6745), .ZN(n6733)
         );
  XNOR2_X1 U8538 ( .A(n6734), .B(n6733), .ZN(n9602) );
  NAND2_X1 U8539 ( .A1(n10087), .A2(n6525), .ZN(n6729) );
  OR2_X1 U8540 ( .A1(n9603), .A2(n6748), .ZN(n6728) );
  NAND2_X1 U8541 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  XNOR2_X1 U8542 ( .A(n6730), .B(n6746), .ZN(n6735) );
  NOR2_X1 U8543 ( .A1(n9603), .A2(n6745), .ZN(n6731) );
  AOI21_X1 U8544 ( .B1(n10087), .B2(n6732), .A(n6731), .ZN(n6736) );
  XNOR2_X1 U8545 ( .A(n6735), .B(n6736), .ZN(n9697) );
  NOR2_X1 U8546 ( .A1(n6734), .A2(n6733), .ZN(n9698) );
  INV_X1 U8547 ( .A(n6735), .ZN(n6738) );
  INV_X1 U8548 ( .A(n6736), .ZN(n6737) );
  NAND2_X1 U8549 ( .A1(n10083), .A2(n6525), .ZN(n6740) );
  OR2_X1 U8550 ( .A1(n9704), .A2(n6748), .ZN(n6739) );
  NAND2_X1 U8551 ( .A1(n6740), .A2(n6739), .ZN(n6741) );
  XNOR2_X1 U8552 ( .A(n6741), .B(n6746), .ZN(n6744) );
  NOR2_X1 U8553 ( .A1(n9704), .A2(n6745), .ZN(n6742) );
  AOI21_X1 U8554 ( .B1(n10083), .B2(n6543), .A(n6742), .ZN(n6743) );
  NAND2_X1 U8555 ( .A1(n6744), .A2(n6743), .ZN(n6774) );
  OAI21_X1 U8556 ( .B1(n6744), .B2(n6743), .A(n6774), .ZN(n8632) );
  OAI22_X1 U8557 ( .A1(n9891), .A2(n6748), .B1(n4609), .B2(n6745), .ZN(n6747)
         );
  XNOR2_X1 U8558 ( .A(n6747), .B(n6746), .ZN(n6750) );
  OAI22_X1 U8559 ( .A1(n9891), .A2(n6542), .B1(n4609), .B2(n6748), .ZN(n6749)
         );
  XNOR2_X1 U8560 ( .A(n6750), .B(n6749), .ZN(n6756) );
  INV_X1 U8561 ( .A(n6756), .ZN(n6775) );
  AND2_X1 U8562 ( .A1(n6751), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6752) );
  OR2_X1 U8563 ( .A1(n10208), .A2(n6752), .ZN(n6753) );
  NAND2_X1 U8564 ( .A1(n6782), .A2(n7449), .ZN(n6763) );
  OR2_X1 U8565 ( .A1(n10490), .A2(n7322), .ZN(n6754) );
  NAND3_X1 U8566 ( .A1(n6775), .A2(n9716), .A3(n6774), .ZN(n6755) );
  NAND3_X1 U8567 ( .A1(n8634), .A2(n6756), .A3(n9716), .ZN(n6780) );
  INV_X1 U8568 ( .A(n9891), .ZN(n6778) );
  OR2_X1 U8569 ( .A1(n7455), .A2(n7023), .ZN(n7952) );
  INV_X1 U8570 ( .A(n7952), .ZN(n6758) );
  NAND2_X1 U8571 ( .A1(n6771), .A2(n6758), .ZN(n6761) );
  NAND2_X1 U8572 ( .A1(n7042), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8315) );
  NAND2_X1 U8573 ( .A1(n10490), .A2(n8315), .ZN(n6762) );
  NAND2_X1 U8574 ( .A1(n6763), .A2(n6762), .ZN(n7535) );
  NOR2_X1 U8575 ( .A1(n6765), .A2(n6764), .ZN(n6766) );
  NAND2_X1 U8576 ( .A1(n7535), .A2(n6766), .ZN(n6767) );
  NAND2_X1 U8577 ( .A1(n6767), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6769) );
  AND2_X1 U8578 ( .A1(n6768), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7047) );
  AOI22_X1 U8579 ( .A1(n9710), .A2(n6772), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6773) );
  OAI21_X1 U8580 ( .B1(n9708), .B2(n9888), .A(n6773), .ZN(n6777) );
  NOR3_X1 U8581 ( .A1(n6775), .A2(n9695), .A3(n6774), .ZN(n6776) );
  AOI211_X1 U8582 ( .C1(n6778), .C2(n9693), .A(n6777), .B(n6776), .ZN(n6779)
         );
  NAND3_X1 U8583 ( .A1(n6781), .A2(n6780), .A3(n6779), .ZN(P1_U3220) );
  NAND2_X1 U8584 ( .A1(n6785), .A2(n6784), .ZN(P1_U3519) );
  INV_X1 U8585 ( .A(n9398), .ZN(n6792) );
  AOI22_X1 U8586 ( .A1(n9233), .A2(n8797), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6789) );
  OAI21_X1 U8587 ( .B1(n8701), .B2(n8782), .A(n6789), .ZN(n6790) );
  AOI21_X1 U8588 ( .B1(n9237), .B2(n8779), .A(n6790), .ZN(n6791) );
  OAI21_X1 U8589 ( .B1(n6792), .B2(n8800), .A(n6791), .ZN(n6793) );
  INV_X1 U8590 ( .A(n6793), .ZN(n6794) );
  INV_X1 U8591 ( .A(n7005), .ZN(n6898) );
  AND2_X1 U8592 ( .A1(n6898), .A2(n6795), .ZN(n7029) );
  NAND2_X1 U8593 ( .A1(n6813), .A2(n6796), .ZN(n6948) );
  OR2_X1 U8594 ( .A1(n6948), .A2(n6797), .ZN(n6902) );
  INV_X1 U8595 ( .A(n7953), .ZN(n7456) );
  NAND2_X1 U8596 ( .A1(n7456), .A2(n7335), .ZN(n6878) );
  AOI21_X1 U8597 ( .B1(n6511), .B2(n10429), .A(n8628), .ZN(n6799) );
  NAND3_X1 U8598 ( .A1(n6800), .A2(n6878), .A3(n6799), .ZN(n6801) );
  NOR2_X1 U8599 ( .A1(n6802), .A2(n6801), .ZN(n6803) );
  OAI21_X1 U8600 ( .B1(n6907), .B2(n6803), .A(n6904), .ZN(n6807) );
  NAND2_X1 U8601 ( .A1(n6804), .A2(n6921), .ZN(n6805) );
  AOI21_X1 U8602 ( .B1(n6807), .B2(n6806), .A(n6805), .ZN(n6808) );
  NAND2_X1 U8603 ( .A1(n6923), .A2(n8413), .ZN(n6930) );
  AND2_X1 U8604 ( .A1(n8518), .A2(n10310), .ZN(n6929) );
  OAI21_X1 U8605 ( .B1(n6808), .B2(n6930), .A(n6929), .ZN(n6809) );
  NAND3_X1 U8606 ( .A1(n6809), .A2(n6924), .A3(n6937), .ZN(n6816) );
  NOR2_X1 U8607 ( .A1(n10147), .A2(n6810), .ZN(n6945) );
  INV_X1 U8608 ( .A(n6945), .ZN(n6811) );
  AND2_X1 U8609 ( .A1(n6811), .A2(n6943), .ZN(n6812) );
  NOR2_X1 U8610 ( .A1(n10143), .A2(n8512), .ZN(n6946) );
  NAND2_X1 U8611 ( .A1(n6813), .A2(n6946), .ZN(n6814) );
  AND2_X1 U8612 ( .A1(n6815), .A2(n6814), .ZN(n6941) );
  OAI211_X1 U8613 ( .C1(n6902), .C2(n6816), .A(n6941), .B(n6940), .ZN(n6820)
         );
  AND2_X1 U8614 ( .A1(n6955), .A2(n6817), .ZN(n6954) );
  INV_X1 U8615 ( .A(n6954), .ZN(n6819) );
  AND2_X1 U8616 ( .A1(n6952), .A2(n6818), .ZN(n6958) );
  OAI21_X1 U8617 ( .B1(n6820), .B2(n6819), .A(n6958), .ZN(n6821) );
  NAND3_X1 U8618 ( .A1(n6821), .A2(n6964), .A3(n6955), .ZN(n6822) );
  AND2_X1 U8619 ( .A1(n6822), .A2(n6961), .ZN(n6841) );
  OR2_X1 U8620 ( .A1(n10108), .A2(n9594), .ZN(n6823) );
  NAND2_X1 U8621 ( .A1(n6825), .A2(n6824), .ZN(n6826) );
  NAND2_X1 U8622 ( .A1(n6826), .A2(n6983), .ZN(n6836) );
  NAND2_X1 U8623 ( .A1(n6966), .A2(n6965), .ZN(n6963) );
  INV_X1 U8624 ( .A(n6963), .ZN(n6828) );
  NAND4_X1 U8625 ( .A1(n6839), .A2(n6992), .A3(n6836), .A4(n6828), .ZN(n7028)
         );
  NAND2_X1 U8626 ( .A1(n9945), .A2(n6831), .ZN(n6977) );
  INV_X1 U8627 ( .A(n6977), .ZN(n6834) );
  NAND2_X1 U8628 ( .A1(n6962), .A2(n6832), .ZN(n6970) );
  AND2_X1 U8629 ( .A1(n6970), .A2(n6966), .ZN(n6972) );
  INV_X1 U8630 ( .A(n6972), .ZN(n6833) );
  NAND3_X1 U8631 ( .A1(n6983), .A2(n6834), .A3(n6833), .ZN(n6835) );
  NAND3_X1 U8632 ( .A1(n6992), .A2(n6836), .A3(n6835), .ZN(n6837) );
  NAND3_X1 U8633 ( .A1(n9905), .A2(n6994), .A3(n6837), .ZN(n6838) );
  NAND2_X1 U8634 ( .A1(n6839), .A2(n6838), .ZN(n6840) );
  AND2_X1 U8635 ( .A1(n7001), .A2(n6840), .ZN(n7032) );
  OAI21_X1 U8636 ( .B1(n6841), .B2(n7028), .A(n7032), .ZN(n6842) );
  NAND2_X1 U8637 ( .A1(n7029), .A2(n6842), .ZN(n6860) );
  INV_X1 U8638 ( .A(n6843), .ZN(n6844) );
  NAND2_X1 U8639 ( .A1(n6844), .A2(SI_29_), .ZN(n6851) );
  NAND2_X1 U8640 ( .A1(n6846), .A2(n6845), .ZN(n6849) );
  NAND3_X1 U8641 ( .A1(n6849), .A2(n6848), .A3(n6847), .ZN(n6850) );
  NAND2_X1 U8642 ( .A1(n6851), .A2(n6850), .ZN(n6858) );
  INV_X1 U8643 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10221) );
  INV_X1 U8644 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6852) );
  MUX2_X1 U8645 ( .A(n10221), .B(n6852), .S(n7290), .Z(n6854) );
  INV_X1 U8646 ( .A(SI_30_), .ZN(n6853) );
  NAND2_X1 U8647 ( .A1(n6854), .A2(n6853), .ZN(n6861) );
  INV_X1 U8648 ( .A(n6854), .ZN(n6855) );
  NAND2_X1 U8649 ( .A1(n6855), .A2(SI_30_), .ZN(n6856) );
  NAND2_X1 U8650 ( .A1(n6861), .A2(n6856), .ZN(n6857) );
  NAND2_X1 U8651 ( .A1(n6858), .A2(n6857), .ZN(n6859) );
  INV_X1 U8652 ( .A(n9727), .ZN(n6874) );
  AND2_X1 U8653 ( .A1(n6860), .A2(n7035), .ZN(n6876) );
  INV_X1 U8654 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10214) );
  INV_X1 U8655 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6863) );
  MUX2_X1 U8656 ( .A(n10214), .B(n6863), .S(n7290), .Z(n6864) );
  XNOR2_X1 U8657 ( .A(n6864), .B(SI_31_), .ZN(n6865) );
  OR2_X1 U8658 ( .A1(n4412), .A2(n10214), .ZN(n6867) );
  INV_X1 U8659 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U8660 ( .A1(n6869), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U8661 ( .A1(n6870), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6871) );
  OAI211_X1 U8662 ( .C1(n6126), .C2(n7676), .A(n6872), .B(n6871), .ZN(n9878)
         );
  INV_X1 U8663 ( .A(n9878), .ZN(n6873) );
  NAND2_X1 U8664 ( .A1(n7013), .A2(n6873), .ZN(n7017) );
  OR2_X1 U8665 ( .A1(n7014), .A2(n6874), .ZN(n6875) );
  NAND2_X1 U8666 ( .A1(n7017), .A2(n6875), .ZN(n6900) );
  OAI21_X1 U8667 ( .B1(n6876), .B2(n6900), .A(n4494), .ZN(n6877) );
  MUX2_X1 U8668 ( .A(n7044), .B(n6515), .S(n6877), .Z(n7049) );
  NOR2_X1 U8669 ( .A1(n8178), .A2(n10406), .ZN(n6882) );
  NOR2_X1 U8670 ( .A1(n10388), .A2(n8093), .ZN(n6881) );
  NAND2_X1 U8671 ( .A1(n7958), .A2(n6878), .ZN(n7480) );
  NOR2_X1 U8672 ( .A1(n7480), .A2(n7959), .ZN(n6880) );
  NOR2_X1 U8673 ( .A1(n8103), .A2(n4966), .ZN(n6879) );
  NAND4_X1 U8674 ( .A1(n6882), .A2(n6881), .A3(n6880), .A4(n6879), .ZN(n6883)
         );
  NOR3_X1 U8675 ( .A1(n6885), .A2(n6884), .A3(n6883), .ZN(n6886) );
  NAND4_X1 U8676 ( .A1(n10318), .A2(n6887), .A3(n8411), .A4(n6886), .ZN(n6888)
         );
  NOR2_X1 U8677 ( .A1(n8522), .A2(n6888), .ZN(n6889) );
  NAND4_X1 U8678 ( .A1(n10063), .A2(n6889), .A3(n8509), .A4(n8598), .ZN(n6890)
         );
  NOR2_X1 U8679 ( .A1(n10018), .A2(n6890), .ZN(n6891) );
  NAND4_X1 U8680 ( .A1(n10004), .A2(n6954), .A3(n6958), .A4(n6891), .ZN(n6892)
         );
  NOR2_X1 U8681 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  NAND4_X1 U8682 ( .A1(n5249), .A2(n6894), .A3(n6973), .A4(n9992), .ZN(n6895)
         );
  OR4_X1 U8683 ( .A1(n9904), .A2(n6895), .A3(n9925), .A4(n9935), .ZN(n6896) );
  NOR2_X1 U8684 ( .A1(n6897), .A2(n6896), .ZN(n6899) );
  NAND4_X1 U8685 ( .A1(n4494), .A2(n7035), .A3(n6899), .A4(n6898), .ZN(n6901)
         );
  NOR2_X1 U8686 ( .A1(n6901), .A2(n6900), .ZN(n7020) );
  NAND3_X1 U8687 ( .A1(n5282), .A2(n8270), .A3(n7020), .ZN(n7052) );
  INV_X1 U8688 ( .A(n6902), .ZN(n6938) );
  INV_X1 U8689 ( .A(n6909), .ZN(n6910) );
  NAND2_X1 U8690 ( .A1(n6910), .A2(n8288), .ZN(n6911) );
  NAND2_X1 U8691 ( .A1(n10344), .A2(n6912), .ZN(n6913) );
  NAND2_X1 U8692 ( .A1(n6913), .A2(n7010), .ZN(n6914) );
  NAND2_X1 U8693 ( .A1(n6927), .A2(n10343), .ZN(n6916) );
  MUX2_X1 U8694 ( .A(n6916), .B(n6915), .S(n7022), .Z(n6917) );
  INV_X1 U8695 ( .A(n6917), .ZN(n6918) );
  NAND2_X1 U8696 ( .A1(n6920), .A2(n8413), .ZN(n6922) );
  NAND3_X1 U8697 ( .A1(n6922), .A2(n6921), .A3(n10310), .ZN(n6925) );
  NAND4_X1 U8698 ( .A1(n6925), .A2(n6924), .A3(n6923), .A4(n7010), .ZN(n6936)
         );
  AOI21_X1 U8699 ( .B1(n6928), .B2(n6927), .A(n6926), .ZN(n6931) );
  OAI211_X1 U8700 ( .C1(n6931), .C2(n6930), .A(n6929), .B(n7022), .ZN(n6935)
         );
  AND2_X1 U8701 ( .A1(n9742), .A2(n7010), .ZN(n6933) );
  OAI21_X1 U8702 ( .B1(n7010), .B2(n9742), .A(n10317), .ZN(n6932) );
  OAI21_X1 U8703 ( .B1(n6933), .B2(n10317), .A(n6932), .ZN(n6934) );
  NAND3_X1 U8704 ( .A1(n6938), .A2(n6944), .A3(n6937), .ZN(n6939) );
  NAND3_X1 U8705 ( .A1(n6941), .A2(n6940), .A3(n6939), .ZN(n6947) );
  INV_X1 U8706 ( .A(n6948), .ZN(n6950) );
  NOR3_X1 U8707 ( .A1(n6950), .A2(n6949), .A3(n7010), .ZN(n6951) );
  NAND3_X1 U8708 ( .A1(n6961), .A2(n7010), .A3(n6952), .ZN(n6953) );
  AOI211_X1 U8709 ( .C1(n6954), .C2(n6957), .A(n6953), .B(n6970), .ZN(n6960)
         );
  NAND3_X1 U8710 ( .A1(n6964), .A2(n7022), .A3(n6955), .ZN(n6956) );
  AOI211_X1 U8711 ( .C1(n6958), .C2(n6957), .A(n6956), .B(n6963), .ZN(n6959)
         );
  NAND2_X1 U8712 ( .A1(n6961), .A2(n7022), .ZN(n6969) );
  NAND3_X1 U8713 ( .A1(n6963), .A2(n6962), .A3(n7022), .ZN(n6968) );
  NAND4_X1 U8714 ( .A1(n6966), .A2(n7010), .A3(n6965), .A4(n6964), .ZN(n6967)
         );
  OAI211_X1 U8715 ( .C1(n6970), .C2(n6969), .A(n6968), .B(n6967), .ZN(n6971)
         );
  AOI21_X1 U8716 ( .B1(n7010), .B2(n6972), .A(n6971), .ZN(n6974) );
  INV_X1 U8717 ( .A(n6978), .ZN(n6979) );
  AOI21_X1 U8718 ( .B1(n6982), .B2(n5289), .A(n6981), .ZN(n6986) );
  INV_X1 U8719 ( .A(n6983), .ZN(n6984) );
  MUX2_X1 U8720 ( .A(n9936), .B(n6984), .S(n7022), .Z(n6985) );
  NOR2_X1 U8721 ( .A1(n6986), .A2(n6985), .ZN(n6993) );
  INV_X1 U8722 ( .A(n6987), .ZN(n6988) );
  AOI21_X1 U8723 ( .B1(n7010), .B2(n6988), .A(n7002), .ZN(n6990) );
  NAND2_X1 U8724 ( .A1(n5127), .A2(n7022), .ZN(n6989) );
  NAND2_X1 U8725 ( .A1(n6997), .A2(n7001), .ZN(n6998) );
  AOI21_X1 U8726 ( .B1(n7002), .B2(n7001), .A(n7000), .ZN(n7003) );
  MUX2_X1 U8727 ( .A(n7006), .B(n7005), .S(n7022), .Z(n7007) );
  AND2_X1 U8728 ( .A1(n9727), .A2(n9878), .ZN(n7034) );
  NAND2_X1 U8729 ( .A1(n7013), .A2(n9727), .ZN(n7016) );
  INV_X1 U8730 ( .A(n7020), .ZN(n7021) );
  NOR4_X1 U8731 ( .A1(n8456), .A2(n7024), .A3(n8628), .A4(n7023), .ZN(n7025)
         );
  OR2_X1 U8732 ( .A1(n7028), .A2(n10005), .ZN(n7031) );
  INV_X1 U8733 ( .A(n7029), .ZN(n7030) );
  AOI21_X1 U8734 ( .B1(n7032), .B2(n7031), .A(n7030), .ZN(n7033) );
  INV_X1 U8735 ( .A(n7033), .ZN(n7036) );
  INV_X1 U8736 ( .A(n7037), .ZN(n7038) );
  OAI211_X1 U8737 ( .C1(n10079), .C2(n9878), .A(n7038), .B(n4494), .ZN(n7041)
         );
  NAND2_X1 U8738 ( .A1(n7322), .A2(n8270), .ZN(n7039) );
  AOI21_X1 U8739 ( .B1(n7043), .B2(n7042), .A(n8456), .ZN(n7050) );
  NOR4_X1 U8740 ( .A1(n7326), .A2(n9701), .A3(n7044), .A4(n6123), .ZN(n7045)
         );
  AOI211_X1 U8741 ( .C1(n7047), .C2(n8438), .A(n7046), .B(n7045), .ZN(n7048)
         );
  AOI21_X1 U8742 ( .B1(n7050), .B2(n7049), .A(n7048), .ZN(n7051) );
  NAND2_X1 U8743 ( .A1(n7529), .A2(n7982), .ZN(n7053) );
  OR2_X1 U8744 ( .A1(n4730), .A2(n4404), .ZN(n7055) );
  NAND2_X1 U8745 ( .A1(n7899), .A2(n7055), .ZN(n10536) );
  NAND2_X1 U8746 ( .A1(n7057), .A2(n4774), .ZN(n8874) );
  NAND2_X1 U8747 ( .A1(n7901), .A2(n4774), .ZN(n7058) );
  NAND2_X1 U8748 ( .A1(n9035), .A2(n7060), .ZN(n7059) );
  NAND2_X1 U8749 ( .A1(n7109), .A2(n10555), .ZN(n7061) );
  OR2_X1 U8750 ( .A1(n9034), .A2(n8147), .ZN(n8136) );
  OAI21_X1 U8751 ( .B1(n4764), .B2(n7110), .A(n8136), .ZN(n7066) );
  NAND2_X1 U8752 ( .A1(n7110), .A2(n8138), .ZN(n7062) );
  NAND2_X1 U8753 ( .A1(n7947), .A2(n7062), .ZN(n7064) );
  AND2_X1 U8754 ( .A1(n9034), .A2(n8138), .ZN(n7063) );
  AOI22_X1 U8755 ( .A1(n7064), .A2(n8147), .B1(n7063), .B2(n7110), .ZN(n7065)
         );
  NAND2_X1 U8756 ( .A1(n7990), .A2(n8059), .ZN(n7067) );
  NAND2_X1 U8757 ( .A1(n8065), .A2(n7067), .ZN(n7069) );
  INV_X1 U8758 ( .A(n8059), .ZN(n9442) );
  NAND2_X1 U8759 ( .A1(n7111), .A2(n9442), .ZN(n7068) );
  NAND2_X1 U8760 ( .A1(n7069), .A2(n7068), .ZN(n8167) );
  OR2_X2 U8761 ( .A1(n9032), .A2(n7070), .ZN(n8854) );
  NAND2_X1 U8762 ( .A1(n7070), .A2(n9032), .ZN(n8851) );
  NAND2_X1 U8763 ( .A1(n8854), .A2(n8851), .ZN(n8165) );
  OR2_X1 U8764 ( .A1(n9033), .A2(n8200), .ZN(n8168) );
  NAND2_X1 U8765 ( .A1(n8167), .A2(n8170), .ZN(n7074) );
  OR2_X1 U8766 ( .A1(n9033), .A2(n8247), .ZN(n8853) );
  NAND2_X1 U8767 ( .A1(n9033), .A2(n8247), .ZN(n8164) );
  NAND2_X1 U8768 ( .A1(n8853), .A2(n8164), .ZN(n8194) );
  NAND3_X1 U8769 ( .A1(n8901), .A2(n8165), .A3(n8168), .ZN(n7072) );
  INV_X1 U8770 ( .A(n7070), .ZN(n8266) );
  AND2_X1 U8771 ( .A1(n8266), .A2(n9032), .ZN(n8278) );
  AOI21_X1 U8772 ( .B1(n9031), .B2(n8611), .A(n8278), .ZN(n7071) );
  AND2_X1 U8773 ( .A1(n7072), .A2(n7071), .ZN(n7073) );
  NAND2_X1 U8774 ( .A1(n7074), .A2(n7073), .ZN(n7076) );
  OR2_X1 U8775 ( .A1(n8611), .A2(n9031), .ZN(n7075) );
  NOR2_X1 U8776 ( .A1(n8485), .A2(n9030), .ZN(n7078) );
  NAND2_X1 U8777 ( .A1(n8485), .A2(n9030), .ZN(n7077) );
  NAND2_X1 U8778 ( .A1(n8921), .A2(n9028), .ZN(n7081) );
  NAND2_X1 U8779 ( .A1(n8926), .A2(n8925), .ZN(n8927) );
  NOR2_X1 U8780 ( .A1(n8934), .A2(n9383), .ZN(n7082) );
  NAND2_X1 U8781 ( .A1(n9521), .A2(n8708), .ZN(n8940) );
  NAND2_X1 U8782 ( .A1(n8942), .A2(n8940), .ZN(n8932) );
  NAND2_X1 U8783 ( .A1(n9521), .A2(n9370), .ZN(n7083) );
  NAND2_X1 U8784 ( .A1(n9514), .A2(n9359), .ZN(n8945) );
  NAND2_X1 U8785 ( .A1(n8948), .A2(n8945), .ZN(n8811) );
  NAND2_X1 U8786 ( .A1(n9514), .A2(n9381), .ZN(n7084) );
  NAND2_X1 U8787 ( .A1(n9363), .A2(n9371), .ZN(n8946) );
  NAND2_X1 U8788 ( .A1(n9431), .A2(n8769), .ZN(n8949) );
  NAND2_X1 U8789 ( .A1(n9431), .A2(n9371), .ZN(n7085) );
  AND2_X1 U8790 ( .A1(n9507), .A2(n9027), .ZN(n7086) );
  OR2_X1 U8791 ( .A1(n9507), .A2(n9027), .ZN(n7087) );
  NAND2_X1 U8792 ( .A1(n9329), .A2(n9345), .ZN(n9314) );
  NAND2_X1 U8793 ( .A1(n8810), .A2(n9314), .ZN(n7091) );
  NAND2_X1 U8794 ( .A1(n9329), .A2(n9318), .ZN(n9311) );
  NAND2_X1 U8795 ( .A1(n9491), .A2(n9317), .ZN(n8963) );
  NAND2_X1 U8796 ( .A1(n8964), .A2(n8963), .ZN(n9302) );
  INV_X1 U8797 ( .A(n9491), .ZN(n8685) );
  OAI21_X1 U8798 ( .B1(n8974), .B2(n9273), .A(n9266), .ZN(n7094) );
  NAND2_X1 U8799 ( .A1(n9469), .A2(n9026), .ZN(n8970) );
  NAND2_X1 U8800 ( .A1(n8975), .A2(n8970), .ZN(n9255) );
  INV_X1 U8801 ( .A(n9469), .ZN(n9260) );
  NAND2_X1 U8802 ( .A1(n7095), .A2(n8701), .ZN(n7097) );
  NAND2_X1 U8803 ( .A1(n9398), .A2(n9249), .ZN(n7128) );
  NAND2_X1 U8804 ( .A1(n7099), .A2(n7098), .ZN(n7103) );
  NAND2_X1 U8805 ( .A1(n9536), .A2(n5624), .ZN(n7101) );
  NAND2_X1 U8806 ( .A1(n5906), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7100) );
  NAND2_X1 U8807 ( .A1(n8646), .A2(n9025), .ZN(n8806) );
  XNOR2_X1 U8808 ( .A(n7103), .B(n7102), .ZN(n7106) );
  NAND2_X1 U8809 ( .A1(n10530), .A2(n4635), .ZN(n10529) );
  OR2_X1 U8810 ( .A1(n7110), .A2(n10560), .ZN(n8886) );
  INV_X1 U8811 ( .A(n9035), .ZN(n7109) );
  NAND2_X1 U8812 ( .A1(n7110), .A2(n10560), .ZN(n8132) );
  INV_X1 U8813 ( .A(n8147), .ZN(n10566) );
  NAND2_X1 U8814 ( .A1(n9034), .A2(n10566), .ZN(n8896) );
  AND2_X1 U8815 ( .A1(n8132), .A2(n8896), .ZN(n8891) );
  AND2_X1 U8816 ( .A1(n9035), .A2(n10555), .ZN(n8889) );
  OR2_X1 U8817 ( .A1(n9034), .A2(n10566), .ZN(n8885) );
  INV_X1 U8818 ( .A(n7990), .ZN(n7111) );
  NAND2_X1 U8819 ( .A1(n7111), .A2(n8059), .ZN(n8897) );
  AND2_X1 U8820 ( .A1(n8851), .A2(n8164), .ZN(n8859) );
  NAND2_X1 U8821 ( .A1(n8485), .A2(n8535), .ZN(n8912) );
  INV_X1 U8822 ( .A(n9029), .ZN(n8689) );
  AND2_X1 U8823 ( .A1(n8530), .A2(n8689), .ZN(n8911) );
  INV_X1 U8824 ( .A(n8911), .ZN(n7115) );
  OR2_X1 U8825 ( .A1(n8530), .A2(n8689), .ZN(n8916) );
  XNOR2_X1 U8826 ( .A(n8921), .B(n9028), .ZN(n8919) );
  NAND2_X1 U8827 ( .A1(n8390), .A2(n8919), .ZN(n8389) );
  INV_X1 U8828 ( .A(n9028), .ZN(n8920) );
  OR2_X1 U8829 ( .A1(n8921), .A2(n8920), .ZN(n8923) );
  NAND2_X1 U8830 ( .A1(n8389), .A2(n8923), .ZN(n8428) );
  NAND2_X1 U8831 ( .A1(n8751), .A2(n8925), .ZN(n7116) );
  NAND2_X1 U8832 ( .A1(n8926), .A2(n8691), .ZN(n7117) );
  XNOR2_X1 U8833 ( .A(n8934), .B(n9383), .ZN(n8827) );
  OR2_X1 U8834 ( .A1(n8934), .A2(n8933), .ZN(n8936) );
  NAND2_X1 U8835 ( .A1(n9377), .A2(n8940), .ZN(n7118) );
  NAND2_X1 U8836 ( .A1(n7118), .A2(n8942), .ZN(n9367) );
  NAND2_X1 U8837 ( .A1(n9367), .A2(n8945), .ZN(n7119) );
  INV_X1 U8838 ( .A(n8849), .ZN(n7120) );
  NAND2_X1 U8839 ( .A1(n9507), .A2(n9358), .ZN(n8950) );
  OAI211_X1 U8840 ( .C1(n7120), .C2(n8950), .A(n8960), .B(n9311), .ZN(n7121)
         );
  INV_X1 U8841 ( .A(n7121), .ZN(n7122) );
  NAND2_X1 U8842 ( .A1(n7123), .A2(n8963), .ZN(n9289) );
  OR2_X1 U8843 ( .A1(n9291), .A2(n8754), .ZN(n7124) );
  NAND2_X1 U8844 ( .A1(n9289), .A2(n7124), .ZN(n7126) );
  NAND2_X1 U8845 ( .A1(n9291), .A2(n8754), .ZN(n7125) );
  NAND2_X1 U8846 ( .A1(n9481), .A2(n9288), .ZN(n8843) );
  NAND2_X1 U8847 ( .A1(n6792), .A2(n9249), .ZN(n7131) );
  NAND2_X1 U8848 ( .A1(n9456), .A2(n8836), .ZN(n7132) );
  AOI21_X1 U8849 ( .B1(n8992), .B2(n8869), .A(n5743), .ZN(n7133) );
  AND2_X1 U8850 ( .A1(n10565), .A2(n7133), .ZN(n7134) );
  INV_X1 U8851 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n7139) );
  NAND2_X1 U8852 ( .A1(n4408), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U8853 ( .A1(n7135), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7136) );
  OAI211_X1 U8854 ( .C1(n7139), .C2(n7138), .A(n7137), .B(n7136), .ZN(n7140)
         );
  INV_X1 U8855 ( .A(n7140), .ZN(n7141) );
  NAND2_X1 U8856 ( .A1(n4746), .A2(P2_B_REG_SCAN_IN), .ZN(n7143) );
  NAND2_X1 U8857 ( .A1(n9380), .A2(n7143), .ZN(n9218) );
  OAI22_X1 U8858 ( .A1(n8836), .A2(n10537), .B1(n8839), .B2(n9218), .ZN(n7144)
         );
  OR2_X1 U8859 ( .A1(n7161), .A2(n9020), .ZN(n8191) );
  OR2_X1 U8860 ( .A1(n7146), .A2(n8191), .ZN(n7147) );
  NAND2_X1 U8861 ( .A1(n7974), .A2(n7148), .ZN(n7149) );
  NAND2_X1 U8862 ( .A1(n7150), .A2(n7149), .ZN(n7154) );
  NAND2_X1 U8863 ( .A1(n7152), .A2(n7151), .ZN(n7153) );
  NAND2_X1 U8864 ( .A1(n7155), .A2(n4523), .ZN(n7156) );
  INV_X1 U8865 ( .A(n8646), .ZN(n7170) );
  NAND2_X1 U8866 ( .A1(n7156), .A2(n5275), .ZN(P2_U3456) );
  AND3_X1 U8867 ( .A1(n7158), .A2(n7314), .A3(n7157), .ZN(n7160) );
  OAI21_X1 U8868 ( .B1(n10565), .B2(n7161), .A(n7972), .ZN(n7163) );
  NAND3_X1 U8869 ( .A1(n8992), .A2(n9020), .A3(n9198), .ZN(n7162) );
  NAND2_X1 U8870 ( .A1(n7163), .A2(n7973), .ZN(n7166) );
  INV_X1 U8871 ( .A(n7973), .ZN(n7164) );
  NAND2_X1 U8872 ( .A1(n7164), .A2(n7969), .ZN(n7165) );
  INV_X1 U8873 ( .A(n10578), .ZN(n7168) );
  INV_X1 U8874 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7167) );
  NAND2_X1 U8875 ( .A1(n7168), .A2(n7167), .ZN(n7169) );
  INV_X1 U8876 ( .A(n7174), .ZN(n8452) );
  NOR2_X1 U8877 ( .A1(n7171), .A2(P1_U3086), .ZN(n7172) );
  NAND2_X1 U8878 ( .A1(n8999), .A2(n7173), .ZN(n7175) );
  NAND2_X1 U8879 ( .A1(n7175), .A2(n7174), .ZN(n7280) );
  NAND2_X1 U8880 ( .A1(n7280), .A2(n4746), .ZN(n7177) );
  NAND2_X1 U8881 ( .A1(n7177), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8882 ( .A(n7259), .ZN(n8111) );
  INV_X1 U8883 ( .A(n7935), .ZN(n7310) );
  INV_X1 U8884 ( .A(n7472), .ZN(n7303) );
  NOR2_X1 U8885 ( .A1(n7224), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7178) );
  OAI21_X1 U8886 ( .B1(n7347), .B2(n7178), .A(n7180), .ZN(n7349) );
  INV_X1 U8887 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U8888 ( .A1(n7350), .A2(n7180), .ZN(n7513) );
  NAND2_X1 U8889 ( .A1(n7514), .A2(n7513), .ZN(n7512) );
  INV_X1 U8890 ( .A(n7520), .ZN(n7292) );
  NAND2_X1 U8891 ( .A1(n7292), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7181) );
  NAND2_X1 U8892 ( .A1(n7420), .A2(n7437), .ZN(n7183) );
  INV_X1 U8893 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n8030) );
  XNOR2_X1 U8894 ( .A(n7431), .B(n8030), .ZN(n7436) );
  NAND2_X1 U8895 ( .A1(n7431), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7184) );
  XNOR2_X1 U8896 ( .A(n7472), .B(n8067), .ZN(n7469) );
  INV_X1 U8897 ( .A(n7187), .ZN(n7925) );
  INV_X1 U8898 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8212) );
  XNOR2_X1 U8899 ( .A(n7935), .B(n8212), .ZN(n7926) );
  XNOR2_X1 U8900 ( .A(n7259), .B(n8375), .ZN(n8113) );
  INV_X1 U8901 ( .A(n7189), .ZN(n7191) );
  INV_X1 U8902 ( .A(n7264), .ZN(n8230) );
  INV_X1 U8903 ( .A(n7194), .ZN(n7190) );
  XNOR2_X1 U8904 ( .A(n9038), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7193) );
  OR3_X1 U8905 ( .A1(n7194), .A2(n7192), .A3(n7193), .ZN(n7195) );
  NOR2_X1 U8906 ( .A1(n7278), .A2(P2_U3151), .ZN(n9541) );
  NAND2_X1 U8907 ( .A1(n7280), .A2(n9541), .ZN(n7505) );
  AOI21_X1 U8908 ( .B1(n9039), .B2(n7195), .A(n9217), .ZN(n7289) );
  NAND2_X1 U8909 ( .A1(n7347), .A2(n7199), .ZN(n7198) );
  NAND2_X1 U8910 ( .A1(n7198), .A2(n7197), .ZN(n7352) );
  NAND2_X1 U8911 ( .A1(n7352), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7200) );
  NAND2_X1 U8912 ( .A1(n7200), .A2(n7199), .ZN(n7516) );
  NAND2_X1 U8913 ( .A1(n7517), .A2(n7516), .ZN(n7515) );
  NAND2_X1 U8914 ( .A1(n7292), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7201) );
  NAND2_X1 U8915 ( .A1(n7421), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7204) );
  NAND2_X1 U8916 ( .A1(n7202), .A2(n7418), .ZN(n7203) );
  NAND2_X1 U8917 ( .A1(n7361), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7208) );
  NAND2_X1 U8918 ( .A1(n7206), .A2(n7296), .ZN(n7207) );
  MUX2_X1 U8919 ( .A(n7242), .B(P2_REG1_REG_6__SCAN_IN), .S(n7472), .Z(n7467)
         );
  OR2_X1 U8920 ( .A1(n7472), .A2(n7242), .ZN(n7209) );
  NAND2_X1 U8921 ( .A1(n7860), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7212) );
  NAND2_X1 U8922 ( .A1(n7210), .A2(n5177), .ZN(n7211) );
  NAND2_X1 U8923 ( .A1(n7310), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7213) );
  NAND2_X1 U8924 ( .A1(n8007), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7216) );
  INV_X1 U8925 ( .A(n8016), .ZN(n7330) );
  NAND2_X1 U8926 ( .A1(n7214), .A2(n7330), .ZN(n7215) );
  NAND2_X1 U8927 ( .A1(n7216), .A2(n7215), .ZN(n8109) );
  XNOR2_X1 U8928 ( .A(n7259), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n8110) );
  NOR2_X1 U8929 ( .A1(n7259), .A2(n8397), .ZN(n7217) );
  AOI21_X1 U8930 ( .B1(n8109), .B2(n8110), .A(n7217), .ZN(n7218) );
  INV_X1 U8931 ( .A(n9038), .ZN(n9057) );
  AOI22_X1 U8932 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n9057), .B1(n9038), .B2(
        n8443), .ZN(n7219) );
  OAI21_X1 U8933 ( .B1(n7220), .B2(n7219), .A(n9058), .ZN(n7221) );
  AND2_X1 U8934 ( .A1(n7221), .A2(n9173), .ZN(n7288) );
  MUX2_X1 U8935 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n5378), .Z(n7226) );
  INV_X1 U8936 ( .A(n7347), .ZN(n7222) );
  MUX2_X1 U8937 ( .A(n7224), .B(n7223), .S(n9181), .Z(n7225) );
  NAND2_X1 U8938 ( .A1(n7346), .A2(n7504), .ZN(n7228) );
  NAND2_X1 U8939 ( .A1(n7226), .A2(n7347), .ZN(n7227) );
  NAND2_X1 U8940 ( .A1(n7228), .A2(n7227), .ZN(n7510) );
  MUX2_X1 U8941 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n9181), .Z(n7229) );
  XNOR2_X1 U8942 ( .A(n7520), .B(n7229), .ZN(n7511) );
  NAND2_X1 U8943 ( .A1(n7510), .A2(n7511), .ZN(n7231) );
  NAND2_X1 U8944 ( .A1(n7229), .A2(n7292), .ZN(n7230) );
  NAND2_X1 U8945 ( .A1(n7231), .A2(n7230), .ZN(n7416) );
  MUX2_X1 U8946 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n4401), .Z(n7233) );
  XNOR2_X1 U8947 ( .A(n7233), .B(n7418), .ZN(n7417) );
  MUX2_X1 U8948 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4402), .Z(n7237) );
  XNOR2_X1 U8949 ( .A(n7237), .B(n7232), .ZN(n7427) );
  INV_X1 U8950 ( .A(n7233), .ZN(n7235) );
  NAND2_X1 U8951 ( .A1(n7235), .A2(n7234), .ZN(n7428) );
  AND2_X1 U8952 ( .A1(n7427), .A2(n7428), .ZN(n7236) );
  NAND2_X1 U8953 ( .A1(n7429), .A2(n7236), .ZN(n7430) );
  NAND2_X1 U8954 ( .A1(n7237), .A2(n7431), .ZN(n7238) );
  NAND2_X1 U8955 ( .A1(n7430), .A2(n7238), .ZN(n7360) );
  MUX2_X1 U8956 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n4402), .Z(n7239) );
  XNOR2_X1 U8957 ( .A(n7239), .B(n4800), .ZN(n7359) );
  NAND2_X1 U8958 ( .A1(n7360), .A2(n7359), .ZN(n7241) );
  NAND2_X1 U8959 ( .A1(n7239), .A2(n7296), .ZN(n7240) );
  NAND2_X1 U8960 ( .A1(n7241), .A2(n7240), .ZN(n7464) );
  MUX2_X1 U8961 ( .A(n8067), .B(n7242), .S(n4402), .Z(n7243) );
  NAND2_X1 U8962 ( .A1(n7243), .A2(n7472), .ZN(n7867) );
  INV_X1 U8963 ( .A(n7243), .ZN(n7244) );
  NAND2_X1 U8964 ( .A1(n7244), .A2(n7303), .ZN(n7245) );
  NAND2_X1 U8965 ( .A1(n7867), .A2(n7245), .ZN(n7463) );
  NAND2_X1 U8966 ( .A1(n7868), .A2(n7867), .ZN(n7249) );
  INV_X1 U8967 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8227) );
  MUX2_X1 U8968 ( .A(n8227), .B(n8245), .S(n4402), .Z(n7246) );
  NAND2_X1 U8969 ( .A1(n7246), .A2(n7862), .ZN(n7932) );
  INV_X1 U8970 ( .A(n7246), .ZN(n7247) );
  NAND2_X1 U8971 ( .A1(n7247), .A2(n5177), .ZN(n7248) );
  AND2_X1 U8972 ( .A1(n7932), .A2(n7248), .ZN(n7865) );
  NAND2_X1 U8973 ( .A1(n7933), .A2(n7932), .ZN(n7253) );
  MUX2_X1 U8974 ( .A(n8212), .B(n8217), .S(n4402), .Z(n7250) );
  NAND2_X1 U8975 ( .A1(n7250), .A2(n7935), .ZN(n8012) );
  INV_X1 U8976 ( .A(n7250), .ZN(n7251) );
  NAND2_X1 U8977 ( .A1(n7251), .A2(n7310), .ZN(n7252) );
  AND2_X1 U8978 ( .A1(n8012), .A2(n7252), .ZN(n7930) );
  NAND2_X1 U8979 ( .A1(n8013), .A2(n8012), .ZN(n7258) );
  MUX2_X1 U8980 ( .A(n7254), .B(n8348), .S(n4402), .Z(n7255) );
  NAND2_X1 U8981 ( .A1(n7255), .A2(n8016), .ZN(n8118) );
  INV_X1 U8982 ( .A(n7255), .ZN(n7256) );
  NAND2_X1 U8983 ( .A1(n7256), .A2(n7330), .ZN(n7257) );
  AND2_X1 U8984 ( .A1(n8118), .A2(n7257), .ZN(n8010) );
  NAND2_X1 U8985 ( .A1(n8117), .A2(n8118), .ZN(n7263) );
  MUX2_X1 U8986 ( .A(n8375), .B(n8397), .S(n4401), .Z(n7260) );
  NAND2_X1 U8987 ( .A1(n7260), .A2(n7259), .ZN(n8233) );
  INV_X1 U8988 ( .A(n7260), .ZN(n7261) );
  NAND2_X1 U8989 ( .A1(n7261), .A2(n8111), .ZN(n7262) );
  AND2_X1 U8990 ( .A1(n8233), .A2(n7262), .ZN(n8119) );
  NAND2_X1 U8991 ( .A1(n8234), .A2(n8233), .ZN(n7268) );
  MUX2_X1 U8992 ( .A(n8384), .B(n8380), .S(n4402), .Z(n7265) );
  NAND2_X1 U8993 ( .A1(n7265), .A2(n7264), .ZN(n7275) );
  INV_X1 U8994 ( .A(n7265), .ZN(n7266) );
  NAND2_X1 U8995 ( .A1(n7266), .A2(n8230), .ZN(n7267) );
  AND2_X1 U8996 ( .A1(n7275), .A2(n7267), .ZN(n8231) );
  NAND2_X1 U8997 ( .A1(n8236), .A2(n7275), .ZN(n7272) );
  MUX2_X1 U8998 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n4402), .Z(n7269) );
  NAND2_X1 U8999 ( .A1(n9057), .A2(n7269), .ZN(n7271) );
  INV_X1 U9000 ( .A(n7269), .ZN(n7270) );
  NAND2_X1 U9001 ( .A1(n7270), .A2(n9038), .ZN(n9052) );
  AND2_X1 U9002 ( .A1(n7271), .A2(n9052), .ZN(n7273) );
  INV_X1 U9003 ( .A(n7273), .ZN(n7274) );
  NAND3_X1 U9004 ( .A1(n8236), .A2(n7275), .A3(n7274), .ZN(n7276) );
  AOI21_X1 U9005 ( .B1(n9053), .B2(n7276), .A(n9159), .ZN(n7287) );
  INV_X1 U9006 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7285) );
  NAND2_X1 U9007 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8688) );
  NOR2_X1 U9008 ( .A1(n4401), .A2(P2_U3151), .ZN(n9544) );
  AND2_X1 U9009 ( .A1(n9544), .A2(n7278), .ZN(n7279) );
  NAND2_X1 U9010 ( .A1(n7280), .A2(n7279), .ZN(n7283) );
  NAND2_X1 U9011 ( .A1(n7281), .A2(n9541), .ZN(n7282) );
  NAND2_X1 U9012 ( .A1(n7283), .A2(n7282), .ZN(n9209) );
  NAND2_X1 U9013 ( .A1(n9209), .A2(n9038), .ZN(n7284) );
  OAI211_X1 U9014 ( .C1(n9171), .C2(n7285), .A(n8688), .B(n7284), .ZN(n7286)
         );
  XNOR2_X1 U9015 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U9016 ( .A1(n7290), .A2(P2_U3151), .ZN(n8451) );
  INV_X2 U9017 ( .A(n8451), .ZN(n9547) );
  NOR2_X1 U9018 ( .A1(n7290), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9545) );
  INV_X2 U9019 ( .A(n9545), .ZN(n9537) );
  OAI222_X1 U9020 ( .A1(n9547), .A2(n7291), .B1(n9537), .B2(n5332), .C1(
        P2_U3151), .C2(n7347), .ZN(P2_U3294) );
  NOR2_X1 U9021 ( .A1(n7290), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10217) );
  INV_X2 U9022 ( .A(n10217), .ZN(n8271) );
  OAI222_X1 U9023 ( .A1(n10224), .A2(n4640), .B1(n8271), .B2(n7291), .C1(n7392), .C2(P1_U3086), .ZN(P1_U3354) );
  OAI222_X1 U9024 ( .A1(n9547), .A2(n7295), .B1(n7418), .B2(P2_U3151), .C1(
        n5410), .C2(n9537), .ZN(P2_U3292) );
  OAI222_X1 U9025 ( .A1(n10224), .A2(n5039), .B1(n8271), .B2(n7293), .C1(
        P1_U3086), .C2(n7839), .ZN(P1_U3353) );
  OAI222_X1 U9026 ( .A1(n9537), .A2(n7294), .B1(n9547), .B2(n7293), .C1(
        P2_U3151), .C2(n7292), .ZN(P2_U3293) );
  OAI222_X1 U9027 ( .A1(P1_U3086), .A2(n7396), .B1(n8271), .B2(n7295), .C1(
        n5409), .C2(n10224), .ZN(P1_U3352) );
  OAI222_X1 U9028 ( .A1(n9547), .A2(n7297), .B1(n7296), .B2(P2_U3151), .C1(
        n4580), .C2(n9537), .ZN(P2_U3290) );
  OAI222_X1 U9029 ( .A1(P1_U3086), .A2(n7400), .B1(n8271), .B2(n7297), .C1(
        n5468), .C2(n10224), .ZN(P1_U3350) );
  OAI222_X1 U9030 ( .A1(n9547), .A2(n7298), .B1(n7431), .B2(P2_U3151), .C1(
        n5001), .C2(n9537), .ZN(P2_U3291) );
  OAI222_X1 U9031 ( .A1(P1_U3086), .A2(n7856), .B1(n8271), .B2(n7298), .C1(
        n5002), .C2(n10224), .ZN(P1_U3351) );
  INV_X1 U9032 ( .A(n7969), .ZN(n7299) );
  NAND2_X1 U9033 ( .A1(n7299), .A2(n7314), .ZN(n7300) );
  OAI21_X1 U9034 ( .B1(n7314), .B2(n5952), .A(n7300), .ZN(P2_U3377) );
  INV_X1 U9035 ( .A(n7301), .ZN(n7307) );
  OAI222_X1 U9036 ( .A1(n9547), .A2(n7307), .B1(n5177), .B2(P2_U3151), .C1(
        n4881), .C2(n9537), .ZN(P2_U3288) );
  INV_X1 U9037 ( .A(n7302), .ZN(n7305) );
  OAI222_X1 U9038 ( .A1(n9537), .A2(n7304), .B1(n9547), .B2(n7305), .C1(
        P2_U3151), .C2(n7303), .ZN(P2_U3289) );
  OAI222_X1 U9039 ( .A1(n10224), .A2(n7306), .B1(n8271), .B2(n7305), .C1(
        P1_U3086), .C2(n9790), .ZN(P1_U3349) );
  OAI222_X1 U9040 ( .A1(n10224), .A2(n4829), .B1(n8271), .B2(n7307), .C1(n9804), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U9041 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7785) );
  INV_X1 U9042 ( .A(n7308), .ZN(n7311) );
  INV_X1 U9043 ( .A(n9821), .ZN(n7309) );
  OAI222_X1 U9044 ( .A1(n10224), .A2(n7785), .B1(n8271), .B2(n7311), .C1(
        P1_U3086), .C2(n7309), .ZN(P1_U3347) );
  INV_X1 U9045 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7625) );
  OAI222_X1 U9046 ( .A1(n9537), .A2(n7625), .B1(n9547), .B2(n7311), .C1(
        P2_U3151), .C2(n7310), .ZN(P2_U3287) );
  INV_X1 U9047 ( .A(n7312), .ZN(n7313) );
  INV_X1 U9048 ( .A(n7315), .ZN(n7316) );
  AOI22_X1 U9049 ( .A1(n7319), .A2(n7318), .B1(n7317), .B2(n7316), .ZN(
        P2_U3376) );
  AND2_X1 U9050 ( .A1(n7319), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U9051 ( .A1(n7319), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U9052 ( .A1(n7319), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U9053 ( .A1(n7319), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U9054 ( .A1(n7319), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U9055 ( .A1(n7319), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U9056 ( .A1(n7319), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U9057 ( .A1(n7319), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U9058 ( .A1(n7319), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U9059 ( .A1(n7319), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U9060 ( .A1(n7319), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U9061 ( .A1(n7319), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U9062 ( .A1(n7319), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U9063 ( .A1(n7319), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U9064 ( .A1(n7319), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U9065 ( .A1(n7319), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U9066 ( .A1(n7319), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U9067 ( .A1(n7319), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U9068 ( .A1(n7319), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U9069 ( .A1(n7319), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U9070 ( .A1(n7319), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U9071 ( .A1(n7319), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U9072 ( .A1(n7319), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U9073 ( .A1(n7319), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U9074 ( .A1(n7319), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U9075 ( .A1(n7319), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U9076 ( .A1(n7319), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U9077 ( .A1(n7319), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U9078 ( .A1(n7319), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U9079 ( .A1(n7319), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U9080 ( .A(n10224), .ZN(n8151) );
  AOI22_X1 U9081 ( .A1(n7884), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n8151), .ZN(n7320) );
  OAI21_X1 U9082 ( .B1(n7321), .B2(n8271), .A(n7320), .ZN(P1_U3345) );
  OAI222_X1 U9083 ( .A1(n9547), .A2(n7321), .B1(n8111), .B2(P2_U3151), .C1(
        n4810), .C2(n9537), .ZN(P2_U3285) );
  NAND2_X1 U9084 ( .A1(n7323), .A2(n7322), .ZN(n7325) );
  AND2_X1 U9085 ( .A1(n7325), .A2(n7324), .ZN(n7387) );
  INV_X1 U9086 ( .A(n7387), .ZN(n7327) );
  NAND2_X1 U9087 ( .A1(n8456), .A2(n7326), .ZN(n7388) );
  NOR2_X1 U9088 ( .A1(n10233), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U9089 ( .A(n7328), .ZN(n7332) );
  OAI222_X1 U9090 ( .A1(n9547), .A2(n7332), .B1(n7330), .B2(P2_U3151), .C1(
        n7329), .C2(n9537), .ZN(P2_U3286) );
  INV_X1 U9091 ( .A(n7491), .ZN(n7331) );
  OAI222_X1 U9092 ( .A1(n10224), .A2(n7787), .B1(n8271), .B2(n7332), .C1(n7331), .C2(P1_U3086), .ZN(P1_U3346) );
  NAND2_X1 U9093 ( .A1(P1_U3973), .A2(n9878), .ZN(n7333) );
  OAI21_X1 U9094 ( .B1(P1_U3973), .B2(n6863), .A(n7333), .ZN(P1_U3585) );
  NAND2_X1 U9095 ( .A1(P1_U3973), .A2(n6511), .ZN(n7334) );
  OAI21_X1 U9096 ( .B1(P1_U3973), .B2(n5332), .A(n7334), .ZN(P1_U3555) );
  INV_X1 U9097 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7727) );
  NAND2_X1 U9098 ( .A1(n7335), .A2(P1_U3973), .ZN(n7336) );
  OAI21_X1 U9099 ( .B1(P1_U3973), .B2(n7727), .A(n7336), .ZN(P1_U3554) );
  INV_X1 U9100 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7793) );
  NAND2_X1 U9101 ( .A1(n8691), .A2(P2_U3893), .ZN(n7337) );
  OAI21_X1 U9102 ( .B1(P2_U3893), .B2(n7793), .A(n7337), .ZN(P2_U3504) );
  INV_X1 U9103 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7796) );
  INV_X1 U9104 ( .A(n7338), .ZN(n7340) );
  INV_X1 U9105 ( .A(n9840), .ZN(n7339) );
  OAI222_X1 U9106 ( .A1(n10224), .A2(n7796), .B1(n8271), .B2(n7340), .C1(
        P1_U3086), .C2(n7339), .ZN(P1_U3344) );
  INV_X1 U9107 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7341) );
  OAI222_X1 U9108 ( .A1(n9537), .A2(n7341), .B1(n9547), .B2(n7340), .C1(
        P2_U3151), .C2(n8230), .ZN(P2_U3284) );
  INV_X1 U9109 ( .A(n7342), .ZN(n7345) );
  AOI22_X1 U9110 ( .A1(n8044), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n8151), .ZN(n7343) );
  OAI21_X1 U9111 ( .B1(n7345), .B2(n8271), .A(n7343), .ZN(P1_U3343) );
  INV_X1 U9112 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7344) );
  OAI222_X1 U9113 ( .A1(n9547), .A2(n7345), .B1(n9057), .B2(P2_U3151), .C1(
        n7344), .C2(n9537), .ZN(P2_U3283) );
  XNOR2_X1 U9114 ( .A(n7346), .B(n7504), .ZN(n7357) );
  OAI22_X1 U9115 ( .A1(n9154), .A2(n7347), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8082), .ZN(n7348) );
  AOI21_X1 U9116 ( .B1(n9210), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n7348), .ZN(
        n7356) );
  INV_X1 U9117 ( .A(n7349), .ZN(n7351) );
  OAI21_X1 U9118 ( .B1(n7351), .B2(P2_REG2_REG_1__SCAN_IN), .A(n7350), .ZN(
        n7354) );
  XNOR2_X1 U9119 ( .A(n7352), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n7353) );
  AOI22_X1 U9120 ( .A1(n9146), .A2(n7354), .B1(n9173), .B2(n7353), .ZN(n7355)
         );
  OAI211_X1 U9121 ( .C1(n9159), .C2(n7357), .A(n7356), .B(n7355), .ZN(P2_U3183) );
  NAND2_X1 U9122 ( .A1(n9738), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7358) );
  OAI21_X1 U9123 ( .B1(n9593), .B2(n9738), .A(n7358), .ZN(P1_U3574) );
  XNOR2_X1 U9124 ( .A(n7360), .B(n7359), .ZN(n7371) );
  XOR2_X1 U9125 ( .A(n7361), .B(n5461), .Z(n7369) );
  INV_X1 U9126 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7367) );
  OAI21_X1 U9127 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n7363), .A(n7362), .ZN(
        n7364) );
  NAND2_X1 U9128 ( .A1(n9146), .A2(n7364), .ZN(n7366) );
  AND2_X1 U9129 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7992) );
  AOI21_X1 U9130 ( .B1(n9209), .B2(n4800), .A(n7992), .ZN(n7365) );
  OAI211_X1 U9131 ( .C1(n9171), .C2(n7367), .A(n7366), .B(n7365), .ZN(n7368)
         );
  AOI21_X1 U9132 ( .B1(n9173), .B2(n7369), .A(n7368), .ZN(n7370) );
  OAI21_X1 U9133 ( .B1(n7371), .B2(n9159), .A(n7370), .ZN(P2_U3187) );
  XNOR2_X1 U9134 ( .A(n7491), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n7386) );
  INV_X1 U9135 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10513) );
  MUX2_X1 U9136 ( .A(n10513), .B(P1_REG1_REG_2__SCAN_IN), .S(n7839), .Z(n7835)
         );
  INV_X1 U9137 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10511) );
  MUX2_X1 U9138 ( .A(n10511), .B(P1_REG1_REG_1__SCAN_IN), .S(n7392), .Z(n9758)
         );
  AND2_X1 U9139 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9757) );
  NAND2_X1 U9140 ( .A1(n9758), .A2(n9757), .ZN(n9756) );
  NAND2_X1 U9141 ( .A1(n9759), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7372) );
  NAND2_X1 U9142 ( .A1(n9756), .A2(n7372), .ZN(n7834) );
  NAND2_X1 U9143 ( .A1(n7835), .A2(n7834), .ZN(n7833) );
  OR2_X1 U9144 ( .A1(n7839), .A2(n10513), .ZN(n7373) );
  NAND2_X1 U9145 ( .A1(n7833), .A2(n7373), .ZN(n9769) );
  XNOR2_X1 U9146 ( .A(n7396), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9770) );
  NAND2_X1 U9147 ( .A1(n9769), .A2(n9770), .ZN(n9768) );
  INV_X1 U9148 ( .A(n7396), .ZN(n9767) );
  NAND2_X1 U9149 ( .A1(n9767), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7374) );
  NAND2_X1 U9150 ( .A1(n9768), .A2(n7374), .ZN(n7848) );
  XNOR2_X1 U9151 ( .A(n7856), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U9152 ( .A1(n7848), .A2(n7849), .ZN(n7847) );
  INV_X1 U9153 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7375) );
  OR2_X1 U9154 ( .A1(n7856), .A2(n7375), .ZN(n7376) );
  NAND2_X1 U9155 ( .A1(n7847), .A2(n7376), .ZN(n9782) );
  XNOR2_X1 U9156 ( .A(n7400), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9783) );
  NAND2_X1 U9157 ( .A1(n9782), .A2(n9783), .ZN(n9781) );
  INV_X1 U9158 ( .A(n7400), .ZN(n9780) );
  NAND2_X1 U9159 ( .A1(n9780), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7377) );
  NAND2_X1 U9160 ( .A1(n9781), .A2(n7377), .ZN(n9796) );
  XNOR2_X1 U9161 ( .A(n9790), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9797) );
  NAND2_X1 U9162 ( .A1(n9796), .A2(n9797), .ZN(n9795) );
  INV_X1 U9163 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7378) );
  OR2_X1 U9164 ( .A1(n9790), .A2(n7378), .ZN(n7379) );
  NAND2_X1 U9165 ( .A1(n9795), .A2(n7379), .ZN(n9813) );
  MUX2_X1 U9166 ( .A(n7380), .B(P1_REG1_REG_7__SCAN_IN), .S(n9804), .Z(n9814)
         );
  OR2_X1 U9167 ( .A1(n9804), .A2(n7380), .ZN(n7381) );
  NAND2_X1 U9168 ( .A1(n9812), .A2(n7381), .ZN(n9827) );
  XNOR2_X1 U9169 ( .A(n9821), .B(n7382), .ZN(n9826) );
  NAND2_X1 U9170 ( .A1(n9827), .A2(n9826), .ZN(n9825) );
  NAND2_X1 U9171 ( .A1(n9821), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7383) );
  NAND2_X1 U9172 ( .A1(n9825), .A2(n7383), .ZN(n7385) );
  INV_X1 U9173 ( .A(n7487), .ZN(n7384) );
  AOI21_X1 U9174 ( .B1(n7386), .B2(n7385), .A(n7384), .ZN(n7414) );
  NAND2_X1 U9175 ( .A1(n7388), .A2(n7387), .ZN(n10235) );
  OR2_X1 U9176 ( .A1(n10235), .A2(n7831), .ZN(n9868) );
  INV_X1 U9177 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7391) );
  NOR2_X1 U9178 ( .A1(n7389), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8568) );
  INV_X1 U9179 ( .A(n8568), .ZN(n7390) );
  OAI21_X1 U9180 ( .B1(n10308), .B2(n7391), .A(n7390), .ZN(n7412) );
  INV_X1 U9181 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7610) );
  AND2_X1 U9182 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9754) );
  NAND2_X1 U9183 ( .A1(n9759), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7393) );
  NAND2_X1 U9184 ( .A1(n9753), .A2(n7393), .ZN(n7837) );
  NAND2_X1 U9185 ( .A1(n7838), .A2(n7837), .ZN(n7836) );
  OR2_X1 U9186 ( .A1(n7839), .A2(n7394), .ZN(n7395) );
  NAND2_X1 U9187 ( .A1(n7836), .A2(n7395), .ZN(n9772) );
  XNOR2_X1 U9188 ( .A(n7396), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9773) );
  NAND2_X1 U9189 ( .A1(n9772), .A2(n9773), .ZN(n9771) );
  NAND2_X1 U9190 ( .A1(n9767), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7397) );
  NAND2_X1 U9191 ( .A1(n9771), .A2(n7397), .ZN(n7853) );
  XNOR2_X1 U9192 ( .A(n7856), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U9193 ( .A1(n7853), .A2(n7854), .ZN(n7852) );
  OR2_X1 U9194 ( .A1(n7856), .A2(n7398), .ZN(n7399) );
  NAND2_X1 U9195 ( .A1(n7852), .A2(n7399), .ZN(n9785) );
  XNOR2_X1 U9196 ( .A(n7400), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9786) );
  NAND2_X1 U9197 ( .A1(n9785), .A2(n9786), .ZN(n9784) );
  NAND2_X1 U9198 ( .A1(n9780), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7401) );
  NAND2_X1 U9199 ( .A1(n9784), .A2(n7401), .ZN(n9799) );
  XNOR2_X1 U9200 ( .A(n9790), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9800) );
  NAND2_X1 U9201 ( .A1(n9799), .A2(n9800), .ZN(n9798) );
  OR2_X1 U9202 ( .A1(n9790), .A2(n7402), .ZN(n7403) );
  NAND2_X1 U9203 ( .A1(n9798), .A2(n7403), .ZN(n9810) );
  MUX2_X1 U9204 ( .A(n7404), .B(P1_REG2_REG_7__SCAN_IN), .S(n9804), .Z(n9811)
         );
  OR2_X1 U9205 ( .A1(n9804), .A2(n7404), .ZN(n7405) );
  NAND2_X1 U9206 ( .A1(n9809), .A2(n7405), .ZN(n9824) );
  XNOR2_X1 U9207 ( .A(n9821), .B(n7563), .ZN(n9823) );
  NAND2_X1 U9208 ( .A1(n9824), .A2(n9823), .ZN(n9822) );
  NAND2_X1 U9209 ( .A1(n9821), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7406) );
  NAND2_X1 U9210 ( .A1(n9822), .A2(n7406), .ZN(n7408) );
  XNOR2_X1 U9211 ( .A(n7491), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7407) );
  NAND2_X1 U9212 ( .A1(n7408), .A2(n7407), .ZN(n7410) );
  OR2_X1 U9213 ( .A1(n6115), .A2(n6123), .ZN(n7409) );
  AOI21_X1 U9214 ( .B1(n7493), .B2(n7410), .A(n10269), .ZN(n7411) );
  AOI211_X1 U9215 ( .C1(n10305), .C2(n7491), .A(n7412), .B(n7411), .ZN(n7413)
         );
  OAI21_X1 U9216 ( .B1(n7414), .B2(n10299), .A(n7413), .ZN(P1_U3252) );
  INV_X1 U9217 ( .A(n7429), .ZN(n7415) );
  AOI21_X1 U9218 ( .B1(n7417), .B2(n7416), .A(n7415), .ZN(n7426) );
  AND2_X1 U9219 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7822) );
  NOR2_X1 U9220 ( .A1(n9154), .A2(n7418), .ZN(n7419) );
  AOI211_X1 U9221 ( .C1(n9210), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n7822), .B(
        n7419), .ZN(n7425) );
  XNOR2_X1 U9222 ( .A(n7421), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n7422) );
  AOI22_X1 U9223 ( .A1(n9146), .A2(n7423), .B1(n9173), .B2(n7422), .ZN(n7424)
         );
  OAI211_X1 U9224 ( .C1(n7426), .C2(n9159), .A(n7425), .B(n7424), .ZN(P2_U3185) );
  AOI21_X1 U9225 ( .B1(n7429), .B2(n7428), .A(n7427), .ZN(n7446) );
  NAND2_X1 U9226 ( .A1(n7430), .A2(n9215), .ZN(n7445) );
  NOR2_X1 U9227 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4833), .ZN(n7949) );
  NOR2_X1 U9228 ( .A1(n9154), .A2(n7431), .ZN(n7432) );
  AOI211_X1 U9229 ( .C1(n9210), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7949), .B(
        n7432), .ZN(n7444) );
  OAI21_X1 U9230 ( .B1(n7435), .B2(n7434), .A(n7433), .ZN(n7442) );
  INV_X1 U9231 ( .A(n7436), .ZN(n7438) );
  NAND3_X1 U9232 ( .A1(n7420), .A2(n7438), .A3(n7437), .ZN(n7439) );
  AOI21_X1 U9233 ( .B1(n7440), .B2(n7439), .A(n9217), .ZN(n7441) );
  AOI21_X1 U9234 ( .B1(n9173), .B2(n7442), .A(n7441), .ZN(n7443) );
  OAI211_X1 U9235 ( .C1(n7446), .C2(n7445), .A(n7444), .B(n7443), .ZN(P2_U3186) );
  INV_X1 U9236 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7447) );
  OAI222_X1 U9237 ( .A1(n9547), .A2(n7527), .B1(n9084), .B2(P2_U3151), .C1(
        n7447), .C2(n9537), .ZN(P2_U3282) );
  NAND3_X1 U9238 ( .A1(n7449), .A2(n7534), .A3(n7448), .ZN(n7458) );
  NAND3_X1 U9239 ( .A1(n7480), .A2(n7450), .A3(n7455), .ZN(n7453) );
  NOR2_X1 U9240 ( .A1(n7451), .A2(n9703), .ZN(n7536) );
  INV_X1 U9241 ( .A(n7536), .ZN(n7452) );
  OAI211_X1 U9242 ( .C1(n10382), .C2(n7454), .A(n7453), .B(n7452), .ZN(n7460)
         );
  INV_X1 U9243 ( .A(n6515), .ZN(n7457) );
  NOR4_X1 U9244 ( .A1(n7458), .A2(n7457), .A3(n7456), .A4(n7455), .ZN(n7459)
         );
  AOI21_X1 U9245 ( .B1(n10324), .B2(n7460), .A(n7459), .ZN(n7461) );
  OAI21_X1 U9246 ( .B1(n7829), .B2(n10324), .A(n7461), .ZN(P1_U3293) );
  INV_X1 U9247 ( .A(n7868), .ZN(n7462) );
  AOI21_X1 U9248 ( .B1(n7464), .B2(n7463), .A(n7462), .ZN(n7479) );
  OAI21_X1 U9249 ( .B1(n7467), .B2(n7466), .A(n7465), .ZN(n7477) );
  INV_X1 U9250 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7475) );
  AND3_X1 U9251 ( .A1(n7362), .A2(n7469), .A3(n7468), .ZN(n7470) );
  OAI21_X1 U9252 ( .B1(n7471), .B2(n7470), .A(n9146), .ZN(n7474) );
  AND2_X1 U9253 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8061) );
  AOI21_X1 U9254 ( .B1(n9209), .B2(n7472), .A(n8061), .ZN(n7473) );
  OAI211_X1 U9255 ( .C1(n9171), .C2(n7475), .A(n7474), .B(n7473), .ZN(n7476)
         );
  AOI21_X1 U9256 ( .B1(n9173), .B2(n7477), .A(n7476), .ZN(n7478) );
  OAI21_X1 U9257 ( .B1(n7479), .B2(n9159), .A(n7478), .ZN(P2_U3188) );
  INV_X1 U9258 ( .A(n7480), .ZN(n7481) );
  AOI21_X1 U9259 ( .B1(n10048), .B2(n10153), .A(n7481), .ZN(n7482) );
  AOI211_X1 U9260 ( .C1(n7483), .C2(n7953), .A(n7536), .B(n7482), .ZN(n10425)
         );
  NAND2_X1 U9261 ( .A1(n10526), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7484) );
  OAI21_X1 U9262 ( .B1(n10425), .B2(n10526), .A(n7484), .ZN(P1_U3522) );
  INV_X1 U9263 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7485) );
  MUX2_X1 U9264 ( .A(n7485), .B(P1_REG1_REG_10__SCAN_IN), .S(n7884), .Z(n7490)
         );
  OR2_X1 U9265 ( .A1(n7491), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7486) );
  INV_X1 U9266 ( .A(n7878), .ZN(n7488) );
  AOI211_X1 U9267 ( .C1(n7490), .C2(n7489), .A(n10299), .B(n7488), .ZN(n7501)
         );
  XNOR2_X1 U9268 ( .A(n7884), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7496) );
  OR2_X1 U9269 ( .A1(n7491), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7492) );
  INV_X1 U9270 ( .A(n7886), .ZN(n7494) );
  AOI211_X1 U9271 ( .C1(n7496), .C2(n7495), .A(n10269), .B(n7494), .ZN(n7500)
         );
  INV_X1 U9272 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7498) );
  NAND2_X1 U9273 ( .A1(n10305), .A2(n7884), .ZN(n7497) );
  NAND2_X1 U9274 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8554) );
  OAI211_X1 U9275 ( .C1(n10308), .C2(n7498), .A(n7497), .B(n8554), .ZN(n7499)
         );
  OR3_X1 U9276 ( .A1(n7501), .A2(n7500), .A3(n7499), .ZN(P1_U3253) );
  INV_X1 U9277 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7509) );
  MUX2_X1 U9278 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n4401), .Z(n7502) );
  NAND2_X1 U9279 ( .A1(n7502), .A2(n5142), .ZN(n7503) );
  AOI22_X1 U9280 ( .A1(n9159), .A2(n7505), .B1(n7504), .B2(n7503), .ZN(n7506)
         );
  AOI21_X1 U9281 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n7506), .ZN(
        n7508) );
  NAND2_X1 U9282 ( .A1(n9209), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7507) );
  OAI211_X1 U9283 ( .C1(n7509), .C2(n9171), .A(n7508), .B(n7507), .ZN(P2_U3182) );
  XOR2_X1 U9284 ( .A(n7510), .B(n7511), .Z(n7525) );
  INV_X1 U9285 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7523) );
  OAI21_X1 U9286 ( .B1(n7514), .B2(n7513), .A(n7512), .ZN(n7519) );
  OAI21_X1 U9287 ( .B1(n7517), .B2(n7516), .A(n7515), .ZN(n7518) );
  AOI22_X1 U9288 ( .A1(n9146), .A2(n7519), .B1(n9173), .B2(n7518), .ZN(n7522)
         );
  AOI22_X1 U9289 ( .A1(n9209), .A2(n7520), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n7521) );
  OAI211_X1 U9290 ( .C1(n7523), .C2(n9171), .A(n7522), .B(n7521), .ZN(n7524)
         );
  AOI21_X1 U9291 ( .B1(n9215), .B2(n7525), .A(n7524), .ZN(n7526) );
  INV_X1 U9292 ( .A(n7526), .ZN(P2_U3184) );
  INV_X1 U9293 ( .A(n9853), .ZN(n7528) );
  OAI222_X1 U9294 ( .A1(P1_U3086), .A2(n7528), .B1(n10224), .B2(n7793), .C1(
        n7527), .C2(n8271), .ZN(P1_U3342) );
  AND2_X1 U9295 ( .A1(n7529), .A2(n7814), .ZN(n8870) );
  OR2_X1 U9296 ( .A1(n8870), .A2(n8867), .ZN(n7975) );
  INV_X1 U9297 ( .A(n7975), .ZN(n8815) );
  NAND2_X1 U9298 ( .A1(n8748), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7549) );
  NAND2_X1 U9299 ( .A1(n7549), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7531) );
  AOI22_X1 U9300 ( .A1(n8779), .A2(n4404), .B1(n8784), .B2(n7982), .ZN(n7530)
         );
  OAI211_X1 U9301 ( .C1(n8786), .C2(n8815), .A(n7531), .B(n7530), .ZN(P2_U3172) );
  XNOR2_X1 U9302 ( .A(n7532), .B(n7533), .ZN(n7828) );
  NAND2_X1 U9303 ( .A1(n9693), .A2(n7953), .ZN(n7538) );
  NAND2_X1 U9304 ( .A1(n7535), .A2(n7534), .ZN(n7919) );
  AOI22_X1 U9305 ( .A1(n9710), .A2(n7536), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n7919), .ZN(n7537) );
  OAI211_X1 U9306 ( .C1(n7828), .C2(n9695), .A(n7538), .B(n7537), .ZN(P1_U3232) );
  XOR2_X1 U9307 ( .A(n7540), .B(n7539), .Z(n7544) );
  AOI22_X1 U9308 ( .A1(n8793), .A2(n4404), .B1(n8779), .B2(n9035), .ZN(n7541)
         );
  OAI21_X1 U9309 ( .B1(n4774), .B2(n8800), .A(n7541), .ZN(n7542) );
  AOI21_X1 U9310 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7549), .A(n7542), .ZN(
        n7543) );
  OAI21_X1 U9311 ( .B1(n7544), .B2(n8786), .A(n7543), .ZN(P2_U3177) );
  XOR2_X1 U9312 ( .A(n7545), .B(n7546), .Z(n7551) );
  AOI22_X1 U9313 ( .A1(n8779), .A2(n7057), .B1(n8793), .B2(n7529), .ZN(n7547)
         );
  OAI21_X1 U9314 ( .B1(n8800), .B2(n8868), .A(n7547), .ZN(n7548) );
  AOI21_X1 U9315 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7549), .A(n7548), .ZN(
        n7550) );
  OAI21_X1 U9316 ( .B1(n8786), .B2(n7551), .A(n7550), .ZN(P2_U3162) );
  OR2_X1 U9317 ( .A1(n7552), .A2(n9701), .ZN(n7554) );
  OR2_X1 U9318 ( .A1(n8100), .A2(n9703), .ZN(n7553) );
  NAND2_X1 U9319 ( .A1(n7554), .A2(n7553), .ZN(n7962) );
  AOI22_X1 U9320 ( .A1(n9710), .A2(n7962), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n7919), .ZN(n7560) );
  OAI21_X1 U9321 ( .B1(n7557), .B2(n7556), .A(n7555), .ZN(n7558) );
  NAND2_X1 U9322 ( .A1(n7558), .A2(n9716), .ZN(n7559) );
  OAI211_X1 U9323 ( .C1(n10429), .C2(n9725), .A(n7560), .B(n7559), .ZN(
        P1_U3222) );
  MUX2_X1 U9324 ( .A(n9664), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9738), .Z(n7812) );
  NOR4_X1 U9325 ( .A1(SI_15_), .A2(P1_REG3_REG_21__SCAN_IN), .A3(
        P2_ADDR_REG_10__SCAN_IN), .A4(n7676), .ZN(n7561) );
  NAND3_X1 U9326 ( .A1(SI_21_), .A2(P1_REG1_REG_25__SCAN_IN), .A3(n7561), .ZN(
        n7572) );
  NAND4_X1 U9327 ( .A1(n7563), .A2(n7562), .A3(P1_REG2_REG_2__SCAN_IN), .A4(
        n10214), .ZN(n7564) );
  NOR3_X1 U9328 ( .A1(n7564), .A2(P1_REG0_REG_15__SCAN_IN), .A3(n7693), .ZN(
        n7570) );
  NAND4_X1 U9329 ( .A1(P2_REG0_REG_3__SCAN_IN), .A2(n6127), .A3(n8671), .A4(
        n9101), .ZN(n7568) );
  NAND4_X1 U9330 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P1_DATAO_REG_23__SCAN_IN), 
        .A3(n7648), .A4(n8067), .ZN(n7567) );
  NAND4_X1 U9331 ( .A1(SI_26_), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P2_ADDR_REG_15__SCAN_IN), .A4(n7670), .ZN(n7566) );
  NAND4_X1 U9332 ( .A1(SI_5_), .A2(P1_REG1_REG_10__SCAN_IN), .A3(
        P2_IR_REG_22__SCAN_IN), .A4(P2_REG0_REG_4__SCAN_IN), .ZN(n7565) );
  NOR4_X1 U9333 ( .A1(n7568), .A2(n7567), .A3(n7566), .A4(n7565), .ZN(n7569)
         );
  NAND4_X1 U9334 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P2_REG0_REG_24__SCAN_IN), 
        .A3(n7570), .A4(n7569), .ZN(n7571) );
  NOR4_X1 U9335 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_REG0_REG_20__SCAN_IN), 
        .A3(n7572), .A4(n7571), .ZN(n7609) );
  INV_X1 U9336 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7709) );
  NAND4_X1 U9337 ( .A1(n7574), .A2(n7573), .A3(P1_ADDR_REG_6__SCAN_IN), .A4(
        n7709), .ZN(n7607) );
  INV_X1 U9338 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10263) );
  NOR4_X1 U9339 ( .A1(P2_REG0_REG_16__SCAN_IN), .A2(P1_REG2_REG_27__SCAN_IN), 
        .A3(n6102), .A4(n10263), .ZN(n7581) );
  INV_X1 U9340 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n7772) );
  NOR4_X1 U9341 ( .A1(P1_REG0_REG_2__SCAN_IN), .A2(P1_REG1_REG_17__SCAN_IN), 
        .A3(P2_WR_REG_SCAN_IN), .A4(n7772), .ZN(n7580) );
  NAND4_X1 U9342 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG0_REG_26__SCAN_IN), 
        .A3(n6377), .A4(n8443), .ZN(n7578) );
  NAND4_X1 U9343 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_REG0_REG_16__SCAN_IN), 
        .A3(P2_D_REG_10__SCAN_IN), .A4(P2_REG3_REG_28__SCAN_IN), .ZN(n7577) );
  NAND4_X1 U9344 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P2_REG2_REG_8__SCAN_IN), 
        .A3(n10179), .A4(n7787), .ZN(n7576) );
  NAND4_X1 U9345 ( .A1(P1_REG0_REG_1__SCAN_IN), .A2(P2_REG0_REG_0__SCAN_IN), 
        .A3(n7793), .A4(n7796), .ZN(n7575) );
  NOR4_X1 U9346 ( .A1(n7578), .A2(n7577), .A3(n7576), .A4(n7575), .ZN(n7579)
         );
  NAND3_X1 U9347 ( .A1(n7581), .A2(n7580), .A3(n7579), .ZN(n7606) );
  NAND4_X1 U9348 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P2_REG1_REG_18__SCAN_IN), 
        .A3(n4833), .A4(n5461), .ZN(n7585) );
  INV_X1 U9349 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8427) );
  INV_X1 U9350 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7708) );
  NAND4_X1 U9351 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_REG2_REG_29__SCAN_IN), 
        .A3(n8427), .A4(n7708), .ZN(n7584) );
  NAND4_X1 U9352 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(P2_DATAO_REG_23__SCAN_IN), .A3(P1_REG1_REG_0__SCAN_IN), .A4(P2_REG1_REG_15__SCAN_IN), .ZN(n7583) );
  NAND4_X1 U9353 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .A3(P2_ADDR_REG_17__SCAN_IN), .A4(n7382), .ZN(n7582) );
  NOR4_X1 U9354 ( .A1(n7585), .A2(n7584), .A3(n7583), .A4(n7582), .ZN(n7604)
         );
  INV_X1 U9355 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n7725) );
  INV_X1 U9356 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7724) );
  NAND4_X1 U9357 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(P1_DATAO_REG_0__SCAN_IN), 
        .A3(n7725), .A4(n7724), .ZN(n7586) );
  NOR3_X1 U9358 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .A3(n7586), .ZN(n7587) );
  NAND3_X1 U9359 ( .A1(n7587), .A2(P1_DATAO_REG_29__SCAN_IN), .A3(
        P2_DATAO_REG_2__SCAN_IN), .ZN(n7590) );
  NAND4_X1 U9360 ( .A1(P2_REG1_REG_27__SCAN_IN), .A2(P1_REG2_REG_30__SCAN_IN), 
        .A3(n6319), .A4(n9373), .ZN(n7589) );
  NAND4_X1 U9361 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P2_DATAO_REG_8__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n7588) );
  NOR3_X1 U9362 ( .A1(n7590), .A2(n7589), .A3(n7588), .ZN(n7603) );
  NAND4_X1 U9363 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .A3(
        P2_DATAO_REG_28__SCAN_IN), .A4(P1_ADDR_REG_13__SCAN_IN), .ZN(n7594) );
  INV_X1 U9364 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7637) );
  INV_X1 U9365 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8758) );
  NAND4_X1 U9366 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P2_REG2_REG_21__SCAN_IN), 
        .A3(n8758), .A4(n8397), .ZN(n7592) );
  INV_X1 U9367 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7624) );
  NAND4_X1 U9368 ( .A1(n7625), .A2(n7404), .A3(n7624), .A4(n6863), .ZN(n7591)
         );
  OR4_X1 U9369 ( .A1(n7637), .A2(n9168), .A3(n7592), .A4(n7591), .ZN(n7593) );
  NOR4_X1 U9370 ( .A1(n7594), .A2(n7593), .A3(P2_IR_REG_14__SCAN_IN), .A4(
        n8582), .ZN(n7602) );
  NAND4_X1 U9371 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(n8129), .ZN(n7600) );
  INV_X1 U9372 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10256) );
  INV_X1 U9373 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7734) );
  NAND4_X1 U9374 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .A3(n10256), .A4(n7734), .ZN(n7597) );
  NAND4_X1 U9375 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .A3(n7595), .A4(n8547), .ZN(n7596) );
  OR4_X1 U9376 ( .A1(n7610), .A2(P2_IR_REG_28__SCAN_IN), .A3(n7597), .A4(n7596), .ZN(n7599) );
  NOR4_X1 U9377 ( .A1(n7600), .A2(n7599), .A3(n7598), .A4(n7611), .ZN(n7601)
         );
  NAND4_X1 U9378 ( .A1(n7604), .A2(n7603), .A3(n7602), .A4(n7601), .ZN(n7605)
         );
  NOR4_X1 U9379 ( .A1(n4841), .A2(n7607), .A3(n7606), .A4(n7605), .ZN(n7608)
         );
  AOI21_X1 U9380 ( .B1(n7609), .B2(n7608), .A(P2_IR_REG_23__SCAN_IN), .ZN(
        n7810) );
  XOR2_X1 U9381 ( .A(n7598), .B(keyinput113), .Z(n7615) );
  XOR2_X1 U9382 ( .A(n7610), .B(keyinput35), .Z(n7614) );
  XNOR2_X1 U9383 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput92), .ZN(n7613) );
  XNOR2_X1 U9384 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput24), .ZN(n7612) );
  NAND4_X1 U9385 ( .A1(n7615), .A2(n7614), .A3(n7613), .A4(n7612), .ZN(n7621)
         );
  XNOR2_X1 U9386 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput9), .ZN(n7619) );
  XNOR2_X1 U9387 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput26), .ZN(n7618) );
  XNOR2_X1 U9388 ( .A(P2_REG0_REG_14__SCAN_IN), .B(keyinput50), .ZN(n7617) );
  XNOR2_X1 U9389 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput67), .ZN(n7616) );
  NAND4_X1 U9390 ( .A1(n7619), .A2(n7618), .A3(n7617), .A4(n7616), .ZN(n7620)
         );
  NOR2_X1 U9391 ( .A1(n7621), .A2(n7620), .ZN(n7658) );
  AOI22_X1 U9392 ( .A1(n8129), .A2(keyinput48), .B1(n6070), .B2(keyinput45), 
        .ZN(n7622) );
  OAI221_X1 U9393 ( .B1(n8129), .B2(keyinput48), .C1(n6070), .C2(keyinput45), 
        .A(n7622), .ZN(n7629) );
  AOI22_X1 U9394 ( .A1(n7625), .A2(keyinput104), .B1(keyinput116), .B2(n7624), 
        .ZN(n7623) );
  OAI221_X1 U9395 ( .B1(n7625), .B2(keyinput104), .C1(n7624), .C2(keyinput116), 
        .A(n7623), .ZN(n7628) );
  XNOR2_X1 U9396 ( .A(n7626), .B(keyinput13), .ZN(n7627) );
  OR3_X1 U9397 ( .A1(n7629), .A2(n7628), .A3(n7627), .ZN(n7634) );
  AOI22_X1 U9398 ( .A1(n7404), .A2(keyinput83), .B1(keyinput94), .B2(n6863), 
        .ZN(n7630) );
  OAI221_X1 U9399 ( .B1(n7404), .B2(keyinput83), .C1(n6863), .C2(keyinput94), 
        .A(n7630), .ZN(n7633) );
  INV_X1 U9400 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n7631) );
  XNOR2_X1 U9401 ( .A(n7631), .B(keyinput7), .ZN(n7632) );
  NOR3_X1 U9402 ( .A1(n7634), .A2(n7633), .A3(n7632), .ZN(n7657) );
  AOI22_X1 U9403 ( .A1(n8758), .A2(keyinput46), .B1(keyinput44), .B2(n9307), 
        .ZN(n7635) );
  OAI221_X1 U9404 ( .B1(n8758), .B2(keyinput46), .C1(n9307), .C2(keyinput44), 
        .A(n7635), .ZN(n7644) );
  AOI22_X1 U9405 ( .A1(n7637), .A2(keyinput53), .B1(keyinput6), .B2(n9168), 
        .ZN(n7636) );
  OAI221_X1 U9406 ( .B1(n7637), .B2(keyinput53), .C1(n9168), .C2(keyinput6), 
        .A(n7636), .ZN(n7643) );
  XNOR2_X1 U9407 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput49), .ZN(n7641) );
  XNOR2_X1 U9408 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput70), .ZN(n7640) );
  XNOR2_X1 U9409 ( .A(P2_REG1_REG_10__SCAN_IN), .B(keyinput31), .ZN(n7639) );
  XNOR2_X1 U9410 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput38), .ZN(n7638) );
  NAND4_X1 U9411 ( .A1(n7641), .A2(n7640), .A3(n7639), .A4(n7638), .ZN(n7642)
         );
  NOR3_X1 U9412 ( .A1(n7644), .A2(n7643), .A3(n7642), .ZN(n7656) );
  AOI22_X1 U9413 ( .A1(n6399), .A2(keyinput76), .B1(P1_U3086), .B2(keyinput117), .ZN(n7645) );
  OAI221_X1 U9414 ( .B1(n6399), .B2(keyinput76), .C1(P1_U3086), .C2(
        keyinput117), .A(n7645), .ZN(n7654) );
  INV_X1 U9415 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n8355) );
  AOI22_X1 U9416 ( .A1(n8355), .A2(keyinput41), .B1(n8640), .B2(keyinput72), 
        .ZN(n7646) );
  OAI221_X1 U9417 ( .B1(n8355), .B2(keyinput41), .C1(n8640), .C2(keyinput72), 
        .A(n7646), .ZN(n7653) );
  AOI22_X1 U9418 ( .A1(n8067), .A2(keyinput105), .B1(n7648), .B2(keyinput86), 
        .ZN(n7647) );
  OAI221_X1 U9419 ( .B1(n8067), .B2(keyinput105), .C1(n7648), .C2(keyinput86), 
        .A(n7647), .ZN(n7652) );
  INV_X1 U9420 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n7650) );
  AOI22_X1 U9421 ( .A1(n7650), .A2(keyinput95), .B1(n8454), .B2(keyinput82), 
        .ZN(n7649) );
  OAI221_X1 U9422 ( .B1(n7650), .B2(keyinput95), .C1(n8454), .C2(keyinput82), 
        .A(n7649), .ZN(n7651) );
  NOR4_X1 U9423 ( .A1(n7654), .A2(n7653), .A3(n7652), .A4(n7651), .ZN(n7655)
         );
  NAND4_X1 U9424 ( .A1(n7658), .A2(n7657), .A3(n7656), .A4(n7655), .ZN(n7808)
         );
  AOI22_X1 U9425 ( .A1(n5425), .A2(keyinput51), .B1(n6127), .B2(keyinput120), 
        .ZN(n7659) );
  OAI221_X1 U9426 ( .B1(n5425), .B2(keyinput51), .C1(n6127), .C2(keyinput120), 
        .A(n7659), .ZN(n7667) );
  AOI22_X1 U9427 ( .A1(n8671), .A2(keyinput57), .B1(keyinput2), .B2(n9101), 
        .ZN(n7660) );
  OAI221_X1 U9428 ( .B1(n8671), .B2(keyinput57), .C1(n9101), .C2(keyinput2), 
        .A(n7660), .ZN(n7666) );
  INV_X1 U9429 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10419) );
  XNOR2_X1 U9430 ( .A(n10419), .B(keyinput110), .ZN(n7665) );
  XOR2_X1 U9431 ( .A(n5448), .B(keyinput22), .Z(n7663) );
  XNOR2_X1 U9432 ( .A(SI_5_), .B(keyinput73), .ZN(n7662) );
  XNOR2_X1 U9433 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput52), .ZN(n7661) );
  NAND3_X1 U9434 ( .A1(n7663), .A2(n7662), .A3(n7661), .ZN(n7664) );
  NOR4_X1 U9435 ( .A1(n7667), .A2(n7666), .A3(n7665), .A4(n7664), .ZN(n7706)
         );
  INV_X1 U9436 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9110) );
  AOI22_X1 U9437 ( .A1(n7485), .A2(keyinput14), .B1(keyinput125), .B2(n9110), 
        .ZN(n7668) );
  OAI221_X1 U9438 ( .B1(n7485), .B2(keyinput14), .C1(n9110), .C2(keyinput125), 
        .A(n7668), .ZN(n7680) );
  INV_X1 U9439 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U9440 ( .A1(n7670), .A2(keyinput32), .B1(n10417), .B2(keyinput58), 
        .ZN(n7669) );
  OAI221_X1 U9441 ( .B1(n7670), .B2(keyinput32), .C1(n10417), .C2(keyinput58), 
        .A(n7669), .ZN(n7679) );
  AOI22_X1 U9442 ( .A1(n7673), .A2(keyinput27), .B1(keyinput118), .B2(n7672), 
        .ZN(n7671) );
  OAI221_X1 U9443 ( .B1(n7673), .B2(keyinput27), .C1(n7672), .C2(keyinput118), 
        .A(n7671), .ZN(n7678) );
  AOI22_X1 U9444 ( .A1(n7676), .A2(keyinput28), .B1(n7675), .B2(keyinput54), 
        .ZN(n7674) );
  OAI221_X1 U9445 ( .B1(n7676), .B2(keyinput28), .C1(n7675), .C2(keyinput54), 
        .A(n7674), .ZN(n7677) );
  NOR4_X1 U9446 ( .A1(n7680), .A2(n7679), .A3(n7678), .A4(n7677), .ZN(n7705)
         );
  INV_X1 U9447 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9596) );
  AOI22_X1 U9448 ( .A1(n9596), .A2(keyinput25), .B1(n6368), .B2(keyinput77), 
        .ZN(n7681) );
  OAI221_X1 U9449 ( .B1(n9596), .B2(keyinput25), .C1(n6368), .C2(keyinput77), 
        .A(n7681), .ZN(n7691) );
  INV_X1 U9450 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7683) );
  AOI22_X1 U9451 ( .A1(n7684), .A2(keyinput20), .B1(keyinput115), .B2(n7683), 
        .ZN(n7682) );
  OAI221_X1 U9452 ( .B1(n7684), .B2(keyinput20), .C1(n7683), .C2(keyinput115), 
        .A(n7682), .ZN(n7690) );
  INV_X1 U9453 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U9454 ( .A1(n10214), .A2(keyinput75), .B1(n10203), .B2(keyinput8), 
        .ZN(n7685) );
  OAI221_X1 U9455 ( .B1(n10214), .B2(keyinput75), .C1(n10203), .C2(keyinput8), 
        .A(n7685), .ZN(n7689) );
  XNOR2_X1 U9456 ( .A(P1_REG0_REG_20__SCAN_IN), .B(keyinput81), .ZN(n7687) );
  XNOR2_X1 U9457 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput16), .ZN(n7686) );
  NAND2_X1 U9458 ( .A1(n7687), .A2(n7686), .ZN(n7688) );
  NOR4_X1 U9459 ( .A1(n7691), .A2(n7690), .A3(n7689), .A4(n7688), .ZN(n7704)
         );
  INV_X1 U9460 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9792) );
  AOI22_X1 U9461 ( .A1(n9792), .A2(keyinput37), .B1(n7693), .B2(keyinput101), 
        .ZN(n7692) );
  OAI221_X1 U9462 ( .B1(n9792), .B2(keyinput37), .C1(n7693), .C2(keyinput101), 
        .A(n7692), .ZN(n7702) );
  AOI22_X1 U9463 ( .A1(n7394), .A2(keyinput55), .B1(n7563), .B2(keyinput119), 
        .ZN(n7694) );
  OAI221_X1 U9464 ( .B1(n7394), .B2(keyinput55), .C1(n7563), .C2(keyinput119), 
        .A(n7694), .ZN(n7701) );
  INV_X1 U9465 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n7696) );
  AOI22_X1 U9466 ( .A1(n7696), .A2(keyinput11), .B1(keyinput97), .B2(n4841), 
        .ZN(n7695) );
  OAI221_X1 U9467 ( .B1(n7696), .B2(keyinput11), .C1(n4841), .C2(keyinput97), 
        .A(n7695), .ZN(n7700) );
  XNOR2_X1 U9468 ( .A(P2_REG0_REG_24__SCAN_IN), .B(keyinput102), .ZN(n7698) );
  XNOR2_X1 U9469 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput103), .ZN(n7697) );
  NAND2_X1 U9470 ( .A1(n7698), .A2(n7697), .ZN(n7699) );
  NOR4_X1 U9471 ( .A1(n7702), .A2(n7701), .A3(n7700), .A4(n7699), .ZN(n7703)
         );
  NAND4_X1 U9472 ( .A1(n7706), .A2(n7705), .A3(n7704), .A4(n7703), .ZN(n7807)
         );
  AOI22_X1 U9473 ( .A1(n7709), .A2(keyinput21), .B1(n7708), .B2(keyinput71), 
        .ZN(n7707) );
  OAI221_X1 U9474 ( .B1(n7709), .B2(keyinput21), .C1(n7708), .C2(keyinput71), 
        .A(n7707), .ZN(n7719) );
  INV_X1 U9475 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n7712) );
  INV_X1 U9476 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n7711) );
  AOI22_X1 U9477 ( .A1(n7712), .A2(keyinput47), .B1(keyinput30), .B2(n7711), 
        .ZN(n7710) );
  OAI221_X1 U9478 ( .B1(n7712), .B2(keyinput47), .C1(n7711), .C2(keyinput30), 
        .A(n7710), .ZN(n7718) );
  AOI22_X1 U9479 ( .A1(n5461), .A2(keyinput63), .B1(n7714), .B2(keyinput74), 
        .ZN(n7713) );
  OAI221_X1 U9480 ( .B1(n5461), .B2(keyinput63), .C1(n7714), .C2(keyinput74), 
        .A(n7713), .ZN(n7717) );
  AOI22_X1 U9481 ( .A1(n8427), .A2(keyinput5), .B1(keyinput121), .B2(n8642), 
        .ZN(n7715) );
  OAI221_X1 U9482 ( .B1(n8427), .B2(keyinput5), .C1(n8642), .C2(keyinput121), 
        .A(n7715), .ZN(n7716) );
  NOR4_X1 U9483 ( .A1(n7719), .A2(n7718), .A3(n7717), .A4(n7716), .ZN(n7757)
         );
  AOI22_X1 U9484 ( .A1(n6319), .A2(keyinput114), .B1(keyinput112), .B2(n7721), 
        .ZN(n7720) );
  OAI221_X1 U9485 ( .B1(n6319), .B2(keyinput114), .C1(n7721), .C2(keyinput112), 
        .A(n7720), .ZN(n7731) );
  INV_X1 U9486 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10420) );
  AOI22_X1 U9487 ( .A1(n10420), .A2(keyinput34), .B1(keyinput106), .B2(n9373), 
        .ZN(n7722) );
  OAI221_X1 U9488 ( .B1(n10420), .B2(keyinput34), .C1(n9373), .C2(keyinput106), 
        .A(n7722), .ZN(n7730) );
  AOI22_X1 U9489 ( .A1(n7725), .A2(keyinput122), .B1(keyinput89), .B2(n7724), 
        .ZN(n7723) );
  OAI221_X1 U9490 ( .B1(n7725), .B2(keyinput122), .C1(n7724), .C2(keyinput89), 
        .A(n7723), .ZN(n7729) );
  AOI22_X1 U9491 ( .A1(n6484), .A2(keyinput90), .B1(n7727), .B2(keyinput79), 
        .ZN(n7726) );
  OAI221_X1 U9492 ( .B1(n6484), .B2(keyinput90), .C1(n7727), .C2(keyinput79), 
        .A(n7726), .ZN(n7728) );
  NOR4_X1 U9493 ( .A1(n7731), .A2(n7730), .A3(n7729), .A4(n7728), .ZN(n7756)
         );
  AOI22_X1 U9494 ( .A1(n4838), .A2(keyinput4), .B1(n10256), .B2(keyinput39), 
        .ZN(n7732) );
  OAI221_X1 U9495 ( .B1(n4838), .B2(keyinput4), .C1(n10256), .C2(keyinput39), 
        .A(n7732), .ZN(n7743) );
  AOI22_X1 U9496 ( .A1(n7734), .A2(keyinput68), .B1(n8317), .B2(keyinput80), 
        .ZN(n7733) );
  OAI221_X1 U9497 ( .B1(n7734), .B2(keyinput68), .C1(n8317), .C2(keyinput80), 
        .A(n7733), .ZN(n7742) );
  INV_X1 U9498 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n7737) );
  AOI22_X1 U9499 ( .A1(n7737), .A2(keyinput43), .B1(n7736), .B2(keyinput88), 
        .ZN(n7735) );
  OAI221_X1 U9500 ( .B1(n7737), .B2(keyinput43), .C1(n7736), .C2(keyinput88), 
        .A(n7735), .ZN(n7741) );
  XNOR2_X1 U9501 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput42), .ZN(n7739) );
  XNOR2_X1 U9502 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput69), .ZN(n7738) );
  NAND2_X1 U9503 ( .A1(n7739), .A2(n7738), .ZN(n7740) );
  NOR4_X1 U9504 ( .A1(n7743), .A2(n7742), .A3(n7741), .A4(n7740), .ZN(n7755)
         );
  INV_X1 U9505 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8351) );
  AOI22_X1 U9506 ( .A1(n8351), .A2(keyinput29), .B1(n9437), .B2(keyinput66), 
        .ZN(n7744) );
  OAI221_X1 U9507 ( .B1(n8351), .B2(keyinput29), .C1(n9437), .C2(keyinput66), 
        .A(n7744), .ZN(n7748) );
  INV_X1 U9508 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10422) );
  XNOR2_X1 U9509 ( .A(n10422), .B(keyinput1), .ZN(n7747) );
  XNOR2_X1 U9510 ( .A(n7745), .B(keyinput64), .ZN(n7746) );
  OR3_X1 U9511 ( .A1(n7748), .A2(n7747), .A3(n7746), .ZN(n7753) );
  AOI22_X1 U9512 ( .A1(n9427), .A2(keyinput59), .B1(n4833), .B2(keyinput126), 
        .ZN(n7749) );
  OAI221_X1 U9513 ( .B1(n9427), .B2(keyinput59), .C1(n4833), .C2(keyinput126), 
        .A(n7749), .ZN(n7752) );
  AOI22_X1 U9514 ( .A1(n7382), .A2(keyinput0), .B1(n8490), .B2(keyinput96), 
        .ZN(n7750) );
  OAI221_X1 U9515 ( .B1(n7382), .B2(keyinput0), .C1(n8490), .C2(keyinput96), 
        .A(n7750), .ZN(n7751) );
  NOR3_X1 U9516 ( .A1(n7753), .A2(n7752), .A3(n7751), .ZN(n7754) );
  NAND4_X1 U9517 ( .A1(n7757), .A2(n7756), .A3(n7755), .A4(n7754), .ZN(n7806)
         );
  INV_X1 U9518 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n7760) );
  INV_X1 U9519 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7759) );
  AOI22_X1 U9520 ( .A1(n7760), .A2(keyinput36), .B1(keyinput93), .B2(n7759), 
        .ZN(n7758) );
  OAI221_X1 U9521 ( .B1(n7760), .B2(keyinput36), .C1(n7759), .C2(keyinput93), 
        .A(n7758), .ZN(n7768) );
  INV_X1 U9522 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10418) );
  AOI22_X1 U9523 ( .A1(n9901), .A2(keyinput84), .B1(n10418), .B2(keyinput60), 
        .ZN(n7761) );
  OAI221_X1 U9524 ( .B1(n9901), .B2(keyinput84), .C1(n10418), .C2(keyinput60), 
        .A(n7761), .ZN(n7767) );
  AOI22_X1 U9525 ( .A1(n8443), .A2(keyinput127), .B1(n7763), .B2(keyinput33), 
        .ZN(n7762) );
  OAI221_X1 U9526 ( .B1(n8443), .B2(keyinput127), .C1(n7763), .C2(keyinput33), 
        .A(n7762), .ZN(n7766) );
  AOI22_X1 U9527 ( .A1(n10199), .A2(keyinput19), .B1(keyinput111), .B2(n9462), 
        .ZN(n7764) );
  OAI221_X1 U9528 ( .B1(n10199), .B2(keyinput19), .C1(n9462), .C2(keyinput111), 
        .A(n7764), .ZN(n7765) );
  NOR4_X1 U9529 ( .A1(n7768), .A2(n7767), .A3(n7766), .A4(n7765), .ZN(n7804)
         );
  INV_X1 U9530 ( .A(keyinput98), .ZN(n7770) );
  XOR2_X1 U9531 ( .A(n6142), .B(keyinput107), .Z(n7769) );
  OAI21_X1 U9532 ( .B1(P2_IR_REG_23__SCAN_IN), .B2(n7770), .A(n7769), .ZN(
        n7779) );
  AOI22_X1 U9533 ( .A1(n10134), .A2(keyinput78), .B1(n7772), .B2(keyinput123), 
        .ZN(n7771) );
  OAI221_X1 U9534 ( .B1(n10134), .B2(keyinput78), .C1(n7772), .C2(keyinput123), 
        .A(n7771), .ZN(n7778) );
  AOI22_X1 U9535 ( .A1(n10263), .A2(keyinput124), .B1(n9513), .B2(keyinput91), 
        .ZN(n7773) );
  OAI221_X1 U9536 ( .B1(n10263), .B2(keyinput124), .C1(n9513), .C2(keyinput91), 
        .A(n7773), .ZN(n7777) );
  INV_X1 U9537 ( .A(P2_WR_REG_SCAN_IN), .ZN(n7775) );
  AOI22_X1 U9538 ( .A1(n7775), .A2(keyinput18), .B1(n6102), .B2(keyinput40), 
        .ZN(n7774) );
  OAI221_X1 U9539 ( .B1(n7775), .B2(keyinput18), .C1(n6102), .C2(keyinput40), 
        .A(n7774), .ZN(n7776) );
  NOR4_X1 U9540 ( .A1(n7779), .A2(n7778), .A3(n7777), .A4(n7776), .ZN(n7803)
         );
  XNOR2_X1 U9541 ( .A(P2_D_REG_23__SCAN_IN), .B(keyinput109), .ZN(n7783) );
  XNOR2_X1 U9542 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(keyinput62), .ZN(n7782) );
  XNOR2_X1 U9543 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput23), .ZN(n7781) );
  XNOR2_X1 U9544 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput61), .ZN(n7780) );
  NAND4_X1 U9545 ( .A1(n7783), .A2(n7782), .A3(n7781), .A4(n7780), .ZN(n7790)
         );
  AOI22_X1 U9546 ( .A1(n6367), .A2(keyinput85), .B1(keyinput17), .B2(n7785), 
        .ZN(n7784) );
  OAI221_X1 U9547 ( .B1(n6367), .B2(keyinput85), .C1(n7785), .C2(keyinput17), 
        .A(n7784), .ZN(n7789) );
  INV_X1 U9548 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8354) );
  AOI22_X1 U9549 ( .A1(n7787), .A2(keyinput15), .B1(keyinput65), .B2(n8354), 
        .ZN(n7786) );
  OAI221_X1 U9550 ( .B1(n7787), .B2(keyinput15), .C1(n8354), .C2(keyinput65), 
        .A(n7786), .ZN(n7788) );
  NOR3_X1 U9551 ( .A1(n7790), .A2(n7789), .A3(n7788), .ZN(n7802) );
  AOI22_X1 U9552 ( .A1(n6112), .A2(keyinput56), .B1(keyinput3), .B2(n5371), 
        .ZN(n7791) );
  OAI221_X1 U9553 ( .B1(n6112), .B2(keyinput56), .C1(n5371), .C2(keyinput3), 
        .A(n7791), .ZN(n7800) );
  AOI22_X1 U9554 ( .A1(n6377), .A2(keyinput12), .B1(keyinput99), .B2(n7793), 
        .ZN(n7792) );
  OAI221_X1 U9555 ( .B1(n6377), .B2(keyinput12), .C1(n7793), .C2(keyinput99), 
        .A(n7792), .ZN(n7799) );
  INV_X1 U9556 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10421) );
  AOI22_X1 U9557 ( .A1(n8212), .A2(keyinput10), .B1(n10421), .B2(keyinput100), 
        .ZN(n7794) );
  OAI221_X1 U9558 ( .B1(n8212), .B2(keyinput10), .C1(n10421), .C2(keyinput100), 
        .A(n7794), .ZN(n7798) );
  AOI22_X1 U9559 ( .A1(n7796), .A2(keyinput87), .B1(keyinput108), .B2(n10179), 
        .ZN(n7795) );
  OAI221_X1 U9560 ( .B1(n7796), .B2(keyinput87), .C1(n10179), .C2(keyinput108), 
        .A(n7795), .ZN(n7797) );
  NOR4_X1 U9561 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n7797), .ZN(n7801)
         );
  NAND4_X1 U9562 ( .A1(n7804), .A2(n7803), .A3(n7802), .A4(n7801), .ZN(n7805)
         );
  NOR4_X1 U9563 ( .A1(n7808), .A2(n7807), .A3(n7806), .A4(n7805), .ZN(n7809)
         );
  OAI21_X1 U9564 ( .B1(keyinput98), .B2(n7810), .A(n7809), .ZN(n7811) );
  XNOR2_X1 U9565 ( .A(n7812), .B(n7811), .ZN(P1_U3575) );
  OAI21_X1 U9566 ( .B1(n10541), .B2(n10562), .A(n7975), .ZN(n7813) );
  NAND2_X1 U9567 ( .A1(n9380), .A2(n4404), .ZN(n7976) );
  OAI211_X1 U9568 ( .C1(n7814), .C2(n10565), .A(n7813), .B(n7976), .ZN(n9447)
         );
  NAND2_X1 U9569 ( .A1(n9447), .A2(n10571), .ZN(n7815) );
  OAI21_X1 U9570 ( .B1(n5371), .B2(n10571), .A(n7815), .ZN(P2_U3390) );
  NAND2_X1 U9571 ( .A1(n9738), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7816) );
  OAI21_X1 U9572 ( .B1(n9663), .B2(n9738), .A(n7816), .ZN(P1_U3577) );
  AOI21_X1 U9573 ( .B1(n7818), .B2(n7817), .A(n8786), .ZN(n7820) );
  NAND2_X1 U9574 ( .A1(n7820), .A2(n7819), .ZN(n7824) );
  INV_X1 U9575 ( .A(n7110), .ZN(n8141) );
  OAI22_X1 U9576 ( .A1(n8800), .A2(n10555), .B1(n8141), .B2(n8795), .ZN(n7821)
         );
  AOI211_X1 U9577 ( .C1(n8793), .C2(n7057), .A(n7822), .B(n7821), .ZN(n7823)
         );
  OAI211_X1 U9578 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8748), .A(n7824), .B(
        n7823), .ZN(P2_U3158) );
  INV_X1 U9579 ( .A(n7825), .ZN(n7875) );
  AOI22_X1 U9580 ( .A1(n10243), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n8151), .ZN(n7826) );
  OAI21_X1 U9581 ( .B1(n7875), .B2(n8271), .A(n7826), .ZN(P1_U3341) );
  NAND2_X1 U9582 ( .A1(n9036), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7827) );
  OAI21_X1 U9583 ( .B1(n9317), .B2(n9036), .A(n7827), .ZN(P2_U3512) );
  MUX2_X1 U9584 ( .A(n7828), .B(n9754), .S(n10230), .Z(n7832) );
  AOI21_X1 U9585 ( .B1(n10230), .B2(n7829), .A(n6115), .ZN(n10229) );
  OAI21_X1 U9586 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n10229), .A(P1_U3973), .ZN(
        n7830) );
  AOI21_X1 U9587 ( .B1(n7832), .B2(n7831), .A(n7830), .ZN(n7859) );
  OAI211_X1 U9588 ( .C1(n7835), .C2(n7834), .A(n10284), .B(n7833), .ZN(n7844)
         );
  OAI211_X1 U9589 ( .C1(n7838), .C2(n7837), .A(n10293), .B(n7836), .ZN(n7843)
         );
  AOI22_X1 U9590 ( .A1(n10233), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n7842) );
  INV_X1 U9591 ( .A(n7839), .ZN(n7840) );
  NAND2_X1 U9592 ( .A1(n10305), .A2(n7840), .ZN(n7841) );
  NAND4_X1 U9593 ( .A1(n7844), .A2(n7843), .A3(n7842), .A4(n7841), .ZN(n7845)
         );
  OR2_X1 U9594 ( .A1(n7859), .A2(n7845), .ZN(P1_U3245) );
  NAND2_X1 U9595 ( .A1(n9305), .A2(P2_U3893), .ZN(n7846) );
  OAI21_X1 U9596 ( .B1(P2_U3893), .B2(n8317), .A(n7846), .ZN(P2_U3511) );
  INV_X1 U9597 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7851) );
  OAI211_X1 U9598 ( .C1(n7849), .C2(n7848), .A(n10284), .B(n7847), .ZN(n7850)
         );
  NAND2_X1 U9599 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n8002) );
  OAI211_X1 U9600 ( .C1(n10308), .C2(n7851), .A(n7850), .B(n8002), .ZN(n7858)
         );
  OAI211_X1 U9601 ( .C1(n7854), .C2(n7853), .A(n10293), .B(n7852), .ZN(n7855)
         );
  OAI21_X1 U9602 ( .B1(n9868), .B2(n7856), .A(n7855), .ZN(n7857) );
  OR3_X1 U9603 ( .A1(n7859), .A2(n7858), .A3(n7857), .ZN(P1_U3247) );
  XNOR2_X1 U9604 ( .A(n7860), .B(n8245), .ZN(n7874) );
  OAI21_X1 U9605 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7861), .A(n7927), .ZN(
        n7872) );
  INV_X1 U9606 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7864) );
  AND2_X1 U9607 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8207) );
  AOI21_X1 U9608 ( .B1(n9209), .B2(n7862), .A(n8207), .ZN(n7863) );
  OAI21_X1 U9609 ( .B1(n9171), .B2(n7864), .A(n7863), .ZN(n7871) );
  INV_X1 U9610 ( .A(n7865), .ZN(n7866) );
  NAND3_X1 U9611 ( .A1(n7868), .A2(n7867), .A3(n7866), .ZN(n7869) );
  AOI21_X1 U9612 ( .B1(n7933), .B2(n7869), .A(n9159), .ZN(n7870) );
  AOI211_X1 U9613 ( .C1(n7872), .C2(n9146), .A(n7871), .B(n7870), .ZN(n7873)
         );
  OAI21_X1 U9614 ( .B1(n7874), .B2(n9213), .A(n7873), .ZN(P2_U3189) );
  INV_X1 U9615 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7876) );
  INV_X1 U9616 ( .A(n9102), .ZN(n9094) );
  OAI222_X1 U9617 ( .A1(n9537), .A2(n7876), .B1(n9547), .B2(n7875), .C1(
        P2_U3151), .C2(n9094), .ZN(P2_U3281) );
  MUX2_X1 U9618 ( .A(n6060), .B(P1_REG1_REG_12__SCAN_IN), .S(n8044), .Z(n7882)
         );
  NAND2_X1 U9619 ( .A1(n7884), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7877) );
  NAND2_X1 U9620 ( .A1(n7878), .A2(n7877), .ZN(n9833) );
  MUX2_X1 U9621 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6211), .S(n9840), .Z(n9832)
         );
  NAND2_X1 U9622 ( .A1(n9833), .A2(n9832), .ZN(n9831) );
  NAND2_X1 U9623 ( .A1(n9840), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7879) );
  NAND2_X1 U9624 ( .A1(n9831), .A2(n7879), .ZN(n7881) );
  INV_X1 U9625 ( .A(n8040), .ZN(n7880) );
  AOI21_X1 U9626 ( .B1(n7882), .B2(n7881), .A(n7880), .ZN(n7895) );
  INV_X1 U9627 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7883) );
  NAND2_X1 U9628 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8497) );
  OAI21_X1 U9629 ( .B1(n10308), .B2(n7883), .A(n8497), .ZN(n7893) );
  NAND2_X1 U9630 ( .A1(n7884), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7885) );
  XNOR2_X1 U9631 ( .A(n9840), .B(n7887), .ZN(n9835) );
  NAND2_X1 U9632 ( .A1(n9836), .A2(n9835), .ZN(n9834) );
  NAND2_X1 U9633 ( .A1(n9840), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7888) );
  NAND2_X1 U9634 ( .A1(n9834), .A2(n7888), .ZN(n7890) );
  XNOR2_X1 U9635 ( .A(n8044), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U9636 ( .A1(n7890), .A2(n7889), .ZN(n7891) );
  AOI21_X1 U9637 ( .B1(n8046), .B2(n7891), .A(n10269), .ZN(n7892) );
  AOI211_X1 U9638 ( .C1(n10305), .C2(n8044), .A(n7893), .B(n7892), .ZN(n7894)
         );
  OAI21_X1 U9639 ( .B1(n7895), .B2(n10299), .A(n7894), .ZN(P1_U3255) );
  OAI21_X1 U9640 ( .B1(n8867), .B2(n7896), .A(n7897), .ZN(n8086) );
  INV_X1 U9641 ( .A(n7529), .ZN(n7902) );
  INV_X1 U9642 ( .A(n10541), .ZN(n9356) );
  NAND3_X1 U9643 ( .A1(n7896), .A2(n7982), .A3(n7529), .ZN(n7898) );
  AND2_X1 U9644 ( .A1(n7899), .A2(n7898), .ZN(n7900) );
  OAI222_X1 U9645 ( .A1(n10537), .A2(n7902), .B1(n10539), .B2(n7901), .C1(
        n9356), .C2(n7900), .ZN(n8083) );
  AOI21_X1 U9646 ( .B1(n10562), .B2(n8086), .A(n8083), .ZN(n7907) );
  OAI22_X1 U9647 ( .A1(n9424), .A2(n8868), .B1(n10578), .B2(n5362), .ZN(n7903)
         );
  INV_X1 U9648 ( .A(n7903), .ZN(n7904) );
  OAI21_X1 U9649 ( .B1(n7907), .B2(n7168), .A(n7904), .ZN(P2_U3460) );
  OAI22_X1 U9650 ( .A1(n8868), .A2(n9500), .B1(n10571), .B2(n5353), .ZN(n7905)
         );
  INV_X1 U9651 ( .A(n7905), .ZN(n7906) );
  OAI21_X1 U9652 ( .B1(n7907), .B2(n10573), .A(n7906), .ZN(P2_U3393) );
  INV_X1 U9653 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7909) );
  INV_X1 U9654 ( .A(n7908), .ZN(n7910) );
  OAI222_X1 U9655 ( .A1(n9537), .A2(n7909), .B1(n9547), .B2(n7910), .C1(
        P2_U3151), .C2(n5173), .ZN(P2_U3280) );
  INV_X1 U9656 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7911) );
  INV_X1 U9657 ( .A(n10260), .ZN(n9858) );
  OAI222_X1 U9658 ( .A1(n10224), .A2(n7911), .B1(n8271), .B2(n7910), .C1(
        P1_U3086), .C2(n9858), .ZN(P1_U3340) );
  INV_X1 U9659 ( .A(n6526), .ZN(n10433) );
  INV_X1 U9660 ( .A(n7555), .ZN(n7915) );
  INV_X1 U9661 ( .A(n7912), .ZN(n7913) );
  NOR3_X1 U9662 ( .A1(n7915), .A2(n7914), .A3(n7913), .ZN(n7916) );
  OAI21_X1 U9663 ( .B1(n7916), .B2(n4527), .A(n9716), .ZN(n7921) );
  OR2_X1 U9664 ( .A1(n7999), .A2(n9703), .ZN(n7918) );
  NAND2_X1 U9665 ( .A1(n9687), .A2(n6511), .ZN(n7917) );
  NAND2_X1 U9666 ( .A1(n7918), .A2(n7917), .ZN(n10398) );
  AOI22_X1 U9667 ( .A1(n9710), .A2(n10398), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n7919), .ZN(n7920) );
  OAI211_X1 U9668 ( .C1(n10433), .C2(n9725), .A(n7921), .B(n7920), .ZN(
        P1_U3237) );
  XOR2_X1 U9669 ( .A(n7922), .B(n7923), .Z(n7942) );
  INV_X1 U9670 ( .A(n7924), .ZN(n7929) );
  NAND3_X1 U9671 ( .A1(n7927), .A2(n7926), .A3(n7925), .ZN(n7928) );
  AOI21_X1 U9672 ( .B1(n7929), .B2(n7928), .A(n9217), .ZN(n7940) );
  INV_X1 U9673 ( .A(n7930), .ZN(n7931) );
  NAND3_X1 U9674 ( .A1(n7933), .A2(n7932), .A3(n7931), .ZN(n7934) );
  AOI21_X1 U9675 ( .B1(n8013), .B2(n7934), .A(n9159), .ZN(n7939) );
  INV_X1 U9676 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U9677 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8261) );
  NAND2_X1 U9678 ( .A1(n9209), .A2(n7935), .ZN(n7936) );
  OAI211_X1 U9679 ( .C1(n9171), .C2(n7937), .A(n8261), .B(n7936), .ZN(n7938)
         );
  NOR3_X1 U9680 ( .A1(n7940), .A2(n7939), .A3(n7938), .ZN(n7941) );
  OAI21_X1 U9681 ( .B1(n7942), .B2(n9213), .A(n7941), .ZN(P2_U3190) );
  OAI21_X1 U9682 ( .B1(n7945), .B2(n7944), .A(n7943), .ZN(n7946) );
  NAND2_X1 U9683 ( .A1(n7946), .A2(n8790), .ZN(n7951) );
  OAI22_X1 U9684 ( .A1(n8800), .A2(n10560), .B1(n7947), .B2(n8795), .ZN(n7948)
         );
  AOI211_X1 U9685 ( .C1(n8793), .C2(n9035), .A(n7949), .B(n7948), .ZN(n7950)
         );
  OAI211_X1 U9686 ( .C1(n8031), .C2(n8748), .A(n7951), .B(n7950), .ZN(P2_U3170) );
  AOI21_X1 U9687 ( .B1(n7953), .B2(n4750), .A(n10407), .ZN(n7954) );
  NAND2_X1 U9688 ( .A1(n7954), .A2(n10408), .ZN(n10427) );
  INV_X1 U9689 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7955) );
  OAI22_X1 U9690 ( .A1(n10411), .A2(n10427), .B1(n7955), .B2(n10382), .ZN(
        n7956) );
  AOI21_X1 U9691 ( .B1(n10332), .B2(n4750), .A(n7956), .ZN(n7968) );
  INV_X1 U9692 ( .A(n8090), .ZN(n8299) );
  XNOR2_X1 U9693 ( .A(n7957), .B(n7959), .ZN(n10426) );
  INV_X1 U9694 ( .A(n8297), .ZN(n10496) );
  NAND2_X1 U9695 ( .A1(n10426), .A2(n10496), .ZN(n7965) );
  NAND2_X1 U9696 ( .A1(n7959), .A2(n7958), .ZN(n7960) );
  NAND2_X1 U9697 ( .A1(n7961), .A2(n7960), .ZN(n7963) );
  AOI21_X1 U9698 ( .B1(n7963), .B2(n10399), .A(n7962), .ZN(n7964) );
  NAND2_X1 U9699 ( .A1(n7965), .A2(n7964), .ZN(n10431) );
  AOI21_X1 U9700 ( .B1(n8299), .B2(n10426), .A(n10431), .ZN(n7966) );
  MUX2_X1 U9701 ( .A(n7610), .B(n7966), .S(n10324), .Z(n7967) );
  NAND2_X1 U9702 ( .A1(n7968), .A2(n7967), .ZN(P1_U3292) );
  NAND2_X1 U9703 ( .A1(n7973), .A2(n7969), .ZN(n7970) );
  OAI211_X1 U9704 ( .C1(n7973), .C2(n7972), .A(n7971), .B(n7970), .ZN(n7979)
         );
  INV_X1 U9705 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7978) );
  NAND3_X1 U9706 ( .A1(n7975), .A2(n10565), .A3(n7974), .ZN(n7977) );
  OAI211_X1 U9707 ( .C1(n7978), .C2(n10533), .A(n7977), .B(n7976), .ZN(n7980)
         );
  MUX2_X1 U9708 ( .A(n7980), .B(P2_REG2_REG_0__SCAN_IN), .S(n10550), .Z(n7981)
         );
  AOI21_X1 U9709 ( .B1(n4398), .B2(n7982), .A(n7981), .ZN(n7983) );
  INV_X1 U9710 ( .A(n7983), .ZN(P2_U3233) );
  NAND2_X1 U9711 ( .A1(n9738), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7984) );
  OAI21_X1 U9712 ( .B1(n9604), .B2(n9738), .A(n7984), .ZN(P1_U3578) );
  INV_X1 U9713 ( .A(n7985), .ZN(n8036) );
  AOI22_X1 U9714 ( .A1(n10274), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n8151), .ZN(n7986) );
  OAI21_X1 U9715 ( .B1(n8036), .B2(n8271), .A(n7986), .ZN(P1_U3339) );
  XNOR2_X1 U9716 ( .A(n7988), .B(n7987), .ZN(n7989) );
  NAND2_X1 U9717 ( .A1(n7989), .A2(n8790), .ZN(n7994) );
  OAI22_X1 U9718 ( .A1(n8800), .A2(n10566), .B1(n7990), .B2(n8795), .ZN(n7991)
         );
  AOI211_X1 U9719 ( .C1(n8793), .C2(n7110), .A(n7992), .B(n7991), .ZN(n7993)
         );
  OAI211_X1 U9720 ( .C1(n8145), .C2(n8748), .A(n7994), .B(n7993), .ZN(P2_U3167) );
  AND2_X1 U9721 ( .A1(n9569), .A2(n7995), .ZN(n7998) );
  OAI211_X1 U9722 ( .C1(n7998), .C2(n7997), .A(n9716), .B(n7996), .ZN(n8006)
         );
  OR2_X1 U9723 ( .A1(n7999), .A2(n9701), .ZN(n8001) );
  OR2_X1 U9724 ( .A1(n8181), .A2(n9703), .ZN(n8000) );
  AND2_X1 U9725 ( .A1(n8001), .A2(n8000), .ZN(n10378) );
  OAI21_X1 U9726 ( .B1(n9719), .B2(n10378), .A(n8002), .ZN(n8003) );
  AOI21_X1 U9727 ( .B1(n9693), .B2(n8004), .A(n8003), .ZN(n8005) );
  OAI211_X1 U9728 ( .C1(n9708), .C2(n10381), .A(n8006), .B(n8005), .ZN(
        P1_U3230) );
  XNOR2_X1 U9729 ( .A(n8007), .B(n8348), .ZN(n8023) );
  OAI21_X1 U9730 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n8009), .A(n8008), .ZN(
        n8021) );
  INV_X1 U9731 ( .A(n8010), .ZN(n8011) );
  NAND3_X1 U9732 ( .A1(n8013), .A2(n8012), .A3(n8011), .ZN(n8014) );
  AOI21_X1 U9733 ( .B1(n8117), .B2(n8014), .A(n9159), .ZN(n8020) );
  INV_X1 U9734 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U9735 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8342) );
  INV_X1 U9736 ( .A(n8342), .ZN(n8015) );
  AOI21_X1 U9737 ( .B1(n9209), .B2(n8016), .A(n8015), .ZN(n8017) );
  OAI21_X1 U9738 ( .B1(n9171), .B2(n8018), .A(n8017), .ZN(n8019) );
  AOI211_X1 U9739 ( .C1(n8021), .C2(n9146), .A(n8020), .B(n8019), .ZN(n8022)
         );
  OAI21_X1 U9740 ( .B1(n8023), .B2(n9213), .A(n8022), .ZN(P2_U3191) );
  AND2_X1 U9741 ( .A1(n8024), .A2(n5967), .ZN(n10547) );
  INV_X1 U9742 ( .A(n10547), .ZN(n8222) );
  NAND2_X1 U9743 ( .A1(n10544), .A2(n8222), .ZN(n8025) );
  INV_X1 U9744 ( .A(n8889), .ZN(n8875) );
  NAND2_X1 U9745 ( .A1(n8026), .A2(n8816), .ZN(n8073) );
  NAND2_X1 U9746 ( .A1(n8073), .A2(n8890), .ZN(n8134) );
  NAND2_X1 U9747 ( .A1(n8886), .A2(n8132), .ZN(n8028) );
  INV_X1 U9748 ( .A(n8028), .ZN(n8882) );
  XNOR2_X1 U9749 ( .A(n8134), .B(n8882), .ZN(n10563) );
  INV_X1 U9750 ( .A(n10563), .ZN(n8035) );
  XNOR2_X1 U9751 ( .A(n8027), .B(n8028), .ZN(n8029) );
  AOI222_X1 U9752 ( .A1(n10541), .A2(n8029), .B1(n9035), .B2(n9382), .C1(n9034), .C2(n9380), .ZN(n10559) );
  MUX2_X1 U9753 ( .A(n8030), .B(n10559), .S(n9385), .Z(n8034) );
  INV_X1 U9754 ( .A(n8031), .ZN(n8032) );
  AOI22_X1 U9755 ( .A1(n4398), .A2(n4764), .B1(n9388), .B2(n8032), .ZN(n8033)
         );
  OAI211_X1 U9756 ( .C1(n9366), .C2(n8035), .A(n8034), .B(n8033), .ZN(P2_U3229) );
  INV_X1 U9757 ( .A(n9148), .ZN(n9142) );
  OAI222_X1 U9758 ( .A1(n9537), .A2(n8037), .B1(P2_U3151), .B2(n9142), .C1(
        n8036), .C2(n9547), .ZN(P2_U3279) );
  MUX2_X1 U9759 ( .A(n8038), .B(P1_REG1_REG_13__SCAN_IN), .S(n9853), .Z(n8043)
         );
  OR2_X1 U9760 ( .A1(n8044), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8039) );
  INV_X1 U9761 ( .A(n9845), .ZN(n8041) );
  AOI211_X1 U9762 ( .C1(n8043), .C2(n8042), .A(n10299), .B(n8041), .ZN(n8053)
         );
  XNOR2_X1 U9763 ( .A(n9853), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n8049) );
  OR2_X1 U9764 ( .A1(n8044), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8045) );
  INV_X1 U9765 ( .A(n9855), .ZN(n8047) );
  AOI211_X1 U9766 ( .C1(n8049), .C2(n8048), .A(n10269), .B(n8047), .ZN(n8052)
         );
  NAND2_X1 U9767 ( .A1(n10305), .A2(n9853), .ZN(n8050) );
  NAND2_X1 U9768 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8586) );
  OAI211_X1 U9769 ( .C1(n10308), .C2(n8355), .A(n8050), .B(n8586), .ZN(n8051)
         );
  OR3_X1 U9770 ( .A1(n8053), .A2(n8052), .A3(n8051), .ZN(P1_U3256) );
  AOI21_X1 U9771 ( .B1(n8054), .B2(n8055), .A(n8786), .ZN(n8057) );
  NAND2_X1 U9772 ( .A1(n8057), .A2(n8056), .ZN(n8063) );
  OAI22_X1 U9773 ( .A1(n8800), .A2(n8059), .B1(n8058), .B2(n8795), .ZN(n8060)
         );
  AOI211_X1 U9774 ( .C1(n8793), .C2(n9034), .A(n8061), .B(n8060), .ZN(n8062)
         );
  OAI211_X1 U9775 ( .C1(n8068), .C2(n8748), .A(n8063), .B(n8062), .ZN(P2_U3179) );
  XNOR2_X1 U9776 ( .A(n8064), .B(n8814), .ZN(n9444) );
  INV_X1 U9777 ( .A(n9444), .ZN(n8072) );
  XNOR2_X1 U9778 ( .A(n8065), .B(n8814), .ZN(n8066) );
  AOI222_X1 U9779 ( .A1(n10541), .A2(n8066), .B1(n9033), .B2(n9380), .C1(n9034), .C2(n9382), .ZN(n9446) );
  MUX2_X1 U9780 ( .A(n8067), .B(n9446), .S(n9385), .Z(n8071) );
  INV_X1 U9781 ( .A(n8068), .ZN(n8069) );
  AOI22_X1 U9782 ( .A1(n4398), .A2(n9442), .B1(n9388), .B2(n8069), .ZN(n8070)
         );
  OAI211_X1 U9783 ( .C1(n9366), .C2(n8072), .A(n8071), .B(n8070), .ZN(P2_U3227) );
  INV_X1 U9784 ( .A(n9366), .ZN(n9295) );
  OAI21_X1 U9785 ( .B1(n8026), .B2(n8816), .A(n8073), .ZN(n10558) );
  INV_X1 U9786 ( .A(n4398), .ZN(n9362) );
  OAI22_X1 U9787 ( .A1(n9362), .A2(n10555), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10533), .ZN(n8080) );
  INV_X1 U9788 ( .A(n8816), .ZN(n8074) );
  XNOR2_X1 U9789 ( .A(n8075), .B(n8074), .ZN(n8076) );
  NAND2_X1 U9790 ( .A1(n8076), .A2(n10541), .ZN(n8078) );
  AOI22_X1 U9791 ( .A1(n9382), .A2(n7057), .B1(n7110), .B2(n9380), .ZN(n8077)
         );
  NAND2_X1 U9792 ( .A1(n8078), .A2(n8077), .ZN(n10556) );
  MUX2_X1 U9793 ( .A(n10556), .B(P2_REG2_REG_3__SCAN_IN), .S(n10550), .Z(n8079) );
  AOI211_X1 U9794 ( .C1(n9295), .C2(n10558), .A(n8080), .B(n8079), .ZN(n8081)
         );
  INV_X1 U9795 ( .A(n8081), .ZN(P2_U3230) );
  INV_X1 U9796 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8082) );
  OAI22_X1 U9797 ( .A1(n9362), .A2(n8868), .B1(n8082), .B2(n10533), .ZN(n8085)
         );
  MUX2_X1 U9798 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n8083), .S(n9385), .Z(n8084)
         );
  AOI211_X1 U9799 ( .C1(n9295), .C2(n8086), .A(n8085), .B(n8084), .ZN(n8087)
         );
  INV_X1 U9800 ( .A(n8087), .ZN(P2_U3232) );
  XOR2_X1 U9801 ( .A(n8088), .B(n8093), .Z(n8089) );
  OAI22_X1 U9802 ( .A1(n9750), .A2(n9701), .B1(n8293), .B2(n9703), .ZN(n8157)
         );
  AOI21_X1 U9803 ( .B1(n8089), .B2(n10399), .A(n8157), .ZN(n10454) );
  AND2_X1 U9804 ( .A1(n8297), .A2(n8090), .ZN(n8091) );
  XNOR2_X1 U9805 ( .A(n8092), .B(n8093), .ZN(n10457) );
  INV_X1 U9806 ( .A(n8094), .ZN(n10453) );
  INV_X2 U9807 ( .A(n10332), .ZN(n10385) );
  AOI211_X1 U9808 ( .C1(n8094), .C2(n10389), .A(n10407), .B(n4438), .ZN(n10451) );
  NAND2_X1 U9809 ( .A1(n10451), .A2(n10393), .ZN(n8096) );
  AOI22_X1 U9810 ( .A1(n10402), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n8160), .B2(
        n10401), .ZN(n8095) );
  OAI211_X1 U9811 ( .C1(n10453), .C2(n10385), .A(n8096), .B(n8095), .ZN(n8097)
         );
  AOI21_X1 U9812 ( .B1(n10394), .B2(n10457), .A(n8097), .ZN(n8098) );
  OAI21_X1 U9813 ( .B1(n10402), .B2(n10454), .A(n8098), .ZN(P1_U3288) );
  XNOR2_X1 U9814 ( .A(n8099), .B(n8103), .ZN(n8101) );
  OAI22_X1 U9815 ( .A1(n8100), .A2(n9701), .B1(n9750), .B2(n9703), .ZN(n9573)
         );
  AOI21_X1 U9816 ( .B1(n8101), .B2(n10399), .A(n9573), .ZN(n10438) );
  XNOR2_X1 U9817 ( .A(n8102), .B(n8103), .ZN(n10444) );
  INV_X1 U9818 ( .A(n6539), .ZN(n10441) );
  AOI211_X1 U9819 ( .C1(n6539), .C2(n10409), .A(n10407), .B(n10391), .ZN(
        n10439) );
  NAND2_X1 U9820 ( .A1(n10439), .A2(n10393), .ZN(n8106) );
  INV_X1 U9821 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8104) );
  AOI22_X1 U9822 ( .A1(n10402), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10401), .B2(
        n8104), .ZN(n8105) );
  OAI211_X1 U9823 ( .C1(n10441), .C2(n10385), .A(n8106), .B(n8105), .ZN(n8107)
         );
  AOI21_X1 U9824 ( .B1(n10394), .B2(n10444), .A(n8107), .ZN(n8108) );
  OAI21_X1 U9825 ( .B1(n10402), .B2(n10438), .A(n8108), .ZN(P1_U3290) );
  XOR2_X1 U9826 ( .A(n8109), .B(n8110), .Z(n8126) );
  NAND2_X1 U9827 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8480) );
  OAI21_X1 U9828 ( .B1(n9154), .B2(n8111), .A(n8480), .ZN(n8116) );
  NAND3_X1 U9829 ( .A1(n8008), .A2(n8113), .A3(n4418), .ZN(n8114) );
  AOI21_X1 U9830 ( .B1(n4762), .B2(n8114), .A(n9217), .ZN(n8115) );
  AOI211_X1 U9831 ( .C1(n9210), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n8116), .B(
        n8115), .ZN(n8125) );
  INV_X1 U9832 ( .A(n8117), .ZN(n8121) );
  INV_X1 U9833 ( .A(n8118), .ZN(n8120) );
  NOR3_X1 U9834 ( .A1(n8121), .A2(n8120), .A3(n8119), .ZN(n8123) );
  INV_X1 U9835 ( .A(n8234), .ZN(n8122) );
  OAI21_X1 U9836 ( .B1(n8123), .B2(n8122), .A(n9215), .ZN(n8124) );
  OAI211_X1 U9837 ( .C1(n8126), .C2(n9213), .A(n8125), .B(n8124), .ZN(P2_U3192) );
  INV_X1 U9838 ( .A(n8127), .ZN(n8130) );
  INV_X1 U9839 ( .A(n10286), .ZN(n8128) );
  OAI222_X1 U9840 ( .A1(n10224), .A2(n8129), .B1(n8271), .B2(n8130), .C1(
        P1_U3086), .C2(n8128), .ZN(P1_U3338) );
  OAI222_X1 U9841 ( .A1(n9537), .A2(n8131), .B1(n9547), .B2(n8130), .C1(
        P2_U3151), .C2(n5166), .ZN(P2_U3278) );
  INV_X1 U9842 ( .A(n8886), .ZN(n8133) );
  OAI21_X1 U9843 ( .B1(n8134), .B2(n8133), .A(n8132), .ZN(n8137) );
  NAND2_X1 U9844 ( .A1(n9034), .A2(n8147), .ZN(n8135) );
  NAND2_X1 U9845 ( .A1(n8136), .A2(n8135), .ZN(n8812) );
  XNOR2_X1 U9846 ( .A(n8137), .B(n8812), .ZN(n10568) );
  INV_X1 U9847 ( .A(n8027), .ZN(n8139) );
  OAI21_X1 U9848 ( .B1(n8139), .B2(n7110), .A(n4764), .ZN(n8140) );
  OAI21_X1 U9849 ( .B1(n8141), .B2(n8027), .A(n8140), .ZN(n8142) );
  XNOR2_X1 U9850 ( .A(n8142), .B(n8812), .ZN(n8143) );
  AOI222_X1 U9851 ( .A1(n10541), .A2(n8143), .B1(n7111), .B2(n9380), .C1(n7110), .C2(n9382), .ZN(n10564) );
  MUX2_X1 U9852 ( .A(n8144), .B(n10564), .S(n9385), .Z(n8149) );
  INV_X1 U9853 ( .A(n8145), .ZN(n8146) );
  AOI22_X1 U9854 ( .A1(n4398), .A2(n8147), .B1(n9388), .B2(n8146), .ZN(n8148)
         );
  OAI211_X1 U9855 ( .C1(n9366), .C2(n10568), .A(n8149), .B(n8148), .ZN(
        P2_U3228) );
  INV_X1 U9856 ( .A(n8150), .ZN(n8210) );
  AOI22_X1 U9857 ( .A1(n10304), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n8151), .ZN(n8152) );
  OAI21_X1 U9858 ( .B1(n8210), .B2(n8271), .A(n8152), .ZN(P1_U3337) );
  NAND2_X1 U9859 ( .A1(n8153), .A2(n8154), .ZN(n8155) );
  XOR2_X1 U9860 ( .A(n8156), .B(n8155), .Z(n8162) );
  AOI22_X1 U9861 ( .A1(n9710), .A2(n8157), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n8158) );
  OAI21_X1 U9862 ( .B1(n10453), .B2(n9725), .A(n8158), .ZN(n8159) );
  AOI21_X1 U9863 ( .B1(n8160), .B2(n9721), .A(n8159), .ZN(n8161) );
  OAI21_X1 U9864 ( .B1(n8162), .B2(n9695), .A(n8161), .ZN(P1_U3227) );
  NAND2_X1 U9865 ( .A1(n8163), .A2(n8164), .ZN(n8166) );
  INV_X1 U9866 ( .A(n8165), .ZN(n8821) );
  XNOR2_X1 U9867 ( .A(n8166), .B(n8821), .ZN(n8220) );
  NAND2_X1 U9868 ( .A1(n8193), .A2(n8168), .ZN(n8169) );
  NAND2_X1 U9869 ( .A1(n8169), .A2(n8821), .ZN(n8171) );
  NAND2_X1 U9870 ( .A1(n8193), .A2(n8170), .ZN(n8280) );
  NAND3_X1 U9871 ( .A1(n8171), .A2(n10541), .A3(n8280), .ZN(n8173) );
  AOI22_X1 U9872 ( .A1(n9382), .A2(n9033), .B1(n9031), .B2(n9380), .ZN(n8172)
         );
  AND2_X1 U9873 ( .A1(n8173), .A2(n8172), .ZN(n8216) );
  INV_X1 U9874 ( .A(n8216), .ZN(n8174) );
  NAND2_X1 U9875 ( .A1(n8174), .A2(n10571), .ZN(n8176) );
  AOI22_X1 U9876 ( .A1(n9520), .A2(n8266), .B1(P2_REG0_REG_8__SCAN_IN), .B2(
        n10573), .ZN(n8175) );
  OAI211_X1 U9877 ( .C1(n8220), .C2(n9524), .A(n8176), .B(n8175), .ZN(P2_U3414) );
  XNOR2_X1 U9878 ( .A(n8177), .B(n8178), .ZN(n10461) );
  INV_X1 U9879 ( .A(n10461), .ZN(n8190) );
  NOR2_X1 U9880 ( .A1(n8179), .A2(n8178), .ZN(n8290) );
  AND2_X1 U9881 ( .A1(n8179), .A2(n8178), .ZN(n8180) );
  OAI21_X1 U9882 ( .B1(n8290), .B2(n8180), .A(n10399), .ZN(n8184) );
  OR2_X1 U9883 ( .A1(n8181), .A2(n9701), .ZN(n8183) );
  OR2_X1 U9884 ( .A1(n8464), .A2(n9703), .ZN(n8182) );
  AND2_X1 U9885 ( .A1(n8183), .A2(n8182), .ZN(n8252) );
  NAND2_X1 U9886 ( .A1(n8184), .A2(n8252), .ZN(n10459) );
  OAI211_X1 U9887 ( .C1(n5079), .C2(n4438), .A(n5080), .B(n10390), .ZN(n10458)
         );
  NOR2_X1 U9888 ( .A1(n10458), .A2(n10411), .ZN(n8188) );
  INV_X1 U9889 ( .A(n8253), .ZN(n8185) );
  AOI22_X1 U9890 ( .A1(n10402), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n8185), .B2(
        n10401), .ZN(n8186) );
  OAI21_X1 U9891 ( .B1(n10385), .B2(n5079), .A(n8186), .ZN(n8187) );
  AOI211_X1 U9892 ( .C1(n10459), .C2(n10324), .A(n8188), .B(n8187), .ZN(n8189)
         );
  OAI21_X1 U9893 ( .B1(n8190), .B2(n10412), .A(n8189), .ZN(P1_U3287) );
  INV_X1 U9894 ( .A(n8191), .ZN(n10554) );
  OAI21_X1 U9895 ( .B1(n8192), .B2(n8901), .A(n8163), .ZN(n8223) );
  INV_X1 U9896 ( .A(n8223), .ZN(n8199) );
  AOI22_X1 U9897 ( .A1(n7111), .A2(n9382), .B1(n9380), .B2(n9032), .ZN(n8198)
         );
  INV_X1 U9898 ( .A(n8167), .ZN(n8195) );
  OAI21_X1 U9899 ( .B1(n8195), .B2(n8194), .A(n8193), .ZN(n8196) );
  NAND2_X1 U9900 ( .A1(n8196), .A2(n10541), .ZN(n8197) );
  OAI211_X1 U9901 ( .C1(n8223), .C2(n10544), .A(n8198), .B(n8197), .ZN(n8225)
         );
  AOI21_X1 U9902 ( .B1(n10554), .B2(n8199), .A(n8225), .ZN(n8244) );
  AOI22_X1 U9903 ( .A1(n9520), .A2(n8200), .B1(P2_REG0_REG_7__SCAN_IN), .B2(
        n10573), .ZN(n8201) );
  OAI21_X1 U9904 ( .B1(n8244), .B2(n10573), .A(n8201), .ZN(P2_U3411) );
  OAI21_X1 U9905 ( .B1(n8203), .B2(n4521), .A(n8202), .ZN(n8204) );
  NAND2_X1 U9906 ( .A1(n8204), .A2(n8790), .ZN(n8209) );
  OAI22_X1 U9907 ( .A1(n8800), .A2(n8247), .B1(n8205), .B2(n8795), .ZN(n8206)
         );
  AOI211_X1 U9908 ( .C1(n8793), .C2(n7111), .A(n8207), .B(n8206), .ZN(n8208)
         );
  OAI211_X1 U9909 ( .C1(n8221), .C2(n8748), .A(n8209), .B(n8208), .ZN(P2_U3153) );
  INV_X1 U9910 ( .A(n9187), .ZN(n9203) );
  OAI222_X1 U9911 ( .A1(n9537), .A2(n8211), .B1(n9203), .B2(P2_U3151), .C1(
        n9547), .C2(n8210), .ZN(P2_U3277) );
  MUX2_X1 U9912 ( .A(n8216), .B(n8212), .S(n10550), .Z(n8215) );
  INV_X1 U9913 ( .A(n8263), .ZN(n8213) );
  AOI22_X1 U9914 ( .A1(n4398), .A2(n8266), .B1(n9388), .B2(n8213), .ZN(n8214)
         );
  OAI211_X1 U9915 ( .C1(n8220), .C2(n9366), .A(n8215), .B(n8214), .ZN(P2_U3225) );
  MUX2_X1 U9916 ( .A(n8217), .B(n8216), .S(n10578), .Z(n8219) );
  NAND2_X1 U9917 ( .A1(n9438), .A2(n8266), .ZN(n8218) );
  OAI211_X1 U9918 ( .C1(n8220), .C2(n9441), .A(n8219), .B(n8218), .ZN(P2_U3467) );
  OAI22_X1 U9919 ( .A1(n8223), .A2(n8222), .B1(n8221), .B2(n10533), .ZN(n8224)
         );
  NOR2_X1 U9920 ( .A1(n8225), .A2(n8224), .ZN(n8226) );
  MUX2_X1 U9921 ( .A(n8227), .B(n8226), .S(n9385), .Z(n8228) );
  OAI21_X1 U9922 ( .B1(n8247), .B2(n9362), .A(n8228), .ZN(P2_U3226) );
  AOI21_X1 U9923 ( .B1(n8384), .B2(n8229), .A(n7192), .ZN(n8243) );
  NAND2_X1 U9924 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8534) );
  OAI21_X1 U9925 ( .B1(n9154), .B2(n8230), .A(n8534), .ZN(n8238) );
  INV_X1 U9926 ( .A(n8231), .ZN(n8232) );
  NAND3_X1 U9927 ( .A1(n8234), .A2(n8233), .A3(n8232), .ZN(n8235) );
  AOI21_X1 U9928 ( .B1(n8236), .B2(n8235), .A(n9159), .ZN(n8237) );
  AOI211_X1 U9929 ( .C1(n9210), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n8238), .B(
        n8237), .ZN(n8242) );
  XNOR2_X1 U9930 ( .A(n8239), .B(n8380), .ZN(n8240) );
  NAND2_X1 U9931 ( .A1(n8240), .A2(n9173), .ZN(n8241) );
  OAI211_X1 U9932 ( .C1(n8243), .C2(n9217), .A(n8242), .B(n8241), .ZN(P2_U3193) );
  MUX2_X1 U9933 ( .A(n8245), .B(n8244), .S(n10578), .Z(n8246) );
  OAI21_X1 U9934 ( .B1(n8247), .B2(n9424), .A(n8246), .ZN(P2_U3466) );
  INV_X1 U9935 ( .A(n8248), .ZN(n8249) );
  AOI21_X1 U9936 ( .B1(n8251), .B2(n8250), .A(n8249), .ZN(n8258) );
  NAND2_X1 U9937 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9791) );
  OAI21_X1 U9938 ( .B1(n9719), .B2(n8252), .A(n9791), .ZN(n8255) );
  NOR2_X1 U9939 ( .A1(n9708), .A2(n8253), .ZN(n8254) );
  AOI211_X1 U9940 ( .C1(n8256), .C2(n9693), .A(n8255), .B(n8254), .ZN(n8257)
         );
  OAI21_X1 U9941 ( .B1(n8258), .B2(n9695), .A(n8257), .ZN(P1_U3239) );
  XOR2_X1 U9942 ( .A(n8259), .B(n8260), .Z(n8268) );
  NAND2_X1 U9943 ( .A1(n8793), .A2(n9033), .ZN(n8262) );
  OAI211_X1 U9944 ( .C1(n8309), .C2(n8795), .A(n8262), .B(n8261), .ZN(n8265)
         );
  NOR2_X1 U9945 ( .A1(n8748), .A2(n8263), .ZN(n8264) );
  AOI211_X1 U9946 ( .C1(n8266), .C2(n8784), .A(n8265), .B(n8264), .ZN(n8267)
         );
  OAI21_X1 U9947 ( .B1(n8268), .B2(n8786), .A(n8267), .ZN(P2_U3161) );
  INV_X1 U9948 ( .A(n8269), .ZN(n8273) );
  OAI222_X1 U9949 ( .A1(n10224), .A2(n8272), .B1(n8271), .B2(n8273), .C1(
        P1_U3086), .C2(n8270), .ZN(P1_U3336) );
  OAI222_X1 U9950 ( .A1(n9537), .A2(n8274), .B1(n9547), .B2(n8273), .C1(
        P2_U3151), .C2(n9198), .ZN(P2_U3276) );
  NAND2_X1 U9951 ( .A1(n8276), .A2(n8819), .ZN(n8277) );
  NAND2_X1 U9952 ( .A1(n8275), .A2(n8277), .ZN(n8613) );
  INV_X1 U9953 ( .A(n8613), .ZN(n8285) );
  INV_X1 U9954 ( .A(n8278), .ZN(n8279) );
  NAND2_X1 U9955 ( .A1(n8280), .A2(n8279), .ZN(n8281) );
  XNOR2_X1 U9956 ( .A(n8281), .B(n8819), .ZN(n8284) );
  OR2_X1 U9957 ( .A1(n8613), .A2(n10544), .ZN(n8283) );
  AOI22_X1 U9958 ( .A1(n9382), .A2(n9032), .B1(n9030), .B2(n9380), .ZN(n8282)
         );
  OAI211_X1 U9959 ( .C1(n9356), .C2(n8284), .A(n8283), .B(n8282), .ZN(n8608)
         );
  AOI21_X1 U9960 ( .B1(n10554), .B2(n8285), .A(n8608), .ZN(n8347) );
  AOI22_X1 U9961 ( .A1(n9520), .A2(n8611), .B1(P2_REG0_REG_9__SCAN_IN), .B2(
        n10573), .ZN(n8286) );
  OAI21_X1 U9962 ( .B1(n8347), .B2(n10573), .A(n8286), .ZN(P2_U3417) );
  XNOR2_X1 U9963 ( .A(n8287), .B(n8288), .ZN(n8298) );
  INV_X1 U9964 ( .A(n8298), .ZN(n10467) );
  OAI21_X1 U9965 ( .B1(n8290), .B2(n8289), .A(n8288), .ZN(n10342) );
  INV_X1 U9966 ( .A(n10342), .ZN(n8292) );
  NOR3_X1 U9967 ( .A1(n8290), .A2(n8289), .A3(n8288), .ZN(n8291) );
  OAI21_X1 U9968 ( .B1(n8292), .B2(n8291), .A(n10399), .ZN(n8296) );
  OR2_X1 U9969 ( .A1(n8293), .A2(n9701), .ZN(n8295) );
  OR2_X1 U9970 ( .A1(n8566), .A2(n9703), .ZN(n8294) );
  AND2_X1 U9971 ( .A1(n8295), .A2(n8294), .ZN(n8328) );
  OAI211_X1 U9972 ( .C1(n8298), .C2(n8297), .A(n8296), .B(n8328), .ZN(n10465)
         );
  AOI21_X1 U9973 ( .B1(n8299), .B2(n10467), .A(n10465), .ZN(n8305) );
  OAI21_X1 U9974 ( .B1(n8300), .B2(n10464), .A(n10390), .ZN(n8301) );
  NOR2_X1 U9975 ( .A1(n8301), .A2(n10373), .ZN(n10462) );
  NOR2_X1 U9976 ( .A1(n10385), .A2(n10464), .ZN(n8303) );
  OAI22_X1 U9977 ( .A1(n10324), .A2(n7404), .B1(n8329), .B2(n10382), .ZN(n8302) );
  AOI211_X1 U9978 ( .C1(n10462), .C2(n10393), .A(n8303), .B(n8302), .ZN(n8304)
         );
  OAI21_X1 U9979 ( .B1(n8305), .B2(n10402), .A(n8304), .ZN(P1_U3286) );
  NAND2_X1 U9980 ( .A1(n8275), .A2(n8306), .ZN(n8307) );
  XNOR2_X1 U9981 ( .A(n8485), .B(n9030), .ZN(n8820) );
  XNOR2_X1 U9982 ( .A(n8307), .B(n8820), .ZN(n8379) );
  INV_X1 U9983 ( .A(n8379), .ZN(n8313) );
  XOR2_X1 U9984 ( .A(n8308), .B(n8820), .Z(n8311) );
  OAI22_X1 U9985 ( .A1(n8309), .A2(n10537), .B1(n8689), .B2(n10539), .ZN(n8310) );
  AOI21_X1 U9986 ( .B1(n8311), .B2(n10541), .A(n8310), .ZN(n8312) );
  OAI21_X1 U9987 ( .B1(n8379), .B2(n10544), .A(n8312), .ZN(n8373) );
  AOI21_X1 U9988 ( .B1(n10554), .B2(n8313), .A(n8373), .ZN(n8396) );
  AOI22_X1 U9989 ( .A1(n9520), .A2(n8485), .B1(P2_REG0_REG_10__SCAN_IN), .B2(
        n10573), .ZN(n8314) );
  OAI21_X1 U9990 ( .B1(n8396), .B2(n10573), .A(n8314), .ZN(P2_U3420) );
  NAND2_X1 U9991 ( .A1(n8335), .A2(n10217), .ZN(n8316) );
  OAI211_X1 U9992 ( .C1(n8317), .C2(n10224), .A(n8316), .B(n8315), .ZN(
        P1_U3335) );
  XOR2_X1 U9993 ( .A(n8318), .B(n8823), .Z(n8388) );
  XNOR2_X1 U9994 ( .A(n8319), .B(n8823), .ZN(n8320) );
  AOI222_X1 U9995 ( .A1(n10541), .A2(n8320), .B1(n9028), .B2(n9380), .C1(n9030), .C2(n9382), .ZN(n8383) );
  INV_X1 U9996 ( .A(n8383), .ZN(n8321) );
  NAND2_X1 U9997 ( .A1(n8321), .A2(n10571), .ZN(n8323) );
  AOI22_X1 U9998 ( .A1(n8530), .A2(n9520), .B1(P2_REG0_REG_11__SCAN_IN), .B2(
        n10573), .ZN(n8322) );
  OAI211_X1 U9999 ( .C1(n8388), .C2(n9524), .A(n8323), .B(n8322), .ZN(P2_U3423) );
  NAND2_X1 U10000 ( .A1(n8325), .A2(n8324), .ZN(n8327) );
  XOR2_X1 U10001 ( .A(n8327), .B(n8326), .Z(n8334) );
  NAND2_X1 U10002 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9805) );
  OAI21_X1 U10003 ( .B1(n9719), .B2(n8328), .A(n9805), .ZN(n8331) );
  NOR2_X1 U10004 ( .A1(n9708), .A2(n8329), .ZN(n8330) );
  OAI21_X1 U10005 ( .B1(n8334), .B2(n9695), .A(n8333), .ZN(P1_U3213) );
  INV_X1 U10006 ( .A(n8335), .ZN(n8337) );
  OAI222_X1 U10007 ( .A1(n9547), .A2(n8337), .B1(n8994), .B2(P2_U3151), .C1(
        n8336), .C2(n9537), .ZN(P2_U3275) );
  INV_X1 U10008 ( .A(n8611), .ZN(n8350) );
  AOI21_X1 U10009 ( .B1(n8339), .B2(n8338), .A(n8786), .ZN(n8341) );
  NAND2_X1 U10010 ( .A1(n8341), .A2(n8340), .ZN(n8346) );
  OAI21_X1 U10011 ( .B1(n8795), .B2(n8535), .A(n8342), .ZN(n8344) );
  NOR2_X1 U10012 ( .A1(n8748), .A2(n8609), .ZN(n8343) );
  AOI211_X1 U10013 ( .C1(n8793), .C2(n9032), .A(n8344), .B(n8343), .ZN(n8345)
         );
  OAI211_X1 U10014 ( .C1(n8350), .C2(n8800), .A(n8346), .B(n8345), .ZN(
        P2_U3171) );
  MUX2_X1 U10015 ( .A(n8348), .B(n8347), .S(n10578), .Z(n8349) );
  OAI21_X1 U10016 ( .B1(n8350), .B2(n9424), .A(n8349), .ZN(P2_U3468) );
  INV_X1 U10017 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10585) );
  INV_X1 U10018 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U10019 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n10292), .B2(n8351), .ZN(n10591) );
  NOR2_X1 U10020 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8352) );
  AOI21_X1 U10021 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n8352), .ZN(n10594) );
  AOI22_X1 U10022 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .B1(n10263), .B2(n9110), .ZN(n10597) );
  NOR2_X1 U10023 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8353) );
  AOI21_X1 U10024 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n8353), .ZN(n10600) );
  AOI22_X1 U10025 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .B1(n8355), .B2(n8354), .ZN(n10603) );
  NOR2_X1 U10026 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8356) );
  AOI21_X1 U10027 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n8356), .ZN(n10606) );
  NOR2_X1 U10028 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8357) );
  AOI21_X1 U10029 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n8357), .ZN(n10609) );
  NOR2_X1 U10030 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8358) );
  AOI21_X1 U10031 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n8358), .ZN(n10612) );
  NOR2_X1 U10032 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n8359) );
  AOI21_X1 U10033 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n8359), .ZN(n10618) );
  NOR2_X1 U10034 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n8360) );
  AOI21_X1 U10035 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n8360), .ZN(n10624) );
  NOR2_X1 U10036 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n8361) );
  AOI21_X1 U10037 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n8361), .ZN(n10621) );
  NOR2_X1 U10038 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n8362) );
  AOI21_X1 U10039 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n8362), .ZN(n10627) );
  NOR2_X1 U10040 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n8363) );
  AOI21_X1 U10041 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n8363), .ZN(n10615) );
  AND2_X1 U10042 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n8364) );
  NOR2_X1 U10043 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n8364), .ZN(n10580) );
  INV_X1 U10044 ( .A(n10580), .ZN(n10581) );
  INV_X1 U10045 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10583) );
  NAND3_X1 U10046 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10582) );
  NAND2_X1 U10047 ( .A1(n10583), .A2(n10582), .ZN(n10579) );
  NAND2_X1 U10048 ( .A1(n10581), .A2(n10579), .ZN(n10630) );
  NAND2_X1 U10049 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n8365) );
  OAI21_X1 U10050 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n8365), .ZN(n10629) );
  NOR2_X1 U10051 ( .A1(n10630), .A2(n10629), .ZN(n10628) );
  AOI21_X1 U10052 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10628), .ZN(n10633) );
  NAND2_X1 U10053 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n8366) );
  OAI21_X1 U10054 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n8366), .ZN(n10632) );
  NOR2_X1 U10055 ( .A1(n10633), .A2(n10632), .ZN(n10631) );
  AOI21_X1 U10056 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10631), .ZN(n10636) );
  NOR2_X1 U10057 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8367) );
  AOI21_X1 U10058 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n8367), .ZN(n10635) );
  NAND2_X1 U10059 ( .A1(n10636), .A2(n10635), .ZN(n10634) );
  OAI21_X1 U10060 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10634), .ZN(n10614) );
  NAND2_X1 U10061 ( .A1(n10615), .A2(n10614), .ZN(n10613) );
  OAI21_X1 U10062 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10613), .ZN(n10626) );
  NAND2_X1 U10063 ( .A1(n10627), .A2(n10626), .ZN(n10625) );
  OAI21_X1 U10064 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10625), .ZN(n10620) );
  NAND2_X1 U10065 ( .A1(n10621), .A2(n10620), .ZN(n10619) );
  OAI21_X1 U10066 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10619), .ZN(n10623) );
  NAND2_X1 U10067 ( .A1(n10624), .A2(n10623), .ZN(n10622) );
  OAI21_X1 U10068 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10622), .ZN(n10617) );
  NAND2_X1 U10069 ( .A1(n10618), .A2(n10617), .ZN(n10616) );
  OAI21_X1 U10070 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10616), .ZN(n10611) );
  NAND2_X1 U10071 ( .A1(n10612), .A2(n10611), .ZN(n10610) );
  OAI21_X1 U10072 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10610), .ZN(n10608) );
  NAND2_X1 U10073 ( .A1(n10609), .A2(n10608), .ZN(n10607) );
  OAI21_X1 U10074 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10607), .ZN(n10605) );
  NAND2_X1 U10075 ( .A1(n10606), .A2(n10605), .ZN(n10604) );
  OAI21_X1 U10076 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10604), .ZN(n10602) );
  NAND2_X1 U10077 ( .A1(n10603), .A2(n10602), .ZN(n10601) );
  OAI21_X1 U10078 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10601), .ZN(n10599) );
  NAND2_X1 U10079 ( .A1(n10600), .A2(n10599), .ZN(n10598) );
  OAI21_X1 U10080 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10598), .ZN(n10596) );
  NAND2_X1 U10081 ( .A1(n10597), .A2(n10596), .ZN(n10595) );
  OAI21_X1 U10082 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10595), .ZN(n10593) );
  NAND2_X1 U10083 ( .A1(n10594), .A2(n10593), .ZN(n10592) );
  OAI21_X1 U10084 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10592), .ZN(n10590) );
  NAND2_X1 U10085 ( .A1(n10591), .A2(n10590), .ZN(n10589) );
  OAI21_X1 U10086 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10589), .ZN(n10586) );
  NAND2_X1 U10087 ( .A1(n10585), .A2(n10586), .ZN(n8368) );
  NOR2_X1 U10088 ( .A1(n10585), .A2(n10586), .ZN(n10584) );
  AOI21_X1 U10089 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n8368), .A(n10584), .ZN(
        n8372) );
  NOR2_X1 U10090 ( .A1(n8370), .A2(n8369), .ZN(n8371) );
  XNOR2_X1 U10091 ( .A(n8372), .B(n8371), .ZN(ADD_1068_U4) );
  NAND2_X1 U10092 ( .A1(n9385), .A2(n10547), .ZN(n8643) );
  INV_X1 U10093 ( .A(n8373), .ZN(n8374) );
  MUX2_X1 U10094 ( .A(n8375), .B(n8374), .S(n9385), .Z(n8378) );
  INV_X1 U10095 ( .A(n8483), .ZN(n8376) );
  AOI22_X1 U10096 ( .A1(n8485), .A2(n4398), .B1(n9388), .B2(n8376), .ZN(n8377)
         );
  OAI211_X1 U10097 ( .C1(n8379), .C2(n8643), .A(n8378), .B(n8377), .ZN(
        P2_U3223) );
  MUX2_X1 U10098 ( .A(n8380), .B(n8383), .S(n10578), .Z(n8382) );
  NAND2_X1 U10099 ( .A1(n8530), .A2(n9438), .ZN(n8381) );
  OAI211_X1 U10100 ( .C1(n8388), .C2(n9441), .A(n8382), .B(n8381), .ZN(
        P2_U3470) );
  MUX2_X1 U10101 ( .A(n8384), .B(n8383), .S(n9385), .Z(n8387) );
  INV_X1 U10102 ( .A(n8536), .ZN(n8385) );
  AOI22_X1 U10103 ( .A1(n8530), .A2(n4398), .B1(n9388), .B2(n8385), .ZN(n8386)
         );
  OAI211_X1 U10104 ( .C1(n8388), .C2(n9366), .A(n8387), .B(n8386), .ZN(
        P2_U3222) );
  OAI21_X1 U10105 ( .B1(n8390), .B2(n8919), .A(n8389), .ZN(n8448) );
  XNOR2_X1 U10106 ( .A(n8391), .B(n8919), .ZN(n8392) );
  OAI222_X1 U10107 ( .A1(n10537), .A2(n8689), .B1(n10539), .B2(n8925), .C1(
        n8392), .C2(n9356), .ZN(n8442) );
  NAND2_X1 U10108 ( .A1(n8442), .A2(n9385), .ZN(n8395) );
  OAI22_X1 U10109 ( .A1(n9385), .A2(n9037), .B1(n8693), .B2(n10533), .ZN(n8393) );
  AOI21_X1 U10110 ( .B1(n8921), .B2(n4398), .A(n8393), .ZN(n8394) );
  OAI211_X1 U10111 ( .C1(n8448), .C2(n9366), .A(n8395), .B(n8394), .ZN(
        P2_U3221) );
  INV_X1 U10112 ( .A(n8485), .ZN(n8399) );
  MUX2_X1 U10113 ( .A(n8397), .B(n8396), .S(n10578), .Z(n8398) );
  OAI21_X1 U10114 ( .B1(n8399), .B2(n9424), .A(n8398), .ZN(P2_U3469) );
  INV_X1 U10115 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8406) );
  INV_X1 U10116 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8400) );
  OR2_X1 U10117 ( .A1(n8401), .A2(n8400), .ZN(n8405) );
  INV_X1 U10118 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8402) );
  OR2_X1 U10119 ( .A1(n8403), .A2(n8402), .ZN(n8404) );
  OAI211_X1 U10120 ( .C1(n7138), .C2(n8406), .A(n8405), .B(n8404), .ZN(n8407)
         );
  INV_X1 U10121 ( .A(n8407), .ZN(n8408) );
  INV_X1 U10122 ( .A(n9219), .ZN(n9011) );
  NAND2_X1 U10123 ( .A1(n9011), .A2(P2_U3893), .ZN(n8410) );
  OAI21_X1 U10124 ( .B1(P2_U3893), .B2(n10214), .A(n8410), .ZN(P2_U3522) );
  XNOR2_X1 U10125 ( .A(n8412), .B(n8411), .ZN(n10493) );
  NAND2_X1 U10126 ( .A1(n10325), .A2(n8413), .ZN(n8415) );
  NAND2_X1 U10127 ( .A1(n8415), .A2(n8414), .ZN(n8416) );
  NAND3_X1 U10128 ( .A1(n8416), .A2(n10311), .A3(n10399), .ZN(n8420) );
  OR2_X1 U10129 ( .A1(n8417), .A2(n9703), .ZN(n8419) );
  NAND2_X1 U10130 ( .A1(n9687), .A2(n9744), .ZN(n8418) );
  AND2_X1 U10131 ( .A1(n8419), .A2(n8418), .ZN(n9679) );
  NAND2_X1 U10132 ( .A1(n8420), .A2(n9679), .ZN(n10488) );
  INV_X1 U10133 ( .A(n8421), .ZN(n10336) );
  AOI211_X1 U10134 ( .C1(n10489), .C2(n10336), .A(n10407), .B(n5279), .ZN(
        n10487) );
  NAND2_X1 U10135 ( .A1(n10487), .A2(n10393), .ZN(n8423) );
  AOI22_X1 U10136 ( .A1(n10402), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9677), 
        .B2(n10401), .ZN(n8422) );
  OAI211_X1 U10137 ( .C1(n6395), .C2(n10385), .A(n8423), .B(n8422), .ZN(n8424)
         );
  AOI21_X1 U10138 ( .B1(n10324), .B2(n10488), .A(n8424), .ZN(n8425) );
  OAI21_X1 U10139 ( .B1(n10493), .B2(n10412), .A(n8425), .ZN(P1_U3282) );
  INV_X1 U10140 ( .A(n8426), .ZN(n8629) );
  OAI222_X1 U10141 ( .A1(n9547), .A2(n8629), .B1(n8863), .B2(P2_U3151), .C1(
        n8427), .C2(n9537), .ZN(P2_U3274) );
  INV_X1 U10142 ( .A(n8928), .ZN(n8429) );
  NAND2_X1 U10143 ( .A1(n8429), .A2(n8927), .ZN(n8825) );
  XNOR2_X1 U10144 ( .A(n8428), .B(n8825), .ZN(n8475) );
  XNOR2_X1 U10145 ( .A(n8430), .B(n8825), .ZN(n8431) );
  NAND2_X1 U10146 ( .A1(n8431), .A2(n10541), .ZN(n8433) );
  AOI22_X1 U10147 ( .A1(n9382), .A2(n9028), .B1(n9383), .B2(n9380), .ZN(n8432)
         );
  NAND2_X1 U10148 ( .A1(n8433), .A2(n8432), .ZN(n8471) );
  OAI22_X1 U10149 ( .A1(n8926), .A2(n10531), .B1(n8749), .B2(n10533), .ZN(
        n8434) );
  OAI21_X1 U10150 ( .B1(n8471), .B2(n8434), .A(n9385), .ZN(n8436) );
  NAND2_X1 U10151 ( .A1(n10550), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8435) );
  OAI211_X1 U10152 ( .C1(n8475), .C2(n9366), .A(n8436), .B(n8435), .ZN(
        P2_U3220) );
  INV_X1 U10153 ( .A(n8437), .ZN(n8440) );
  OAI222_X1 U10154 ( .A1(n10224), .A2(n8439), .B1(n8271), .B2(n8440), .C1(
        P1_U3086), .C2(n8438), .ZN(P1_U3333) );
  OAI222_X1 U10155 ( .A1(n9537), .A2(n8441), .B1(n9547), .B2(n8440), .C1(
        P2_U3151), .C2(n8869), .ZN(P2_U3273) );
  AOI21_X1 U10156 ( .B1(n9443), .B2(n8921), .A(n8442), .ZN(n8445) );
  MUX2_X1 U10157 ( .A(n8443), .B(n8445), .S(n10578), .Z(n8444) );
  OAI21_X1 U10158 ( .B1(n9441), .B2(n8448), .A(n8444), .ZN(P2_U3471) );
  INV_X1 U10159 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8446) );
  MUX2_X1 U10160 ( .A(n8446), .B(n8445), .S(n10571), .Z(n8447) );
  OAI21_X1 U10161 ( .B1(n8448), .B2(n9524), .A(n8447), .ZN(P2_U3426) );
  MUX2_X1 U10162 ( .A(n8471), .B(P2_REG0_REG_13__SCAN_IN), .S(n10573), .Z(
        n8450) );
  OAI22_X1 U10163 ( .A1(n8475), .A2(n9524), .B1(n8926), .B2(n9500), .ZN(n8449)
         );
  OR2_X1 U10164 ( .A1(n8450), .A2(n8449), .ZN(P2_U3429) );
  NAND2_X1 U10165 ( .A1(n8455), .A2(n8451), .ZN(n8453) );
  NAND2_X1 U10166 ( .A1(n8452), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9022) );
  OAI211_X1 U10167 ( .C1(n8454), .C2(n9537), .A(n8453), .B(n9022), .ZN(
        P2_U3272) );
  NAND2_X1 U10168 ( .A1(n8455), .A2(n10217), .ZN(n8457) );
  OAI211_X1 U10169 ( .C1(n8458), .C2(n10224), .A(n8457), .B(n8456), .ZN(
        P1_U3332) );
  XNOR2_X1 U10170 ( .A(n8459), .B(n8460), .ZN(n8461) );
  NAND2_X1 U10171 ( .A1(n8461), .A2(n8462), .ZN(n8559) );
  OAI21_X1 U10172 ( .B1(n8462), .B2(n8461), .A(n8559), .ZN(n8463) );
  NAND2_X1 U10173 ( .A1(n8463), .A2(n9716), .ZN(n8470) );
  OR2_X1 U10174 ( .A1(n8464), .A2(n9701), .ZN(n8466) );
  OR2_X1 U10175 ( .A1(n8553), .A2(n9703), .ZN(n8465) );
  AND2_X1 U10176 ( .A1(n8466), .A2(n8465), .ZN(n10363) );
  NAND2_X1 U10177 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9818) );
  OAI21_X1 U10178 ( .B1(n9719), .B2(n10363), .A(n9818), .ZN(n8467) );
  AOI21_X1 U10179 ( .B1(n9693), .B2(n8468), .A(n8467), .ZN(n8469) );
  OAI211_X1 U10180 ( .C1(n9708), .C2(n10366), .A(n8470), .B(n8469), .ZN(
        P1_U3221) );
  INV_X1 U10181 ( .A(n8471), .ZN(n8472) );
  MUX2_X1 U10182 ( .A(n8472), .B(n9044), .S(n7168), .Z(n8474) );
  NAND2_X1 U10183 ( .A1(n8751), .A2(n9438), .ZN(n8473) );
  OAI211_X1 U10184 ( .C1(n9441), .C2(n8475), .A(n8474), .B(n8473), .ZN(
        P2_U3472) );
  NAND2_X1 U10185 ( .A1(n8477), .A2(n8476), .ZN(n8478) );
  XOR2_X1 U10186 ( .A(n8479), .B(n8478), .Z(n8487) );
  OAI21_X1 U10187 ( .B1(n8795), .B2(n8689), .A(n8480), .ZN(n8481) );
  AOI21_X1 U10188 ( .B1(n8793), .B2(n9031), .A(n8481), .ZN(n8482) );
  OAI21_X1 U10189 ( .B1(n8483), .B2(n8748), .A(n8482), .ZN(n8484) );
  AOI21_X1 U10190 ( .B1(n8485), .B2(n8784), .A(n8484), .ZN(n8486) );
  OAI21_X1 U10191 ( .B1(n8487), .B2(n8786), .A(n8486), .ZN(P2_U3157) );
  INV_X1 U10192 ( .A(n8488), .ZN(n8492) );
  OAI222_X1 U10193 ( .A1(n10224), .A2(n8490), .B1(n8271), .B2(n8492), .C1(
        n8489), .C2(P1_U3086), .ZN(P1_U3331) );
  OAI222_X1 U10194 ( .A1(n9537), .A2(n8493), .B1(n9547), .B2(n8492), .C1(n8491), .C2(P2_U3151), .ZN(P2_U3271) );
  XOR2_X1 U10195 ( .A(n8495), .B(n8494), .Z(n8501) );
  INV_X1 U10196 ( .A(n8496), .ZN(n9743) );
  AOI22_X1 U10197 ( .A1(n9649), .A2(n9741), .B1(n9743), .B2(n9687), .ZN(n10314) );
  NAND2_X1 U10198 ( .A1(n9721), .A2(n10316), .ZN(n8498) );
  OAI211_X1 U10199 ( .C1(n9719), .C2(n10314), .A(n8498), .B(n8497), .ZN(n8499)
         );
  AOI21_X1 U10200 ( .B1(n10317), .B2(n9693), .A(n8499), .ZN(n8500) );
  OAI21_X1 U10201 ( .B1(n8501), .B2(n9695), .A(n8500), .ZN(P1_U3224) );
  XNOR2_X1 U10202 ( .A(n8503), .B(n8502), .ZN(n10150) );
  INV_X1 U10203 ( .A(n8504), .ZN(n8505) );
  AOI211_X1 U10204 ( .C1(n10147), .C2(n4437), .A(n10407), .B(n8505), .ZN(
        n10146) );
  INV_X1 U10205 ( .A(n9555), .ZN(n8506) );
  AOI22_X1 U10206 ( .A1(n10402), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8506), 
        .B2(n10401), .ZN(n8507) );
  OAI21_X1 U10207 ( .B1(n8508), .B2(n10385), .A(n8507), .ZN(n8515) );
  XNOR2_X1 U10208 ( .A(n8510), .B(n8509), .ZN(n8513) );
  OAI22_X1 U10209 ( .A1(n8512), .A2(n9703), .B1(n8511), .B2(n9701), .ZN(n9553)
         );
  AOI21_X1 U10210 ( .B1(n8513), .B2(n10399), .A(n9553), .ZN(n10149) );
  NOR2_X1 U10211 ( .A1(n10149), .A2(n10402), .ZN(n8514) );
  AOI211_X1 U10212 ( .C1(n10146), .C2(n10393), .A(n8515), .B(n8514), .ZN(n8516) );
  OAI21_X1 U10213 ( .B1(n10150), .B2(n10412), .A(n8516), .ZN(P1_U3279) );
  XNOR2_X1 U10214 ( .A(n8517), .B(n8522), .ZN(n10508) );
  INV_X1 U10215 ( .A(n10508), .ZN(n8529) );
  NAND2_X1 U10216 ( .A1(n10313), .A2(n8518), .ZN(n8521) );
  INV_X1 U10217 ( .A(n8519), .ZN(n8520) );
  AOI21_X1 U10218 ( .B1(n8522), .B2(n8521), .A(n8520), .ZN(n8523) );
  AOI22_X1 U10219 ( .A1(n9649), .A2(n9740), .B1(n9742), .B2(n9687), .ZN(n8588)
         );
  OAI21_X1 U10220 ( .B1(n8523), .B2(n10048), .A(n8588), .ZN(n10506) );
  OAI211_X1 U10221 ( .C1(n10504), .C2(n8524), .A(n4437), .B(n10390), .ZN(
        n10502) );
  NOR2_X1 U10222 ( .A1(n10502), .A2(n10411), .ZN(n8527) );
  AOI22_X1 U10223 ( .A1(n10402), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8585), 
        .B2(n10401), .ZN(n8525) );
  OAI21_X1 U10224 ( .B1(n10504), .B2(n10385), .A(n8525), .ZN(n8526) );
  AOI211_X1 U10225 ( .C1(n10506), .C2(n10324), .A(n8527), .B(n8526), .ZN(n8528) );
  OAI21_X1 U10226 ( .B1(n8529), .B2(n10412), .A(n8528), .ZN(P1_U3280) );
  INV_X1 U10227 ( .A(n8530), .ZN(n8541) );
  OAI211_X1 U10228 ( .C1(n8533), .C2(n8532), .A(n8531), .B(n8790), .ZN(n8540)
         );
  OAI21_X1 U10229 ( .B1(n8782), .B2(n8535), .A(n8534), .ZN(n8538) );
  NOR2_X1 U10230 ( .A1(n8748), .A2(n8536), .ZN(n8537) );
  AOI211_X1 U10231 ( .C1(n8779), .C2(n9028), .A(n8538), .B(n8537), .ZN(n8539)
         );
  OAI211_X1 U10232 ( .C1(n8541), .C2(n8800), .A(n8540), .B(n8539), .ZN(
        P2_U3176) );
  XNOR2_X1 U10233 ( .A(n8542), .B(n8827), .ZN(n8576) );
  INV_X1 U10234 ( .A(n8827), .ZN(n8938) );
  XNOR2_X1 U10235 ( .A(n8543), .B(n8938), .ZN(n8544) );
  AOI222_X1 U10236 ( .A1(n10541), .A2(n8544), .B1(n8691), .B2(n9382), .C1(
        n9370), .C2(n9380), .ZN(n8571) );
  MUX2_X1 U10237 ( .A(n9101), .B(n8571), .S(n10578), .Z(n8546) );
  NAND2_X1 U10238 ( .A1(n8934), .A2(n9438), .ZN(n8545) );
  OAI211_X1 U10239 ( .C1(n9441), .C2(n8576), .A(n8546), .B(n8545), .ZN(
        P2_U3473) );
  MUX2_X1 U10240 ( .A(n8547), .B(n8571), .S(n10571), .Z(n8549) );
  NAND2_X1 U10241 ( .A1(n8934), .A2(n9520), .ZN(n8548) );
  OAI211_X1 U10242 ( .C1(n8576), .C2(n9524), .A(n8549), .B(n8548), .ZN(
        P2_U3432) );
  XNOR2_X1 U10243 ( .A(n8550), .B(n9672), .ZN(n8551) );
  NOR2_X1 U10244 ( .A1(n8551), .A2(n8552), .ZN(n9671) );
  AOI21_X1 U10245 ( .B1(n8552), .B2(n8551), .A(n9671), .ZN(n8558) );
  INV_X1 U10246 ( .A(n8553), .ZN(n9745) );
  AOI22_X1 U10247 ( .A1(n9649), .A2(n9743), .B1(n9745), .B2(n9687), .ZN(n10327) );
  OAI21_X1 U10248 ( .B1(n9719), .B2(n10327), .A(n8554), .ZN(n8556) );
  NOR2_X1 U10249 ( .A1(n9708), .A2(n10330), .ZN(n8555) );
  AOI211_X1 U10250 ( .C1(n10335), .C2(n9693), .A(n8556), .B(n8555), .ZN(n8557)
         );
  OAI21_X1 U10251 ( .B1(n8558), .B2(n9695), .A(n8557), .ZN(P1_U3217) );
  OAI21_X1 U10252 ( .B1(n8560), .B2(n8459), .A(n8559), .ZN(n8564) );
  XNOR2_X1 U10253 ( .A(n8562), .B(n8561), .ZN(n8563) );
  XNOR2_X1 U10254 ( .A(n8564), .B(n8563), .ZN(n8565) );
  NAND2_X1 U10255 ( .A1(n8565), .A2(n9716), .ZN(n8570) );
  OR2_X1 U10256 ( .A1(n8566), .A2(n9701), .ZN(n10347) );
  NAND2_X1 U10257 ( .A1(n9744), .A2(n9649), .ZN(n10356) );
  AOI21_X1 U10258 ( .B1(n10347), .B2(n10356), .A(n9719), .ZN(n8567) );
  AOI211_X1 U10259 ( .C1(n6101), .C2(n9693), .A(n8568), .B(n8567), .ZN(n8569)
         );
  OAI211_X1 U10260 ( .C1(n9708), .C2(n10350), .A(n8570), .B(n8569), .ZN(
        P1_U3231) );
  INV_X1 U10261 ( .A(n8934), .ZN(n8572) );
  OAI21_X1 U10262 ( .B1(n8572), .B2(n10531), .A(n8571), .ZN(n8573) );
  NAND2_X1 U10263 ( .A1(n8573), .A2(n9385), .ZN(n8575) );
  AOI22_X1 U10264 ( .A1(n10550), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n9388), 
        .B2(n8655), .ZN(n8574) );
  OAI211_X1 U10265 ( .C1(n8576), .C2(n9366), .A(n8575), .B(n8574), .ZN(
        P2_U3219) );
  INV_X1 U10266 ( .A(n8577), .ZN(n8581) );
  OAI222_X1 U10267 ( .A1(n9537), .A2(n8579), .B1(n9547), .B2(n8581), .C1(n8578), .C2(P2_U3151), .ZN(P2_U3270) );
  OAI222_X1 U10268 ( .A1(n10224), .A2(n8582), .B1(n8271), .B2(n8581), .C1(
        n8580), .C2(P1_U3086), .ZN(P1_U3330) );
  XOR2_X1 U10269 ( .A(n8584), .B(n8583), .Z(n8592) );
  NAND2_X1 U10270 ( .A1(n9721), .A2(n8585), .ZN(n8587) );
  OAI211_X1 U10271 ( .C1(n9719), .C2(n8588), .A(n8587), .B(n8586), .ZN(n8589)
         );
  AOI21_X1 U10272 ( .B1(n8590), .B2(n9693), .A(n8589), .ZN(n8591) );
  OAI21_X1 U10273 ( .B1(n8592), .B2(n9695), .A(n8591), .ZN(P1_U3234) );
  INV_X1 U10274 ( .A(n8593), .ZN(n10226) );
  OAI222_X1 U10275 ( .A1(n9547), .A2(n10226), .B1(P2_U3151), .B2(n8595), .C1(
        n8594), .C2(n9537), .ZN(P2_U3269) );
  XNOR2_X1 U10276 ( .A(n8596), .B(n8598), .ZN(n10206) );
  XNOR2_X1 U10277 ( .A(n8597), .B(n8598), .ZN(n8599) );
  NAND2_X1 U10278 ( .A1(n8599), .A2(n10399), .ZN(n8601) );
  AND2_X1 U10279 ( .A1(n9740), .A2(n9687), .ZN(n8600) );
  AOI21_X1 U10280 ( .B1(n9737), .B2(n9649), .A(n8600), .ZN(n9718) );
  NAND2_X1 U10281 ( .A1(n8601), .A2(n9718), .ZN(n10142) );
  INV_X1 U10282 ( .A(n10068), .ZN(n8602) );
  AOI211_X1 U10283 ( .C1(n10143), .C2(n8504), .A(n10407), .B(n8602), .ZN(
        n10141) );
  NAND2_X1 U10284 ( .A1(n10141), .A2(n10393), .ZN(n8605) );
  INV_X1 U10285 ( .A(n8603), .ZN(n9722) );
  AOI22_X1 U10286 ( .A1(n10402), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9722), 
        .B2(n10401), .ZN(n8604) );
  OAI211_X1 U10287 ( .C1(n9726), .C2(n10385), .A(n8605), .B(n8604), .ZN(n8606)
         );
  AOI21_X1 U10288 ( .B1(n10324), .B2(n10142), .A(n8606), .ZN(n8607) );
  OAI21_X1 U10289 ( .B1(n10206), .B2(n10412), .A(n8607), .ZN(P1_U3278) );
  MUX2_X1 U10290 ( .A(n8608), .B(P2_REG2_REG_9__SCAN_IN), .S(n10550), .Z(n8615) );
  NOR2_X1 U10291 ( .A1(n10533), .A2(n8609), .ZN(n8610) );
  AOI21_X1 U10292 ( .B1(n4398), .B2(n8611), .A(n8610), .ZN(n8612) );
  OAI21_X1 U10293 ( .B1(n8613), .B2(n8643), .A(n8612), .ZN(n8614) );
  OR2_X1 U10294 ( .A1(n8615), .A2(n8614), .ZN(P2_U3224) );
  NAND2_X1 U10295 ( .A1(n8617), .A2(n10394), .ZN(n8625) );
  NOR2_X1 U10296 ( .A1(n8618), .A2(n10385), .ZN(n8622) );
  OAI22_X1 U10297 ( .A1(n10324), .A2(n8620), .B1(n8619), .B2(n10382), .ZN(
        n8621) );
  AOI211_X1 U10298 ( .C1(n8623), .C2(n10393), .A(n8622), .B(n8621), .ZN(n8624)
         );
  OAI211_X1 U10299 ( .C1(n8616), .C2(n10402), .A(n8625), .B(n8624), .ZN(
        P1_U3356) );
  INV_X1 U10300 ( .A(n8626), .ZN(n9548) );
  OAI222_X1 U10301 ( .A1(n10224), .A2(n8627), .B1(n8271), .B2(n9548), .C1(
        n6123), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U10302 ( .A1(n10224), .A2(n8630), .B1(n8271), .B2(n8629), .C1(
        n8628), .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U10303 ( .A(n9910), .ZN(n8637) );
  AOI22_X1 U10304 ( .A1(n9731), .A2(n9687), .B1(n9649), .B2(n9729), .ZN(n9908)
         );
  OAI22_X1 U10305 ( .A1(n9719), .A2(n9908), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8635), .ZN(n8636) );
  AOI21_X1 U10306 ( .B1(n8637), .B2(n9721), .A(n8636), .ZN(n8638) );
  INV_X1 U10307 ( .A(n8639), .ZN(n9543) );
  OAI222_X1 U10308 ( .A1(n10224), .A2(n8640), .B1(n8271), .B2(n9543), .C1(
        n6115), .C2(P1_U3086), .ZN(P1_U3327) );
  NAND2_X1 U10309 ( .A1(n8641), .A2(n9388), .ZN(n9220) );
  OAI21_X1 U10310 ( .B1(n9385), .B2(n8642), .A(n9220), .ZN(n8645) );
  NOR2_X1 U10311 ( .A1(n7146), .A2(n8643), .ZN(n8644) );
  AOI211_X1 U10312 ( .C1(n4398), .C2(n8646), .A(n8645), .B(n8644), .ZN(n8647)
         );
  OAI21_X1 U10313 ( .B1(n8648), .B2(n10550), .A(n8647), .ZN(P2_U3204) );
  INV_X1 U10314 ( .A(n8650), .ZN(n8651) );
  AOI21_X1 U10315 ( .B1(n8652), .B2(n8649), .A(n8651), .ZN(n8658) );
  NAND2_X1 U10316 ( .A1(n8793), .A2(n8691), .ZN(n8653) );
  NAND2_X1 U10317 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9070) );
  OAI211_X1 U10318 ( .C1(n8708), .C2(n8795), .A(n8653), .B(n9070), .ZN(n8654)
         );
  AOI21_X1 U10319 ( .B1(n8655), .B2(n8797), .A(n8654), .ZN(n8657) );
  NAND2_X1 U10320 ( .A1(n8934), .A2(n8784), .ZN(n8656) );
  OAI211_X1 U10321 ( .C1(n8658), .C2(n8786), .A(n8657), .B(n8656), .ZN(
        P2_U3155) );
  XNOR2_X1 U10322 ( .A(n8724), .B(n9288), .ZN(n8664) );
  AOI22_X1 U10323 ( .A1(n9283), .A2(n8797), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8661) );
  NAND2_X1 U10324 ( .A1(n9304), .A2(n8793), .ZN(n8660) );
  OAI211_X1 U10325 ( .C1(n8974), .C2(n8795), .A(n8661), .B(n8660), .ZN(n8662)
         );
  AOI21_X1 U10326 ( .B1(n9481), .B2(n8784), .A(n8662), .ZN(n8663) );
  OAI21_X1 U10327 ( .B1(n8664), .B2(n8786), .A(n8663), .ZN(P2_U3156) );
  INV_X1 U10328 ( .A(n9329), .ZN(n9501) );
  NAND2_X1 U10329 ( .A1(n8713), .A2(n8665), .ZN(n8765) );
  XNOR2_X1 U10330 ( .A(n8666), .B(n9027), .ZN(n8766) );
  NAND2_X1 U10331 ( .A1(n8765), .A2(n8766), .ZN(n8764) );
  AND2_X1 U10332 ( .A1(n8764), .A2(n8668), .ZN(n8670) );
  XNOR2_X1 U10333 ( .A(n8667), .B(n9318), .ZN(n8669) );
  NAND3_X1 U10334 ( .A1(n8764), .A2(n8669), .A3(n8668), .ZN(n8733) );
  OAI211_X1 U10335 ( .C1(n8670), .C2(n8669), .A(n8790), .B(n8733), .ZN(n8675)
         );
  NOR2_X1 U10336 ( .A1(n8671), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9208) );
  AOI21_X1 U10337 ( .B1(n9027), .B2(n8793), .A(n9208), .ZN(n8672) );
  OAI21_X1 U10338 ( .B1(n9333), .B2(n8795), .A(n8672), .ZN(n8673) );
  AOI21_X1 U10339 ( .B1(n9337), .B2(n8797), .A(n8673), .ZN(n8674) );
  OAI211_X1 U10340 ( .C1(n9501), .C2(n8800), .A(n8675), .B(n8674), .ZN(
        P2_U3159) );
  OAI21_X1 U10341 ( .B1(n8678), .B2(n8677), .A(n8676), .ZN(n8679) );
  NAND2_X1 U10342 ( .A1(n8679), .A2(n8790), .ZN(n8684) );
  INV_X1 U10343 ( .A(n9308), .ZN(n8681) );
  AOI22_X1 U10344 ( .A1(n9305), .A2(n8793), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8680) );
  OAI21_X1 U10345 ( .B1(n8681), .B2(n8748), .A(n8680), .ZN(n8682) );
  AOI21_X1 U10346 ( .B1(n8779), .B2(n9304), .A(n8682), .ZN(n8683) );
  OAI211_X1 U10347 ( .C1(n8685), .C2(n8800), .A(n8684), .B(n8683), .ZN(
        P2_U3163) );
  XNOR2_X1 U10348 ( .A(n8686), .B(n8920), .ZN(n8687) );
  XNOR2_X1 U10349 ( .A(n4765), .B(n8687), .ZN(n8696) );
  OAI21_X1 U10350 ( .B1(n8782), .B2(n8689), .A(n8688), .ZN(n8690) );
  AOI21_X1 U10351 ( .B1(n8779), .B2(n8691), .A(n8690), .ZN(n8692) );
  OAI21_X1 U10352 ( .B1(n8693), .B2(n8748), .A(n8692), .ZN(n8694) );
  AOI21_X1 U10353 ( .B1(n8921), .B2(n8784), .A(n8694), .ZN(n8695) );
  OAI21_X1 U10354 ( .B1(n8696), .B2(n8786), .A(n8695), .ZN(P2_U3164) );
  XOR2_X1 U10355 ( .A(n8698), .B(n8697), .Z(n8704) );
  AOI22_X1 U10356 ( .A1(n9258), .A2(n8797), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8700) );
  NAND2_X1 U10357 ( .A1(n5874), .A2(n8793), .ZN(n8699) );
  OAI211_X1 U10358 ( .C1(n8701), .C2(n8795), .A(n8700), .B(n8699), .ZN(n8702)
         );
  AOI21_X1 U10359 ( .B1(n9469), .B2(n8784), .A(n8702), .ZN(n8703) );
  OAI21_X1 U10360 ( .B1(n8704), .B2(n8786), .A(n8703), .ZN(P2_U3165) );
  XNOR2_X1 U10361 ( .A(n8706), .B(n8705), .ZN(n8712) );
  NAND2_X1 U10362 ( .A1(n9371), .A2(n8779), .ZN(n8707) );
  NAND2_X1 U10363 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9131) );
  OAI211_X1 U10364 ( .C1(n8708), .C2(n8782), .A(n8707), .B(n9131), .ZN(n8709)
         );
  AOI21_X1 U10365 ( .B1(n9374), .B2(n8797), .A(n8709), .ZN(n8711) );
  NAND2_X1 U10366 ( .A1(n9514), .A2(n8784), .ZN(n8710) );
  OAI211_X1 U10367 ( .C1(n8712), .C2(n8786), .A(n8711), .B(n8710), .ZN(
        P2_U3166) );
  INV_X1 U10368 ( .A(n8713), .ZN(n8714) );
  AOI21_X1 U10369 ( .B1(n8716), .B2(n8715), .A(n8714), .ZN(n8721) );
  NAND2_X1 U10370 ( .A1(n9027), .A2(n8779), .ZN(n8717) );
  NAND2_X1 U10371 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9152) );
  OAI211_X1 U10372 ( .C1(n9359), .C2(n8782), .A(n8717), .B(n9152), .ZN(n8719)
         );
  NOR2_X1 U10373 ( .A1(n9363), .A2(n8800), .ZN(n8718) );
  AOI211_X1 U10374 ( .C1(n9360), .C2(n8797), .A(n8719), .B(n8718), .ZN(n8720)
         );
  OAI21_X1 U10375 ( .B1(n8721), .B2(n8786), .A(n8720), .ZN(P2_U3168) );
  XNOR2_X1 U10376 ( .A(n8725), .B(n8974), .ZN(n8726) );
  XNOR2_X1 U10377 ( .A(n8727), .B(n8726), .ZN(n8732) );
  NOR2_X1 U10378 ( .A1(n9026), .A2(n8795), .ZN(n8730) );
  AOI22_X1 U10379 ( .A1(n9271), .A2(n8797), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8728) );
  OAI21_X1 U10380 ( .B1(n9288), .B2(n8782), .A(n8728), .ZN(n8729) );
  AOI211_X1 U10381 ( .C1(n9475), .C2(n8784), .A(n8730), .B(n8729), .ZN(n8731)
         );
  OAI21_X1 U10382 ( .B1(n8732), .B2(n8786), .A(n8731), .ZN(P2_U3169) );
  OAI21_X1 U10383 ( .B1(n9318), .B2(n8734), .A(n8733), .ZN(n8738) );
  INV_X1 U10384 ( .A(n8735), .ZN(n8736) );
  AOI21_X1 U10385 ( .B1(n8738), .B2(n8737), .A(n8736), .ZN(n8743) );
  AOI22_X1 U10386 ( .A1(n9345), .A2(n8793), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8740) );
  NAND2_X1 U10387 ( .A1(n9319), .A2(n8797), .ZN(n8739) );
  OAI211_X1 U10388 ( .C1(n9317), .C2(n8795), .A(n8740), .B(n8739), .ZN(n8741)
         );
  AOI21_X1 U10389 ( .B1(n7088), .B2(n8784), .A(n8741), .ZN(n8742) );
  OAI21_X1 U10390 ( .B1(n8743), .B2(n8786), .A(n8742), .ZN(P2_U3173) );
  XNOR2_X1 U10391 ( .A(n8745), .B(n8744), .ZN(n8753) );
  NAND2_X1 U10392 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9043) );
  OAI21_X1 U10393 ( .B1(n8795), .B2(n8933), .A(n9043), .ZN(n8746) );
  AOI21_X1 U10394 ( .B1(n8793), .B2(n9028), .A(n8746), .ZN(n8747) );
  OAI21_X1 U10395 ( .B1(n8749), .B2(n8748), .A(n8747), .ZN(n8750) );
  AOI21_X1 U10396 ( .B1(n8751), .B2(n8784), .A(n8750), .ZN(n8752) );
  OAI21_X1 U10397 ( .B1(n8753), .B2(n8786), .A(n8752), .ZN(P2_U3174) );
  XNOR2_X1 U10398 ( .A(n8755), .B(n8754), .ZN(n8756) );
  XNOR2_X1 U10399 ( .A(n8757), .B(n8756), .ZN(n8763) );
  OAI22_X1 U10400 ( .A1(n9317), .A2(n8782), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8758), .ZN(n8759) );
  AOI21_X1 U10401 ( .B1(n9292), .B2(n8797), .A(n8759), .ZN(n8760) );
  OAI21_X1 U10402 ( .B1(n9288), .B2(n8795), .A(n8760), .ZN(n8761) );
  AOI21_X1 U10403 ( .B1(n9291), .B2(n8784), .A(n8761), .ZN(n8762) );
  OAI21_X1 U10404 ( .B1(n8763), .B2(n8786), .A(n8762), .ZN(P2_U3175) );
  INV_X1 U10405 ( .A(n9507), .ZN(n8773) );
  OAI21_X1 U10406 ( .B1(n8766), .B2(n8765), .A(n8764), .ZN(n8767) );
  NAND2_X1 U10407 ( .A1(n8767), .A2(n8790), .ZN(n8772) );
  NAND2_X1 U10408 ( .A1(n9345), .A2(n8779), .ZN(n8768) );
  NAND2_X1 U10409 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9170) );
  OAI211_X1 U10410 ( .C1(n8769), .C2(n8782), .A(n8768), .B(n9170), .ZN(n8770)
         );
  AOI21_X1 U10411 ( .B1(n9348), .B2(n8797), .A(n8770), .ZN(n8771) );
  OAI211_X1 U10412 ( .C1(n8773), .C2(n8800), .A(n8772), .B(n8771), .ZN(
        P2_U3178) );
  NAND2_X1 U10413 ( .A1(n8775), .A2(n8774), .ZN(n8778) );
  XNOR2_X1 U10414 ( .A(n8776), .B(n4907), .ZN(n8777) );
  XNOR2_X1 U10415 ( .A(n8778), .B(n8777), .ZN(n8787) );
  NAND2_X1 U10416 ( .A1(n9249), .A2(n8779), .ZN(n8781) );
  AOI22_X1 U10417 ( .A1(n9251), .A2(n8797), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8780) );
  OAI211_X1 U10418 ( .C1(n9026), .C2(n8782), .A(n8781), .B(n8780), .ZN(n8783)
         );
  AOI21_X1 U10419 ( .B1(n9463), .B2(n8784), .A(n8783), .ZN(n8785) );
  OAI21_X1 U10420 ( .B1(n8787), .B2(n8786), .A(n8785), .ZN(P2_U3180) );
  INV_X1 U10421 ( .A(n9521), .ZN(n8801) );
  AND2_X1 U10422 ( .A1(n8650), .A2(n8788), .ZN(n8792) );
  OAI211_X1 U10423 ( .C1(n8792), .C2(n8791), .A(n8790), .B(n8789), .ZN(n8799)
         );
  NAND2_X1 U10424 ( .A1(n8793), .A2(n9383), .ZN(n8794) );
  NAND2_X1 U10425 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9105) );
  OAI211_X1 U10426 ( .C1(n9359), .C2(n8795), .A(n8794), .B(n9105), .ZN(n8796)
         );
  AOI21_X1 U10427 ( .B1(n9387), .B2(n8797), .A(n8796), .ZN(n8798) );
  OAI211_X1 U10428 ( .C1(n8801), .C2(n8800), .A(n8799), .B(n8798), .ZN(
        P2_U3181) );
  NAND2_X1 U10429 ( .A1(n9527), .A2(n5624), .ZN(n8803) );
  NAND2_X1 U10430 ( .A1(n5757), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8802) );
  OR2_X1 U10431 ( .A1(n9010), .A2(n9219), .ZN(n8993) );
  NAND2_X1 U10432 ( .A1(n9533), .A2(n5624), .ZN(n8805) );
  NAND2_X1 U10433 ( .A1(n5906), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8804) );
  NAND2_X1 U10434 ( .A1(n8840), .A2(n8839), .ZN(n8807) );
  AND2_X1 U10435 ( .A1(n8807), .A2(n8806), .ZN(n9004) );
  INV_X1 U10436 ( .A(n8839), .ZN(n9024) );
  INV_X1 U10437 ( .A(n9009), .ZN(n8835) );
  INV_X1 U10438 ( .A(n8981), .ZN(n8808) );
  INV_X1 U10439 ( .A(n8847), .ZN(n8809) );
  NAND2_X1 U10440 ( .A1(n8845), .A2(n8843), .ZN(n9280) );
  INV_X1 U10441 ( .A(n8810), .ZN(n8831) );
  INV_X1 U10442 ( .A(n8811), .ZN(n9369) );
  NAND4_X1 U10443 ( .A1(n8815), .A2(n8814), .A3(n8813), .A4(n8812), .ZN(n8818)
         );
  NAND4_X1 U10444 ( .A1(n8816), .A2(n8882), .A3(n4635), .A4(n8901), .ZN(n8817)
         );
  NOR2_X1 U10445 ( .A1(n8818), .A2(n8817), .ZN(n8822) );
  AND4_X1 U10446 ( .A1(n8822), .A2(n7113), .A3(n8821), .A4(n8820), .ZN(n8824)
         );
  NAND4_X1 U10447 ( .A1(n8825), .A2(n8824), .A3(n8823), .A4(n8919), .ZN(n8826)
         );
  NOR2_X1 U10448 ( .A1(n8932), .A2(n8826), .ZN(n8828) );
  NAND3_X1 U10449 ( .A1(n9369), .A2(n8828), .A3(n8827), .ZN(n8829) );
  NOR2_X1 U10450 ( .A1(n9355), .A2(n8829), .ZN(n8830) );
  NAND4_X1 U10451 ( .A1(n8831), .A2(n9343), .A3(n9330), .A4(n8830), .ZN(n8832)
         );
  NOR3_X1 U10452 ( .A1(n9280), .A2(n9302), .A3(n8832), .ZN(n8833) );
  NAND3_X1 U10453 ( .A1(n9267), .A2(n8833), .A3(n9290), .ZN(n8834) );
  AND4_X1 U10454 ( .A1(n8835), .A2(n4495), .A3(n9007), .A4(n9234), .ZN(n8838)
         );
  NAND4_X1 U10455 ( .A1(n8993), .A2(n9004), .A3(n8838), .A4(n9225), .ZN(n8842)
         );
  NAND3_X1 U10456 ( .A1(n8840), .A2(n8839), .A3(n8991), .ZN(n8841) );
  NAND3_X1 U10457 ( .A1(n8842), .A2(n7104), .A3(n8841), .ZN(n8998) );
  MUX2_X1 U10458 ( .A(n9237), .B(n9456), .S(n8999), .Z(n8986) );
  OR2_X1 U10459 ( .A1(n8970), .A2(n8999), .ZN(n8973) );
  OR2_X1 U10460 ( .A1(n8843), .A2(n8999), .ZN(n8844) );
  OAI21_X1 U10461 ( .B1(n8845), .B2(n8991), .A(n8844), .ZN(n8846) );
  NOR2_X1 U10462 ( .A1(n8847), .A2(n8846), .ZN(n8848) );
  NAND4_X1 U10463 ( .A1(n8973), .A2(n8848), .A3(n8975), .A4(n8971), .ZN(n8969)
         );
  NAND2_X1 U10464 ( .A1(n8849), .A2(n8999), .ZN(n8850) );
  NOR2_X1 U10465 ( .A1(n8810), .A2(n8850), .ZN(n8959) );
  MUX2_X1 U10466 ( .A(n8854), .B(n8851), .S(n8991), .Z(n8852) );
  NAND2_X1 U10467 ( .A1(n8852), .A2(n7113), .ZN(n8884) );
  AND2_X1 U10468 ( .A1(n8854), .A2(n8853), .ZN(n8856) );
  OAI211_X1 U10469 ( .C1(n8884), .C2(n8856), .A(n8855), .B(n8912), .ZN(n8857)
         );
  NAND2_X1 U10470 ( .A1(n8857), .A2(n8991), .ZN(n8862) );
  OAI21_X1 U10471 ( .B1(n8884), .B2(n8859), .A(n8858), .ZN(n8860) );
  NAND2_X1 U10472 ( .A1(n8860), .A2(n8999), .ZN(n8861) );
  AND2_X1 U10473 ( .A1(n8861), .A2(n8862), .ZN(n8910) );
  NAND2_X1 U10474 ( .A1(n7107), .A2(n8863), .ZN(n8866) );
  INV_X1 U10475 ( .A(n8870), .ZN(n8864) );
  NAND3_X1 U10476 ( .A1(n8864), .A2(n8991), .A3(n7896), .ZN(n8865) );
  OAI21_X1 U10477 ( .B1(n8867), .B2(n8866), .A(n8865), .ZN(n8881) );
  AOI21_X1 U10478 ( .B1(n4404), .B2(n8999), .A(n4730), .ZN(n8873) );
  AOI21_X1 U10479 ( .B1(n10538), .B2(n8991), .A(n8868), .ZN(n8872) );
  NAND3_X1 U10480 ( .A1(n8870), .A2(n8869), .A3(n7107), .ZN(n8871) );
  OAI211_X1 U10481 ( .C1(n8873), .C2(n8872), .A(n4635), .B(n8871), .ZN(n8880)
         );
  NAND2_X1 U10482 ( .A1(n8890), .A2(n7108), .ZN(n8877) );
  NAND2_X1 U10483 ( .A1(n8875), .A2(n8874), .ZN(n8876) );
  MUX2_X1 U10484 ( .A(n8877), .B(n8876), .S(n8991), .Z(n8878) );
  INV_X1 U10485 ( .A(n8878), .ZN(n8879) );
  OAI21_X1 U10486 ( .B1(n8881), .B2(n8880), .A(n8879), .ZN(n8883) );
  NAND2_X1 U10487 ( .A1(n8883), .A2(n8882), .ZN(n8894) );
  INV_X1 U10488 ( .A(n8884), .ZN(n8906) );
  NAND2_X1 U10489 ( .A1(n8895), .A2(n8885), .ZN(n8902) );
  INV_X1 U10490 ( .A(n8902), .ZN(n8887) );
  AND4_X1 U10491 ( .A1(n8901), .A2(n8887), .A3(n8999), .A4(n8886), .ZN(n8888)
         );
  OAI211_X1 U10492 ( .C1(n8894), .C2(n8889), .A(n8906), .B(n8888), .ZN(n8909)
         );
  INV_X1 U10493 ( .A(n8890), .ZN(n8893) );
  AND4_X1 U10494 ( .A1(n8901), .A2(n8991), .A3(n8891), .A4(n8897), .ZN(n8892)
         );
  OAI211_X1 U10495 ( .C1(n8894), .C2(n8893), .A(n8906), .B(n8892), .ZN(n8908)
         );
  NAND2_X1 U10496 ( .A1(n7112), .A2(n8999), .ZN(n8900) );
  NAND3_X1 U10497 ( .A1(n8897), .A2(n8896), .A3(n8999), .ZN(n8899) );
  OR2_X1 U10498 ( .A1(n8897), .A2(n8999), .ZN(n8898) );
  NAND4_X1 U10499 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n8898), .ZN(n8904)
         );
  NOR2_X1 U10500 ( .A1(n8902), .A2(n8999), .ZN(n8903) );
  NOR2_X1 U10501 ( .A1(n8904), .A2(n8903), .ZN(n8905) );
  NAND2_X1 U10502 ( .A1(n8906), .A2(n8905), .ZN(n8907) );
  NAND4_X1 U10503 ( .A1(n8910), .A2(n8909), .A3(n8908), .A4(n8907), .ZN(n8915)
         );
  NAND3_X1 U10504 ( .A1(n8915), .A2(n8912), .A3(n7115), .ZN(n8913) );
  NAND2_X1 U10505 ( .A1(n8915), .A2(n8914), .ZN(n8918) );
  INV_X1 U10506 ( .A(n8916), .ZN(n8917) );
  NAND2_X1 U10507 ( .A1(n8921), .A2(n8920), .ZN(n8922) );
  MUX2_X1 U10508 ( .A(n8923), .B(n8922), .S(n8999), .Z(n8924) );
  MUX2_X1 U10509 ( .A(n8926), .B(n8925), .S(n8991), .Z(n8929) );
  NAND2_X1 U10510 ( .A1(n8929), .A2(n8927), .ZN(n8931) );
  NOR2_X1 U10511 ( .A1(n8929), .A2(n8928), .ZN(n8930) );
  INV_X1 U10512 ( .A(n8932), .ZN(n9378) );
  NAND2_X1 U10513 ( .A1(n8934), .A2(n8933), .ZN(n8935) );
  MUX2_X1 U10514 ( .A(n8936), .B(n8935), .S(n8999), .Z(n8937) );
  OAI211_X1 U10515 ( .C1(n8939), .C2(n8938), .A(n9378), .B(n8937), .ZN(n8944)
         );
  AND2_X1 U10516 ( .A1(n8945), .A2(n8940), .ZN(n8941) );
  MUX2_X1 U10517 ( .A(n8942), .B(n8941), .S(n8991), .Z(n8943) );
  INV_X1 U10518 ( .A(n9355), .ZN(n9353) );
  INV_X1 U10519 ( .A(n8945), .ZN(n8947) );
  INV_X1 U10520 ( .A(n8948), .ZN(n8954) );
  NAND2_X1 U10521 ( .A1(n9311), .A2(n8991), .ZN(n8956) );
  NAND2_X1 U10522 ( .A1(n8950), .A2(n8949), .ZN(n8951) );
  NOR2_X1 U10523 ( .A1(n8956), .A2(n8951), .ZN(n8952) );
  INV_X1 U10524 ( .A(n8955), .ZN(n8958) );
  INV_X1 U10525 ( .A(n8956), .ZN(n8957) );
  NAND2_X1 U10526 ( .A1(n8963), .A2(n8960), .ZN(n8961) );
  NAND2_X1 U10527 ( .A1(n8961), .A2(n8999), .ZN(n8962) );
  MUX2_X1 U10528 ( .A(n8964), .B(n8963), .S(n8991), .Z(n8965) );
  NAND2_X1 U10529 ( .A1(n9291), .A2(n9304), .ZN(n8967) );
  MUX2_X1 U10530 ( .A(n9304), .B(n9291), .S(n8991), .Z(n8966) );
  OAI21_X1 U10531 ( .B1(n8999), .B2(n8971), .A(n8970), .ZN(n8972) );
  NAND2_X1 U10532 ( .A1(n8973), .A2(n8972), .ZN(n8978) );
  NAND4_X1 U10533 ( .A1(n8975), .A2(n8974), .A3(n8999), .A4(n9475), .ZN(n8977)
         );
  OR2_X1 U10534 ( .A1(n8975), .A2(n8999), .ZN(n8976) );
  INV_X1 U10535 ( .A(n8979), .ZN(n8980) );
  MUX2_X1 U10536 ( .A(n8981), .B(n8980), .S(n8999), .Z(n8982) );
  MUX2_X1 U10537 ( .A(n9249), .B(n9398), .S(n8999), .Z(n8983) );
  OR2_X1 U10538 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  OAI21_X1 U10539 ( .B1(n9003), .B2(n9237), .A(n9004), .ZN(n8990) );
  NOR3_X1 U10540 ( .A1(n8988), .A2(n4836), .A3(n8987), .ZN(n8989) );
  INV_X1 U10541 ( .A(n8993), .ZN(n8995) );
  INV_X1 U10542 ( .A(n9007), .ZN(n9000) );
  NOR3_X1 U10543 ( .A1(n9009), .A2(n9000), .A3(n8999), .ZN(n9001) );
  OAI211_X1 U10544 ( .C1(n9456), .C2(n9003), .A(n9002), .B(n9001), .ZN(n9014)
         );
  INV_X1 U10545 ( .A(n9004), .ZN(n9006) );
  AOI21_X1 U10546 ( .B1(n9453), .B2(n9219), .A(n9010), .ZN(n9005) );
  OAI22_X1 U10547 ( .A1(n9012), .A2(n7104), .B1(n9450), .B2(n9011), .ZN(n9013)
         );
  AOI21_X1 U10548 ( .B1(n9015), .B2(n9014), .A(n9013), .ZN(n9016) );
  XNOR2_X1 U10549 ( .A(n9016), .B(n5743), .ZN(n9023) );
  NAND3_X1 U10550 ( .A1(n9018), .A2(n9017), .A3(n4402), .ZN(n9019) );
  OAI211_X1 U10551 ( .C1(n9020), .C2(n9022), .A(n9019), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9021) );
  OAI21_X1 U10552 ( .B1(n9023), .B2(n9022), .A(n9021), .ZN(P2_U3296) );
  MUX2_X1 U10553 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9024), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10554 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n9227), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10555 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9237), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10556 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9249), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10557 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n4907), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10558 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9268), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10559 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n5874), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10560 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n9269), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10561 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9304), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10562 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9345), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10563 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9027), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10564 ( .A(n9371), .B(P2_DATAO_REG_17__SCAN_IN), .S(n9036), .Z(
        P2_U3508) );
  MUX2_X1 U10565 ( .A(n9381), .B(P2_DATAO_REG_16__SCAN_IN), .S(n9036), .Z(
        P2_U3507) );
  MUX2_X1 U10566 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9370), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10567 ( .A(n9383), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9036), .Z(
        P2_U3505) );
  MUX2_X1 U10568 ( .A(n9028), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9036), .Z(
        P2_U3503) );
  MUX2_X1 U10569 ( .A(n9029), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9036), .Z(
        P2_U3502) );
  MUX2_X1 U10570 ( .A(n9030), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9036), .Z(
        P2_U3501) );
  MUX2_X1 U10571 ( .A(n9031), .B(P2_DATAO_REG_9__SCAN_IN), .S(n9036), .Z(
        P2_U3500) );
  MUX2_X1 U10572 ( .A(n9032), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9036), .Z(
        P2_U3499) );
  MUX2_X1 U10573 ( .A(n9033), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9036), .Z(
        P2_U3498) );
  MUX2_X1 U10574 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n7111), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10575 ( .A(n9034), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9036), .Z(
        P2_U3496) );
  MUX2_X1 U10576 ( .A(n7110), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9036), .Z(
        P2_U3495) );
  MUX2_X1 U10577 ( .A(n9035), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9036), .Z(
        P2_U3494) );
  MUX2_X1 U10578 ( .A(n7057), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9036), .Z(
        P2_U3493) );
  MUX2_X1 U10579 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n4404), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10580 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n7529), .S(P2_U3893), .Z(
        P2_U3491) );
  INV_X1 U10581 ( .A(n9066), .ZN(n9041) );
  AOI21_X1 U10582 ( .B1(n9045), .B2(n9042), .A(n9041), .ZN(n9065) );
  OAI21_X1 U10583 ( .B1(n9154), .B2(n9084), .A(n9043), .ZN(n9056) );
  NAND2_X1 U10584 ( .A1(n9053), .A2(n9052), .ZN(n9049) );
  MUX2_X1 U10585 ( .A(n9045), .B(n9044), .S(n4401), .Z(n9046) );
  NAND2_X1 U10586 ( .A1(n9046), .A2(n9060), .ZN(n9078) );
  INV_X1 U10587 ( .A(n9046), .ZN(n9047) );
  NAND2_X1 U10588 ( .A1(n9047), .A2(n9084), .ZN(n9048) );
  AND2_X1 U10589 ( .A1(n9078), .A2(n9048), .ZN(n9050) );
  INV_X1 U10590 ( .A(n9050), .ZN(n9051) );
  NAND3_X1 U10591 ( .A1(n9053), .A2(n9052), .A3(n9051), .ZN(n9054) );
  AOI21_X1 U10592 ( .B1(n9079), .B2(n9054), .A(n9159), .ZN(n9055) );
  AOI211_X1 U10593 ( .C1(n9210), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n9056), .B(
        n9055), .ZN(n9064) );
  NAND2_X1 U10594 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n9057), .ZN(n9059) );
  NAND2_X1 U10595 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9061), .ZN(n9085) );
  OAI21_X1 U10596 ( .B1(n9061), .B2(P2_REG1_REG_13__SCAN_IN), .A(n9085), .ZN(
        n9062) );
  NAND2_X1 U10597 ( .A1(n9062), .A2(n9173), .ZN(n9063) );
  OAI211_X1 U10598 ( .C1(n9065), .C2(n9217), .A(n9064), .B(n9063), .ZN(
        P2_U3195) );
  XNOR2_X1 U10599 ( .A(n9102), .B(n9071), .ZN(n9068) );
  AND3_X1 U10600 ( .A1(n9066), .A2(n9068), .A3(n9067), .ZN(n9069) );
  OAI21_X1 U10601 ( .B1(n9093), .B2(n9069), .A(n9146), .ZN(n9092) );
  OAI21_X1 U10602 ( .B1(n9154), .B2(n9094), .A(n9070), .ZN(n9082) );
  NAND2_X1 U10603 ( .A1(n9079), .A2(n9078), .ZN(n9075) );
  MUX2_X1 U10604 ( .A(n9071), .B(n9101), .S(n4402), .Z(n9072) );
  NAND2_X1 U10605 ( .A1(n9072), .A2(n9102), .ZN(n9096) );
  INV_X1 U10606 ( .A(n9072), .ZN(n9073) );
  NAND2_X1 U10607 ( .A1(n9073), .A2(n9094), .ZN(n9074) );
  AND2_X1 U10608 ( .A1(n9096), .A2(n9074), .ZN(n9076) );
  INV_X1 U10609 ( .A(n9076), .ZN(n9077) );
  NAND3_X1 U10610 ( .A1(n9079), .A2(n9078), .A3(n9077), .ZN(n9080) );
  AOI21_X1 U10611 ( .B1(n9097), .B2(n9080), .A(n9159), .ZN(n9081) );
  AOI211_X1 U10612 ( .C1(n9210), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n9082), .B(
        n9081), .ZN(n9091) );
  NAND2_X1 U10613 ( .A1(n9084), .A2(n9083), .ZN(n9086) );
  XNOR2_X1 U10614 ( .A(n9102), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n9087) );
  OAI21_X1 U10615 ( .B1(n9088), .B2(n9087), .A(n9103), .ZN(n9089) );
  NAND2_X1 U10616 ( .A1(n9089), .A2(n9173), .ZN(n9090) );
  NAND3_X1 U10617 ( .A1(n9092), .A2(n9091), .A3(n9090), .ZN(P2_U3196) );
  OAI21_X1 U10618 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n9095), .A(n9122), .ZN(
        n9112) );
  MUX2_X1 U10619 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n4402), .Z(n9114) );
  XNOR2_X1 U10620 ( .A(n9114), .B(n9115), .ZN(n9098) );
  NAND2_X1 U10621 ( .A1(n9099), .A2(n9098), .ZN(n9118) );
  OAI21_X1 U10622 ( .B1(n9099), .B2(n9098), .A(n9118), .ZN(n9100) );
  NAND2_X1 U10623 ( .A1(n9100), .A2(n9215), .ZN(n9109) );
  OR2_X1 U10624 ( .A1(n9102), .A2(n9101), .ZN(n9104) );
  XNOR2_X1 U10625 ( .A(n9127), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n9107) );
  OAI21_X1 U10626 ( .B1(n9154), .B2(n5173), .A(n9105), .ZN(n9106) );
  AOI21_X1 U10627 ( .B1(n9173), .B2(n9107), .A(n9106), .ZN(n9108) );
  OAI211_X1 U10628 ( .C1(n9171), .C2(n9110), .A(n9109), .B(n9108), .ZN(n9111)
         );
  AOI21_X1 U10629 ( .B1(n9112), .B2(n9146), .A(n9111), .ZN(n9113) );
  INV_X1 U10630 ( .A(n9113), .ZN(P2_U3197) );
  INV_X1 U10631 ( .A(n9114), .ZN(n9116) );
  NAND2_X1 U10632 ( .A1(n9116), .A2(n9115), .ZN(n9117) );
  MUX2_X1 U10633 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n4402), .Z(n9120) );
  INV_X1 U10634 ( .A(n9120), .ZN(n9119) );
  NAND2_X1 U10635 ( .A1(n9119), .A2(n9148), .ZN(n9140) );
  NAND2_X1 U10636 ( .A1(n9120), .A2(n9142), .ZN(n9138) );
  NAND2_X1 U10637 ( .A1(n9140), .A2(n9138), .ZN(n9121) );
  XNOR2_X1 U10638 ( .A(n9139), .B(n9121), .ZN(n9137) );
  NAND2_X1 U10639 ( .A1(n9122), .A2(n4465), .ZN(n9124) );
  XNOR2_X1 U10640 ( .A(n9148), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n9123) );
  NOR2_X1 U10641 ( .A1(n9124), .A2(n9123), .ZN(n9125) );
  OAI21_X1 U10642 ( .B1(n9126), .B2(n9125), .A(n9146), .ZN(n9136) );
  NAND2_X1 U10643 ( .A1(n9127), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9130) );
  NAND2_X1 U10644 ( .A1(n5173), .A2(n9128), .ZN(n9129) );
  XNOR2_X1 U10645 ( .A(n9148), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n9150) );
  XNOR2_X1 U10646 ( .A(n9151), .B(n9150), .ZN(n9134) );
  NAND2_X1 U10647 ( .A1(n9210), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n9132) );
  OAI211_X1 U10648 ( .C1(n9142), .C2(n9154), .A(n9132), .B(n9131), .ZN(n9133)
         );
  AOI21_X1 U10649 ( .B1(n9173), .B2(n9134), .A(n9133), .ZN(n9135) );
  OAI211_X1 U10650 ( .C1(n9159), .C2(n9137), .A(n9136), .B(n9135), .ZN(
        P2_U3198) );
  MUX2_X1 U10651 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n4402), .Z(n9175) );
  XNOR2_X1 U10652 ( .A(n9175), .B(n9176), .ZN(n9179) );
  NAND2_X1 U10653 ( .A1(n9139), .A2(n9138), .ZN(n9141) );
  NAND2_X1 U10654 ( .A1(n9141), .A2(n9140), .ZN(n9180) );
  XOR2_X1 U10655 ( .A(n9179), .B(n9180), .Z(n9160) );
  NAND2_X1 U10656 ( .A1(n9145), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9165) );
  OAI21_X1 U10657 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n9145), .A(n9165), .ZN(
        n9147) );
  NAND2_X1 U10658 ( .A1(n9147), .A2(n9146), .ZN(n9158) );
  INV_X1 U10659 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9434) );
  NOR2_X1 U10660 ( .A1(n9148), .A2(n9434), .ZN(n9149) );
  XOR2_X1 U10661 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9169), .Z(n9156) );
  NAND2_X1 U10662 ( .A1(n9210), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n9153) );
  OAI211_X1 U10663 ( .C1(n9154), .C2(n5166), .A(n9153), .B(n9152), .ZN(n9155)
         );
  AOI21_X1 U10664 ( .B1(n9173), .B2(n9156), .A(n9155), .ZN(n9157) );
  OAI211_X1 U10665 ( .C1(n9160), .C2(n9159), .A(n9158), .B(n9157), .ZN(
        P2_U3199) );
  INV_X1 U10666 ( .A(n9161), .ZN(n9164) );
  INV_X1 U10667 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9347) );
  OR2_X1 U10668 ( .A1(n9187), .A2(n9347), .ZN(n9192) );
  NAND2_X1 U10669 ( .A1(n9187), .A2(n9347), .ZN(n9162) );
  NAND2_X1 U10670 ( .A1(n9192), .A2(n9162), .ZN(n9163) );
  AND3_X1 U10671 ( .A1(n9165), .A2(n9164), .A3(n9163), .ZN(n9166) );
  OAI22_X1 U10672 ( .A1(n9169), .A2(n9168), .B1(n9176), .B2(n9167), .ZN(n9205)
         );
  XNOR2_X1 U10673 ( .A(n9187), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n9204) );
  XNOR2_X1 U10674 ( .A(n9205), .B(n9204), .ZN(n9174) );
  INV_X1 U10675 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10587) );
  OAI21_X1 U10676 ( .B1(n9171), .B2(n10587), .A(n9170), .ZN(n9172) );
  AOI21_X1 U10677 ( .B1(n9174), .B2(n9173), .A(n9172), .ZN(n9191) );
  INV_X1 U10678 ( .A(n9175), .ZN(n9177) );
  AND2_X1 U10679 ( .A1(n9177), .A2(n9176), .ZN(n9178) );
  MUX2_X1 U10680 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n4402), .Z(n9183) );
  AND2_X1 U10681 ( .A1(n9182), .A2(n9183), .ZN(n9195) );
  INV_X1 U10682 ( .A(n9196), .ZN(n9184) );
  INV_X1 U10683 ( .A(n9186), .ZN(n9185) );
  NAND2_X1 U10684 ( .A1(n9185), .A2(n9215), .ZN(n9189) );
  INV_X1 U10685 ( .A(n9192), .ZN(n9193) );
  XNOR2_X1 U10686 ( .A(n5743), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n9200) );
  AOI21_X1 U10687 ( .B1(n9203), .B2(n9196), .A(n9195), .ZN(n9202) );
  MUX2_X1 U10688 ( .A(n9206), .B(n9200), .S(n9199), .Z(n9201) );
  XNOR2_X1 U10689 ( .A(n9202), .B(n9201), .ZN(n9216) );
  XNOR2_X1 U10690 ( .A(n9207), .B(n9206), .ZN(n9214) );
  AOI21_X1 U10691 ( .B1(n9209), .B2(n5743), .A(n9208), .ZN(n9212) );
  NAND2_X1 U10692 ( .A1(n9210), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n9211) );
  AOI21_X1 U10693 ( .B1(n9448), .B2(n9220), .A(n10550), .ZN(n9222) );
  AOI21_X1 U10694 ( .B1(n10550), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9222), .ZN(
        n9221) );
  OAI21_X1 U10695 ( .B1(n9450), .B2(n9362), .A(n9221), .ZN(P2_U3202) );
  AOI21_X1 U10696 ( .B1(n10550), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9222), .ZN(
        n9223) );
  OAI21_X1 U10697 ( .B1(n9453), .B2(n9362), .A(n9223), .ZN(P2_U3203) );
  XNOR2_X1 U10698 ( .A(n9224), .B(n9225), .ZN(n9459) );
  INV_X1 U10699 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9228) );
  AOI22_X1 U10700 ( .A1(n9456), .A2(n4398), .B1(n9388), .B2(n9229), .ZN(n9230)
         );
  OAI21_X1 U10701 ( .B1(n9232), .B2(n9234), .A(n9231), .ZN(n9401) );
  INV_X1 U10702 ( .A(n9233), .ZN(n9242) );
  XNOR2_X1 U10703 ( .A(n9236), .B(n9235), .ZN(n9241) );
  AOI21_X2 U10704 ( .B1(n9241), .B2(n10541), .A(n9240), .ZN(n9400) );
  OAI21_X1 U10705 ( .B1(n9242), .B2(n10533), .A(n9400), .ZN(n9243) );
  NAND2_X1 U10706 ( .A1(n9243), .A2(n9385), .ZN(n9245) );
  AOI22_X1 U10707 ( .A1(n9398), .A2(n4398), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n10550), .ZN(n9244) );
  OAI211_X1 U10708 ( .C1(n9401), .C2(n9366), .A(n9245), .B(n9244), .ZN(
        P2_U3206) );
  XNOR2_X1 U10709 ( .A(n9246), .B(n9248), .ZN(n9466) );
  INV_X1 U10710 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9250) );
  MUX2_X1 U10711 ( .A(n9250), .B(n9461), .S(n9385), .Z(n9253) );
  AOI22_X1 U10712 ( .A1(n9463), .A2(n4398), .B1(n9388), .B2(n9251), .ZN(n9252)
         );
  OAI211_X1 U10713 ( .C1(n9466), .C2(n9366), .A(n9253), .B(n9252), .ZN(
        P2_U3207) );
  XOR2_X1 U10714 ( .A(n9254), .B(n9255), .Z(n9472) );
  XNOR2_X1 U10715 ( .A(n9256), .B(n9255), .ZN(n9257) );
  AOI222_X1 U10716 ( .A1(n10541), .A2(n9257), .B1(n5874), .B2(n9382), .C1(
        n4907), .C2(n9380), .ZN(n9467) );
  INV_X1 U10717 ( .A(n9467), .ZN(n9262) );
  INV_X1 U10718 ( .A(n9258), .ZN(n9259) );
  OAI22_X1 U10719 ( .A1(n9260), .A2(n10531), .B1(n9259), .B2(n10533), .ZN(
        n9261) );
  OAI21_X1 U10720 ( .B1(n9262), .B2(n9261), .A(n9385), .ZN(n9264) );
  NAND2_X1 U10721 ( .A1(n10550), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9263) );
  OAI211_X1 U10722 ( .C1(n9472), .C2(n9366), .A(n9264), .B(n9263), .ZN(
        P2_U3208) );
  XOR2_X1 U10723 ( .A(n9265), .B(n9267), .Z(n9478) );
  XOR2_X1 U10724 ( .A(n9267), .B(n9266), .Z(n9270) );
  AOI222_X1 U10725 ( .A1(n10541), .A2(n9270), .B1(n9269), .B2(n9382), .C1(
        n9268), .C2(n9380), .ZN(n9473) );
  INV_X1 U10726 ( .A(n9473), .ZN(n9275) );
  INV_X1 U10727 ( .A(n9271), .ZN(n9272) );
  OAI22_X1 U10728 ( .A1(n9273), .A2(n10531), .B1(n9272), .B2(n10533), .ZN(
        n9274) );
  OAI21_X1 U10729 ( .B1(n9275), .B2(n9274), .A(n9385), .ZN(n9277) );
  NAND2_X1 U10730 ( .A1(n10550), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9276) );
  OAI211_X1 U10731 ( .C1(n9478), .C2(n9366), .A(n9277), .B(n9276), .ZN(
        P2_U3209) );
  XNOR2_X1 U10732 ( .A(n9278), .B(n9280), .ZN(n9484) );
  INV_X1 U10733 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9282) );
  XNOR2_X1 U10734 ( .A(n9279), .B(n9280), .ZN(n9281) );
  AOI222_X1 U10735 ( .A1(n10541), .A2(n9281), .B1(n9304), .B2(n9382), .C1(
        n5874), .C2(n9380), .ZN(n9479) );
  MUX2_X1 U10736 ( .A(n9282), .B(n9479), .S(n9385), .Z(n9285) );
  AOI22_X1 U10737 ( .A1(n9481), .A2(n4398), .B1(n9388), .B2(n9283), .ZN(n9284)
         );
  OAI211_X1 U10738 ( .C1(n9484), .C2(n9366), .A(n9285), .B(n9284), .ZN(
        P2_U3210) );
  XOR2_X1 U10739 ( .A(n9290), .B(n9286), .Z(n9287) );
  OAI222_X1 U10740 ( .A1(n10539), .A2(n9288), .B1(n10537), .B2(n9317), .C1(
        n9287), .C2(n9356), .ZN(n9414) );
  INV_X1 U10741 ( .A(n9414), .ZN(n9297) );
  XNOR2_X1 U10742 ( .A(n9289), .B(n9290), .ZN(n9415) );
  INV_X1 U10743 ( .A(n9291), .ZN(n9488) );
  AOI22_X1 U10744 ( .A1(n9292), .A2(n9388), .B1(P2_REG2_REG_22__SCAN_IN), .B2(
        n10550), .ZN(n9293) );
  OAI21_X1 U10745 ( .B1(n9488), .B2(n9362), .A(n9293), .ZN(n9294) );
  AOI21_X1 U10746 ( .B1(n9415), .B2(n9295), .A(n9294), .ZN(n9296) );
  OAI21_X1 U10747 ( .B1(n9297), .B2(n10550), .A(n9296), .ZN(P2_U3211) );
  NAND2_X1 U10748 ( .A1(n9299), .A2(n9298), .ZN(n9300) );
  XOR2_X1 U10749 ( .A(n9302), .B(n9300), .Z(n9494) );
  XNOR2_X1 U10750 ( .A(n9303), .B(n9302), .ZN(n9306) );
  AOI222_X1 U10751 ( .A1(n10541), .A2(n9306), .B1(n9305), .B2(n9382), .C1(
        n9304), .C2(n9380), .ZN(n9489) );
  MUX2_X1 U10752 ( .A(n9307), .B(n9489), .S(n9385), .Z(n9310) );
  AOI22_X1 U10753 ( .A1(n9491), .A2(n4398), .B1(n9388), .B2(n9308), .ZN(n9309)
         );
  OAI211_X1 U10754 ( .C1(n9494), .C2(n9366), .A(n9310), .B(n9309), .ZN(
        P2_U3212) );
  NAND2_X1 U10755 ( .A1(n4442), .A2(n9343), .ZN(n9342) );
  NAND3_X1 U10756 ( .A1(n9342), .A2(n9330), .A3(n9326), .ZN(n9325) );
  NAND2_X1 U10757 ( .A1(n9325), .A2(n9311), .ZN(n9312) );
  XNOR2_X1 U10758 ( .A(n9312), .B(n8810), .ZN(n9498) );
  NAND2_X1 U10759 ( .A1(n9332), .A2(n9314), .ZN(n9315) );
  XNOR2_X1 U10760 ( .A(n9315), .B(n8810), .ZN(n9316) );
  OAI222_X1 U10761 ( .A1(n10537), .A2(n9318), .B1(n10539), .B2(n9317), .C1(
        n9316), .C2(n9356), .ZN(n9421) );
  NAND2_X1 U10762 ( .A1(n9421), .A2(n9385), .ZN(n9324) );
  INV_X1 U10763 ( .A(n9319), .ZN(n9321) );
  INV_X1 U10764 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9320) );
  OAI22_X1 U10765 ( .A1(n9321), .A2(n10533), .B1(n9385), .B2(n9320), .ZN(n9322) );
  AOI21_X1 U10766 ( .B1(n7088), .B2(n4398), .A(n9322), .ZN(n9323) );
  OAI211_X1 U10767 ( .C1(n9498), .C2(n9366), .A(n9324), .B(n9323), .ZN(
        P2_U3213) );
  INV_X1 U10768 ( .A(n9325), .ZN(n9328) );
  AOI21_X1 U10769 ( .B1(n9342), .B2(n9326), .A(n9330), .ZN(n9327) );
  NOR2_X1 U10770 ( .A1(n9328), .A2(n9327), .ZN(n9502) );
  AOI22_X1 U10771 ( .A1(n9329), .A2(n4398), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n10550), .ZN(n9341) );
  NAND2_X1 U10772 ( .A1(n9313), .A2(n9330), .ZN(n9331) );
  NAND3_X1 U10773 ( .A1(n9332), .A2(n10541), .A3(n9331), .ZN(n9336) );
  OAI22_X1 U10774 ( .A1(n9333), .A2(n10539), .B1(n9358), .B2(n10537), .ZN(
        n9334) );
  INV_X1 U10775 ( .A(n9334), .ZN(n9335) );
  NAND2_X1 U10776 ( .A1(n9336), .A2(n9335), .ZN(n9499) );
  INV_X1 U10777 ( .A(n9337), .ZN(n9338) );
  NOR2_X1 U10778 ( .A1(n9338), .A2(n10533), .ZN(n9339) );
  OAI21_X1 U10779 ( .B1(n9499), .B2(n9339), .A(n9385), .ZN(n9340) );
  OAI211_X1 U10780 ( .C1(n9502), .C2(n9366), .A(n9341), .B(n9340), .ZN(
        P2_U3214) );
  OAI21_X1 U10781 ( .B1(n4442), .B2(n9343), .A(n9342), .ZN(n9510) );
  XNOR2_X1 U10782 ( .A(n9344), .B(n9343), .ZN(n9346) );
  AOI222_X1 U10783 ( .A1(n10541), .A2(n9346), .B1(n9371), .B2(n9382), .C1(
        n9345), .C2(n9380), .ZN(n9505) );
  MUX2_X1 U10784 ( .A(n9347), .B(n9505), .S(n9385), .Z(n9350) );
  AOI22_X1 U10785 ( .A1(n9507), .A2(n4398), .B1(n9388), .B2(n9348), .ZN(n9349)
         );
  OAI211_X1 U10786 ( .C1(n9510), .C2(n9366), .A(n9350), .B(n9349), .ZN(
        P2_U3215) );
  XNOR2_X1 U10787 ( .A(n9352), .B(n9353), .ZN(n9433) );
  XNOR2_X1 U10788 ( .A(n9354), .B(n9355), .ZN(n9357) );
  OAI222_X1 U10789 ( .A1(n10537), .A2(n9359), .B1(n10539), .B2(n9358), .C1(
        n9357), .C2(n9356), .ZN(n9430) );
  AOI22_X1 U10790 ( .A1(n10550), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9388), 
        .B2(n9360), .ZN(n9361) );
  OAI21_X1 U10791 ( .B1(n9363), .B2(n9362), .A(n9361), .ZN(n9364) );
  AOI21_X1 U10792 ( .B1(n9430), .B2(n9385), .A(n9364), .ZN(n9365) );
  OAI21_X1 U10793 ( .B1(n9433), .B2(n9366), .A(n9365), .ZN(P2_U3216) );
  XNOR2_X1 U10794 ( .A(n9367), .B(n9369), .ZN(n9517) );
  XNOR2_X1 U10795 ( .A(n9368), .B(n9369), .ZN(n9372) );
  AOI222_X1 U10796 ( .A1(n10541), .A2(n9372), .B1(n9371), .B2(n9380), .C1(
        n9370), .C2(n9382), .ZN(n9512) );
  MUX2_X1 U10797 ( .A(n9373), .B(n9512), .S(n9385), .Z(n9376) );
  AOI22_X1 U10798 ( .A1(n9514), .A2(n4398), .B1(n9388), .B2(n9374), .ZN(n9375)
         );
  OAI211_X1 U10799 ( .C1(n9517), .C2(n9366), .A(n9376), .B(n9375), .ZN(
        P2_U3217) );
  XNOR2_X1 U10800 ( .A(n9377), .B(n9378), .ZN(n9525) );
  INV_X1 U10801 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9386) );
  XNOR2_X1 U10802 ( .A(n9379), .B(n9378), .ZN(n9384) );
  AOI222_X1 U10803 ( .A1(n10541), .A2(n9384), .B1(n9383), .B2(n9382), .C1(
        n9381), .C2(n9380), .ZN(n9518) );
  MUX2_X1 U10804 ( .A(n9386), .B(n9518), .S(n9385), .Z(n9391) );
  AOI22_X1 U10805 ( .A1(n9521), .A2(n4398), .B1(n9388), .B2(n9387), .ZN(n9390)
         );
  OAI211_X1 U10806 ( .C1(n9525), .C2(n9366), .A(n9391), .B(n9390), .ZN(
        P2_U3218) );
  NOR2_X1 U10807 ( .A1(n9448), .A2(n7168), .ZN(n9393) );
  AOI21_X1 U10808 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n7168), .A(n9393), .ZN(
        n9392) );
  OAI21_X1 U10809 ( .B1(n9450), .B2(n9424), .A(n9392), .ZN(P2_U3490) );
  AOI21_X1 U10810 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n7168), .A(n9393), .ZN(
        n9394) );
  OAI21_X1 U10811 ( .B1(n9453), .B2(n9424), .A(n9394), .ZN(P2_U3489) );
  NAND2_X1 U10812 ( .A1(n9456), .A2(n9438), .ZN(n9396) );
  OAI211_X1 U10813 ( .C1(n9459), .C2(n9441), .A(n9397), .B(n9396), .ZN(
        P2_U3487) );
  NAND2_X1 U10814 ( .A1(n9398), .A2(n9443), .ZN(n9399) );
  OAI211_X1 U10815 ( .C1(n10567), .C2(n9401), .A(n9400), .B(n9399), .ZN(n9460)
         );
  MUX2_X1 U10816 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9460), .S(n10578), .Z(
        P2_U3486) );
  INV_X1 U10817 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9402) );
  MUX2_X1 U10818 ( .A(n9402), .B(n9461), .S(n10578), .Z(n9404) );
  NAND2_X1 U10819 ( .A1(n9463), .A2(n9438), .ZN(n9403) );
  OAI211_X1 U10820 ( .C1(n9441), .C2(n9466), .A(n9404), .B(n9403), .ZN(
        P2_U3485) );
  MUX2_X1 U10821 ( .A(n9405), .B(n9467), .S(n10578), .Z(n9407) );
  NAND2_X1 U10822 ( .A1(n9469), .A2(n9438), .ZN(n9406) );
  OAI211_X1 U10823 ( .C1(n9472), .C2(n9441), .A(n9407), .B(n9406), .ZN(
        P2_U3484) );
  INV_X1 U10824 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9408) );
  MUX2_X1 U10825 ( .A(n9408), .B(n9473), .S(n10578), .Z(n9410) );
  NAND2_X1 U10826 ( .A1(n9475), .A2(n9438), .ZN(n9409) );
  OAI211_X1 U10827 ( .C1(n9441), .C2(n9478), .A(n9410), .B(n9409), .ZN(
        P2_U3483) );
  MUX2_X1 U10828 ( .A(n9411), .B(n9479), .S(n10578), .Z(n9413) );
  NAND2_X1 U10829 ( .A1(n9481), .A2(n9438), .ZN(n9412) );
  OAI211_X1 U10830 ( .C1(n9441), .C2(n9484), .A(n9413), .B(n9412), .ZN(
        P2_U3482) );
  AOI21_X1 U10831 ( .B1(n10562), .B2(n9415), .A(n9414), .ZN(n9485) );
  MUX2_X1 U10832 ( .A(n9416), .B(n9485), .S(n10578), .Z(n9417) );
  OAI21_X1 U10833 ( .B1(n9488), .B2(n9424), .A(n9417), .ZN(P2_U3481) );
  INV_X1 U10834 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9418) );
  MUX2_X1 U10835 ( .A(n9418), .B(n9489), .S(n10578), .Z(n9420) );
  NAND2_X1 U10836 ( .A1(n9491), .A2(n9438), .ZN(n9419) );
  OAI211_X1 U10837 ( .C1(n9494), .C2(n9441), .A(n9420), .B(n9419), .ZN(
        P2_U3480) );
  AOI21_X1 U10838 ( .B1(n9443), .B2(n7088), .A(n9421), .ZN(n9495) );
  MUX2_X1 U10839 ( .A(n9422), .B(n9495), .S(n10578), .Z(n9423) );
  OAI21_X1 U10840 ( .B1(n9441), .B2(n9498), .A(n9423), .ZN(P2_U3479) );
  MUX2_X1 U10841 ( .A(n9499), .B(P2_REG1_REG_19__SCAN_IN), .S(n7168), .Z(n9426) );
  OAI22_X1 U10842 ( .A1(n9502), .A2(n9441), .B1(n9501), .B2(n9424), .ZN(n9425)
         );
  OR2_X1 U10843 ( .A1(n9426), .A2(n9425), .ZN(P2_U3478) );
  MUX2_X1 U10844 ( .A(n9427), .B(n9505), .S(n10578), .Z(n9429) );
  NAND2_X1 U10845 ( .A1(n9507), .A2(n9438), .ZN(n9428) );
  OAI211_X1 U10846 ( .C1(n9441), .C2(n9510), .A(n9429), .B(n9428), .ZN(
        P2_U3477) );
  AOI21_X1 U10847 ( .B1(n9443), .B2(n9431), .A(n9430), .ZN(n9432) );
  OAI21_X1 U10848 ( .B1(n10567), .B2(n9433), .A(n9432), .ZN(n9511) );
  MUX2_X1 U10849 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9511), .S(n10578), .Z(
        P2_U3476) );
  MUX2_X1 U10850 ( .A(n9434), .B(n9512), .S(n10578), .Z(n9436) );
  NAND2_X1 U10851 ( .A1(n9514), .A2(n9438), .ZN(n9435) );
  OAI211_X1 U10852 ( .C1(n9517), .C2(n9441), .A(n9436), .B(n9435), .ZN(
        P2_U3475) );
  MUX2_X1 U10853 ( .A(n9437), .B(n9518), .S(n10578), .Z(n9440) );
  NAND2_X1 U10854 ( .A1(n9521), .A2(n9438), .ZN(n9439) );
  OAI211_X1 U10855 ( .C1(n9525), .C2(n9441), .A(n9440), .B(n9439), .ZN(
        P2_U3474) );
  AOI22_X1 U10856 ( .A1(n9444), .A2(n10562), .B1(n9443), .B2(n9442), .ZN(n9445) );
  NAND2_X1 U10857 ( .A1(n9446), .A2(n9445), .ZN(n9526) );
  MUX2_X1 U10858 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9526), .S(n10578), .Z(
        P2_U3465) );
  MUX2_X1 U10859 ( .A(n9447), .B(P2_REG1_REG_0__SCAN_IN), .S(n7168), .Z(
        P2_U3459) );
  NOR2_X1 U10860 ( .A1(n9448), .A2(n10573), .ZN(n9451) );
  AOI21_X1 U10861 ( .B1(n10573), .B2(P2_REG0_REG_31__SCAN_IN), .A(n9451), .ZN(
        n9449) );
  OAI21_X1 U10862 ( .B1(n9450), .B2(n9500), .A(n9449), .ZN(P2_U3458) );
  AOI21_X1 U10863 ( .B1(n10573), .B2(P2_REG0_REG_30__SCAN_IN), .A(n9451), .ZN(
        n9452) );
  OAI21_X1 U10864 ( .B1(n9453), .B2(n9500), .A(n9452), .ZN(P2_U3457) );
  INV_X1 U10865 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U10866 ( .A1(n9456), .A2(n9520), .ZN(n9457) );
  OAI211_X1 U10867 ( .C1(n9459), .C2(n9524), .A(n9458), .B(n9457), .ZN(
        P2_U3455) );
  MUX2_X1 U10868 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9460), .S(n10571), .Z(
        P2_U3454) );
  MUX2_X1 U10869 ( .A(n9462), .B(n9461), .S(n10571), .Z(n9465) );
  NAND2_X1 U10870 ( .A1(n9463), .A2(n9520), .ZN(n9464) );
  OAI211_X1 U10871 ( .C1(n9466), .C2(n9524), .A(n9465), .B(n9464), .ZN(
        P2_U3453) );
  INV_X1 U10872 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9468) );
  MUX2_X1 U10873 ( .A(n9468), .B(n9467), .S(n10571), .Z(n9471) );
  NAND2_X1 U10874 ( .A1(n9469), .A2(n9520), .ZN(n9470) );
  OAI211_X1 U10875 ( .C1(n9472), .C2(n9524), .A(n9471), .B(n9470), .ZN(
        P2_U3452) );
  MUX2_X1 U10876 ( .A(n9474), .B(n9473), .S(n10571), .Z(n9477) );
  NAND2_X1 U10877 ( .A1(n9475), .A2(n9520), .ZN(n9476) );
  OAI211_X1 U10878 ( .C1(n9478), .C2(n9524), .A(n9477), .B(n9476), .ZN(
        P2_U3451) );
  INV_X1 U10879 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9480) );
  MUX2_X1 U10880 ( .A(n9480), .B(n9479), .S(n10571), .Z(n9483) );
  NAND2_X1 U10881 ( .A1(n9481), .A2(n9520), .ZN(n9482) );
  OAI211_X1 U10882 ( .C1(n9484), .C2(n9524), .A(n9483), .B(n9482), .ZN(
        P2_U3450) );
  INV_X1 U10883 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9486) );
  MUX2_X1 U10884 ( .A(n9486), .B(n9485), .S(n10571), .Z(n9487) );
  OAI21_X1 U10885 ( .B1(n9488), .B2(n9500), .A(n9487), .ZN(P2_U3449) );
  INV_X1 U10886 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9490) );
  MUX2_X1 U10887 ( .A(n9490), .B(n9489), .S(n10571), .Z(n9493) );
  NAND2_X1 U10888 ( .A1(n9491), .A2(n9520), .ZN(n9492) );
  OAI211_X1 U10889 ( .C1(n9494), .C2(n9524), .A(n9493), .B(n9492), .ZN(
        P2_U3448) );
  INV_X1 U10890 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9496) );
  MUX2_X1 U10891 ( .A(n9496), .B(n9495), .S(n10571), .Z(n9497) );
  OAI21_X1 U10892 ( .B1(n9498), .B2(n9524), .A(n9497), .ZN(P2_U3447) );
  MUX2_X1 U10893 ( .A(n9499), .B(P2_REG0_REG_19__SCAN_IN), .S(n10573), .Z(
        n9504) );
  OAI22_X1 U10894 ( .A1(n9502), .A2(n9524), .B1(n9501), .B2(n9500), .ZN(n9503)
         );
  OR2_X1 U10895 ( .A1(n9504), .A2(n9503), .ZN(P2_U3446) );
  INV_X1 U10896 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9506) );
  MUX2_X1 U10897 ( .A(n9506), .B(n9505), .S(n10571), .Z(n9509) );
  NAND2_X1 U10898 ( .A1(n9507), .A2(n9520), .ZN(n9508) );
  OAI211_X1 U10899 ( .C1(n9510), .C2(n9524), .A(n9509), .B(n9508), .ZN(
        P2_U3444) );
  MUX2_X1 U10900 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9511), .S(n10571), .Z(
        P2_U3441) );
  MUX2_X1 U10901 ( .A(n9513), .B(n9512), .S(n10571), .Z(n9516) );
  NAND2_X1 U10902 ( .A1(n9514), .A2(n9520), .ZN(n9515) );
  OAI211_X1 U10903 ( .C1(n9517), .C2(n9524), .A(n9516), .B(n9515), .ZN(
        P2_U3438) );
  INV_X1 U10904 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9519) );
  MUX2_X1 U10905 ( .A(n9519), .B(n9518), .S(n10571), .Z(n9523) );
  NAND2_X1 U10906 ( .A1(n9521), .A2(n9520), .ZN(n9522) );
  OAI211_X1 U10907 ( .C1(n9525), .C2(n9524), .A(n9523), .B(n9522), .ZN(
        P2_U3435) );
  MUX2_X1 U10908 ( .A(P2_REG0_REG_6__SCAN_IN), .B(n9526), .S(n10571), .Z(
        P2_U3408) );
  INV_X1 U10909 ( .A(n9527), .ZN(n9532) );
  NOR4_X1 U10910 ( .A1(n9529), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9528), .ZN(n9530) );
  AOI21_X1 U10911 ( .B1(n9545), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9530), .ZN(
        n9531) );
  OAI21_X1 U10912 ( .B1(n9532), .B2(n9547), .A(n9531), .ZN(P2_U3264) );
  INV_X1 U10913 ( .A(n9533), .ZN(n10220) );
  AOI22_X1 U10914 ( .A1(n9534), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9545), .ZN(n9535) );
  OAI21_X1 U10915 ( .B1(n10220), .B2(n9547), .A(n9535), .ZN(P2_U3265) );
  INV_X1 U10916 ( .A(n9536), .ZN(n10222) );
  INV_X1 U10917 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9538) );
  OAI222_X1 U10918 ( .A1(n9547), .A2(n10222), .B1(n9540), .B2(P2_U3151), .C1(
        n9538), .C2(n9537), .ZN(P2_U3266) );
  AOI21_X1 U10919 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9545), .A(n9541), .ZN(
        n9542) );
  OAI21_X1 U10920 ( .B1(n9543), .B2(n9547), .A(n9542), .ZN(P2_U3267) );
  AOI21_X1 U10921 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9545), .A(n9544), .ZN(
        n9546) );
  OAI21_X1 U10922 ( .B1(n9548), .B2(n9547), .A(n9546), .ZN(P2_U3268) );
  MUX2_X1 U10923 ( .A(n9549), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  XNOR2_X1 U10924 ( .A(n9550), .B(n9610), .ZN(n9551) );
  NOR2_X1 U10925 ( .A1(n9551), .A2(n9552), .ZN(n9609) );
  AOI21_X1 U10926 ( .B1(n9552), .B2(n9551), .A(n9609), .ZN(n9558) );
  NAND2_X1 U10927 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10249)
         );
  NAND2_X1 U10928 ( .A1(n9710), .A2(n9553), .ZN(n9554) );
  OAI211_X1 U10929 ( .C1(n9708), .C2(n9555), .A(n10249), .B(n9554), .ZN(n9556)
         );
  AOI21_X1 U10930 ( .B1(n10147), .B2(n9693), .A(n9556), .ZN(n9557) );
  OAI21_X1 U10931 ( .B1(n9558), .B2(n9695), .A(n9557), .ZN(P1_U3215) );
  INV_X1 U10932 ( .A(n9634), .ZN(n9561) );
  NOR3_X1 U10933 ( .A1(n4751), .A2(n9660), .A3(n9559), .ZN(n9560) );
  OAI21_X1 U10934 ( .B1(n9561), .B2(n9560), .A(n9716), .ZN(n9568) );
  OR2_X1 U10935 ( .A1(n9604), .A2(n9703), .ZN(n9563) );
  NAND2_X1 U10936 ( .A1(n9733), .A2(n9687), .ZN(n9562) );
  NAND2_X1 U10937 ( .A1(n9563), .A2(n9562), .ZN(n10101) );
  INV_X1 U10938 ( .A(n9966), .ZN(n9565) );
  OAI22_X1 U10939 ( .A1(n9565), .A2(n9708), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9564), .ZN(n9566) );
  AOI21_X1 U10940 ( .B1(n10101), .B2(n9710), .A(n9566), .ZN(n9567) );
  OAI211_X1 U10941 ( .C1(n9968), .C2(n9725), .A(n9568), .B(n9567), .ZN(
        P1_U3216) );
  OAI21_X1 U10942 ( .B1(n9571), .B2(n9570), .A(n9569), .ZN(n9572) );
  NAND2_X1 U10943 ( .A1(n9572), .A2(n9716), .ZN(n9577) );
  AOI22_X1 U10944 ( .A1(n9710), .A2(n9573), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n9576) );
  NAND2_X1 U10945 ( .A1(n9721), .A2(n8104), .ZN(n9575) );
  NAND2_X1 U10946 ( .A1(n9693), .A2(n6539), .ZN(n9574) );
  NAND4_X1 U10947 ( .A1(n9577), .A2(n9576), .A3(n9575), .A4(n9574), .ZN(
        P1_U3218) );
  XNOR2_X1 U10948 ( .A(n9578), .B(n9579), .ZN(n9684) );
  NOR2_X1 U10949 ( .A1(n9684), .A2(n9685), .ZN(n9683) );
  AOI21_X1 U10950 ( .B1(n9578), .B2(n9579), .A(n9683), .ZN(n9583) );
  XNOR2_X1 U10951 ( .A(n9581), .B(n9580), .ZN(n9582) );
  XNOR2_X1 U10952 ( .A(n9583), .B(n9582), .ZN(n9590) );
  OR2_X1 U10953 ( .A1(n9593), .A2(n9703), .ZN(n9586) );
  OR2_X1 U10954 ( .A1(n9584), .A2(n9701), .ZN(n9585) );
  AND2_X1 U10955 ( .A1(n9586), .A2(n9585), .ZN(n10020) );
  NAND2_X1 U10956 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U10957 ( .A1(n9721), .A2(n10024), .ZN(n9587) );
  OAI211_X1 U10958 ( .C1(n10020), .C2(n9719), .A(n9875), .B(n9587), .ZN(n9588)
         );
  AOI21_X1 U10959 ( .B1(n10123), .B2(n9693), .A(n9588), .ZN(n9589) );
  OAI21_X1 U10960 ( .B1(n9590), .B2(n9695), .A(n9589), .ZN(P1_U3219) );
  XOR2_X1 U10961 ( .A(n9592), .B(n9591), .Z(n9600) );
  OAI22_X1 U10962 ( .A1(n9594), .A2(n9703), .B1(n9593), .B2(n9701), .ZN(n9595)
         );
  INV_X1 U10963 ( .A(n9595), .ZN(n9994) );
  OAI22_X1 U10964 ( .A1(n9994), .A2(n9719), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9596), .ZN(n9598) );
  NOR2_X1 U10965 ( .A1(n5075), .A2(n9725), .ZN(n9597) );
  AOI211_X1 U10966 ( .C1(n9997), .C2(n9721), .A(n9598), .B(n9597), .ZN(n9599)
         );
  OAI21_X1 U10967 ( .B1(n9600), .B2(n9695), .A(n9599), .ZN(P1_U3223) );
  AOI21_X1 U10968 ( .B1(n9602), .B2(n9601), .A(n9699), .ZN(n9608) );
  OAI22_X1 U10969 ( .A1(n9604), .A2(n9701), .B1(n9603), .B2(n9703), .ZN(n9940)
         );
  AOI22_X1 U10970 ( .A1(n9931), .A2(n9721), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9605) );
  OAI21_X1 U10971 ( .B1(n4549), .B2(n9719), .A(n9605), .ZN(n9606) );
  AOI21_X1 U10972 ( .B1(n10091), .B2(n9693), .A(n9606), .ZN(n9607) );
  OAI21_X1 U10973 ( .B1(n9608), .B2(n9695), .A(n9607), .ZN(P1_U3225) );
  AOI21_X1 U10974 ( .B1(n9610), .B2(n9550), .A(n9609), .ZN(n9613) );
  XNOR2_X1 U10975 ( .A(n9613), .B(n9611), .ZN(n9714) );
  INV_X1 U10976 ( .A(n9612), .ZN(n9715) );
  NAND2_X1 U10977 ( .A1(n9714), .A2(n9715), .ZN(n9713) );
  OAI21_X1 U10978 ( .B1(n9614), .B2(n9613), .A(n9713), .ZN(n9619) );
  OAI21_X1 U10979 ( .B1(n9617), .B2(n9616), .A(n9615), .ZN(n9618) );
  XNOR2_X1 U10980 ( .A(n9619), .B(n9618), .ZN(n9623) );
  NOR2_X1 U10981 ( .A1(n9708), .A2(n10069), .ZN(n9621) );
  AOI22_X1 U10982 ( .A1(n9736), .A2(n9649), .B1(n9687), .B2(n9739), .ZN(n10065) );
  NAND2_X1 U10983 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10275)
         );
  OAI21_X1 U10984 ( .B1(n9719), .B2(n10065), .A(n10275), .ZN(n9620) );
  AOI211_X1 U10985 ( .C1(n10138), .C2(n9693), .A(n9621), .B(n9620), .ZN(n9622)
         );
  OAI21_X1 U10986 ( .B1(n9623), .B2(n9695), .A(n9622), .ZN(P1_U3226) );
  NAND2_X1 U10987 ( .A1(n9625), .A2(n9624), .ZN(n9626) );
  XNOR2_X1 U10988 ( .A(n9627), .B(n9626), .ZN(n9631) );
  AOI22_X1 U10989 ( .A1(n9735), .A2(n9649), .B1(n9687), .B2(n9737), .ZN(n10047) );
  NAND2_X1 U10990 ( .A1(n9721), .A2(n10051), .ZN(n9628) );
  NAND2_X1 U10991 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10290)
         );
  OAI211_X1 U10992 ( .C1(n10047), .C2(n9719), .A(n9628), .B(n10290), .ZN(n9629) );
  AOI21_X1 U10993 ( .B1(n10133), .B2(n9693), .A(n9629), .ZN(n9630) );
  OAI21_X1 U10994 ( .B1(n9631), .B2(n9695), .A(n9630), .ZN(P1_U3228) );
  AND3_X1 U10995 ( .A1(n9634), .A2(n9633), .A3(n9632), .ZN(n9635) );
  OAI21_X1 U10996 ( .B1(n9636), .B2(n9635), .A(n9716), .ZN(n9644) );
  OR2_X1 U10997 ( .A1(n9702), .A2(n9703), .ZN(n9638) );
  OR2_X1 U10998 ( .A1(n9663), .A2(n9701), .ZN(n9637) );
  AND2_X1 U10999 ( .A1(n9638), .A2(n9637), .ZN(n9946) );
  INV_X1 U11000 ( .A(n9946), .ZN(n9642) );
  OAI22_X1 U11001 ( .A1(n9640), .A2(n9708), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9639), .ZN(n9641) );
  AOI21_X1 U11002 ( .B1(n9642), .B2(n9710), .A(n9641), .ZN(n9643) );
  OAI211_X1 U11003 ( .C1(n9955), .C2(n9725), .A(n9644), .B(n9643), .ZN(
        P1_U3229) );
  XNOR2_X1 U11004 ( .A(n9646), .B(n9645), .ZN(n9647) );
  XNOR2_X1 U11005 ( .A(n9648), .B(n9647), .ZN(n9655) );
  AOI22_X1 U11006 ( .A1(n9664), .A2(n9649), .B1(n9687), .B2(n9734), .ZN(n10006) );
  INV_X1 U11007 ( .A(n10006), .ZN(n9650) );
  AOI22_X1 U11008 ( .A1(n9650), .A2(n9710), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9651) );
  OAI21_X1 U11009 ( .B1(n9708), .B2(n9652), .A(n9651), .ZN(n9653) );
  AOI21_X1 U11010 ( .B1(n10118), .B2(n9693), .A(n9653), .ZN(n9654) );
  OAI21_X1 U11011 ( .B1(n9655), .B2(n9695), .A(n9654), .ZN(P1_U3233) );
  OAI21_X1 U11012 ( .B1(n9658), .B2(n9660), .A(n9657), .ZN(n9659) );
  OAI21_X1 U11013 ( .B1(n4593), .B2(n9660), .A(n9659), .ZN(n9661) );
  NAND2_X1 U11014 ( .A1(n9661), .A2(n9716), .ZN(n9670) );
  INV_X1 U11015 ( .A(n9662), .ZN(n9985) );
  OR2_X1 U11016 ( .A1(n9663), .A2(n9703), .ZN(n9666) );
  NAND2_X1 U11017 ( .A1(n9664), .A2(n9687), .ZN(n9665) );
  AND2_X1 U11018 ( .A1(n9666), .A2(n9665), .ZN(n9982) );
  OAI22_X1 U11019 ( .A1(n9982), .A2(n9719), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9667), .ZN(n9668) );
  AOI21_X1 U11020 ( .B1(n9985), .B2(n9721), .A(n9668), .ZN(n9669) );
  OAI211_X1 U11021 ( .C1(n9988), .C2(n9725), .A(n9670), .B(n9669), .ZN(
        P1_U3235) );
  AOI21_X1 U11022 ( .B1(n8550), .B2(n9672), .A(n9671), .ZN(n9676) );
  XNOR2_X1 U11023 ( .A(n9674), .B(n9673), .ZN(n9675) );
  XNOR2_X1 U11024 ( .A(n9676), .B(n9675), .ZN(n9682) );
  NAND2_X1 U11025 ( .A1(n9721), .A2(n9677), .ZN(n9678) );
  NAND2_X1 U11026 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9837) );
  OAI211_X1 U11027 ( .C1(n9719), .C2(n9679), .A(n9678), .B(n9837), .ZN(n9680)
         );
  AOI21_X1 U11028 ( .B1(n10489), .B2(n9693), .A(n9680), .ZN(n9681) );
  OAI21_X1 U11029 ( .B1(n9682), .B2(n9695), .A(n9681), .ZN(P1_U3236) );
  AOI21_X1 U11030 ( .B1(n9685), .B2(n9684), .A(n9683), .ZN(n9696) );
  OR2_X1 U11031 ( .A1(n9686), .A2(n9703), .ZN(n9689) );
  NAND2_X1 U11032 ( .A1(n9736), .A2(n9687), .ZN(n9688) );
  NAND2_X1 U11033 ( .A1(n9689), .A2(n9688), .ZN(n10033) );
  NAND2_X1 U11034 ( .A1(n10033), .A2(n9710), .ZN(n9690) );
  NAND2_X1 U11035 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10306)
         );
  OAI211_X1 U11036 ( .C1(n9708), .C2(n9691), .A(n9690), .B(n10306), .ZN(n9692)
         );
  AOI21_X1 U11037 ( .B1(n10128), .B2(n9693), .A(n9692), .ZN(n9694) );
  OAI21_X1 U11038 ( .B1(n9696), .B2(n9695), .A(n9694), .ZN(P1_U3238) );
  OR2_X1 U11039 ( .A1(n9702), .A2(n9701), .ZN(n9706) );
  OR2_X1 U11040 ( .A1(n9704), .A2(n9703), .ZN(n9705) );
  AND2_X1 U11041 ( .A1(n9706), .A2(n9705), .ZN(n9926) );
  INV_X1 U11042 ( .A(n9926), .ZN(n9711) );
  INV_X1 U11043 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9707) );
  OAI22_X1 U11044 ( .A1(n9708), .A2(n9920), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9707), .ZN(n9709) );
  AOI21_X1 U11045 ( .B1(n9711), .B2(n9710), .A(n9709), .ZN(n9712) );
  OAI21_X1 U11046 ( .B1(n9715), .B2(n9714), .A(n9713), .ZN(n9717) );
  NAND2_X1 U11047 ( .A1(n9717), .A2(n9716), .ZN(n9724) );
  NAND2_X1 U11048 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10261)
         );
  OAI21_X1 U11049 ( .B1(n9719), .B2(n9718), .A(n10261), .ZN(n9720) );
  AOI21_X1 U11050 ( .B1(n9722), .B2(n9721), .A(n9720), .ZN(n9723) );
  OAI211_X1 U11051 ( .C1(n9726), .C2(n9725), .A(n9724), .B(n9723), .ZN(
        P1_U3241) );
  MUX2_X1 U11052 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9727), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U11053 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9728), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U11054 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9729), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U11055 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9730), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U11056 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9731), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U11057 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9732), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U11058 ( .A(n9733), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9738), .Z(
        P1_U3576) );
  MUX2_X1 U11059 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9734), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U11060 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9735), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U11061 ( .A(n9736), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9738), .Z(
        P1_U3571) );
  MUX2_X1 U11062 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9737), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U11063 ( .A(n9739), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9738), .Z(
        P1_U3569) );
  MUX2_X1 U11064 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9740), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U11065 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9741), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U11066 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9742), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U11067 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9743), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U11068 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9744), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U11069 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9745), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U11070 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9746), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U11071 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9747), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U11072 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9748), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U11073 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9749), .S(P1_U3973), .Z(
        P1_U3559) );
  INV_X1 U11074 ( .A(n9750), .ZN(n9751) );
  MUX2_X1 U11075 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9751), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U11076 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9752), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U11077 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n4735), .S(P1_U3973), .Z(
        P1_U3556) );
  OAI211_X1 U11078 ( .C1(n9755), .C2(n9754), .A(n10293), .B(n9753), .ZN(n9763)
         );
  OAI211_X1 U11079 ( .C1(n9758), .C2(n9757), .A(n10284), .B(n9756), .ZN(n9762)
         );
  AOI22_X1 U11080 ( .A1(n10233), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9761) );
  NAND2_X1 U11081 ( .A1(n10305), .A2(n9759), .ZN(n9760) );
  NAND4_X1 U11082 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(
        P1_U3244) );
  INV_X1 U11083 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9765) );
  NAND2_X1 U11084 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9764) );
  OAI21_X1 U11085 ( .B1(n10308), .B2(n9765), .A(n9764), .ZN(n9766) );
  AOI21_X1 U11086 ( .B1(n9767), .B2(n10305), .A(n9766), .ZN(n9776) );
  OAI211_X1 U11087 ( .C1(n9770), .C2(n9769), .A(n10284), .B(n9768), .ZN(n9775)
         );
  OAI211_X1 U11088 ( .C1(n9773), .C2(n9772), .A(n10293), .B(n9771), .ZN(n9774)
         );
  NAND3_X1 U11089 ( .A1(n9776), .A2(n9775), .A3(n9774), .ZN(P1_U3246) );
  INV_X1 U11090 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U11091 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9777) );
  OAI21_X1 U11092 ( .B1(n10308), .B2(n9778), .A(n9777), .ZN(n9779) );
  AOI21_X1 U11093 ( .B1(n9780), .B2(n10305), .A(n9779), .ZN(n9789) );
  OAI211_X1 U11094 ( .C1(n9783), .C2(n9782), .A(n10284), .B(n9781), .ZN(n9788)
         );
  OAI211_X1 U11095 ( .C1(n9786), .C2(n9785), .A(n10293), .B(n9784), .ZN(n9787)
         );
  NAND3_X1 U11096 ( .A1(n9789), .A2(n9788), .A3(n9787), .ZN(P1_U3248) );
  INV_X1 U11097 ( .A(n9790), .ZN(n9794) );
  OAI21_X1 U11098 ( .B1(n10308), .B2(n9792), .A(n9791), .ZN(n9793) );
  AOI21_X1 U11099 ( .B1(n9794), .B2(n10305), .A(n9793), .ZN(n9803) );
  OAI211_X1 U11100 ( .C1(n9797), .C2(n9796), .A(n10284), .B(n9795), .ZN(n9802)
         );
  OAI211_X1 U11101 ( .C1(n9800), .C2(n9799), .A(n10293), .B(n9798), .ZN(n9801)
         );
  NAND3_X1 U11102 ( .A1(n9803), .A2(n9802), .A3(n9801), .ZN(P1_U3249) );
  INV_X1 U11103 ( .A(n9804), .ZN(n9808) );
  INV_X1 U11104 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9806) );
  OAI21_X1 U11105 ( .B1(n10308), .B2(n9806), .A(n9805), .ZN(n9807) );
  AOI21_X1 U11106 ( .B1(n9808), .B2(n10305), .A(n9807), .ZN(n9817) );
  OAI211_X1 U11107 ( .C1(n9811), .C2(n9810), .A(n10293), .B(n9809), .ZN(n9816)
         );
  OAI211_X1 U11108 ( .C1(n9814), .C2(n9813), .A(n10284), .B(n9812), .ZN(n9815)
         );
  NAND3_X1 U11109 ( .A1(n9817), .A2(n9816), .A3(n9815), .ZN(P1_U3250) );
  INV_X1 U11110 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9819) );
  OAI21_X1 U11111 ( .B1(n10308), .B2(n9819), .A(n9818), .ZN(n9820) );
  AOI21_X1 U11112 ( .B1(n9821), .B2(n10305), .A(n9820), .ZN(n9830) );
  OAI211_X1 U11113 ( .C1(n9824), .C2(n9823), .A(n9822), .B(n10293), .ZN(n9829)
         );
  OAI211_X1 U11114 ( .C1(n9827), .C2(n9826), .A(n9825), .B(n10284), .ZN(n9828)
         );
  NAND3_X1 U11115 ( .A1(n9830), .A2(n9829), .A3(n9828), .ZN(P1_U3251) );
  OAI211_X1 U11116 ( .C1(n9833), .C2(n9832), .A(n9831), .B(n10284), .ZN(n9843)
         );
  OAI211_X1 U11117 ( .C1(n9836), .C2(n9835), .A(n9834), .B(n10293), .ZN(n9842)
         );
  INV_X1 U11118 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9838) );
  OAI21_X1 U11119 ( .B1(n10308), .B2(n9838), .A(n9837), .ZN(n9839) );
  AOI21_X1 U11120 ( .B1(n9840), .B2(n10305), .A(n9839), .ZN(n9841) );
  NAND3_X1 U11121 ( .A1(n9843), .A2(n9842), .A3(n9841), .ZN(P1_U3254) );
  INV_X1 U11122 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U11123 ( .A1(n9853), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9844) );
  NAND2_X1 U11124 ( .A1(n9845), .A2(n9844), .ZN(n10238) );
  INV_X1 U11125 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9846) );
  XNOR2_X1 U11126 ( .A(n10243), .B(n9846), .ZN(n10237) );
  NOR2_X1 U11127 ( .A1(n9847), .A2(n9858), .ZN(n9848) );
  INV_X1 U11128 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10253) );
  XNOR2_X1 U11129 ( .A(n9858), .B(n9847), .ZN(n10254) );
  NOR2_X1 U11130 ( .A1(n10253), .A2(n10254), .ZN(n10252) );
  INV_X1 U11131 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10139) );
  XNOR2_X1 U11132 ( .A(n10274), .B(n10139), .ZN(n10265) );
  NOR2_X1 U11133 ( .A1(n10274), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9849) );
  AOI21_X1 U11134 ( .B1(n10264), .B2(n10265), .A(n9849), .ZN(n10283) );
  XNOR2_X1 U11135 ( .A(n10286), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10282) );
  OAI22_X1 U11136 ( .A1(n10283), .A2(n10282), .B1(P1_REG1_REG_17__SCAN_IN), 
        .B2(n10286), .ZN(n10301) );
  NAND2_X1 U11137 ( .A1(n10304), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9850) );
  OAI21_X1 U11138 ( .B1(n10304), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9850), .ZN(
        n10300) );
  NOR2_X1 U11139 ( .A1(n10301), .A2(n10300), .ZN(n10298) );
  INV_X1 U11140 ( .A(n9850), .ZN(n9851) );
  NOR2_X1 U11141 ( .A1(n10298), .A2(n9851), .ZN(n9852) );
  XNOR2_X1 U11142 ( .A(n9852), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9869) );
  NAND2_X1 U11143 ( .A1(n9853), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U11144 ( .A1(n9855), .A2(n9854), .ZN(n10240) );
  OR2_X1 U11145 ( .A1(n10243), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9857) );
  NAND2_X1 U11146 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n10243), .ZN(n9856) );
  AND2_X1 U11147 ( .A1(n9857), .A2(n9856), .ZN(n10239) );
  NOR2_X1 U11148 ( .A1(n9859), .A2(n9858), .ZN(n9860) );
  XOR2_X1 U11149 ( .A(n10260), .B(n9859), .Z(n10257) );
  NOR2_X1 U11150 ( .A1(n10256), .A2(n10257), .ZN(n10255) );
  XNOR2_X1 U11151 ( .A(n10274), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n10270) );
  NAND2_X1 U11152 ( .A1(n10274), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9861) );
  INV_X1 U11153 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9862) );
  XNOR2_X1 U11154 ( .A(n10286), .B(n9862), .ZN(n10280) );
  NAND2_X1 U11155 ( .A1(n10279), .A2(n10280), .ZN(n10278) );
  OR2_X1 U11156 ( .A1(n10286), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9863) );
  NAND2_X1 U11157 ( .A1(n10304), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9865) );
  OR2_X1 U11158 ( .A1(n10304), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9864) );
  AND2_X1 U11159 ( .A1(n9865), .A2(n9864), .ZN(n10295) );
  NAND2_X1 U11160 ( .A1(n10294), .A2(n9865), .ZN(n9866) );
  INV_X1 U11161 ( .A(n9871), .ZN(n9867) );
  OAI21_X1 U11162 ( .B1(n9869), .B2(n10299), .A(n9868), .ZN(n9870) );
  AOI21_X1 U11163 ( .B1(n10293), .B2(n9871), .A(n9870), .ZN(n9873) );
  NAND2_X1 U11164 ( .A1(n9883), .A2(n10079), .ZN(n9882) );
  XNOR2_X1 U11165 ( .A(n10076), .B(n9882), .ZN(n9877) );
  NAND2_X1 U11166 ( .A1(n9877), .A2(n10390), .ZN(n10075) );
  NAND2_X1 U11167 ( .A1(n9879), .A2(n9878), .ZN(n10077) );
  NOR2_X1 U11168 ( .A1(n10402), .A2(n10077), .ZN(n9885) );
  NOR2_X1 U11169 ( .A1(n10076), .A2(n10385), .ZN(n9880) );
  AOI211_X1 U11170 ( .C1(n10402), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9885), .B(
        n9880), .ZN(n9881) );
  OAI21_X1 U11171 ( .B1(n10075), .B2(n10411), .A(n9881), .ZN(P1_U3263) );
  OAI211_X1 U11172 ( .C1(n9883), .C2(n10079), .A(n10390), .B(n9882), .ZN(
        n10078) );
  NOR2_X1 U11173 ( .A1(n10079), .A2(n10385), .ZN(n9884) );
  AOI211_X1 U11174 ( .C1(n10402), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9885), .B(
        n9884), .ZN(n9886) );
  OAI21_X1 U11175 ( .B1(n10411), .B2(n10078), .A(n9886), .ZN(P1_U3264) );
  INV_X1 U11176 ( .A(n10158), .ZN(n9896) );
  NOR2_X1 U11177 ( .A1(n9887), .A2(n10411), .ZN(n9893) );
  NOR2_X1 U11178 ( .A1(n10382), .A2(n9888), .ZN(n9889) );
  AOI21_X1 U11179 ( .B1(n10402), .B2(P1_REG2_REG_28__SCAN_IN), .A(n9889), .ZN(
        n9890) );
  OAI21_X1 U11180 ( .B1(n9891), .B2(n10385), .A(n9890), .ZN(n9892) );
  AOI211_X1 U11181 ( .C1(n9894), .C2(n10324), .A(n9893), .B(n9892), .ZN(n9895)
         );
  OAI21_X1 U11182 ( .B1(n9896), .B2(n10412), .A(n9895), .ZN(P1_U3265) );
  AOI211_X1 U11183 ( .C1(n10083), .C2(n9918), .A(n10407), .B(n9900), .ZN(
        n10082) );
  OAI22_X1 U11184 ( .A1(n9902), .A2(n10385), .B1(n9901), .B2(n10324), .ZN(
        n9903) );
  AOI21_X1 U11185 ( .B1(n10082), .B2(n10393), .A(n9903), .ZN(n9913) );
  OAI21_X1 U11186 ( .B1(n9907), .B2(n9906), .A(n10399), .ZN(n9909) );
  NOR2_X1 U11187 ( .A1(n10382), .A2(n9910), .ZN(n9911) );
  OAI21_X1 U11188 ( .B1(n10081), .B2(n9911), .A(n10324), .ZN(n9912) );
  OAI211_X1 U11189 ( .C1(n10163), .C2(n10412), .A(n9913), .B(n9912), .ZN(
        P1_U3266) );
  INV_X1 U11190 ( .A(n9914), .ZN(n9917) );
  INV_X1 U11191 ( .A(n9915), .ZN(n9916) );
  INV_X1 U11192 ( .A(n9918), .ZN(n9919) );
  AOI211_X1 U11193 ( .C1(n10087), .C2(n9930), .A(n10407), .B(n9919), .ZN(
        n10085) );
  NOR2_X1 U11194 ( .A1(n5084), .A2(n10385), .ZN(n9923) );
  OAI22_X1 U11195 ( .A1(n10324), .A2(n9921), .B1(n9920), .B2(n10382), .ZN(
        n9922) );
  AOI211_X1 U11196 ( .C1(n10085), .C2(n10393), .A(n9923), .B(n9922), .ZN(n9928) );
  NAND2_X1 U11197 ( .A1(n10086), .A2(n10324), .ZN(n9927) );
  OAI211_X1 U11198 ( .C1(n10167), .C2(n10412), .A(n9928), .B(n9927), .ZN(
        P1_U3267) );
  XNOR2_X1 U11199 ( .A(n9929), .B(n9935), .ZN(n10094) );
  AOI211_X1 U11200 ( .C1(n10091), .C2(n9949), .A(n10407), .B(n5085), .ZN(
        n10090) );
  AOI22_X1 U11201 ( .A1(n9931), .A2(n10401), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10402), .ZN(n9932) );
  OAI21_X1 U11202 ( .B1(n9933), .B2(n10385), .A(n9932), .ZN(n9941) );
  OAI21_X1 U11203 ( .B1(n9937), .B2(n9936), .A(n9935), .ZN(n9939) );
  OAI21_X1 U11204 ( .B1(n10094), .B2(n10412), .A(n9942), .ZN(P1_U3268) );
  XNOR2_X1 U11205 ( .A(n9943), .B(n9944), .ZN(n10172) );
  NAND2_X1 U11206 ( .A1(n9934), .A2(n10399), .ZN(n9948) );
  AOI21_X1 U11207 ( .B1(n9969), .B2(n9945), .A(n5249), .ZN(n9947) );
  OAI21_X1 U11208 ( .B1(n9948), .B2(n9947), .A(n9946), .ZN(n10096) );
  INV_X1 U11209 ( .A(n9964), .ZN(n9951) );
  INV_X1 U11210 ( .A(n9949), .ZN(n9950) );
  AOI211_X1 U11211 ( .C1(n10097), .C2(n9951), .A(n10407), .B(n9950), .ZN(
        n10095) );
  NAND2_X1 U11212 ( .A1(n10095), .A2(n10393), .ZN(n9954) );
  AOI22_X1 U11213 ( .A1(n9952), .A2(n10401), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10402), .ZN(n9953) );
  OAI211_X1 U11214 ( .C1(n9955), .C2(n10385), .A(n9954), .B(n9953), .ZN(n9956)
         );
  AOI21_X1 U11215 ( .B1(n10324), .B2(n10096), .A(n9956), .ZN(n9957) );
  OAI21_X1 U11216 ( .B1(n10172), .B2(n10412), .A(n9957), .ZN(P1_U3269) );
  INV_X1 U11217 ( .A(n9958), .ZN(n9959) );
  NAND2_X1 U11218 ( .A1(n9960), .A2(n9959), .ZN(n9978) );
  NOR2_X1 U11219 ( .A1(n9977), .A2(n9961), .ZN(n9962) );
  XNOR2_X1 U11220 ( .A(n9962), .B(n9971), .ZN(n10105) );
  INV_X1 U11221 ( .A(n9963), .ZN(n9965) );
  AOI211_X1 U11222 ( .C1(n10102), .C2(n9965), .A(n10407), .B(n9964), .ZN(
        n10100) );
  AOI22_X1 U11223 ( .A1(n9966), .A2(n10401), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10402), .ZN(n9967) );
  OAI21_X1 U11224 ( .B1(n9968), .B2(n10385), .A(n9967), .ZN(n9975) );
  OAI21_X1 U11225 ( .B1(n9971), .B2(n9970), .A(n9969), .ZN(n9972) );
  NAND2_X1 U11226 ( .A1(n9972), .A2(n10399), .ZN(n10103) );
  INV_X1 U11227 ( .A(n10101), .ZN(n9973) );
  AOI21_X1 U11228 ( .B1(n10103), .B2(n9973), .A(n10402), .ZN(n9974) );
  AOI211_X1 U11229 ( .C1(n10100), .C2(n10393), .A(n9975), .B(n9974), .ZN(n9976) );
  OAI21_X1 U11230 ( .B1(n10105), .B2(n10412), .A(n9976), .ZN(P1_U3270) );
  AOI21_X1 U11231 ( .B1(n6973), .B2(n9978), .A(n9977), .ZN(n9979) );
  INV_X1 U11232 ( .A(n9979), .ZN(n10177) );
  XNOR2_X1 U11233 ( .A(n9981), .B(n9980), .ZN(n9983) );
  OAI21_X1 U11234 ( .B1(n9983), .B2(n10048), .A(n9982), .ZN(n10106) );
  INV_X1 U11235 ( .A(n9996), .ZN(n9984) );
  AOI211_X1 U11236 ( .C1(n10108), .C2(n9984), .A(n10407), .B(n9963), .ZN(
        n10107) );
  NAND2_X1 U11237 ( .A1(n10107), .A2(n10393), .ZN(n9987) );
  AOI22_X1 U11238 ( .A1(n9985), .A2(n10401), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10402), .ZN(n9986) );
  OAI211_X1 U11239 ( .C1(n9988), .C2(n10385), .A(n9987), .B(n9986), .ZN(n9989)
         );
  AOI21_X1 U11240 ( .B1(n10324), .B2(n10106), .A(n9989), .ZN(n9990) );
  OAI21_X1 U11241 ( .B1(n10177), .B2(n10412), .A(n9990), .ZN(P1_U3271) );
  XNOR2_X1 U11242 ( .A(n9991), .B(n9992), .ZN(n10181) );
  XNOR2_X1 U11243 ( .A(n9993), .B(n9992), .ZN(n9995) );
  OAI21_X1 U11244 ( .B1(n9995), .B2(n10048), .A(n9994), .ZN(n10111) );
  AOI211_X1 U11245 ( .C1(n10113), .C2(n10008), .A(n10407), .B(n9996), .ZN(
        n10112) );
  NAND2_X1 U11246 ( .A1(n10112), .A2(n10393), .ZN(n9999) );
  AOI22_X1 U11247 ( .A1(n9997), .A2(n10401), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n10402), .ZN(n9998) );
  OAI211_X1 U11248 ( .C1(n5075), .C2(n10385), .A(n9999), .B(n9998), .ZN(n10000) );
  AOI21_X1 U11249 ( .B1(n10324), .B2(n10111), .A(n10000), .ZN(n10001) );
  OAI21_X1 U11250 ( .B1(n10181), .B2(n10412), .A(n10001), .ZN(P1_U3272) );
  XOR2_X1 U11251 ( .A(n10004), .B(n10002), .Z(n10185) );
  OAI211_X1 U11252 ( .C1(n10005), .C2(n10004), .A(n10003), .B(n10399), .ZN(
        n10007) );
  NAND2_X1 U11253 ( .A1(n10007), .A2(n10006), .ZN(n10117) );
  INV_X1 U11254 ( .A(n10008), .ZN(n10009) );
  AOI211_X1 U11255 ( .C1(n10118), .C2(n4457), .A(n10407), .B(n10009), .ZN(
        n10116) );
  NAND2_X1 U11256 ( .A1(n10116), .A2(n10393), .ZN(n10012) );
  AOI22_X1 U11257 ( .A1(n10010), .A2(n10401), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n10402), .ZN(n10011) );
  OAI211_X1 U11258 ( .C1(n10013), .C2(n10385), .A(n10012), .B(n10011), .ZN(
        n10014) );
  AOI21_X1 U11259 ( .B1(n10324), .B2(n10117), .A(n10014), .ZN(n10015) );
  OAI21_X1 U11260 ( .B1(n10185), .B2(n10412), .A(n10015), .ZN(P1_U3273) );
  XNOR2_X1 U11261 ( .A(n10017), .B(n10016), .ZN(n10189) );
  XNOR2_X1 U11262 ( .A(n10019), .B(n10018), .ZN(n10021) );
  OAI21_X1 U11263 ( .B1(n10021), .B2(n10048), .A(n10020), .ZN(n10121) );
  INV_X1 U11264 ( .A(n4457), .ZN(n10023) );
  AOI211_X1 U11265 ( .C1(n10123), .C2(n10022), .A(n10407), .B(n10023), .ZN(
        n10122) );
  NAND2_X1 U11266 ( .A1(n10122), .A2(n10393), .ZN(n10026) );
  AOI22_X1 U11267 ( .A1(n10024), .A2(n10401), .B1(n10402), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n10025) );
  OAI211_X1 U11268 ( .C1(n10027), .C2(n10385), .A(n10026), .B(n10025), .ZN(
        n10028) );
  AOI21_X1 U11269 ( .B1(n10324), .B2(n10121), .A(n10028), .ZN(n10029) );
  OAI21_X1 U11270 ( .B1(n10189), .B2(n10412), .A(n10029), .ZN(P1_U3274) );
  XOR2_X1 U11271 ( .A(n10031), .B(n10030), .Z(n10193) );
  XOR2_X1 U11272 ( .A(n10032), .B(n10031), .Z(n10035) );
  INV_X1 U11273 ( .A(n10033), .ZN(n10034) );
  OAI21_X1 U11274 ( .B1(n10035), .B2(n10048), .A(n10034), .ZN(n10126) );
  INV_X1 U11275 ( .A(n10036), .ZN(n10038) );
  INV_X1 U11276 ( .A(n10022), .ZN(n10037) );
  AOI211_X1 U11277 ( .C1(n10128), .C2(n10038), .A(n10407), .B(n10037), .ZN(
        n10127) );
  NAND2_X1 U11278 ( .A1(n10127), .A2(n10393), .ZN(n10041) );
  AOI22_X1 U11279 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n10402), .B1(n10039), 
        .B2(n10401), .ZN(n10040) );
  OAI211_X1 U11280 ( .C1(n10042), .C2(n10385), .A(n10041), .B(n10040), .ZN(
        n10043) );
  AOI21_X1 U11281 ( .B1(n10324), .B2(n10126), .A(n10043), .ZN(n10044) );
  OAI21_X1 U11282 ( .B1(n10193), .B2(n10412), .A(n10044), .ZN(P1_U3275) );
  XNOR2_X1 U11283 ( .A(n4516), .B(n10046), .ZN(n10197) );
  XOR2_X1 U11284 ( .A(n10045), .B(n10046), .Z(n10049) );
  OAI21_X1 U11285 ( .B1(n10049), .B2(n10048), .A(n10047), .ZN(n10131) );
  INV_X1 U11286 ( .A(n10067), .ZN(n10050) );
  AOI211_X1 U11287 ( .C1(n10133), .C2(n10050), .A(n10407), .B(n10036), .ZN(
        n10132) );
  NAND2_X1 U11288 ( .A1(n10132), .A2(n10393), .ZN(n10053) );
  AOI22_X1 U11289 ( .A1(n10402), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10051), 
        .B2(n10401), .ZN(n10052) );
  OAI211_X1 U11290 ( .C1(n10054), .C2(n10385), .A(n10053), .B(n10052), .ZN(
        n10055) );
  AOI21_X1 U11291 ( .B1(n10324), .B2(n10131), .A(n10055), .ZN(n10056) );
  OAI21_X1 U11292 ( .B1(n10197), .B2(n10412), .A(n10056), .ZN(P1_U3276) );
  INV_X1 U11293 ( .A(n10057), .ZN(n10058) );
  AOI21_X1 U11294 ( .B1(n10063), .B2(n10059), .A(n10058), .ZN(n10060) );
  INV_X1 U11295 ( .A(n10060), .ZN(n10201) );
  OAI21_X1 U11296 ( .B1(n10063), .B2(n10061), .A(n10062), .ZN(n10064) );
  NAND2_X1 U11297 ( .A1(n10064), .A2(n10399), .ZN(n10066) );
  NAND2_X1 U11298 ( .A1(n10066), .A2(n10065), .ZN(n10137) );
  AOI211_X1 U11299 ( .C1(n10138), .C2(n10068), .A(n10407), .B(n10067), .ZN(
        n10136) );
  NAND2_X1 U11300 ( .A1(n10136), .A2(n10393), .ZN(n10072) );
  INV_X1 U11301 ( .A(n10069), .ZN(n10070) );
  AOI22_X1 U11302 ( .A1(n10402), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10070), 
        .B2(n10401), .ZN(n10071) );
  OAI211_X1 U11303 ( .C1(n6250), .C2(n10385), .A(n10072), .B(n10071), .ZN(
        n10073) );
  AOI21_X1 U11304 ( .B1(n10324), .B2(n10137), .A(n10073), .ZN(n10074) );
  OAI21_X1 U11305 ( .B1(n10201), .B2(n10412), .A(n10074), .ZN(P1_U3277) );
  OAI211_X1 U11306 ( .C1(n10079), .C2(n10503), .A(n10078), .B(n10077), .ZN(
        n10152) );
  MUX2_X1 U11307 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10152), .S(n10528), .Z(
        P1_U3552) );
  INV_X1 U11308 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10084) );
  INV_X1 U11309 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10088) );
  MUX2_X1 U11310 ( .A(n10088), .B(n10164), .S(n10528), .Z(n10089) );
  OAI21_X1 U11311 ( .B1(n10167), .B2(n10145), .A(n10089), .ZN(P1_U3548) );
  AOI21_X1 U11312 ( .B1(n10490), .B2(n10091), .A(n10090), .ZN(n10092) );
  OAI211_X1 U11313 ( .C1(n10094), .C2(n10153), .A(n10093), .B(n10092), .ZN(
        n10168) );
  MUX2_X1 U11314 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10168), .S(n10528), .Z(
        P1_U3547) );
  AOI211_X1 U11315 ( .C1(n10490), .C2(n10097), .A(n10096), .B(n10095), .ZN(
        n10169) );
  MUX2_X1 U11316 ( .A(n10098), .B(n10169), .S(n10528), .Z(n10099) );
  OAI21_X1 U11317 ( .B1(n10172), .B2(n10145), .A(n10099), .ZN(P1_U3546) );
  AOI211_X1 U11318 ( .C1(n10490), .C2(n10102), .A(n10101), .B(n10100), .ZN(
        n10104) );
  AOI211_X1 U11319 ( .C1(n10490), .C2(n10108), .A(n10107), .B(n10106), .ZN(
        n10174) );
  MUX2_X1 U11320 ( .A(n10109), .B(n10174), .S(n10528), .Z(n10110) );
  OAI21_X1 U11321 ( .B1(n10177), .B2(n10145), .A(n10110), .ZN(P1_U3544) );
  INV_X1 U11322 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10114) );
  AOI211_X1 U11323 ( .C1(n10490), .C2(n10113), .A(n10112), .B(n10111), .ZN(
        n10178) );
  MUX2_X1 U11324 ( .A(n10114), .B(n10178), .S(n10528), .Z(n10115) );
  OAI21_X1 U11325 ( .B1(n10181), .B2(n10145), .A(n10115), .ZN(P1_U3543) );
  INV_X1 U11326 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10119) );
  AOI211_X1 U11327 ( .C1(n10490), .C2(n10118), .A(n10117), .B(n10116), .ZN(
        n10182) );
  MUX2_X1 U11328 ( .A(n10119), .B(n10182), .S(n10528), .Z(n10120) );
  OAI21_X1 U11329 ( .B1(n10185), .B2(n10145), .A(n10120), .ZN(P1_U3542) );
  AOI211_X1 U11330 ( .C1(n10490), .C2(n10123), .A(n10122), .B(n10121), .ZN(
        n10186) );
  MUX2_X1 U11331 ( .A(n10124), .B(n10186), .S(n10528), .Z(n10125) );
  OAI21_X1 U11332 ( .B1(n10189), .B2(n10145), .A(n10125), .ZN(P1_U3541) );
  AOI211_X1 U11333 ( .C1(n10490), .C2(n10128), .A(n10127), .B(n10126), .ZN(
        n10190) );
  MUX2_X1 U11334 ( .A(n10129), .B(n10190), .S(n10528), .Z(n10130) );
  OAI21_X1 U11335 ( .B1(n10193), .B2(n10145), .A(n10130), .ZN(P1_U3540) );
  AOI211_X1 U11336 ( .C1(n10490), .C2(n10133), .A(n10132), .B(n10131), .ZN(
        n10194) );
  MUX2_X1 U11337 ( .A(n10134), .B(n10194), .S(n10528), .Z(n10135) );
  OAI21_X1 U11338 ( .B1(n10197), .B2(n10145), .A(n10135), .ZN(P1_U3539) );
  AOI211_X1 U11339 ( .C1(n10490), .C2(n10138), .A(n10137), .B(n10136), .ZN(
        n10198) );
  MUX2_X1 U11340 ( .A(n10139), .B(n10198), .S(n10528), .Z(n10140) );
  OAI21_X1 U11341 ( .B1(n10201), .B2(n10145), .A(n10140), .ZN(P1_U3538) );
  AOI211_X1 U11342 ( .C1(n10490), .C2(n10143), .A(n10142), .B(n10141), .ZN(
        n10202) );
  MUX2_X1 U11343 ( .A(n10253), .B(n10202), .S(n10528), .Z(n10144) );
  OAI21_X1 U11344 ( .B1(n10206), .B2(n10145), .A(n10144), .ZN(P1_U3537) );
  AOI21_X1 U11345 ( .B1(n10490), .B2(n10147), .A(n10146), .ZN(n10148) );
  OAI211_X1 U11346 ( .C1(n10150), .C2(n10153), .A(n10149), .B(n10148), .ZN(
        n10207) );
  MUX2_X1 U11347 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10207), .S(n10528), .Z(
        P1_U3536) );
  MUX2_X1 U11348 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10151), .S(n10510), .Z(
        P1_U3521) );
  MUX2_X1 U11349 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10152), .S(n10510), .Z(
        P1_U3520) );
  NOR2_X1 U11350 ( .A1(n10509), .A2(n10153), .ZN(n10160) );
  NAND2_X1 U11351 ( .A1(n10509), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n10155) );
  NAND2_X1 U11352 ( .A1(n10156), .A2(n10155), .ZN(n10157) );
  AOI21_X1 U11353 ( .B1(n10158), .B2(n10160), .A(n10157), .ZN(n10159) );
  INV_X1 U11354 ( .A(n10159), .ZN(P1_U3518) );
  MUX2_X1 U11355 ( .A(n10165), .B(n10164), .S(n10510), .Z(n10166) );
  OAI21_X1 U11356 ( .B1(n10167), .B2(n10205), .A(n10166), .ZN(P1_U3516) );
  MUX2_X1 U11357 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10168), .S(n10510), .Z(
        P1_U3515) );
  INV_X1 U11358 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10170) );
  MUX2_X1 U11359 ( .A(n10170), .B(n10169), .S(n10510), .Z(n10171) );
  OAI21_X1 U11360 ( .B1(n10172), .B2(n10205), .A(n10171), .ZN(P1_U3514) );
  MUX2_X1 U11361 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10173), .S(n10510), .Z(
        P1_U3513) );
  INV_X1 U11362 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10175) );
  MUX2_X1 U11363 ( .A(n10175), .B(n10174), .S(n10510), .Z(n10176) );
  OAI21_X1 U11364 ( .B1(n10177), .B2(n10205), .A(n10176), .ZN(P1_U3512) );
  MUX2_X1 U11365 ( .A(n10179), .B(n10178), .S(n10510), .Z(n10180) );
  OAI21_X1 U11366 ( .B1(n10181), .B2(n10205), .A(n10180), .ZN(P1_U3511) );
  MUX2_X1 U11367 ( .A(n10183), .B(n10182), .S(n10510), .Z(n10184) );
  OAI21_X1 U11368 ( .B1(n10185), .B2(n10205), .A(n10184), .ZN(P1_U3510) );
  INV_X1 U11369 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10187) );
  MUX2_X1 U11370 ( .A(n10187), .B(n10186), .S(n10510), .Z(n10188) );
  OAI21_X1 U11371 ( .B1(n10189), .B2(n10205), .A(n10188), .ZN(P1_U3509) );
  INV_X1 U11372 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10191) );
  MUX2_X1 U11373 ( .A(n10191), .B(n10190), .S(n10510), .Z(n10192) );
  OAI21_X1 U11374 ( .B1(n10193), .B2(n10205), .A(n10192), .ZN(P1_U3507) );
  INV_X1 U11375 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10195) );
  MUX2_X1 U11376 ( .A(n10195), .B(n10194), .S(n10510), .Z(n10196) );
  OAI21_X1 U11377 ( .B1(n10197), .B2(n10205), .A(n10196), .ZN(P1_U3504) );
  MUX2_X1 U11378 ( .A(n10199), .B(n10198), .S(n10510), .Z(n10200) );
  OAI21_X1 U11379 ( .B1(n10201), .B2(n10205), .A(n10200), .ZN(P1_U3501) );
  MUX2_X1 U11380 ( .A(n10203), .B(n10202), .S(n10510), .Z(n10204) );
  OAI21_X1 U11381 ( .B1(n10206), .B2(n10205), .A(n10204), .ZN(P1_U3498) );
  MUX2_X1 U11382 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10207), .S(n10510), .Z(
        P1_U3495) );
  MUX2_X1 U11383 ( .A(P1_D_REG_1__SCAN_IN), .B(n10210), .S(n10423), .Z(
        P1_U3440) );
  MUX2_X1 U11384 ( .A(P1_D_REG_0__SCAN_IN), .B(n10211), .S(n10423), .Z(
        P1_U3439) );
  INV_X1 U11385 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10213) );
  NAND3_X1 U11386 ( .A1(n10213), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n10215) );
  OAI22_X1 U11387 ( .A1(n10212), .A2(n10215), .B1(n10214), .B2(n10224), .ZN(
        n10216) );
  AOI21_X1 U11388 ( .B1(n9527), .B2(n10217), .A(n10216), .ZN(n10218) );
  INV_X1 U11389 ( .A(n10218), .ZN(P1_U3324) );
  OAI222_X1 U11390 ( .A1(n10224), .A2(n10221), .B1(n8271), .B2(n10220), .C1(
        P1_U3086), .C2(n10219), .ZN(P1_U3325) );
  OAI222_X1 U11391 ( .A1(n10224), .A2(n10223), .B1(n8271), .B2(n10222), .C1(
        n6049), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U11392 ( .A1(n10227), .A2(P1_U3086), .B1(n8271), .B2(n10226), .C1(
        n10225), .C2(n10224), .ZN(P1_U3329) );
  MUX2_X1 U11393 ( .A(n10228), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U11394 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  OAI21_X1 U11395 ( .B1(n10230), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10229), .ZN(
        n10231) );
  XOR2_X1 U11396 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10231), .Z(n10236) );
  AOI22_X1 U11397 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10233), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10234) );
  OAI21_X1 U11398 ( .B1(n10236), .B2(n10235), .A(n10234), .ZN(P1_U3243) );
  INV_X1 U11399 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10251) );
  OAI21_X1 U11400 ( .B1(n10238), .B2(n10237), .A(n10284), .ZN(n10246) );
  OAI21_X1 U11401 ( .B1(n10240), .B2(n10239), .A(n10293), .ZN(n10241) );
  OR2_X1 U11402 ( .A1(n10242), .A2(n10241), .ZN(n10245) );
  NAND2_X1 U11403 ( .A1(n10305), .A2(n10243), .ZN(n10244) );
  OAI211_X1 U11404 ( .C1(n10247), .C2(n10246), .A(n10245), .B(n10244), .ZN(
        n10248) );
  INV_X1 U11405 ( .A(n10248), .ZN(n10250) );
  OAI211_X1 U11406 ( .C1(n10308), .C2(n10251), .A(n10250), .B(n10249), .ZN(
        P1_U3257) );
  AOI211_X1 U11407 ( .C1(n10254), .C2(n10253), .A(n10252), .B(n10299), .ZN(
        n10259) );
  AOI211_X1 U11408 ( .C1(n10257), .C2(n10256), .A(n10255), .B(n10269), .ZN(
        n10258) );
  AOI211_X1 U11409 ( .C1(n10305), .C2(n10260), .A(n10259), .B(n10258), .ZN(
        n10262) );
  OAI211_X1 U11410 ( .C1(n10308), .C2(n10263), .A(n10262), .B(n10261), .ZN(
        P1_U3258) );
  INV_X1 U11411 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10277) );
  XOR2_X1 U11412 ( .A(n10265), .B(n10264), .Z(n10266) );
  NOR2_X1 U11413 ( .A1(n10266), .A2(n10299), .ZN(n10273) );
  INV_X1 U11414 ( .A(n10267), .ZN(n10268) );
  AOI211_X1 U11415 ( .C1(n10271), .C2(n10270), .A(n10269), .B(n10268), .ZN(
        n10272) );
  AOI211_X1 U11416 ( .C1(n10305), .C2(n10274), .A(n10273), .B(n10272), .ZN(
        n10276) );
  OAI211_X1 U11417 ( .C1(n10308), .C2(n10277), .A(n10276), .B(n10275), .ZN(
        P1_U3259) );
  OAI21_X1 U11418 ( .B1(n10280), .B2(n10279), .A(n10278), .ZN(n10281) );
  NAND2_X1 U11419 ( .A1(n10281), .A2(n10293), .ZN(n10289) );
  XNOR2_X1 U11420 ( .A(n10283), .B(n10282), .ZN(n10285) );
  NAND2_X1 U11421 ( .A1(n10285), .A2(n10284), .ZN(n10288) );
  NAND2_X1 U11422 ( .A1(n10305), .A2(n10286), .ZN(n10287) );
  AND3_X1 U11423 ( .A1(n10289), .A2(n10288), .A3(n10287), .ZN(n10291) );
  OAI211_X1 U11424 ( .C1(n10308), .C2(n10292), .A(n10291), .B(n10290), .ZN(
        P1_U3260) );
  OAI211_X1 U11425 ( .C1(n10296), .C2(n10295), .A(n10294), .B(n10293), .ZN(
        n10297) );
  INV_X1 U11426 ( .A(n10297), .ZN(n10303) );
  AOI211_X1 U11427 ( .C1(n10301), .C2(n10300), .A(n10299), .B(n10298), .ZN(
        n10302) );
  AOI211_X1 U11428 ( .C1(n10305), .C2(n10304), .A(n10303), .B(n10302), .ZN(
        n10307) );
  OAI211_X1 U11429 ( .C1(n10308), .C2(n10585), .A(n10307), .B(n10306), .ZN(
        P1_U3261) );
  INV_X1 U11430 ( .A(n10318), .ZN(n10309) );
  NAND3_X1 U11431 ( .A1(n10311), .A2(n10310), .A3(n10309), .ZN(n10312) );
  NAND3_X1 U11432 ( .A1(n10313), .A2(n10399), .A3(n10312), .ZN(n10315) );
  AOI222_X1 U11433 ( .A1(n10317), .A2(n10332), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10402), .C1(n10316), .C2(n10401), .ZN(n10323) );
  XNOR2_X1 U11434 ( .A(n10319), .B(n10318), .ZN(n10501) );
  INV_X1 U11435 ( .A(n8524), .ZN(n10320) );
  OAI211_X1 U11436 ( .C1(n10499), .C2(n5279), .A(n10320), .B(n10390), .ZN(
        n10497) );
  INV_X1 U11437 ( .A(n10497), .ZN(n10321) );
  AOI22_X1 U11438 ( .A1(n10501), .A2(n10394), .B1(n10393), .B2(n10321), .ZN(
        n10322) );
  OAI211_X1 U11439 ( .C1(n10402), .C2(n10498), .A(n10323), .B(n10322), .ZN(
        P1_U3281) );
  OAI21_X1 U11440 ( .B1(n10333), .B2(n10326), .A(n10325), .ZN(n10329) );
  INV_X1 U11441 ( .A(n10327), .ZN(n10328) );
  AOI21_X1 U11442 ( .B1(n10329), .B2(n10399), .A(n10328), .ZN(n10483) );
  INV_X1 U11443 ( .A(n10330), .ZN(n10331) );
  AOI222_X1 U11444 ( .A1(n10335), .A2(n10332), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n10402), .C1(n10331), .C2(n10401), .ZN(n10340) );
  XNOR2_X1 U11445 ( .A(n10334), .B(n10333), .ZN(n10486) );
  OAI21_X1 U11446 ( .B1(n10372), .B2(n6101), .A(n10335), .ZN(n10337) );
  NAND3_X1 U11447 ( .A1(n10337), .A2(n10390), .A3(n10336), .ZN(n10482) );
  INV_X1 U11448 ( .A(n10482), .ZN(n10338) );
  AOI22_X1 U11449 ( .A1(n10486), .A2(n10394), .B1(n10393), .B2(n10338), .ZN(
        n10339) );
  OAI211_X1 U11450 ( .C1(n10402), .C2(n10483), .A(n10340), .B(n10339), .ZN(
        P1_U3283) );
  NAND2_X1 U11451 ( .A1(n10342), .A2(n10341), .ZN(n10362) );
  INV_X1 U11452 ( .A(n10343), .ZN(n10345) );
  OAI21_X1 U11453 ( .B1(n10362), .B2(n10345), .A(n10344), .ZN(n10346) );
  XNOR2_X1 U11454 ( .A(n10346), .B(n10354), .ZN(n10349) );
  INV_X1 U11455 ( .A(n10347), .ZN(n10348) );
  AOI21_X1 U11456 ( .B1(n10349), .B2(n10399), .A(n10348), .ZN(n10477) );
  NOR2_X1 U11457 ( .A1(n10382), .A2(n10350), .ZN(n10351) );
  AOI21_X1 U11458 ( .B1(n10402), .B2(P1_REG2_REG_9__SCAN_IN), .A(n10351), .ZN(
        n10352) );
  OAI21_X1 U11459 ( .B1(n10385), .B2(n6393), .A(n10352), .ZN(n10353) );
  INV_X1 U11460 ( .A(n10353), .ZN(n10361) );
  XNOR2_X1 U11461 ( .A(n10355), .B(n10354), .ZN(n10480) );
  XNOR2_X1 U11462 ( .A(n10372), .B(n6393), .ZN(n10358) );
  INV_X1 U11463 ( .A(n10356), .ZN(n10357) );
  AOI21_X1 U11464 ( .B1(n10358), .B2(n10390), .A(n10357), .ZN(n10476) );
  INV_X1 U11465 ( .A(n10476), .ZN(n10359) );
  AOI22_X1 U11466 ( .A1(n10480), .A2(n10394), .B1(n10393), .B2(n10359), .ZN(
        n10360) );
  OAI211_X1 U11467 ( .C1(n10402), .C2(n10477), .A(n10361), .B(n10360), .ZN(
        P1_U3284) );
  XNOR2_X1 U11468 ( .A(n10362), .B(n10370), .ZN(n10365) );
  INV_X1 U11469 ( .A(n10363), .ZN(n10364) );
  AOI21_X1 U11470 ( .B1(n10365), .B2(n10399), .A(n10364), .ZN(n10471) );
  NOR2_X1 U11471 ( .A1(n10382), .A2(n10366), .ZN(n10367) );
  AOI21_X1 U11472 ( .B1(n10402), .B2(P1_REG2_REG_8__SCAN_IN), .A(n10367), .ZN(
        n10368) );
  OAI21_X1 U11473 ( .B1(n10385), .B2(n4697), .A(n10368), .ZN(n10369) );
  INV_X1 U11474 ( .A(n10369), .ZN(n10376) );
  XNOR2_X1 U11475 ( .A(n10371), .B(n10370), .ZN(n10474) );
  OAI211_X1 U11476 ( .C1(n10373), .C2(n4697), .A(n10372), .B(n10390), .ZN(
        n10470) );
  INV_X1 U11477 ( .A(n10470), .ZN(n10374) );
  AOI22_X1 U11478 ( .A1(n10474), .A2(n10394), .B1(n10393), .B2(n10374), .ZN(
        n10375) );
  OAI211_X1 U11479 ( .C1(n10402), .C2(n10471), .A(n10376), .B(n10375), .ZN(
        P1_U3285) );
  XNOR2_X1 U11480 ( .A(n10377), .B(n10388), .ZN(n10380) );
  INV_X1 U11481 ( .A(n10378), .ZN(n10379) );
  AOI21_X1 U11482 ( .B1(n10380), .B2(n10399), .A(n10379), .ZN(n10447) );
  NOR2_X1 U11483 ( .A1(n10382), .A2(n10381), .ZN(n10383) );
  AOI21_X1 U11484 ( .B1(n10402), .B2(P1_REG2_REG_4__SCAN_IN), .A(n10383), .ZN(
        n10384) );
  OAI21_X1 U11485 ( .B1(n10385), .B2(n10446), .A(n10384), .ZN(n10386) );
  INV_X1 U11486 ( .A(n10386), .ZN(n10396) );
  XNOR2_X1 U11487 ( .A(n10388), .B(n10387), .ZN(n10450) );
  OAI211_X1 U11488 ( .C1(n10391), .C2(n10446), .A(n10390), .B(n10389), .ZN(
        n10445) );
  INV_X1 U11489 ( .A(n10445), .ZN(n10392) );
  AOI22_X1 U11490 ( .A1(n10450), .A2(n10394), .B1(n10393), .B2(n10392), .ZN(
        n10395) );
  OAI211_X1 U11491 ( .C1(n10402), .C2(n10447), .A(n10396), .B(n10395), .ZN(
        P1_U3289) );
  XOR2_X1 U11492 ( .A(n10406), .B(n10397), .Z(n10400) );
  AOI21_X1 U11493 ( .B1(n10400), .B2(n10399), .A(n10398), .ZN(n10434) );
  AOI22_X1 U11494 ( .A1(n10402), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10401), .ZN(n10403) );
  OAI21_X1 U11495 ( .B1(n10385), .B2(n10433), .A(n10403), .ZN(n10404) );
  INV_X1 U11496 ( .A(n10404), .ZN(n10416) );
  XNOR2_X1 U11497 ( .A(n10405), .B(n10406), .ZN(n10437) );
  INV_X1 U11498 ( .A(n10437), .ZN(n10413) );
  AOI21_X1 U11499 ( .B1(n10408), .B2(n6526), .A(n10407), .ZN(n10410) );
  NAND2_X1 U11500 ( .A1(n10410), .A2(n10409), .ZN(n10432) );
  OAI22_X1 U11501 ( .A1(n10413), .A2(n10412), .B1(n10411), .B2(n10432), .ZN(
        n10414) );
  INV_X1 U11502 ( .A(n10414), .ZN(n10415) );
  OAI211_X1 U11503 ( .C1(n10402), .C2(n10434), .A(n10416), .B(n10415), .ZN(
        P1_U3291) );
  AND2_X1 U11504 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10424), .ZN(P1_U3294) );
  NOR2_X1 U11505 ( .A1(n10423), .A2(n10417), .ZN(P1_U3295) );
  AND2_X1 U11506 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10424), .ZN(P1_U3296) );
  AND2_X1 U11507 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10424), .ZN(P1_U3297) );
  AND2_X1 U11508 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10424), .ZN(P1_U3298) );
  AND2_X1 U11509 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10424), .ZN(P1_U3299) );
  AND2_X1 U11510 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10424), .ZN(P1_U3300) );
  NOR2_X1 U11511 ( .A1(n10423), .A2(n10418), .ZN(P1_U3301) );
  NOR2_X1 U11512 ( .A1(n10423), .A2(n10419), .ZN(P1_U3302) );
  AND2_X1 U11513 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10424), .ZN(P1_U3303) );
  AND2_X1 U11514 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10424), .ZN(P1_U3304) );
  NOR2_X1 U11515 ( .A1(n10423), .A2(n10420), .ZN(P1_U3305) );
  AND2_X1 U11516 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10424), .ZN(P1_U3306) );
  AND2_X1 U11517 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10424), .ZN(P1_U3307) );
  AND2_X1 U11518 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10424), .ZN(P1_U3308) );
  AND2_X1 U11519 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10424), .ZN(P1_U3309) );
  NOR2_X1 U11520 ( .A1(n10423), .A2(n10421), .ZN(P1_U3310) );
  AND2_X1 U11521 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10424), .ZN(P1_U3311) );
  AND2_X1 U11522 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10424), .ZN(P1_U3312) );
  AND2_X1 U11523 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10424), .ZN(P1_U3313) );
  AND2_X1 U11524 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10424), .ZN(P1_U3314) );
  AND2_X1 U11525 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10424), .ZN(P1_U3315) );
  NOR2_X1 U11526 ( .A1(n10423), .A2(n10422), .ZN(P1_U3316) );
  AND2_X1 U11527 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10424), .ZN(P1_U3317) );
  AND2_X1 U11528 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10424), .ZN(P1_U3318) );
  AND2_X1 U11529 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10424), .ZN(P1_U3319) );
  AND2_X1 U11530 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10424), .ZN(P1_U3320) );
  AND2_X1 U11531 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10424), .ZN(P1_U3321) );
  AND2_X1 U11532 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10424), .ZN(P1_U3322) );
  AND2_X1 U11533 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10424), .ZN(P1_U3323) );
  AOI22_X1 U11534 ( .A1(n10510), .A2(n10425), .B1(n6127), .B2(n10509), .ZN(
        P1_U3453) );
  INV_X1 U11535 ( .A(n10492), .ZN(n10468) );
  NAND2_X1 U11536 ( .A1(n10426), .A2(n10468), .ZN(n10428) );
  OAI211_X1 U11537 ( .C1(n10429), .C2(n10503), .A(n10428), .B(n10427), .ZN(
        n10430) );
  NOR2_X1 U11538 ( .A1(n10431), .A2(n10430), .ZN(n10512) );
  AOI22_X1 U11539 ( .A1(n10510), .A2(n10512), .B1(n6112), .B2(n10509), .ZN(
        P1_U3456) );
  OAI21_X1 U11540 ( .B1(n10433), .B2(n10503), .A(n10432), .ZN(n10436) );
  INV_X1 U11541 ( .A(n10434), .ZN(n10435) );
  AOI211_X1 U11542 ( .C1(n10437), .C2(n10507), .A(n10436), .B(n10435), .ZN(
        n10514) );
  AOI22_X1 U11543 ( .A1(n10510), .A2(n10514), .B1(n6142), .B2(n10509), .ZN(
        P1_U3459) );
  INV_X1 U11544 ( .A(n10438), .ZN(n10443) );
  INV_X1 U11545 ( .A(n10439), .ZN(n10440) );
  OAI21_X1 U11546 ( .B1(n10441), .B2(n10503), .A(n10440), .ZN(n10442) );
  AOI211_X1 U11547 ( .C1(n10507), .C2(n10444), .A(n10443), .B(n10442), .ZN(
        n10516) );
  AOI22_X1 U11548 ( .A1(n10510), .A2(n10516), .B1(n6154), .B2(n10509), .ZN(
        P1_U3462) );
  OAI21_X1 U11549 ( .B1(n10446), .B2(n10503), .A(n10445), .ZN(n10449) );
  INV_X1 U11550 ( .A(n10447), .ZN(n10448) );
  AOI211_X1 U11551 ( .C1(n10507), .C2(n10450), .A(n10449), .B(n10448), .ZN(
        n10517) );
  AOI22_X1 U11552 ( .A1(n10510), .A2(n10517), .B1(n6166), .B2(n10509), .ZN(
        P1_U3465) );
  INV_X1 U11553 ( .A(n10451), .ZN(n10452) );
  OAI21_X1 U11554 ( .B1(n10453), .B2(n10503), .A(n10452), .ZN(n10456) );
  INV_X1 U11555 ( .A(n10454), .ZN(n10455) );
  AOI211_X1 U11556 ( .C1(n10507), .C2(n10457), .A(n10456), .B(n10455), .ZN(
        n10518) );
  AOI22_X1 U11557 ( .A1(n10510), .A2(n10518), .B1(n6181), .B2(n10509), .ZN(
        P1_U3468) );
  OAI21_X1 U11558 ( .B1(n5079), .B2(n10503), .A(n10458), .ZN(n10460) );
  AOI211_X1 U11559 ( .C1(n10507), .C2(n10461), .A(n10460), .B(n10459), .ZN(
        n10519) );
  AOI22_X1 U11560 ( .A1(n10510), .A2(n10519), .B1(n6107), .B2(n10509), .ZN(
        P1_U3471) );
  INV_X1 U11561 ( .A(n10462), .ZN(n10463) );
  OAI21_X1 U11562 ( .B1(n10464), .B2(n10503), .A(n10463), .ZN(n10466) );
  AOI211_X1 U11563 ( .C1(n10468), .C2(n10467), .A(n10466), .B(n10465), .ZN(
        n10520) );
  INV_X1 U11564 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U11565 ( .A1(n10510), .A2(n10520), .B1(n10469), .B2(n10509), .ZN(
        P1_U3474) );
  OAI21_X1 U11566 ( .B1(n4697), .B2(n10503), .A(n10470), .ZN(n10473) );
  INV_X1 U11567 ( .A(n10471), .ZN(n10472) );
  AOI211_X1 U11568 ( .C1(n10507), .C2(n10474), .A(n10473), .B(n10472), .ZN(
        n10521) );
  INV_X1 U11569 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U11570 ( .A1(n10510), .A2(n10521), .B1(n10475), .B2(n10509), .ZN(
        P1_U3477) );
  OAI21_X1 U11571 ( .B1(n6393), .B2(n10503), .A(n10476), .ZN(n10479) );
  INV_X1 U11572 ( .A(n10477), .ZN(n10478) );
  AOI211_X1 U11573 ( .C1(n10507), .C2(n10480), .A(n10479), .B(n10478), .ZN(
        n10522) );
  INV_X1 U11574 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U11575 ( .A1(n10510), .A2(n10522), .B1(n10481), .B2(n10509), .ZN(
        P1_U3480) );
  OAI211_X1 U11576 ( .C1(n10484), .C2(n10503), .A(n10483), .B(n10482), .ZN(
        n10485) );
  AOI21_X1 U11577 ( .B1(n10486), .B2(n10507), .A(n10485), .ZN(n10523) );
  AOI22_X1 U11578 ( .A1(n10510), .A2(n10523), .B1(n6194), .B2(n10509), .ZN(
        P1_U3483) );
  INV_X1 U11579 ( .A(n10493), .ZN(n10495) );
  AOI211_X1 U11580 ( .C1(n10490), .C2(n10489), .A(n10488), .B(n10487), .ZN(
        n10491) );
  OAI21_X1 U11581 ( .B1(n10493), .B2(n10492), .A(n10491), .ZN(n10494) );
  AOI21_X1 U11582 ( .B1(n10496), .B2(n10495), .A(n10494), .ZN(n10524) );
  AOI22_X1 U11583 ( .A1(n10510), .A2(n10524), .B1(n6212), .B2(n10509), .ZN(
        P1_U3486) );
  OAI211_X1 U11584 ( .C1(n10499), .C2(n10503), .A(n10498), .B(n10497), .ZN(
        n10500) );
  AOI21_X1 U11585 ( .B1(n10501), .B2(n10507), .A(n10500), .ZN(n10525) );
  AOI22_X1 U11586 ( .A1(n10510), .A2(n10525), .B1(n6061), .B2(n10509), .ZN(
        P1_U3489) );
  OAI21_X1 U11587 ( .B1(n10504), .B2(n10503), .A(n10502), .ZN(n10505) );
  AOI211_X1 U11588 ( .C1(n10508), .C2(n10507), .A(n10506), .B(n10505), .ZN(
        n10527) );
  AOI22_X1 U11589 ( .A1(n10510), .A2(n10527), .B1(n6050), .B2(n10509), .ZN(
        P1_U3492) );
  AOI22_X1 U11590 ( .A1(n10528), .A2(n10512), .B1(n10511), .B2(n10526), .ZN(
        P1_U3523) );
  AOI22_X1 U11591 ( .A1(n10528), .A2(n10514), .B1(n10513), .B2(n10526), .ZN(
        P1_U3524) );
  INV_X1 U11592 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U11593 ( .A1(n10528), .A2(n10516), .B1(n10515), .B2(n10526), .ZN(
        P1_U3525) );
  AOI22_X1 U11594 ( .A1(n10528), .A2(n10517), .B1(n7375), .B2(n10526), .ZN(
        P1_U3526) );
  AOI22_X1 U11595 ( .A1(n10528), .A2(n10518), .B1(n6179), .B2(n10526), .ZN(
        P1_U3527) );
  AOI22_X1 U11596 ( .A1(n10528), .A2(n10519), .B1(n7378), .B2(n10526), .ZN(
        P1_U3528) );
  AOI22_X1 U11597 ( .A1(n10528), .A2(n10520), .B1(n7380), .B2(n10526), .ZN(
        P1_U3529) );
  AOI22_X1 U11598 ( .A1(n10528), .A2(n10521), .B1(n7382), .B2(n10526), .ZN(
        P1_U3530) );
  AOI22_X1 U11599 ( .A1(n10528), .A2(n10522), .B1(n6075), .B2(n10526), .ZN(
        P1_U3531) );
  AOI22_X1 U11600 ( .A1(n10528), .A2(n10523), .B1(n7485), .B2(n10526), .ZN(
        P1_U3532) );
  AOI22_X1 U11601 ( .A1(n10528), .A2(n10524), .B1(n6211), .B2(n10526), .ZN(
        P1_U3533) );
  AOI22_X1 U11602 ( .A1(n10528), .A2(n10525), .B1(n6060), .B2(n10526), .ZN(
        P1_U3534) );
  AOI22_X1 U11603 ( .A1(n10528), .A2(n10527), .B1(n8038), .B2(n10526), .ZN(
        P1_U3535) );
  OAI21_X1 U11604 ( .B1(n10530), .B2(n4635), .A(n10529), .ZN(n10553) );
  INV_X1 U11605 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10532) );
  OAI22_X1 U11606 ( .A1(n10533), .A2(n10532), .B1(n4774), .B2(n10531), .ZN(
        n10546) );
  INV_X1 U11607 ( .A(n10553), .ZN(n10545) );
  OAI21_X1 U11608 ( .B1(n10536), .B2(n10535), .A(n10534), .ZN(n10542) );
  OAI22_X1 U11609 ( .A1(n7109), .A2(n10539), .B1(n10538), .B2(n10537), .ZN(
        n10540) );
  AOI21_X1 U11610 ( .B1(n10542), .B2(n10541), .A(n10540), .ZN(n10543) );
  OAI21_X1 U11611 ( .B1(n10545), .B2(n10544), .A(n10543), .ZN(n10551) );
  AOI211_X1 U11612 ( .C1(n10547), .C2(n10553), .A(n10546), .B(n10551), .ZN(
        n10548) );
  AOI22_X1 U11613 ( .A1(n10550), .A2(n10549), .B1(n10548), .B2(n9385), .ZN(
        P2_U3231) );
  NOR2_X1 U11614 ( .A1(n4774), .A2(n10565), .ZN(n10552) );
  AOI211_X1 U11615 ( .C1(n10554), .C2(n10553), .A(n10552), .B(n10551), .ZN(
        n10574) );
  AOI22_X1 U11616 ( .A1(n10573), .A2(n5392), .B1(n10574), .B2(n10571), .ZN(
        P2_U3396) );
  NOR2_X1 U11617 ( .A1(n10555), .A2(n10565), .ZN(n10557) );
  AOI211_X1 U11618 ( .C1(n10562), .C2(n10558), .A(n10557), .B(n10556), .ZN(
        n10575) );
  AOI22_X1 U11619 ( .A1(n10573), .A2(n5425), .B1(n10575), .B2(n10571), .ZN(
        P2_U3399) );
  OAI21_X1 U11620 ( .B1(n10560), .B2(n10565), .A(n10559), .ZN(n10561) );
  AOI21_X1 U11621 ( .B1(n10563), .B2(n10562), .A(n10561), .ZN(n10576) );
  AOI22_X1 U11622 ( .A1(n10573), .A2(n5448), .B1(n10576), .B2(n10571), .ZN(
        P2_U3402) );
  INV_X1 U11623 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10572) );
  INV_X1 U11624 ( .A(n10564), .ZN(n10570) );
  OAI22_X1 U11625 ( .A1(n10568), .A2(n10567), .B1(n10566), .B2(n10565), .ZN(
        n10569) );
  NOR2_X1 U11626 ( .A1(n10570), .A2(n10569), .ZN(n10577) );
  AOI22_X1 U11627 ( .A1(n10573), .A2(n10572), .B1(n10577), .B2(n10571), .ZN(
        P2_U3405) );
  AOI22_X1 U11628 ( .A1(n10578), .A2(n10574), .B1(n7196), .B2(n7168), .ZN(
        P2_U3461) );
  AOI22_X1 U11629 ( .A1(n10578), .A2(n10575), .B1(n5424), .B2(n7168), .ZN(
        P2_U3462) );
  AOI22_X1 U11630 ( .A1(n10578), .A2(n10576), .B1(n7205), .B2(n7168), .ZN(
        P2_U3463) );
  AOI22_X1 U11631 ( .A1(n10578), .A2(n10577), .B1(n5461), .B2(n7168), .ZN(
        P2_U3464) );
  OAI222_X1 U11632 ( .A1(n10583), .A2(n10582), .B1(n10583), .B2(n10581), .C1(
        n10580), .C2(n10579), .ZN(ADD_1068_U5) );
  XOR2_X1 U11633 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11634 ( .B1(n10586), .B2(n10585), .A(n10584), .ZN(n10588) );
  XNOR2_X1 U11635 ( .A(n10588), .B(n10587), .ZN(ADD_1068_U55) );
  OAI21_X1 U11636 ( .B1(n10591), .B2(n10590), .A(n10589), .ZN(ADD_1068_U56) );
  OAI21_X1 U11637 ( .B1(n10594), .B2(n10593), .A(n10592), .ZN(ADD_1068_U57) );
  OAI21_X1 U11638 ( .B1(n10597), .B2(n10596), .A(n10595), .ZN(ADD_1068_U58) );
  OAI21_X1 U11639 ( .B1(n10600), .B2(n10599), .A(n10598), .ZN(ADD_1068_U59) );
  OAI21_X1 U11640 ( .B1(n10603), .B2(n10602), .A(n10601), .ZN(ADD_1068_U60) );
  OAI21_X1 U11641 ( .B1(n10606), .B2(n10605), .A(n10604), .ZN(ADD_1068_U61) );
  OAI21_X1 U11642 ( .B1(n10609), .B2(n10608), .A(n10607), .ZN(ADD_1068_U62) );
  OAI21_X1 U11643 ( .B1(n10612), .B2(n10611), .A(n10610), .ZN(ADD_1068_U63) );
  OAI21_X1 U11644 ( .B1(n10615), .B2(n10614), .A(n10613), .ZN(ADD_1068_U51) );
  OAI21_X1 U11645 ( .B1(n10618), .B2(n10617), .A(n10616), .ZN(ADD_1068_U47) );
  OAI21_X1 U11646 ( .B1(n10621), .B2(n10620), .A(n10619), .ZN(ADD_1068_U49) );
  OAI21_X1 U11647 ( .B1(n10624), .B2(n10623), .A(n10622), .ZN(ADD_1068_U48) );
  OAI21_X1 U11648 ( .B1(n10627), .B2(n10626), .A(n10625), .ZN(ADD_1068_U50) );
  AOI21_X1 U11649 ( .B1(n10630), .B2(n10629), .A(n10628), .ZN(ADD_1068_U54) );
  AOI21_X1 U11650 ( .B1(n10633), .B2(n10632), .A(n10631), .ZN(ADD_1068_U53) );
  OAI21_X1 U11651 ( .B1(n10636), .B2(n10635), .A(n10634), .ZN(ADD_1068_U52) );
  INV_X1 U6188 ( .A(n6543), .ZN(n6538) );
  CLKBUF_X2 U5181 ( .A(n6150), .Z(n4412) );
  NAND2_X1 U5353 ( .A1(n4779), .A2(n6392), .ZN(n10372) );
  CLKBUF_X1 U6677 ( .A(n5660), .Z(n5986) );
  CLKBUF_X2 U7085 ( .A(n5372), .Z(n9540) );
endmodule

