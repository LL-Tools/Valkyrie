

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1,
         READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,
         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,
         n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
         n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
         n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168,
         n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176,
         n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
         n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192,
         n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200,
         n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
         n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216,
         n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224,
         n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232,
         n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240,
         n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
         n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256,
         n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264,
         n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
         n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
         n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288,
         n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296,
         n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304,
         n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
         n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,
         n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
         n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336,
         n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,
         n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
         n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360,
         n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368,
         n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
         n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
         n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,
         n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,
         n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408,
         n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,
         n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
         n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432,
         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,
         n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480,
         n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,
         n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
         n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504,
         n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512,
         n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520,
         n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528,
         n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536,
         n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544,
         n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552,
         n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560,
         n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
         n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576,
         n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584,
         n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592,
         n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600,
         n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608,
         n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616,
         n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624,
         n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
         n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
         n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648,
         n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656,
         n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664,
         n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672,
         n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680,
         n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688,
         n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696,
         n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,
         n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,
         n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720,
         n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728,
         n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736,
         n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744,
         n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752,
         n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,
         n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768,
         n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,
         n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
         n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792,
         n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800,
         n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808,
         n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,
         n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,
         n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
         n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840,
         n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,
         n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
         n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864,
         n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872,
         n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,
         n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888,
         n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,
         n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904,
         n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912,
         n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920,
         n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,
         n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936,
         n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944,
         n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
         n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960,
         n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,
         n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976,
         n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984,
         n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992,
         n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,
         n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008,
         n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016,
         n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
         n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032,
         n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040,
         n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048,
         n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056,
         n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,
         n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,
         n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080,
         n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088,
         n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
         n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104,
         n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,
         n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120,
         n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128,
         n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,
         n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
         n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152,
         n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160,
         n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
         n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176,
         n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184,
         n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192,
         n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200,
         n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208,
         n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
         n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224,
         n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232,
         n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
         n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248,
         n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256,
         n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,
         n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,
         n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280,
         n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
         n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296,
         n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304,
         n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
         n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320,
         n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
         n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,
         n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
         n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,
         n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
         n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368,
         n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
         n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,
         n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392,
         n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,
         n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,
         n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,
         n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424,
         n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432,
         n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440,
         n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448,
         n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456,
         n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464,
         n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472,
         n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480,
         n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488,
         n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496,
         n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504,
         n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512,
         n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520,
         n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528,
         n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536,
         n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544,
         n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552,
         n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560,
         n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568,
         n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576,
         n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584,
         n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592,
         n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600,
         n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608,
         n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616,
         n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624,
         n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632,
         n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640,
         n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648,
         n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656,
         n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664,
         n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672,
         n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680,
         n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688,
         n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696,
         n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704,
         n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712,
         n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,
         n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728,
         n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,
         n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744,
         n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752,
         n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760,
         n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768,
         n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776,
         n22777, n22778, n22779, n22780, n22781, n22782;

  INV_X2 U11255 ( .A(n17281), .ZN(n14651) );
  XNOR2_X1 U11256 ( .A(n17288), .B(n17087), .ZN(n16359) );
  INV_X1 U11257 ( .A(n21269), .ZN(n21232) );
  AND2_X1 U11258 ( .A1(n15835), .A2(n15766), .ZN(n15836) );
  CLKBUF_X1 U11259 ( .A(n12809), .Z(n13518) );
  INV_X1 U11260 ( .A(n20850), .ZN(n21279) );
  NAND2_X2 U11261 ( .A1(n15564), .A2(n12895), .ZN(n16178) );
  OR3_X1 U11262 ( .A1(n15439), .A2(n17172), .A3(n13858), .ZN(n19930) );
  NAND2_X1 U11263 ( .A1(n13853), .A2(n17172), .ZN(n19904) );
  NAND2_X2 U11264 ( .A1(n12993), .A2(n12992), .ZN(n13640) );
  CLKBUF_X2 U11265 ( .A(n11720), .Z(n11843) );
  INV_X2 U11266 ( .A(n12523), .ZN(n12577) );
  CLKBUF_X2 U11267 ( .A(n12576), .Z(n18416) );
  BUF_X2 U11268 ( .A(n12490), .Z(n18467) );
  CLKBUF_X2 U11269 ( .A(n12524), .Z(n18465) );
  CLKBUF_X2 U11270 ( .A(n12521), .Z(n18469) );
  CLKBUF_X2 U11271 ( .A(n12473), .Z(n18474) );
  AND2_X1 U11272 ( .A1(n14617), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12205) );
  CLKBUF_X2 U11273 ( .A(n12936), .Z(n13523) );
  BUF_X1 U11274 ( .A(n12902), .Z(n17039) );
  CLKBUF_X2 U11275 ( .A(n14120), .Z(n20262) );
  INV_X2 U11276 ( .A(n12891), .ZN(n12888) );
  OR2_X1 U11277 ( .A1(n12828), .A2(n12827), .ZN(n15384) );
  AND4_X1 U11278 ( .A1(n12874), .A2(n12873), .A3(n12872), .A4(n12871), .ZN(
        n12880) );
  INV_X1 U11279 ( .A(n12883), .ZN(n15598) );
  NOR2_X1 U11280 ( .A1(n11184), .A2(n11234), .ZN(n11314) );
  CLKBUF_X2 U11281 ( .A(n14633), .Z(n14627) );
  OAI21_X1 U11282 ( .B1(n11935), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11435), .ZN(n11983) );
  AND2_X4 U11283 ( .A1(n12765), .A2(n15430), .ZN(n12803) );
  AND2_X1 U11284 ( .A1(n12762), .A2(n15429), .ZN(n12817) );
  AND2_X1 U11285 ( .A1(n15353), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12763) );
  CLKBUF_X1 U11286 ( .A(n18732), .Z(n11148) );
  NOR3_X1 U11287 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n18840), .A3(n21481), 
        .ZN(n18732) );
  OAI22_X1 U11288 ( .A1(n15561), .A2(n15596), .B1(n20751), .B2(n15595), .ZN(
        n22597) );
  NAND2_X2 U11289 ( .A1(n16731), .A2(n20689), .ZN(n15595) );
  INV_X1 U11290 ( .A(n17839), .ZN(n11149) );
  INV_X1 U11291 ( .A(n11149), .ZN(n11150) );
  INV_X1 U11292 ( .A(n11149), .ZN(n11151) );
  NOR2_X2 U11294 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12765) );
  AND4_X1 U11295 ( .A1(n12798), .A2(n12797), .A3(n12796), .A4(n12795), .ZN(
        n12799) );
  CLKBUF_X2 U11296 ( .A(n11937), .Z(n14617) );
  OR3_X1 U11297 ( .A1(n15439), .A2(n17172), .A3(n13824), .ZN(n13940) );
  INV_X1 U11298 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11936) );
  INV_X1 U11299 ( .A(n18475), .ZN(n18322) );
  AND2_X1 U11300 ( .A1(n12886), .A2(n15330), .ZN(n13659) );
  AND2_X2 U11301 ( .A1(n17059), .A2(n15429), .ZN(n17061) );
  INV_X1 U11302 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12757) );
  OR2_X1 U11303 ( .A1(n17216), .A2(n17215), .ZN(n11594) );
  OR2_X1 U11304 ( .A1(n13829), .A2(n15439), .ZN(n19942) );
  OR2_X1 U11305 ( .A1(n13843), .A2(n17188), .ZN(n19886) );
  AND3_X1 U11306 ( .A1(n12853), .A2(n11319), .A3(n11316), .ZN(n11315) );
  INV_X1 U11308 ( .A(n11670), .ZN(n11667) );
  AND2_X1 U11309 ( .A1(n12895), .A2(n12891), .ZN(n16419) );
  AND2_X2 U11310 ( .A1(n12782), .A2(n12781), .ZN(n15583) );
  NAND2_X1 U11311 ( .A1(n11778), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11785) );
  AOI221_X1 U11312 ( .B1(n11152), .B2(n12520), .C1(n12720), .C2(n21615), .A(
        n12719), .ZN(n18867) );
  INV_X1 U11313 ( .A(n21762), .ZN(n18793) );
  NAND2_X1 U11314 ( .A1(n21279), .A2(n21843), .ZN(n21792) );
  INV_X1 U11315 ( .A(n11166), .ZN(n16400) );
  INV_X1 U11316 ( .A(n22093), .ZN(n22102) );
  BUF_X1 U11317 ( .A(n19178), .Z(n11173) );
  INV_X2 U11318 ( .A(n14120), .ZN(n11354) );
  OAI211_X1 U11319 ( .C1(n17396), .C2(n17395), .A(n17394), .B(n17408), .ZN(
        n17400) );
  NOR2_X1 U11320 ( .A1(n21371), .A2(n18370), .ZN(n18377) );
  INV_X1 U11321 ( .A(n18840), .ZN(n18887) );
  INV_X1 U11322 ( .A(n21792), .ZN(n21898) );
  INV_X1 U11323 ( .A(n22216), .ZN(n22244) );
  NAND2_X1 U11324 ( .A1(n17288), .A2(n17287), .ZN(n19223) );
  INV_X1 U11325 ( .A(n11171), .ZN(n17188) );
  INV_X2 U11326 ( .A(n21868), .ZN(n21886) );
  NAND2_X2 U11327 ( .A1(n12911), .A2(n12907), .ZN(n12982) );
  INV_X1 U11329 ( .A(n14120), .ZN(n11153) );
  OR2_X2 U11330 ( .A1(n17307), .A2(n17308), .ZN(n11209) );
  NOR2_X2 U11331 ( .A1(n16883), .A2(n13784), .ZN(n11405) );
  AOI211_X2 U11332 ( .C1(n20694), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n22031), .B(n20659), .ZN(n20660) );
  NAND2_X2 U11333 ( .A1(n11953), .A2(n11952), .ZN(n14353) );
  AND2_X1 U11334 ( .A1(n17051), .A2(n17059), .ZN(n11154) );
  AND2_X2 U11335 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11792) );
  XNOR2_X2 U11336 ( .A(n14101), .B(n11431), .ZN(n11574) );
  NAND2_X2 U11337 ( .A1(n11347), .A2(n11346), .ZN(n16031) );
  AND2_X4 U11338 ( .A1(n15678), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11975) );
  NAND2_X1 U11339 ( .A1(n12520), .A2(n21330), .ZN(n12717) );
  NAND4_X2 U11340 ( .A1(n12497), .A2(n12496), .A3(n12495), .A4(n11211), .ZN(
        n12520) );
  XNOR2_X2 U11341 ( .A(n12060), .B(n12059), .ZN(n13807) );
  NOR2_X2 U11342 ( .A1(n15953), .A2(n15954), .ZN(n15883) );
  NAND3_X4 U11343 ( .A1(n12637), .A2(n12636), .A3(n12635), .ZN(n21371) );
  XNOR2_X2 U11344 ( .A(n13081), .B(n13080), .ZN(n13696) );
  NAND2_X2 U11345 ( .A1(n12969), .A2(n12968), .ZN(n13081) );
  AOI211_X1 U11346 ( .C1(n22097), .C2(n22118), .A(n22096), .B(n22095), .ZN(
        n22101) );
  NAND2_X1 U11347 ( .A1(n20647), .A2(n13772), .ZN(n16903) );
  AOI221_X1 U11348 ( .B1(P3_REIP_REG_29__SCAN_IN), .B2(n21801), .C1(n21740), 
        .C2(n21868), .A(n21739), .ZN(n21741) );
  AND2_X1 U11349 ( .A1(n17085), .A2(n12190), .ZN(n16323) );
  INV_X1 U11350 ( .A(n18388), .ZN(n18378) );
  INV_X1 U11351 ( .A(n17793), .ZN(n13945) );
  NAND2_X1 U11352 ( .A1(n11692), .A2(n12062), .ZN(n11352) );
  OAI21_X1 U11353 ( .B1(n13808), .B2(n13814), .A(n13815), .ZN(n12048) );
  CLKBUF_X2 U11354 ( .A(n15262), .Z(n15313) );
  NOR2_X1 U11355 ( .A1(n18864), .A2(n12538), .ZN(n12539) );
  INV_X1 U11356 ( .A(n12520), .ZN(n21451) );
  INV_X2 U11357 ( .A(n21371), .ZN(n21438) );
  INV_X1 U11358 ( .A(n14353), .ZN(n11997) );
  CLKBUF_X3 U11359 ( .A(n12205), .Z(n11174) );
  CLKBUF_X2 U11360 ( .A(n13018), .Z(n13574) );
  BUF_X2 U11361 ( .A(n12817), .Z(n13568) );
  BUF_X2 U11362 ( .A(n12818), .Z(n13576) );
  BUF_X2 U11363 ( .A(n13260), .Z(n13569) );
  AND2_X2 U11364 ( .A1(n14630), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11819) );
  BUF_X2 U11365 ( .A(n12955), .Z(n13550) );
  BUF_X2 U11366 ( .A(n12924), .Z(n13567) );
  CLKBUF_X2 U11367 ( .A(n12994), .Z(n13575) );
  CLKBUF_X2 U11368 ( .A(n20521), .Z(n21955) );
  CLKBUF_X2 U11369 ( .A(n12956), .Z(n13577) );
  INV_X2 U11370 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11761) );
  NOR2_X1 U11371 ( .A1(n17470), .A2(n11216), .ZN(n17474) );
  NAND2_X1 U11372 ( .A1(n11407), .A2(n11196), .ZN(n13803) );
  OAI21_X1 U11373 ( .B1(n17499), .B2(n17485), .A(n17498), .ZN(n17486) );
  AOI21_X1 U11374 ( .B1(n16465), .B2(n16462), .A(n16464), .ZN(n16795) );
  AOI211_X1 U11375 ( .C1(n16323), .C2(n17998), .A(n16322), .B(n16321), .ZN(
        n16324) );
  NAND2_X1 U11376 ( .A1(n14319), .A2(n14318), .ZN(n17409) );
  XNOR2_X1 U11377 ( .A(n16330), .B(n13600), .ZN(n16378) );
  NOR2_X1 U11378 ( .A1(n17421), .A2(n14263), .ZN(n14314) );
  NOR2_X1 U11379 ( .A1(n17494), .A2(n17633), .ZN(n17488) );
  NOR2_X1 U11380 ( .A1(n19246), .A2(n17972), .ZN(n17971) );
  NAND2_X1 U11381 ( .A1(n17475), .A2(n11432), .ZN(n17411) );
  AND2_X1 U11382 ( .A1(n17521), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n19274) );
  NAND2_X1 U11383 ( .A1(n11357), .A2(n11355), .ZN(n18006) );
  AND2_X1 U11384 ( .A1(n17716), .A2(n14116), .ZN(n17521) );
  OR2_X1 U11385 ( .A1(n20648), .A2(n16917), .ZN(n20656) );
  NAND2_X1 U11386 ( .A1(n16990), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16827) );
  NAND2_X1 U11387 ( .A1(n11669), .A2(n11665), .ZN(n16990) );
  NAND2_X1 U11388 ( .A1(n16250), .A2(n16249), .ZN(n20647) );
  NAND2_X1 U11389 ( .A1(n17224), .A2(n17226), .ZN(n17225) );
  OAI21_X1 U11390 ( .B1(n13994), .B2(n11454), .A(n11260), .ZN(n11453) );
  NAND2_X1 U11391 ( .A1(n11660), .A2(n11662), .ZN(n16250) );
  XOR2_X1 U11392 ( .A(n17086), .B(n17085), .Z(n17544) );
  AND2_X1 U11393 ( .A1(n14087), .A2(n13989), .ZN(n14106) );
  OR2_X1 U11394 ( .A1(n14104), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16154) );
  OAI211_X1 U11395 ( .C1(n11440), .C2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11439), .B(n11437), .ZN(n17919) );
  AND2_X1 U11396 ( .A1(n17123), .A2(n11609), .ZN(n17199) );
  XNOR2_X1 U11397 ( .A(n13963), .B(n13964), .ZN(n14104) );
  AND2_X1 U11398 ( .A1(n15880), .A2(n11289), .ZN(n16232) );
  OR2_X1 U11399 ( .A1(n12568), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n21765) );
  OR3_X1 U11400 ( .A1(n16909), .A2(n16905), .A3(n16908), .ZN(n20671) );
  NOR2_X2 U11401 ( .A1(n15777), .A2(n15957), .ZN(n15880) );
  NAND2_X1 U11402 ( .A1(n18631), .A2(n21705), .ZN(n21719) );
  OAI21_X1 U11403 ( .B1(n13740), .B2(n13250), .A(n13059), .ZN(n15835) );
  AND2_X1 U11404 ( .A1(n17255), .A2(n11269), .ZN(n17245) );
  OR2_X1 U11405 ( .A1(n13786), .A2(n13773), .ZN(n20670) );
  NAND2_X1 U11406 ( .A1(n11210), .A2(n13131), .ZN(n13744) );
  XNOR2_X1 U11407 ( .A(n13765), .B(n13135), .ZN(n13752) );
  NOR2_X1 U11408 ( .A1(n17278), .A2(n15098), .ZN(n17264) );
  NAND2_X2 U11409 ( .A1(n13765), .A2(n13764), .ZN(n13786) );
  NAND2_X1 U11410 ( .A1(n13039), .A2(n11198), .ZN(n13765) );
  OAI21_X1 U11411 ( .B1(n15962), .B2(n13250), .A(n13101), .ZN(n15606) );
  NAND2_X1 U11412 ( .A1(n18729), .A2(n21762), .ZN(n18596) );
  NAND2_X1 U11413 ( .A1(n13103), .A2(n13093), .ZN(n15962) );
  NAND2_X1 U11414 ( .A1(n13027), .A2(n15539), .ZN(n13103) );
  NAND2_X1 U11415 ( .A1(n13079), .A2(n13078), .ZN(n15444) );
  NOR2_X1 U11416 ( .A1(n21431), .A2(n21430), .ZN(n21429) );
  NOR2_X1 U11417 ( .A1(n19917), .A2(n13844), .ZN(n13849) );
  AND2_X1 U11418 ( .A1(n16552), .A2(n16538), .ZN(n16540) );
  NAND2_X2 U11419 ( .A1(n13071), .A2(n13074), .ZN(n16347) );
  NAND2_X1 U11420 ( .A1(n13820), .A2(n11171), .ZN(n13947) );
  NAND2_X1 U11421 ( .A1(n11723), .A2(n15439), .ZN(n19864) );
  AND2_X1 U11422 ( .A1(n13832), .A2(n13831), .ZN(n17793) );
  NOR2_X1 U11423 ( .A1(n16565), .A2(n16550), .ZN(n16552) );
  OR2_X1 U11424 ( .A1(n13842), .A2(n17172), .ZN(n13931) );
  AND2_X1 U11425 ( .A1(n11555), .A2(n11556), .ZN(n18553) );
  CLKBUF_X1 U11426 ( .A(n13676), .Z(n16779) );
  NAND2_X1 U11427 ( .A1(n14366), .A2(n14361), .ZN(n15066) );
  NAND2_X1 U11428 ( .A1(n14365), .A2(n14364), .ZN(n15065) );
  NAND2_X1 U11429 ( .A1(n14371), .A2(n14370), .ZN(n14374) );
  NAND2_X1 U11430 ( .A1(n13026), .A2(n13025), .ZN(n15539) );
  CLKBUF_X3 U11431 ( .A(n14362), .Z(n11171) );
  NOR2_X1 U11432 ( .A1(n21102), .A2(n18447), .ZN(n18462) );
  AND2_X1 U11433 ( .A1(n11621), .A2(n11620), .ZN(n11619) );
  XNOR2_X1 U11434 ( .A(n13823), .B(n13819), .ZN(n14362) );
  OR2_X1 U11435 ( .A1(n13697), .A2(n12950), .ZN(n12976) );
  NAND2_X2 U11436 ( .A1(n15798), .A2(n15797), .ZN(n22190) );
  NAND2_X1 U11437 ( .A1(n11335), .A2(n13807), .ZN(n11692) );
  CLKBUF_X1 U11438 ( .A(n16723), .Z(n20623) );
  NAND2_X1 U11439 ( .A1(n12048), .A2(n12047), .ZN(n11335) );
  NAND2_X1 U11440 ( .A1(n13818), .A2(n13813), .ZN(n19023) );
  NAND2_X1 U11441 ( .A1(n21894), .A2(n11323), .ZN(n12740) );
  CLKBUF_X1 U11442 ( .A(n14117), .Z(n18010) );
  XNOR2_X1 U11443 ( .A(n13817), .B(n13816), .ZN(n13823) );
  NAND2_X2 U11444 ( .A1(n17879), .A2(n15370), .ZN(n20696) );
  INV_X2 U11445 ( .A(n20790), .ZN(n20844) );
  NOR2_X2 U11446 ( .A1(n20259), .A2(n20205), .ZN(n20206) );
  NOR2_X2 U11447 ( .A1(n20259), .A2(n20258), .ZN(n20260) );
  NOR2_X2 U11448 ( .A1(n20259), .A2(n20163), .ZN(n16029) );
  NOR2_X2 U11449 ( .A1(n20259), .A2(n20069), .ZN(n20070) );
  NOR2_X2 U11450 ( .A1(n20259), .A2(n20110), .ZN(n20111) );
  NOR2_X2 U11451 ( .A1(n20259), .A2(n20022), .ZN(n20023) );
  NOR2_X2 U11452 ( .A1(n16371), .A2(n22265), .ZN(n15370) );
  XNOR2_X1 U11453 ( .A(n12543), .B(n12544), .ZN(n18832) );
  NOR2_X2 U11454 ( .A1(n20259), .A2(n19833), .ZN(n19834) );
  INV_X1 U11455 ( .A(n13815), .ZN(n13816) );
  XNOR2_X1 U11456 ( .A(n12072), .B(n12074), .ZN(n13806) );
  AND2_X1 U11457 ( .A1(n21893), .A2(n11324), .ZN(n11323) );
  NAND2_X1 U11458 ( .A1(n11322), .A2(n13655), .ZN(n16371) );
  NAND2_X1 U11459 ( .A1(n21279), .A2(n12702), .ZN(n21927) );
  NAND2_X1 U11460 ( .A1(n12058), .A2(n12057), .ZN(n12059) );
  NAND2_X1 U11461 ( .A1(n15215), .A2(n15214), .ZN(n15213) );
  AND3_X1 U11462 ( .A1(n12043), .A2(n12042), .A3(n12041), .ZN(n13814) );
  OAI21_X1 U11463 ( .B1(n13653), .B2(n11285), .A(n13654), .ZN(n11322) );
  AND2_X1 U11464 ( .A1(n12410), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12414) );
  NAND2_X1 U11465 ( .A1(n15701), .A2(n12039), .ZN(n14180) );
  INV_X1 U11466 ( .A(n18490), .ZN(n18489) );
  AND2_X1 U11467 ( .A1(n12038), .A2(n11608), .ZN(n15701) );
  NAND2_X1 U11468 ( .A1(n11397), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12911) );
  XNOR2_X1 U11469 ( .A(n12539), .B(n21564), .ZN(n18856) );
  NOR2_X1 U11470 ( .A1(n15464), .A2(n15465), .ZN(n15825) );
  INV_X2 U11471 ( .A(n12069), .ZN(n12160) );
  INV_X1 U11472 ( .A(n12033), .ZN(n15644) );
  AOI21_X1 U11473 ( .B1(n18109), .B2(n18108), .A(n21948), .ZN(n21277) );
  NOR2_X1 U11474 ( .A1(n11546), .A2(n12746), .ZN(n11545) );
  OR2_X1 U11475 ( .A1(n12051), .A2(n11814), .ZN(n12045) );
  INV_X1 U11476 ( .A(n18844), .ZN(n11562) );
  OR2_X1 U11477 ( .A1(n21472), .A2(n21470), .ZN(n12746) );
  AND4_X1 U11478 ( .A1(n12233), .A2(n12232), .A3(n12231), .A4(n12230), .ZN(
        n16057) );
  NOR2_X1 U11479 ( .A1(n21335), .A2(n19470), .ZN(n12692) );
  AND3_X1 U11480 ( .A1(n11997), .A2(n12004), .A3(n11998), .ZN(n15157) );
  NAND2_X1 U11481 ( .A1(n13640), .A2(n13623), .ZN(n13655) );
  AND2_X1 U11482 ( .A1(n12917), .A2(n15319), .ZN(n12904) );
  NAND2_X1 U11483 ( .A1(n12021), .A2(n11988), .ZN(n15707) );
  OR2_X1 U11484 ( .A1(n13686), .A2(n16435), .ZN(n12917) );
  AND2_X1 U11485 ( .A1(n11607), .A2(n14152), .ZN(n12021) );
  OR2_X1 U11486 ( .A1(n13660), .A2(n12884), .ZN(n15382) );
  AND2_X1 U11487 ( .A1(n11343), .A2(n11341), .ZN(n12004) );
  NAND4_X1 U11488 ( .A1(n20112), .A2(n19835), .A3(n11720), .A4(n11997), .ZN(
        n14195) );
  INV_X1 U11489 ( .A(n14146), .ZN(n20207) );
  OR2_X1 U11490 ( .A1(n11825), .A2(n11824), .ZN(n14093) );
  INV_X1 U11491 ( .A(n12006), .ZN(n19835) );
  AND2_X1 U11492 ( .A1(n12017), .A2(n12010), .ZN(n14156) );
  CLKBUF_X2 U11493 ( .A(n16435), .Z(n11166) );
  NAND2_X1 U11494 ( .A1(n11345), .A2(n11344), .ZN(n14146) );
  NOR2_X1 U11495 ( .A1(n12006), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12192) );
  NAND2_X1 U11496 ( .A1(n13915), .A2(n12215), .ZN(n12334) );
  AND2_X2 U11497 ( .A1(n12888), .A2(n12895), .ZN(n21956) );
  AND2_X2 U11498 ( .A1(n12006), .A2(n12009), .ZN(n15161) );
  NAND2_X1 U11499 ( .A1(n11552), .A2(n11373), .ZN(n21330) );
  NAND2_X1 U11500 ( .A1(n11721), .A2(n14353), .ZN(n12014) );
  NOR2_X2 U11501 ( .A1(n12883), .A2(n15384), .ZN(n17062) );
  INV_X1 U11502 ( .A(n12009), .ZN(n11721) );
  CLKBUF_X1 U11503 ( .A(n12894), .Z(n15381) );
  INV_X1 U11504 ( .A(n12894), .ZN(n15570) );
  INV_X1 U11505 ( .A(n11983), .ZN(n14149) );
  INV_X1 U11506 ( .A(n12885), .ZN(n16726) );
  NAND2_X1 U11507 ( .A1(n11813), .A2(n11812), .ZN(n12009) );
  NAND4_X2 U11508 ( .A1(n12802), .A2(n12801), .A3(n12800), .A4(n12799), .ZN(
        n12894) );
  INV_X2 U11509 ( .A(U212), .ZN(n11155) );
  INV_X2 U11510 ( .A(n14154), .ZN(n11156) );
  AND2_X1 U11511 ( .A1(n12862), .A2(n12850), .ZN(n11313) );
  NAND2_X2 U11512 ( .A1(U214), .A2(n20711), .ZN(n20777) );
  NAND2_X1 U11513 ( .A1(n11229), .A2(n11436), .ZN(n11435) );
  AOI21_X1 U11514 ( .B1(n12818), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n12764), .ZN(n12767) );
  AND4_X1 U11515 ( .A1(n12866), .A2(n12865), .A3(n12864), .A4(n12863), .ZN(
        n12882) );
  AND4_X1 U11516 ( .A1(n12794), .A2(n12793), .A3(n12792), .A4(n12791), .ZN(
        n12800) );
  AND4_X1 U11517 ( .A1(n12858), .A2(n12857), .A3(n12856), .A4(n12855), .ZN(
        n12862) );
  AND4_X1 U11518 ( .A1(n12790), .A2(n12789), .A3(n12788), .A4(n12787), .ZN(
        n12801) );
  AND4_X1 U11519 ( .A1(n11944), .A2(n11943), .A3(n11942), .A4(n11936), .ZN(
        n11946) );
  AND4_X1 U11520 ( .A1(n12775), .A2(n12774), .A3(n12773), .A4(n12772), .ZN(
        n12782) );
  AND4_X1 U11521 ( .A1(n11805), .A2(n11804), .A3(n11803), .A4(n11802), .ZN(
        n11806) );
  AND4_X1 U11522 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n11778) );
  AND4_X1 U11523 ( .A1(n12878), .A2(n12877), .A3(n12876), .A4(n12875), .ZN(
        n12879) );
  BUF_X2 U11524 ( .A(n12521), .Z(n11167) );
  INV_X2 U11525 ( .A(n20544), .ZN(n11157) );
  INV_X2 U11526 ( .A(n15643), .ZN(n11786) );
  CLKBUF_X2 U11527 ( .A(n11960), .Z(n14613) );
  NAND2_X2 U11528 ( .A1(n22306), .A2(n22320), .ZN(n18099) );
  NAND2_X2 U11529 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n22306), .ZN(n18096) );
  BUF_X2 U11530 ( .A(n12475), .Z(n18476) );
  NOR2_X1 U11531 ( .A1(n20000), .A2(n19845), .ZN(n20325) );
  AND2_X1 U11532 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12764) );
  BUF_X2 U11533 ( .A(n12803), .Z(n13413) );
  CLKBUF_X3 U11534 ( .A(n12476), .Z(n18454) );
  INV_X1 U11535 ( .A(n22276), .ZN(n17839) );
  BUF_X4 U11536 ( .A(n12498), .Z(n11158) );
  NOR2_X1 U11537 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14497) );
  BUF_X2 U11538 ( .A(n11773), .Z(n14636) );
  BUF_X4 U11539 ( .A(n11773), .Z(n14630) );
  NAND2_X1 U11540 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21492), .ZN(
        n12443) );
  NAND3_X2 U11541 ( .A1(n21939), .A2(n20846), .A3(n21937), .ZN(n21868) );
  NAND2_X1 U11542 ( .A1(n20877), .A2(n21491), .ZN(n12445) );
  NAND2_X1 U11543 ( .A1(n21460), .A2(n21492), .ZN(n20849) );
  NAND2_X1 U11544 ( .A1(n20877), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12444) );
  INV_X1 U11545 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11762) );
  INV_X2 U11546 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21492) );
  AND2_X2 U11547 ( .A1(n11170), .A2(n11936), .ZN(n14479) );
  AND2_X1 U11548 ( .A1(n17905), .A2(n13838), .ZN(n11723) );
  AND2_X1 U11549 ( .A1(n16474), .A2(n11688), .ZN(n16330) );
  NAND2_X2 U11550 ( .A1(n15875), .A2(n12991), .ZN(n16674) );
  XNOR2_X1 U11551 ( .A(n12912), .B(n12978), .ZN(n15609) );
  NOR2_X2 U11552 ( .A1(n16716), .A2(n16715), .ZN(n16714) );
  NAND3_X4 U11553 ( .A1(n11313), .A2(n11314), .A3(n11315), .ZN(n12895) );
  NOR2_X1 U11554 ( .A1(n18491), .A2(n18378), .ZN(n11159) );
  OR2_X2 U11555 ( .A1(n17343), .A2(n17137), .ZN(n17139) );
  NAND2_X2 U11556 ( .A1(n15491), .A2(n15503), .ZN(n17689) );
  CLKBUF_X1 U11557 ( .A(n15981), .Z(n11160) );
  CLKBUF_X1 U11558 ( .A(n16013), .Z(n11161) );
  AND2_X1 U11559 ( .A1(n16835), .A2(n20676), .ZN(n11162) );
  NOR2_X1 U11560 ( .A1(n11162), .A2(n16834), .ZN(n16836) );
  CLKBUF_X1 U11561 ( .A(n15359), .Z(n11163) );
  INV_X1 U11562 ( .A(n17885), .ZN(n11164) );
  XNOR2_X1 U11563 ( .A(n20628), .B(n13703), .ZN(n15359) );
  OAI21_X2 U11564 ( .B1(n17915), .B2(n14099), .A(n17913), .ZN(n14101) );
  AND2_X2 U11565 ( .A1(n17054), .A2(n12763), .ZN(n13260) );
  INV_X1 U11566 ( .A(n12911), .ZN(n12978) );
  NOR2_X4 U11567 ( .A1(n16712), .A2(n11679), .ZN(n16578) );
  NAND2_X2 U11568 ( .A1(n11406), .A2(n11405), .ZN(n16876) );
  XNOR2_X2 U11569 ( .A(n20658), .B(n20657), .ZN(n22029) );
  NAND2_X2 U11570 ( .A1(n16819), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16821) );
  OAI21_X2 U11571 ( .B1(n13792), .B2(n11667), .A(n13791), .ZN(n16819) );
  NAND2_X1 U11572 ( .A1(n12891), .A2(n15384), .ZN(n16435) );
  BUF_X1 U11573 ( .A(n12890), .Z(n12914) );
  NOR2_X2 U11574 ( .A1(n16139), .A2(n11214), .ZN(n15424) );
  AND2_X2 U11575 ( .A1(n15191), .A2(n12244), .ZN(n16139) );
  XNOR2_X1 U11576 ( .A(n13724), .B(n13719), .ZN(n15818) );
  NAND2_X1 U11577 ( .A1(n13718), .A2(n13717), .ZN(n13724) );
  OAI21_X2 U11578 ( .B1(n13696), .B2(n13762), .A(n13695), .ZN(n20627) );
  NAND2_X2 U11579 ( .A1(n20627), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20628) );
  NOR2_X2 U11580 ( .A1(n15492), .A2(n15493), .ZN(n15491) );
  AND2_X2 U11581 ( .A1(n16484), .A2(n16485), .ZN(n16474) );
  NOR2_X2 U11582 ( .A1(n16497), .A2(n16499), .ZN(n16484) );
  AND2_X1 U11583 ( .A1(n17051), .A2(n17059), .ZN(n11168) );
  AND2_X1 U11584 ( .A1(n17051), .A2(n17059), .ZN(n12809) );
  BUF_X4 U11585 ( .A(n12609), .Z(n18329) );
  AND2_X1 U11586 ( .A1(n15678), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11169) );
  AND2_X4 U11587 ( .A1(n15678), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11170) );
  NOR2_X4 U11588 ( .A1(n16566), .A2(n16568), .ZN(n16547) );
  AND2_X4 U11589 ( .A1(n11786), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14460) );
  NAND2_X2 U11590 ( .A1(n13273), .A2(n13272), .ZN(n16712) );
  OAI22_X1 U11592 ( .A1(n17403), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n17901), 
        .B2(n17083), .ZN(n19178) );
  AND2_X4 U11593 ( .A1(n15161), .A2(n12215), .ZN(n12321) );
  AND2_X1 U11594 ( .A1(n14120), .A2(n14346), .ZN(n12215) );
  AND2_X2 U11595 ( .A1(n16225), .A2(n11685), .ZN(n16647) );
  NOR2_X4 U11596 ( .A1(n16224), .A2(n16223), .ZN(n16225) );
  AND2_X1 U11597 ( .A1(n17059), .A2(n15429), .ZN(n11175) );
  AND2_X2 U11598 ( .A1(n17059), .A2(n15429), .ZN(n11176) );
  INV_X1 U11599 ( .A(n16031), .ZN(n11343) );
  OAI21_X1 U11600 ( .B1(n11221), .B2(n13786), .A(n16821), .ZN(n11407) );
  AND2_X1 U11601 ( .A1(n13786), .A2(n16965), .ZN(n11408) );
  NAND2_X1 U11602 ( .A1(n14175), .A2(n19341), .ZN(n14215) );
  AND4_X1 U11603 ( .A1(n14172), .A2(n15658), .A3(n14171), .A4(n14170), .ZN(
        n14173) );
  NAND2_X1 U11604 ( .A1(n11325), .A2(n21919), .ZN(n21894) );
  NAND2_X1 U11605 ( .A1(n21927), .A2(n12701), .ZN(n11325) );
  AOI21_X1 U11606 ( .B1(n14749), .B2(n14750), .A(n11280), .ZN(n11483) );
  NAND2_X1 U11607 ( .A1(n12005), .A2(n11233), .ZN(n11363) );
  NOR2_X1 U11608 ( .A1(n12050), .A2(n17901), .ZN(n11364) );
  NAND2_X1 U11609 ( .A1(n11841), .A2(n11840), .ZN(n11858) );
  NAND2_X1 U11610 ( .A1(n12894), .A2(n12842), .ZN(n12843) );
  AND4_X1 U11611 ( .A1(n13861), .A2(n11354), .A3(n13860), .A4(n13859), .ZN(
        n13862) );
  AND2_X1 U11612 ( .A1(n16031), .A2(n12006), .ZN(n14152) );
  NOR2_X1 U11613 ( .A1(n21326), .A2(n12717), .ZN(n12519) );
  NAND2_X1 U11614 ( .A1(n11588), .A2(n11587), .ZN(n12716) );
  INV_X1 U11615 ( .A(n21330), .ZN(n11587) );
  NAND2_X1 U11616 ( .A1(n12520), .A2(n11152), .ZN(n11588) );
  INV_X1 U11617 ( .A(n19592), .ZN(n11334) );
  NOR2_X1 U11618 ( .A1(n17039), .A2(n22256), .ZN(n13561) );
  NAND2_X1 U11619 ( .A1(n16619), .A2(n11684), .ZN(n11683) );
  INV_X1 U11620 ( .A(n16713), .ZN(n11684) );
  OR2_X1 U11621 ( .A1(n12842), .A2(n22489), .ZN(n13065) );
  NAND2_X1 U11622 ( .A1(n13777), .A2(n11236), .ZN(n11673) );
  OAI21_X1 U11623 ( .B1(n15964), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12935), 
        .ZN(n13697) );
  NAND2_X1 U11624 ( .A1(n22384), .A2(n22256), .ZN(n13026) );
  NOR2_X1 U11625 ( .A1(n14055), .A2(n14054), .ZN(n14053) );
  INV_X1 U11626 ( .A(n11342), .ZN(n11341) );
  NOR2_X1 U11627 ( .A1(n17104), .A2(n14324), .ZN(n14315) );
  NAND2_X1 U11628 ( .A1(n14269), .A2(n11704), .ZN(n11702) );
  AND2_X1 U11629 ( .A1(n12002), .A2(n11354), .ZN(n12183) );
  NOR2_X1 U11630 ( .A1(n17703), .A2(n11735), .ZN(n11734) );
  INV_X1 U11631 ( .A(n17704), .ZN(n11733) );
  INV_X2 U11632 ( .A(n12066), .ZN(n12181) );
  NAND2_X1 U11633 ( .A1(n11718), .A2(n11717), .ZN(n11722) );
  AOI21_X1 U11634 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n17832), .A(
        n12664), .ZN(n12672) );
  OR2_X1 U11635 ( .A1(n18771), .A2(n21829), .ZN(n12558) );
  OAI21_X1 U11636 ( .B1(n18811), .B2(n18810), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12733) );
  NAND2_X1 U11637 ( .A1(n12535), .A2(n12717), .ZN(n12537) );
  NOR2_X1 U11638 ( .A1(n11380), .A2(n21459), .ZN(n12687) );
  NOR2_X1 U11639 ( .A1(n11382), .A2(n11381), .ZN(n11380) );
  NAND2_X1 U11640 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16298) );
  INV_X1 U11641 ( .A(n13065), .ZN(n13599) );
  AND2_X1 U11642 ( .A1(n11690), .A2(n11689), .ZN(n11688) );
  INV_X1 U11643 ( .A(n16331), .ZN(n11689) );
  NOR2_X1 U11644 ( .A1(n16347), .A2(n15614), .ZN(n22380) );
  OR2_X1 U11645 ( .A1(n16347), .A2(n13696), .ZN(n22486) );
  NOR2_X1 U11646 ( .A1(n15707), .A2(n15129), .ZN(n12002) );
  NAND2_X1 U11647 ( .A1(n14251), .A2(n14252), .ZN(n14261) );
  AND2_X1 U11648 ( .A1(n14382), .A2(n15882), .ZN(n11579) );
  NAND2_X1 U11649 ( .A1(n12707), .A2(n12702), .ZN(n21893) );
  NAND2_X1 U11650 ( .A1(n18642), .A2(n11746), .ZN(n18653) );
  NAND3_X1 U11651 ( .A1(n12647), .A2(n12646), .A3(n12645), .ZN(n20850) );
  AOI211_X1 U11652 ( .C1(n18477), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n12644), .B(n12643), .ZN(n12645) );
  AND2_X1 U11653 ( .A1(n12568), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18662) );
  AOI21_X1 U11654 ( .B1(n18771), .B2(n11563), .A(n18793), .ZN(n12560) );
  NOR2_X1 U11655 ( .A1(n11564), .A2(n11565), .ZN(n11563) );
  INV_X1 U11656 ( .A(n12551), .ZN(n11564) );
  NAND2_X1 U11657 ( .A1(n11566), .A2(n12554), .ZN(n11565) );
  INV_X1 U11658 ( .A(n21925), .ZN(n21912) );
  AND2_X1 U11659 ( .A1(n21924), .A2(n11386), .ZN(n11385) );
  AND2_X1 U11660 ( .A1(n21923), .A2(n21922), .ZN(n11386) );
  AND2_X1 U11661 ( .A1(n22190), .A2(n15799), .ZN(n22215) );
  OAI21_X1 U11662 ( .B1(n17544), .B2(n19285), .A(n11641), .ZN(n11640) );
  NOR2_X1 U11663 ( .A1(n11253), .A2(n11642), .ZN(n11641) );
  OAI21_X1 U11664 ( .B1(n14334), .B2(n17083), .A(n17543), .ZN(n11642) );
  XNOR2_X1 U11665 ( .A(n15066), .B(n15065), .ZN(n19860) );
  NAND2_X1 U11666 ( .A1(n11504), .A2(n11503), .ZN(n11502) );
  AND2_X1 U11667 ( .A1(n14664), .A2(n14663), .ZN(n11503) );
  OAI21_X1 U11668 ( .B1(n11506), .B2(n11505), .A(n14665), .ZN(n11504) );
  XNOR2_X1 U11669 ( .A(n14661), .B(DATAI_27_), .ZN(n14664) );
  AOI22_X1 U11670 ( .A1(n15597), .A2(n14666), .B1(keyinput_134), .B2(DATAI_26_), .ZN(n11501) );
  NAND2_X1 U11671 ( .A1(n11500), .A2(n11499), .ZN(n11498) );
  NAND2_X1 U11672 ( .A1(keyinput_135), .A2(DATAI_25_), .ZN(n11499) );
  NAND2_X1 U11673 ( .A1(n15588), .A2(n14667), .ZN(n11500) );
  NAND2_X1 U11674 ( .A1(n11531), .A2(n14680), .ZN(n11530) );
  NAND2_X1 U11675 ( .A1(n14676), .A2(n14675), .ZN(n11531) );
  INV_X1 U11676 ( .A(n14679), .ZN(n11529) );
  NAND2_X1 U11677 ( .A1(n22779), .A2(keyinput_169), .ZN(n11534) );
  NAND2_X1 U11678 ( .A1(n14729), .A2(P1_M_IO_N_REG_SCAN_IN), .ZN(n11533) );
  NAND2_X1 U11679 ( .A1(n14723), .A2(n14722), .ZN(n11537) );
  AND2_X1 U11680 ( .A1(n14728), .A2(n11288), .ZN(n11535) );
  NAND2_X1 U11681 ( .A1(keyinput_167), .A2(P1_ADS_N_REG_SCAN_IN), .ZN(n11536)
         );
  NAND2_X1 U11682 ( .A1(n11514), .A2(n11513), .ZN(n14746) );
  AND2_X1 U11683 ( .A1(n14739), .A2(n14738), .ZN(n11513) );
  OAI21_X1 U11684 ( .B1(n11519), .B2(n11516), .A(n11515), .ZN(n11514) );
  NAND2_X1 U11685 ( .A1(n11483), .A2(n11481), .ZN(n11480) );
  INV_X1 U11686 ( .A(n14768), .ZN(n11488) );
  NAND2_X1 U11687 ( .A1(keyinput_201), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(
        n11491) );
  NAND2_X1 U11688 ( .A1(n17793), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13833) );
  OAI21_X1 U11689 ( .B1(n14813), .B2(n14812), .A(n11497), .ZN(n11496) );
  AND2_X1 U11690 ( .A1(n14811), .A2(n14810), .ZN(n11497) );
  AND2_X1 U11691 ( .A1(n11976), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11923) );
  BUF_X1 U11692 ( .A(n12848), .Z(n13548) );
  NAND2_X1 U11693 ( .A1(n12841), .A2(n12840), .ZN(n12845) );
  NAND2_X1 U11694 ( .A1(n12952), .A2(n12953), .ZN(n12923) );
  AND2_X1 U11695 ( .A1(n14027), .A2(n11424), .ZN(n14043) );
  AND2_X1 U11696 ( .A1(n11426), .A2(n11425), .ZN(n11424) );
  INV_X1 U11697 ( .A(n14044), .ZN(n11425) );
  AND2_X1 U11698 ( .A1(n11254), .A2(n14038), .ZN(n11426) );
  AOI21_X1 U11699 ( .B1(n14195), .B2(n11343), .A(n14154), .ZN(n12012) );
  AND2_X1 U11700 ( .A1(n14231), .A2(n11359), .ZN(n11358) );
  NAND2_X1 U11701 ( .A1(n11731), .A2(n17685), .ZN(n11359) );
  INV_X1 U11702 ( .A(n14235), .ZN(n11356) );
  NOR2_X1 U11703 ( .A1(n11737), .A2(n17703), .ZN(n11736) );
  INV_X1 U11704 ( .A(n14016), .ZN(n11737) );
  AND2_X1 U11705 ( .A1(n13985), .A2(n13984), .ZN(n14108) );
  NAND2_X1 U11706 ( .A1(n11366), .A2(n14089), .ZN(n13963) );
  INV_X1 U11707 ( .A(n14088), .ZN(n11366) );
  AOI21_X1 U11708 ( .B1(n12071), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n12046), .ZN(n13815) );
  AND2_X1 U11709 ( .A1(n14120), .A2(n14353), .ZN(n11719) );
  NAND2_X1 U11710 ( .A1(n11985), .A2(n11984), .ZN(n12018) );
  NOR2_X1 U11711 ( .A1(n13426), .A2(n13398), .ZN(n11675) );
  INV_X1 U11712 ( .A(n16580), .ZN(n13361) );
  NOR2_X1 U11713 ( .A1(n11682), .A2(n11683), .ZN(n11681) );
  INV_X1 U11714 ( .A(n16608), .ZN(n11682) );
  NOR2_X1 U11715 ( .A1(n11637), .A2(n16501), .ZN(n11636) );
  INV_X1 U11716 ( .A(n11638), .ZN(n11637) );
  NOR2_X1 U11717 ( .A1(n11626), .A2(n16596), .ZN(n11625) );
  INV_X1 U11718 ( .A(n11627), .ZN(n11626) );
  OR2_X1 U11719 ( .A1(n16257), .A2(n11633), .ZN(n11632) );
  INV_X1 U11720 ( .A(n16721), .ZN(n11633) );
  NOR2_X1 U11721 ( .A1(n11661), .A2(n11659), .ZN(n11658) );
  INV_X1 U11722 ( .A(n16202), .ZN(n11661) );
  INV_X1 U11723 ( .A(n16169), .ZN(n11659) );
  AND2_X1 U11724 ( .A1(n16182), .A2(n16181), .ZN(n16183) );
  NAND2_X1 U11725 ( .A1(n16419), .A2(n11165), .ZN(n16430) );
  INV_X1 U11726 ( .A(n13708), .ZN(n13698) );
  AND2_X1 U11727 ( .A1(n15936), .A2(n13009), .ZN(n22446) );
  AND2_X1 U11728 ( .A1(n14163), .A2(n14162), .ZN(n14184) );
  NOR2_X1 U11729 ( .A1(n11421), .A2(n11277), .ZN(n11420) );
  NAND2_X1 U11730 ( .A1(n14043), .A2(n14047), .ZN(n14055) );
  NAND2_X1 U11731 ( .A1(n14027), .A2(n11426), .ZN(n14045) );
  NOR2_X1 U11732 ( .A1(n13995), .A2(n11275), .ZN(n11418) );
  NOR2_X1 U11733 ( .A1(n17221), .A2(n11613), .ZN(n11612) );
  INV_X1 U11734 ( .A(n17227), .ZN(n11613) );
  OAI21_X1 U11735 ( .B1(n12051), .B2(n12028), .A(n12027), .ZN(n12029) );
  NAND2_X1 U11736 ( .A1(n17225), .A2(n11215), .ZN(n14569) );
  NOR2_X1 U11737 ( .A1(n11581), .A2(n11583), .ZN(n11580) );
  INV_X1 U11738 ( .A(n17241), .ZN(n11581) );
  AND3_X1 U11739 ( .A1(n14353), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11354), 
        .ZN(n14588) );
  AND2_X1 U11740 ( .A1(n11612), .A2(n11611), .ZN(n11610) );
  INV_X1 U11741 ( .A(n14299), .ZN(n11611) );
  AND2_X1 U11742 ( .A1(n11228), .A2(n15487), .ZN(n11621) );
  NAND2_X1 U11743 ( .A1(n11706), .A2(n13896), .ZN(n13900) );
  NAND3_X1 U11744 ( .A1(n11706), .A2(n13867), .A3(n11705), .ZN(n14088) );
  AND2_X1 U11745 ( .A1(n13866), .A2(n13896), .ZN(n11705) );
  INV_X1 U11746 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11428) );
  AND4_X1 U11747 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11898) );
  AND4_X1 U11748 ( .A1(n11887), .A2(n11886), .A3(n11885), .A4(n11884), .ZN(
        n11899) );
  AND4_X1 U11749 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11897) );
  INV_X1 U11750 ( .A(n17440), .ZN(n11711) );
  OR2_X1 U11751 ( .A1(n17122), .A2(n14324), .ZN(n14256) );
  INV_X1 U11752 ( .A(n17153), .ZN(n11618) );
  NAND2_X1 U11753 ( .A1(n17966), .A2(n11736), .ZN(n11726) );
  INV_X1 U11754 ( .A(n16229), .ZN(n11614) );
  NOR2_X1 U11755 ( .A1(n16035), .A2(n11616), .ZN(n11615) );
  INV_X1 U11756 ( .A(n15884), .ZN(n11616) );
  INV_X1 U11757 ( .A(n13998), .ZN(n11708) );
  NAND2_X1 U11758 ( .A1(n11646), .A2(n15234), .ZN(n11645) );
  INV_X1 U11759 ( .A(n16138), .ZN(n11646) );
  NOR2_X1 U11760 ( .A1(n16153), .A2(n14108), .ZN(n11576) );
  NAND3_X1 U11761 ( .A1(n13901), .A2(n14088), .A3(n14324), .ZN(n11440) );
  NAND2_X1 U11762 ( .A1(n11915), .A2(n11914), .ZN(n14137) );
  NOR2_X1 U11763 ( .A1(n14146), .A2(n14149), .ZN(n11607) );
  NOR2_X1 U11764 ( .A1(n11542), .A2(n11540), .ZN(n11539) );
  INV_X1 U11765 ( .A(n12617), .ZN(n11542) );
  NAND2_X1 U11766 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20878), .ZN(
        n12523) );
  OR2_X1 U11767 ( .A1(n20849), .A2(n12445), .ZN(n18172) );
  NOR2_X1 U11768 ( .A1(n21123), .A2(n11466), .ZN(n11465) );
  INV_X1 U11769 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11466) );
  NOR2_X1 U11770 ( .A1(n18575), .A2(n21783), .ZN(n12563) );
  AND2_X1 U11771 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12547), .ZN(
        n12548) );
  AND2_X1 U11772 ( .A1(n11558), .A2(n11242), .ZN(n12543) );
  OR2_X1 U11773 ( .A1(n18856), .A2(n11560), .ZN(n11558) );
  NAND2_X1 U11774 ( .A1(n11562), .A2(n11561), .ZN(n11560) );
  INV_X1 U11775 ( .A(n18855), .ZN(n11561) );
  NAND2_X1 U11776 ( .A1(n18858), .A2(n12723), .ZN(n12724) );
  INV_X1 U11777 ( .A(n12716), .ZN(n12714) );
  NAND2_X1 U11778 ( .A1(n11589), .A2(n12716), .ZN(n12718) );
  NAND2_X1 U11779 ( .A1(n11152), .A2(n11590), .ZN(n11589) );
  INV_X1 U11780 ( .A(n12717), .ZN(n11590) );
  INV_X1 U11781 ( .A(n11331), .ZN(n12698) );
  OAI21_X1 U11782 ( .B1(n12687), .B2(n11379), .A(n11332), .ZN(n11331) );
  INV_X1 U11783 ( .A(n21894), .ZN(n16301) );
  NAND2_X1 U11784 ( .A1(n22190), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15815) );
  AND2_X1 U11785 ( .A1(n22489), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13598) );
  AOI21_X1 U11786 ( .B1(n13515), .B2(n13514), .A(n13513), .ZN(n16485) );
  AND2_X1 U11787 ( .A1(n16817), .A2(n13469), .ZN(n13513) );
  OR2_X1 U11788 ( .A1(n13496), .A2(n13495), .ZN(n16499) );
  NOR2_X1 U11789 ( .A1(n13322), .A2(n13321), .ZN(n13323) );
  INV_X1 U11790 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U11791 ( .A1(n13323), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13357) );
  OAI21_X1 U11792 ( .B1(n22245), .B2(n13589), .A(n13290), .ZN(n16713) );
  NOR2_X1 U11793 ( .A1(n11686), .A2(n13235), .ZN(n11685) );
  NOR2_X1 U11794 ( .A1(n11281), .A2(n11687), .ZN(n11686) );
  INV_X1 U11795 ( .A(n16419), .ZN(n16439) );
  NOR2_X1 U11796 ( .A1(n16477), .A2(n16467), .ZN(n16466) );
  OAI21_X1 U11797 ( .B1(n16821), .B2(n16965), .A(n13786), .ZN(n16327) );
  NAND2_X1 U11798 ( .A1(n16488), .A2(n16478), .ZN(n16477) );
  INV_X1 U11799 ( .A(n11666), .ZN(n11665) );
  NAND2_X1 U11800 ( .A1(n13787), .A2(n11670), .ZN(n16991) );
  NAND2_X1 U11801 ( .A1(n11404), .A2(n11401), .ZN(n13787) );
  NOR2_X1 U11802 ( .A1(n13785), .A2(n11402), .ZN(n11401) );
  OR2_X1 U11803 ( .A1(n11180), .A2(n16391), .ZN(n16716) );
  OR2_X1 U11804 ( .A1(n15894), .A2(n15893), .ZN(n15898) );
  NAND2_X1 U11805 ( .A1(n16178), .A2(n11166), .ZN(n16440) );
  NAND2_X1 U11806 ( .A1(n15372), .A2(n15371), .ZN(n15395) );
  NAND2_X1 U11807 ( .A1(n13092), .A2(n15506), .ZN(n13093) );
  AND2_X1 U11808 ( .A1(n15962), .A2(n15961), .ZN(n22417) );
  NOR2_X1 U11809 ( .A1(n15962), .A2(n15732), .ZN(n15841) );
  INV_X1 U11810 ( .A(n15961), .ZN(n15732) );
  NOR2_X1 U11811 ( .A1(n22503), .A2(n22388), .ZN(n22465) );
  INV_X1 U11812 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22487) );
  NOR2_X1 U11813 ( .A1(n22459), .A2(n22388), .ZN(n22512) );
  INV_X1 U11814 ( .A(n22493), .ZN(n15913) );
  OR2_X1 U11815 ( .A1(n11207), .A2(n14270), .ZN(n14272) );
  NOR2_X1 U11816 ( .A1(n14249), .A2(n11905), .ZN(n14251) );
  NAND2_X1 U11817 ( .A1(n14027), .A2(n14028), .ZN(n14032) );
  OR2_X1 U11818 ( .A1(n14018), .A2(n11903), .ZN(n14022) );
  AND2_X1 U11819 ( .A1(n11843), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n14008) );
  NAND2_X1 U11820 ( .A1(n13904), .A2(n13905), .ZN(n13908) );
  NAND2_X1 U11821 ( .A1(n14378), .A2(n11339), .ZN(n11338) );
  NOR2_X1 U11822 ( .A1(n14380), .A2(n11340), .ZN(n11339) );
  INV_X1 U11823 ( .A(n14377), .ZN(n11340) );
  AND2_X1 U11824 ( .A1(n14379), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14380) );
  INV_X1 U11826 ( .A(n11655), .ZN(n11652) );
  NAND2_X1 U11827 ( .A1(n11200), .A2(n11602), .ZN(n11601) );
  INV_X1 U11828 ( .A(n17261), .ZN(n11602) );
  AND3_X1 U11829 ( .A1(n12349), .A2(n12348), .A3(n12347), .ZN(n16210) );
  AND2_X1 U11830 ( .A1(n14588), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n16066) );
  NAND2_X1 U11831 ( .A1(n14379), .A2(n14355), .ZN(n16068) );
  CLKBUF_X1 U11832 ( .A(n16354), .Z(n15306) );
  NAND2_X1 U11833 ( .A1(n11156), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15129) );
  NAND2_X1 U11834 ( .A1(n15128), .A2(n15127), .ZN(n18048) );
  INV_X1 U11835 ( .A(n16354), .ZN(n16353) );
  AND2_X1 U11836 ( .A1(n12151), .A2(n12150), .ZN(n17242) );
  AND2_X1 U11837 ( .A1(n12090), .A2(n12089), .ZN(n15530) );
  CLKBUF_X1 U11838 ( .A(n13902), .Z(n14067) );
  AND2_X1 U11839 ( .A1(n11433), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11432) );
  NOR2_X1 U11840 ( .A1(n14269), .A2(n11704), .ZN(n11703) );
  INV_X1 U11841 ( .A(n11715), .ZN(n11714) );
  OAI21_X1 U11842 ( .B1(n11716), .B2(n14244), .A(n17449), .ZN(n11715) );
  INV_X1 U11843 ( .A(n11728), .ZN(n11727) );
  OAI21_X1 U11844 ( .B1(n14240), .B2(n11729), .A(n11749), .ZN(n11728) );
  NAND2_X1 U11845 ( .A1(n15424), .A2(n15425), .ZN(n15492) );
  AND2_X1 U11846 ( .A1(n11287), .A2(n11643), .ZN(n16078) );
  AND2_X1 U11847 ( .A1(n19860), .A2(n18018), .ZN(n19924) );
  NAND2_X1 U11848 ( .A1(n14140), .A2(n14139), .ZN(n19932) );
  NAND2_X1 U11849 ( .A1(n17803), .A2(n17901), .ZN(n14140) );
  INV_X1 U11850 ( .A(n19932), .ZN(n20259) );
  INV_X1 U11851 ( .A(n21897), .ZN(n21921) );
  NAND2_X1 U11852 ( .A1(n21114), .A2(n11459), .ZN(n11458) );
  INV_X1 U11853 ( .A(n21180), .ZN(n11459) );
  OR2_X1 U11854 ( .A1(n21167), .A2(n11284), .ZN(n11457) );
  OR2_X1 U11855 ( .A1(n21167), .A2(n21168), .ZN(n11460) );
  NOR2_X1 U11856 ( .A1(n21114), .A2(n11455), .ZN(n21117) );
  AND2_X1 U11857 ( .A1(n21116), .A2(n21115), .ZN(n11455) );
  INV_X1 U11858 ( .A(n17836), .ZN(n20848) );
  NOR2_X1 U11859 ( .A1(n20848), .A2(n21278), .ZN(n20853) );
  INV_X2 U11860 ( .A(n18322), .ZN(n18198) );
  INV_X1 U11861 ( .A(n12477), .ZN(n11554) );
  NAND2_X1 U11862 ( .A1(n12482), .A2(n11375), .ZN(n11374) );
  NAND2_X1 U11863 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11375) );
  AOI21_X1 U11864 ( .B1(n12486), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n12488), .ZN(n12496) );
  NOR2_X1 U11865 ( .A1(n21335), .A2(n21336), .ZN(n21459) );
  AND2_X1 U11866 ( .A1(n11392), .A2(n11391), .ZN(n12592) );
  NOR2_X1 U11867 ( .A1(n21492), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11392) );
  INV_X1 U11868 ( .A(n12445), .ZN(n11391) );
  AND2_X1 U11869 ( .A1(n21892), .A2(n21893), .ZN(n21282) );
  INV_X1 U11870 ( .A(n21617), .ZN(n21511) );
  NOR2_X1 U11871 ( .A1(n18824), .A2(n20922), .ZN(n18795) );
  NAND2_X1 U11872 ( .A1(n18822), .A2(n12730), .ZN(n18811) );
  OR2_X1 U11873 ( .A1(n18808), .A2(n21589), .ZN(n11557) );
  NAND2_X1 U11874 ( .A1(n21753), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21731) );
  NOR2_X1 U11875 ( .A1(n12744), .A2(n21707), .ZN(n21753) );
  NAND2_X1 U11876 ( .A1(n12689), .A2(n11186), .ZN(n11324) );
  NOR3_X1 U11877 ( .A1(n12560), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n11192), .ZN(n11371) );
  NAND2_X1 U11878 ( .A1(n12558), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12559) );
  NOR2_X1 U11879 ( .A1(n18793), .A2(n21600), .ZN(n11376) );
  AOI21_X1 U11880 ( .B1(n12679), .B2(n12678), .A(n12677), .ZN(n21901) );
  NAND2_X1 U11881 ( .A1(n21471), .A2(n11546), .ZN(n21892) );
  NOR2_X1 U11882 ( .A1(n21808), .A2(n21929), .ZN(n21926) );
  INV_X1 U11883 ( .A(n21953), .ZN(n15798) );
  NAND2_X1 U11884 ( .A1(n13664), .A2(n13663), .ZN(n16789) );
  NOR2_X1 U11885 ( .A1(n13691), .A2(n16333), .ZN(n13692) );
  NAND2_X1 U11886 ( .A1(n20696), .A2(n13688), .ZN(n20646) );
  INV_X1 U11887 ( .A(n20646), .ZN(n20694) );
  OAI211_X1 U11888 ( .C1(n13803), .C2(n13802), .A(n13801), .B(n13800), .ZN(
        n16943) );
  INV_X1 U11889 ( .A(n22016), .ZN(n21980) );
  NAND2_X1 U11890 ( .A1(n12976), .A2(n12951), .ZN(n13073) );
  CLKBUF_X1 U11891 ( .A(n15964), .Z(n15965) );
  BUF_X1 U11892 ( .A(n15435), .Z(n15961) );
  NOR2_X2 U11893 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22497) );
  INV_X1 U11894 ( .A(n16233), .ZN(n11578) );
  NAND2_X1 U11895 ( .A1(n15159), .A2(n19341), .ZN(n20313) );
  OR2_X1 U11896 ( .A1(n15661), .A2(n15158), .ZN(n15159) );
  AND2_X1 U11897 ( .A1(n17901), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16306) );
  NOR2_X1 U11898 ( .A1(n11209), .A2(n11653), .ZN(n17089) );
  NAND2_X1 U11899 ( .A1(n11655), .A2(n11654), .ZN(n11653) );
  XNOR2_X1 U11900 ( .A(n11694), .B(n14313), .ZN(n16346) );
  AOI21_X1 U11901 ( .B1(n11701), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14310), .ZN(n11696) );
  OR2_X1 U11902 ( .A1(n14215), .A2(n14181), .ZN(n19285) );
  NOR2_X2 U11903 ( .A1(n14178), .A2(n15708), .ZN(n19271) );
  INV_X1 U11904 ( .A(n19327), .ZN(n19281) );
  OR2_X1 U11905 ( .A1(n14215), .A2(n14214), .ZN(n19327) );
  INV_X1 U11906 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20000) );
  INV_X1 U11907 ( .A(n19027), .ZN(n18018) );
  INV_X1 U11908 ( .A(n20200), .ZN(n18023) );
  NOR2_X1 U11909 ( .A1(n19952), .A2(n19910), .ZN(n20373) );
  AND2_X1 U11910 ( .A1(n19882), .A2(n19962), .ZN(n20172) );
  AND2_X1 U11911 ( .A1(n19844), .A2(n19936), .ZN(n20331) );
  NAND2_X1 U11912 ( .A1(n11475), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n11474) );
  OR2_X1 U11913 ( .A1(n21256), .A2(n21253), .ZN(n11475) );
  OR2_X1 U11914 ( .A1(n21249), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n11473) );
  XNOR2_X1 U11915 ( .A(n11477), .B(n21258), .ZN(n11476) );
  NOR2_X1 U11916 ( .A1(n21259), .A2(n21114), .ZN(n11477) );
  NOR2_X1 U11917 ( .A1(n21198), .A2(n21197), .ZN(n21205) );
  INV_X1 U11918 ( .A(n21267), .ZN(n21235) );
  INV_X1 U11919 ( .A(n21272), .ZN(n21193) );
  NAND2_X1 U11920 ( .A1(n21388), .A2(n11279), .ZN(n11328) );
  OR2_X1 U11921 ( .A1(n21390), .A2(n21389), .ZN(n21388) );
  NOR2_X1 U11922 ( .A1(n21397), .A2(n21391), .ZN(n21390) );
  NAND2_X1 U11923 ( .A1(n21398), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n21397) );
  INV_X1 U11924 ( .A(n21402), .ZN(n21419) );
  NAND2_X1 U11925 ( .A1(n21456), .A2(P3_EAX_REG_8__SCAN_IN), .ZN(n21436) );
  NOR2_X1 U11926 ( .A1(n12452), .A2(n12451), .ZN(n21751) );
  NAND2_X1 U11927 ( .A1(n21371), .A2(n21456), .ZN(n21447) );
  OAI21_X1 U11928 ( .B1(n18724), .B2(n11148), .A(n21239), .ZN(n11571) );
  NOR2_X1 U11929 ( .A1(n11570), .A2(n11569), .ZN(n11568) );
  NOR2_X1 U11930 ( .A1(n21868), .A2(n21230), .ZN(n11569) );
  INV_X1 U11931 ( .A(n18727), .ZN(n11570) );
  INV_X1 U11932 ( .A(n18756), .ZN(n18803) );
  NOR2_X2 U11933 ( .A1(n21751), .A2(n18891), .ZN(n18802) );
  INV_X1 U11934 ( .A(n18892), .ZN(n18878) );
  XNOR2_X1 U11935 ( .A(n18721), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21742) );
  NOR2_X2 U11936 ( .A1(n21751), .A2(n21559), .ZN(n21885) );
  NAND2_X1 U11937 ( .A1(n21856), .A2(n21895), .ZN(n21559) );
  AND2_X1 U11938 ( .A1(n11389), .A2(n11265), .ZN(n21947) );
  OAI22_X1 U11939 ( .A1(n11390), .A2(n21917), .B1(n21918), .B2(n21915), .ZN(
        n11389) );
  NAND2_X1 U11940 ( .A1(n21925), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11388) );
  INV_X1 U11941 ( .A(keyinput_133), .ZN(n14661) );
  XNOR2_X1 U11942 ( .A(n14657), .B(DATAI_30_), .ZN(n14658) );
  INV_X1 U11943 ( .A(keyinput_130), .ZN(n14657) );
  OAI22_X1 U11944 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_128), .B1(
        DATAI_31_), .B2(keyinput_129), .ZN(n11505) );
  INV_X1 U11945 ( .A(n14660), .ZN(n11506) );
  INV_X1 U11946 ( .A(keyinput_132), .ZN(n14662) );
  AOI21_X1 U11947 ( .B1(n11502), .B2(n11501), .A(n11498), .ZN(n14672) );
  AOI21_X1 U11948 ( .B1(n11528), .B2(n11527), .A(n11258), .ZN(n14698) );
  AOI22_X1 U11949 ( .A1(n14682), .A2(n14681), .B1(keyinput_145), .B2(DATAI_15_), .ZN(n11527) );
  NAND2_X1 U11950 ( .A1(n11530), .A2(n11529), .ZN(n11528) );
  AOI21_X1 U11951 ( .B1(n11537), .B2(n11535), .A(n11532), .ZN(n14730) );
  NAND2_X1 U11952 ( .A1(n11534), .A2(n11533), .ZN(n11532) );
  NAND2_X1 U11953 ( .A1(n11526), .A2(n11525), .ZN(n11524) );
  NAND2_X1 U11954 ( .A1(n14733), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n11525) );
  NAND2_X1 U11955 ( .A1(n21963), .A2(keyinput_171), .ZN(n11526) );
  NAND2_X1 U11956 ( .A1(n22268), .A2(keyinput_172), .ZN(n11522) );
  NOR2_X1 U11957 ( .A1(n11523), .A2(n11520), .ZN(n11519) );
  NAND2_X1 U11958 ( .A1(n11522), .A2(n11521), .ZN(n11520) );
  NOR2_X1 U11959 ( .A1(n14732), .A2(n11524), .ZN(n11523) );
  NAND2_X1 U11960 ( .A1(n14734), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11521) );
  INV_X1 U11961 ( .A(n14740), .ZN(n11515) );
  NAND2_X1 U11962 ( .A1(n11518), .A2(n11517), .ZN(n11516) );
  NAND2_X1 U11963 ( .A1(n14735), .A2(P1_MORE_REG_SCAN_IN), .ZN(n11517) );
  NAND2_X1 U11964 ( .A1(n17878), .A2(keyinput_173), .ZN(n11518) );
  INV_X1 U11965 ( .A(n14749), .ZN(n11481) );
  AOI21_X1 U11966 ( .B1(n14746), .B2(n14745), .A(n14744), .ZN(n14751) );
  AOI21_X1 U11967 ( .B1(n11201), .B2(n11482), .A(n11286), .ZN(n11479) );
  INV_X1 U11968 ( .A(n11483), .ZN(n11482) );
  NAND2_X1 U11969 ( .A1(n11489), .A2(n11292), .ZN(n11486) );
  AND2_X1 U11970 ( .A1(n14769), .A2(n11490), .ZN(n11489) );
  INV_X1 U11971 ( .A(n14774), .ZN(n11490) );
  OAI21_X1 U11972 ( .B1(n11492), .B2(n11487), .A(n11292), .ZN(n11485) );
  NOR2_X1 U11973 ( .A1(n11488), .A2(n14774), .ZN(n11487) );
  NAND2_X1 U11974 ( .A1(n11512), .A2(n14802), .ZN(n11511) );
  NAND2_X1 U11975 ( .A1(n14799), .A2(n14798), .ZN(n11512) );
  NOR2_X1 U11976 ( .A1(n14801), .A2(n11300), .ZN(n11510) );
  AOI21_X1 U11977 ( .B1(n11509), .B2(n11508), .A(n11507), .ZN(n14805) );
  XNOR2_X1 U11978 ( .A(P1_EBX_REG_24__SCAN_IN), .B(keyinput_219), .ZN(n11507)
         );
  INV_X1 U11979 ( .A(n14804), .ZN(n11508) );
  NAND2_X1 U11980 ( .A1(n11511), .A2(n11510), .ZN(n11509) );
  CLKBUF_X1 U11981 ( .A(n13566), .Z(n13543) );
  INV_X1 U11982 ( .A(n11495), .ZN(n11494) );
  OAI22_X1 U11983 ( .A1(n22234), .A2(n14814), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(keyinput_227), .ZN(n11495) );
  AND2_X1 U11984 ( .A1(n11938), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11436) );
  AOI22_X1 U11985 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11934) );
  OR2_X1 U11986 ( .A1(n12669), .A2(n12670), .ZN(n12662) );
  INV_X1 U11987 ( .A(n13050), .ZN(n11409) );
  INV_X1 U11988 ( .A(n13762), .ZN(n13751) );
  OR2_X1 U11989 ( .A1(n13037), .A2(n13036), .ZN(n13734) );
  OR2_X1 U11990 ( .A1(n13049), .A2(n13048), .ZN(n13737) );
  OR2_X1 U11991 ( .A1(n12934), .A2(n12933), .ZN(n13709) );
  OR2_X1 U11992 ( .A1(n13004), .A2(n13003), .ZN(n13707) );
  INV_X1 U11993 ( .A(n12847), .ZN(n13686) );
  AND3_X1 U11994 ( .A1(n15381), .A2(n12895), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n13642) );
  AOI22_X1 U11995 ( .A1(n13387), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U11996 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12924), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U11997 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12817), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12768) );
  OR2_X1 U11998 ( .A1(n15381), .A2(n22256), .ZN(n12992) );
  NAND2_X1 U11999 ( .A1(n15813), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12993) );
  NOR2_X1 U12000 ( .A1(n16376), .A2(n13628), .ZN(n13645) );
  AND2_X1 U12001 ( .A1(n13751), .A2(n13642), .ZN(n13651) );
  AOI22_X1 U12002 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11802) );
  NAND2_X1 U12003 ( .A1(n12063), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12058) );
  AOI21_X1 U12004 ( .B1(n12071), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n12056), .ZN(n12060) );
  OAI22_X1 U12005 ( .A1(n11363), .A2(n14195), .B1(n12049), .B2(n12085), .ZN(
        n12052) );
  NAND2_X1 U12006 ( .A1(n14238), .A2(n11450), .ZN(n11449) );
  INV_X1 U12007 ( .A(n17503), .ZN(n11450) );
  AND2_X1 U12008 ( .A1(n13958), .A2(n13957), .ZN(n13964) );
  NOR2_X1 U12009 ( .A1(n20262), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12191) );
  OR2_X1 U12010 ( .A1(n11798), .A2(n11797), .ZN(n13865) );
  NAND2_X1 U12011 ( .A1(n14149), .A2(n12006), .ZN(n11994) );
  NAND2_X1 U12012 ( .A1(n14157), .A2(n12011), .ZN(n14190) );
  AND2_X1 U12013 ( .A1(n14160), .A2(n12006), .ZN(n12011) );
  NOR2_X1 U12014 ( .A1(n11493), .A2(n14816), .ZN(n14822) );
  AOI21_X1 U12015 ( .B1(n11496), .B2(n11494), .A(n14656), .ZN(n11493) );
  NAND2_X1 U12016 ( .A1(n11982), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11344) );
  NAND2_X1 U12017 ( .A1(n11974), .A2(n11936), .ZN(n11345) );
  AND2_X1 U12018 ( .A1(n11976), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11756) );
  AOI21_X1 U12019 ( .B1(n11937), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n11923), .ZN(n11925) );
  AOI21_X1 U12020 ( .B1(n11858), .B2(n11857), .A(n11856), .ZN(n11913) );
  AOI21_X1 U12021 ( .B1(n19403), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12661), .ZN(n12670) );
  AND2_X1 U12022 ( .A1(n12671), .A2(n12675), .ZN(n12661) );
  NAND2_X1 U12023 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11541) );
  NOR2_X1 U12024 ( .A1(n21317), .A2(n12542), .ZN(n12546) );
  NOR2_X1 U12025 ( .A1(n11230), .A2(n11320), .ZN(n11319) );
  NAND2_X1 U12026 ( .A1(n12861), .A2(n12859), .ZN(n11320) );
  NOR2_X1 U12027 ( .A1(n11318), .A2(n11317), .ZN(n11316) );
  NAND2_X1 U12028 ( .A1(n12852), .A2(n12849), .ZN(n11317) );
  NOR2_X1 U12029 ( .A1(n16465), .A2(n11691), .ZN(n11690) );
  INV_X1 U12030 ( .A(n16475), .ZN(n11691) );
  NAND2_X1 U12031 ( .A1(n16895), .A2(n13782), .ZN(n16883) );
  AND2_X1 U12032 ( .A1(n16269), .A2(n13191), .ZN(n11687) );
  AND2_X1 U12033 ( .A1(n13064), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13100) );
  NOR2_X1 U12034 ( .A1(n16516), .A2(n11639), .ZN(n11638) );
  INV_X1 U12035 ( .A(n16527), .ZN(n11639) );
  OAI21_X1 U12036 ( .B1(n11405), .B2(n11668), .A(n11667), .ZN(n11666) );
  NAND2_X1 U12037 ( .A1(n11671), .A2(n13788), .ZN(n11668) );
  NAND2_X1 U12038 ( .A1(n22048), .A2(n11403), .ZN(n11402) );
  NOR2_X1 U12039 ( .A1(n11628), .A2(n16613), .ZN(n11627) );
  INV_X1 U12040 ( .A(n16623), .ZN(n11628) );
  NAND2_X1 U12041 ( .A1(n16419), .A2(n22129), .ZN(n11624) );
  NAND2_X1 U12042 ( .A1(n12885), .A2(n12891), .ZN(n13762) );
  NAND2_X1 U12043 ( .A1(n12901), .A2(n12900), .ZN(n15323) );
  OR2_X1 U12044 ( .A1(n12966), .A2(n12965), .ZN(n13708) );
  OR2_X1 U12045 ( .A1(n12946), .A2(n12945), .ZN(n13766) );
  INV_X1 U12046 ( .A(n13642), .ZN(n13624) );
  NAND2_X1 U12047 ( .A1(n12975), .A2(n12951), .ZN(n11400) );
  INV_X1 U12048 ( .A(n13092), .ZN(n13027) );
  NAND2_X1 U12049 ( .A1(n12899), .A2(n12816), .ZN(n12902) );
  INV_X1 U12050 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22476) );
  AND2_X1 U12051 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12983) );
  OR2_X1 U12052 ( .A1(n13611), .A2(n13607), .ZN(n13608) );
  INV_X1 U12053 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22408) );
  INV_X1 U12054 ( .A(n14272), .ZN(n14321) );
  INV_X1 U12055 ( .A(n14024), .ZN(n11427) );
  OR2_X1 U12056 ( .A1(n13996), .A2(n11417), .ZN(n14005) );
  NAND2_X1 U12057 ( .A1(n11418), .A2(n14002), .ZN(n11417) );
  AND3_X1 U12058 ( .A1(n13920), .A2(n11871), .A3(n11411), .ZN(n11410) );
  NOR2_X1 U12059 ( .A1(n13908), .A2(n11413), .ZN(n11412) );
  MUX2_X1 U12060 ( .A(n12050), .B(n14077), .S(n13915), .Z(n13904) );
  NAND2_X1 U12061 ( .A1(n13810), .A2(n13809), .ZN(n13808) );
  NOR2_X1 U12062 ( .A1(n11740), .A2(n11283), .ZN(n11593) );
  NOR2_X1 U12063 ( .A1(n11599), .A2(n17210), .ZN(n11598) );
  NAND2_X1 U12064 ( .A1(n11584), .A2(n11755), .ZN(n11583) );
  INV_X1 U12065 ( .A(n17248), .ZN(n11584) );
  INV_X1 U12066 ( .A(n16244), .ZN(n11603) );
  NOR2_X1 U12067 ( .A1(n11881), .A2(n11880), .ZN(n13983) );
  OR2_X1 U12068 ( .A1(n11836), .A2(n11835), .ZN(n13894) );
  INV_X1 U12069 ( .A(n14195), .ZN(n11362) );
  AND2_X1 U12070 ( .A1(n12004), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11361) );
  AND2_X1 U12071 ( .A1(n12426), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12387) );
  AND2_X1 U12072 ( .A1(n14312), .A2(n14313), .ZN(n11744) );
  AND2_X1 U12073 ( .A1(n11298), .A2(n17565), .ZN(n11433) );
  NAND2_X1 U12074 ( .A1(n11730), .A2(n11732), .ZN(n11729) );
  INV_X1 U12075 ( .A(n11736), .ZN(n11730) );
  NOR2_X1 U12076 ( .A1(n11185), .A2(n17719), .ZN(n11725) );
  INV_X1 U12077 ( .A(n14238), .ZN(n11451) );
  NAND2_X1 U12078 ( .A1(n11446), .A2(n11448), .ZN(n11443) );
  NAND2_X1 U12079 ( .A1(n11208), .A2(n11451), .ZN(n11444) );
  AOI21_X1 U12080 ( .B1(n11447), .B2(n11451), .A(n14234), .ZN(n11446) );
  AOI21_X1 U12081 ( .B1(n11358), .B2(n11360), .A(n11356), .ZN(n11355) );
  NAND2_X1 U12082 ( .A1(n11726), .A2(n11358), .ZN(n11357) );
  INV_X1 U12083 ( .A(n17685), .ZN(n11360) );
  AND2_X1 U12084 ( .A1(n12127), .A2(n12126), .ZN(n17275) );
  OR2_X1 U12085 ( .A1(n11650), .A2(n16210), .ZN(n11649) );
  AND2_X1 U12086 ( .A1(n12122), .A2(n12121), .ZN(n16215) );
  OR2_X1 U12087 ( .A1(n16214), .A2(n16215), .ZN(n17276) );
  NAND2_X1 U12088 ( .A1(n11651), .A2(n15790), .ZN(n11650) );
  INV_X1 U12089 ( .A(n17690), .ZN(n11651) );
  INV_X1 U12090 ( .A(n12334), .ZN(n12346) );
  NAND2_X1 U12091 ( .A1(n11369), .A2(n11368), .ZN(n14007) );
  NAND2_X1 U12092 ( .A1(n11453), .A2(n11194), .ZN(n11369) );
  AND2_X1 U12093 ( .A1(n11194), .A2(n17937), .ZN(n11367) );
  NAND2_X1 U12094 ( .A1(n17531), .A2(n13994), .ZN(n17938) );
  OR2_X1 U12095 ( .A1(n11855), .A2(n11854), .ZN(n14089) );
  INV_X1 U12096 ( .A(n16057), .ZN(n11644) );
  XNOR2_X1 U12097 ( .A(n14088), .B(n14089), .ZN(n14100) );
  CLKBUF_X1 U12098 ( .A(n14070), .Z(n14071) );
  NAND2_X2 U12099 ( .A1(n11772), .A2(n11353), .ZN(n14154) );
  AND2_X1 U12100 ( .A1(n19967), .A2(n19846), .ZN(n15080) );
  NAND2_X1 U12101 ( .A1(n13822), .A2(n13839), .ZN(n13842) );
  NOR2_X1 U12102 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21460), .ZN(
        n12671) );
  NOR2_X1 U12103 ( .A1(n11377), .A2(n20877), .ZN(n12473) );
  NOR2_X1 U12104 ( .A1(n12443), .A2(n12446), .ZN(n12490) );
  NOR2_X1 U12105 ( .A1(n12446), .A2(n21485), .ZN(n12524) );
  NAND2_X1 U12106 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21491), .ZN(
        n12446) );
  INV_X1 U12107 ( .A(n21020), .ZN(n11467) );
  NOR2_X1 U12108 ( .A1(n20974), .A2(n11470), .ZN(n11469) );
  INV_X1 U12109 ( .A(n21765), .ZN(n18663) );
  NAND2_X1 U12110 ( .A1(n18514), .A2(n11747), .ZN(n18575) );
  OR2_X1 U12111 ( .A1(n18511), .A2(n18539), .ZN(n18515) );
  INV_X1 U12112 ( .A(n12553), .ZN(n11566) );
  NAND2_X1 U12113 ( .A1(n18771), .A2(n12551), .ZN(n18552) );
  AND2_X1 U12114 ( .A1(n12546), .A2(n12709), .ZN(n12549) );
  INV_X1 U12115 ( .A(n21751), .ZN(n18501) );
  NAND2_X1 U12116 ( .A1(n18828), .A2(n12727), .ZN(n12729) );
  OR3_X1 U12117 ( .A1(n12740), .A2(n21503), .A3(n11546), .ZN(n21495) );
  NOR3_X1 U12118 ( .A1(n21460), .A2(n21492), .A3(n21491), .ZN(n20878) );
  NOR2_X1 U12119 ( .A1(n16472), .A2(n20576), .ZN(n16446) );
  NOR3_X1 U12120 ( .A1(n22197), .A2(n16569), .A3(n20559), .ZN(n16556) );
  INV_X1 U12121 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n22175) );
  AND2_X1 U12122 ( .A1(n16415), .A2(n16414), .ZN(n16550) );
  AND2_X1 U12123 ( .A1(n16044), .A2(n16043), .ZN(n16176) );
  CLKBUF_X1 U12124 ( .A(n16510), .Z(n16511) );
  AND2_X1 U12125 ( .A1(n15170), .A2(n15169), .ZN(n20504) );
  INV_X1 U12126 ( .A(n22373), .ZN(n15254) );
  AND2_X1 U12127 ( .A1(n15370), .A2(n15121), .ZN(n15136) );
  OR2_X1 U12128 ( .A1(n13595), .A2(n16796), .ZN(n13691) );
  AND2_X1 U12129 ( .A1(n13536), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13537) );
  NAND2_X1 U12130 ( .A1(n13537), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13595) );
  NOR2_X1 U12131 ( .A1(n13491), .A2(n16833), .ZN(n13492) );
  NAND2_X1 U12132 ( .A1(n13492), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13535) );
  AND2_X1 U12133 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n13445), .ZN(
        n13446) );
  INV_X1 U12134 ( .A(n13444), .ZN(n13445) );
  NAND2_X1 U12135 ( .A1(n13446), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13491) );
  AND2_X1 U12136 ( .A1(n13469), .A2(n16855), .ZN(n13423) );
  NOR2_X1 U12137 ( .A1(n13379), .A2(n13378), .ZN(n13380) );
  NAND2_X1 U12138 ( .A1(n13380), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13444) );
  NOR2_X1 U12139 ( .A1(n13357), .A2(n13356), .ZN(n13358) );
  INV_X1 U12140 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n13356) );
  CLKBUF_X1 U12141 ( .A(n16566), .Z(n16567) );
  NAND2_X1 U12142 ( .A1(n11681), .A2(n11680), .ZN(n11679) );
  INV_X1 U12143 ( .A(n16594), .ZN(n11680) );
  AND2_X1 U12144 ( .A1(n13325), .A2(n13324), .ZN(n16608) );
  INV_X1 U12145 ( .A(n16712), .ZN(n11678) );
  NOR2_X1 U12146 ( .A1(n13274), .A2(n13255), .ZN(n13275) );
  NAND2_X1 U12147 ( .A1(n13275), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13322) );
  NAND2_X1 U12148 ( .A1(n13254), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13274) );
  AND2_X1 U12149 ( .A1(n13236), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13254) );
  NOR2_X1 U12150 ( .A1(n13230), .A2(n13204), .ZN(n13236) );
  AND2_X1 U12151 ( .A1(n13188), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13189) );
  NOR2_X1 U12152 ( .A1(n16046), .A2(n16190), .ZN(n11676) );
  INV_X1 U12153 ( .A(n15862), .ZN(n11677) );
  AOI21_X1 U12154 ( .B1(n22178), .B2(n13469), .A(n13170), .ZN(n16223) );
  NOR2_X1 U12155 ( .A1(n13136), .A2(n20645), .ZN(n13156) );
  CLKBUF_X1 U12156 ( .A(n15862), .Z(n15863) );
  NOR2_X1 U12157 ( .A1(n13106), .A2(n20640), .ZN(n13125) );
  NAND2_X1 U12158 ( .A1(n13125), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13136) );
  NOR2_X1 U12159 ( .A1(n11748), .A2(n13058), .ZN(n13059) );
  CLKBUF_X1 U12160 ( .A(n15836), .Z(n15837) );
  NAND2_X1 U12161 ( .A1(n13107), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13106) );
  NOR2_X1 U12162 ( .A1(n13094), .A2(n13054), .ZN(n13107) );
  INV_X1 U12163 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13054) );
  NAND2_X1 U12164 ( .A1(n15511), .A2(n13091), .ZN(n15607) );
  AND2_X1 U12165 ( .A1(n16540), .A2(n11276), .ZN(n16488) );
  INV_X1 U12166 ( .A(n16489), .ZN(n11635) );
  NAND2_X1 U12167 ( .A1(n16540), .A2(n11636), .ZN(n16503) );
  NAND2_X1 U12168 ( .A1(n16540), .A2(n11638), .ZN(n16514) );
  NAND2_X1 U12169 ( .A1(n16540), .A2(n16527), .ZN(n16529) );
  NAND2_X1 U12170 ( .A1(n16714), .A2(n11197), .ZN(n16581) );
  OR2_X1 U12171 ( .A1(n16581), .A2(n16563), .ZN(n16565) );
  INV_X1 U12172 ( .A(n11673), .ZN(n11672) );
  NAND2_X1 U12173 ( .A1(n16714), .A2(n11627), .ZN(n16615) );
  NAND2_X1 U12174 ( .A1(n16714), .A2(n16623), .ZN(n16624) );
  AND2_X1 U12175 ( .A1(n16394), .A2(n16393), .ZN(n16715) );
  NAND2_X1 U12176 ( .A1(n16903), .A2(n13777), .ZN(n16896) );
  NAND2_X1 U12177 ( .A1(n11631), .A2(n11634), .ZN(n11630) );
  INV_X1 U12178 ( .A(n16668), .ZN(n11634) );
  INV_X1 U12179 ( .A(n11632), .ZN(n11631) );
  NOR3_X1 U12180 ( .A1(n16258), .A2(n11245), .A3(n16257), .ZN(n16722) );
  OR2_X1 U12181 ( .A1(n16184), .A2(n16183), .ZN(n16258) );
  NOR2_X1 U12182 ( .A1(n16258), .A2(n16257), .ZN(n20609) );
  AOI21_X1 U12183 ( .B1(n16169), .B2(n11663), .A(n11237), .ZN(n11662) );
  INV_X1 U12184 ( .A(n13761), .ZN(n11663) );
  AND2_X1 U12185 ( .A1(n22018), .A2(n22112), .ZN(n17025) );
  AND2_X1 U12186 ( .A1(n15947), .A2(n15946), .ZN(n15948) );
  NOR2_X1 U12187 ( .A1(n15949), .A2(n15948), .ZN(n16177) );
  OR2_X1 U12188 ( .A1(n15898), .A2(n15897), .ZN(n15949) );
  AND2_X1 U12189 ( .A1(n15772), .A2(n15771), .ZN(n15893) );
  NAND2_X1 U12190 ( .A1(n12982), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11674) );
  INV_X1 U12191 ( .A(n11400), .ZN(n11399) );
  NAND2_X1 U12192 ( .A1(n12981), .A2(n15842), .ZN(n15964) );
  NAND2_X1 U12193 ( .A1(n13013), .A2(n13012), .ZN(n15874) );
  INV_X1 U12194 ( .A(n15841), .ZN(n15846) );
  INV_X1 U12195 ( .A(n22380), .ZN(n22470) );
  OR3_X1 U12196 ( .A1(n22452), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n15551), 
        .ZN(n15599) );
  AND2_X1 U12197 ( .A1(n16347), .A2(n15614), .ZN(n15963) );
  NOR2_X1 U12198 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15551), .ZN(n15593) );
  NAND2_X1 U12199 ( .A1(n14184), .A2(n14183), .ZN(n15650) );
  NAND2_X1 U12200 ( .A1(n14053), .A2(n11278), .ZN(n14249) );
  INV_X1 U12201 ( .A(n14241), .ZN(n11419) );
  NAND2_X1 U12202 ( .A1(n14053), .A2(n14064), .ZN(n14228) );
  NAND2_X1 U12203 ( .A1(n14053), .A2(n11420), .ZN(n14242) );
  AND2_X1 U12204 ( .A1(n12356), .A2(n12355), .ZN(n17363) );
  INV_X1 U12205 ( .A(n12414), .ZN(n12395) );
  NOR2_X1 U12206 ( .A1(n14022), .A2(n11904), .ZN(n14027) );
  NAND2_X1 U12207 ( .A1(n11902), .A2(n11901), .ZN(n14018) );
  INV_X1 U12208 ( .A(n14008), .ZN(n11901) );
  INV_X1 U12209 ( .A(n11418), .ZN(n11416) );
  AND2_X1 U12210 ( .A1(n12170), .A2(n12169), .ZN(n14299) );
  NAND2_X1 U12211 ( .A1(n17123), .A2(n11612), .ZN(n17219) );
  NAND2_X1 U12212 ( .A1(n12005), .A2(n12004), .ZN(n11365) );
  NAND2_X1 U12213 ( .A1(n11592), .A2(n11596), .ZN(n17197) );
  NOR2_X1 U12214 ( .A1(n11598), .A2(n11597), .ZN(n11596) );
  NAND2_X1 U12215 ( .A1(n11594), .A2(n11593), .ZN(n11592) );
  INV_X1 U12216 ( .A(n17204), .ZN(n11597) );
  AND2_X1 U12217 ( .A1(n14286), .A2(n14287), .ZN(n17286) );
  NAND2_X1 U12218 ( .A1(n11600), .A2(n11599), .ZN(n17209) );
  XNOR2_X1 U12219 ( .A(n14569), .B(n11296), .ZN(n17216) );
  AND2_X1 U12220 ( .A1(n12366), .A2(n12365), .ZN(n17127) );
  NAND2_X1 U12221 ( .A1(n11580), .A2(n11349), .ZN(n11348) );
  INV_X1 U12222 ( .A(n17237), .ZN(n11349) );
  NAND2_X1 U12223 ( .A1(n17231), .A2(n17233), .ZN(n17232) );
  OR2_X1 U12224 ( .A1(n17341), .A2(n17340), .ZN(n17343) );
  NAND2_X1 U12225 ( .A1(n17156), .A2(n17157), .ZN(n17341) );
  OR2_X1 U12226 ( .A1(n17689), .A2(n11647), .ZN(n15099) );
  NAND2_X1 U12227 ( .A1(n11648), .A2(n19116), .ZN(n11647) );
  INV_X1 U12228 ( .A(n11649), .ZN(n11648) );
  AND2_X1 U12229 ( .A1(n12354), .A2(n12353), .ZN(n15100) );
  AND2_X1 U12230 ( .A1(n12246), .A2(n12245), .ZN(n16138) );
  NOR2_X1 U12231 ( .A1(n20313), .A2(n15163), .ZN(n16355) );
  NAND2_X1 U12232 ( .A1(n12321), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12200) );
  AND2_X1 U12233 ( .A1(n11610), .A2(n14284), .ZN(n11609) );
  INV_X1 U12234 ( .A(n12424), .ZN(n12390) );
  AND2_X1 U12235 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n12390), .ZN(
        n12426) );
  NAND2_X1 U12236 ( .A1(n12425), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12424) );
  NOR2_X1 U12237 ( .A1(n11206), .A2(n19183), .ZN(n12425) );
  NAND2_X1 U12238 ( .A1(n12419), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12421) );
  INV_X1 U12239 ( .A(n17242), .ZN(n11617) );
  NOR2_X1 U12240 ( .A1(n12417), .A2(n12418), .ZN(n12419) );
  NAND2_X1 U12241 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n12416), .ZN(
        n12415) );
  NAND2_X1 U12242 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12386), .ZN(
        n12417) );
  INV_X1 U12243 ( .A(n12415), .ZN(n12386) );
  NAND2_X1 U12244 ( .A1(n12414), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12413) );
  NOR2_X1 U12245 ( .A1(n12413), .A2(n17489), .ZN(n12416) );
  INV_X1 U12246 ( .A(n12396), .ZN(n12411) );
  NOR2_X1 U12247 ( .A1(n12408), .A2(n17523), .ZN(n12396) );
  NAND2_X1 U12248 ( .A1(n12409), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12408) );
  NOR2_X1 U12249 ( .A1(n12406), .A2(n17988), .ZN(n12409) );
  AND2_X1 U12250 ( .A1(n12109), .A2(n12108), .ZN(n16035) );
  NAND2_X1 U12251 ( .A1(n15883), .A2(n15884), .ZN(n16036) );
  NOR2_X1 U12252 ( .A1(n12100), .A2(n12404), .ZN(n12407) );
  NAND2_X1 U12253 ( .A1(n12405), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12404) );
  AND2_X1 U12254 ( .A1(n12099), .A2(n12098), .ZN(n15954) );
  NOR2_X1 U12255 ( .A1(n12402), .A2(n17958), .ZN(n12405) );
  NAND2_X1 U12256 ( .A1(n12403), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12402) );
  INV_X1 U12257 ( .A(n15530), .ZN(n11620) );
  NAND2_X1 U12258 ( .A1(n16094), .A2(n11621), .ZN(n15529) );
  NOR2_X1 U12259 ( .A1(n12400), .A2(n16143), .ZN(n12403) );
  NAND2_X1 U12260 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n12401), .ZN(
        n12400) );
  NAND2_X1 U12261 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12399), .ZN(
        n12398) );
  NAND2_X1 U12262 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12397) );
  NOR2_X1 U12263 ( .A1(n12397), .A2(n17923), .ZN(n12399) );
  NOR2_X1 U12264 ( .A1(n11656), .A2(n11657), .ZN(n11655) );
  INV_X1 U12265 ( .A(n17285), .ZN(n11656) );
  NOR2_X1 U12266 ( .A1(n14301), .A2(n17087), .ZN(n11654) );
  NAND2_X1 U12267 ( .A1(n14310), .A2(n11702), .ZN(n11701) );
  NOR2_X1 U12268 ( .A1(n11699), .A2(n14311), .ZN(n11695) );
  NOR2_X1 U12269 ( .A1(n11703), .A2(n11700), .ZN(n11699) );
  AOI21_X1 U12270 ( .B1(n11177), .B2(n11716), .A(n11255), .ZN(n11710) );
  OR3_X1 U12271 ( .A1(n14264), .A2(n14324), .A3(n17567), .ZN(n17434) );
  AND2_X1 U12272 ( .A1(n12147), .A2(n12146), .ZN(n17153) );
  NAND2_X1 U12273 ( .A1(n17255), .A2(n11248), .ZN(n17243) );
  NAND2_X1 U12274 ( .A1(n17255), .A2(n11247), .ZN(n17154) );
  OAI211_X1 U12275 ( .C1(n17505), .C2(n11445), .A(n11442), .B(n11370), .ZN(
        n14069) );
  INV_X1 U12276 ( .A(n11446), .ZN(n11445) );
  AND2_X1 U12277 ( .A1(n11444), .A2(n11443), .ZN(n11442) );
  NAND2_X1 U12278 ( .A1(n17505), .A2(n11208), .ZN(n11370) );
  AND2_X1 U12279 ( .A1(n17255), .A2(n17256), .ZN(n17258) );
  INV_X1 U12280 ( .A(n17485), .ZN(n14062) );
  AND2_X1 U12281 ( .A1(n17508), .A2(n17504), .ZN(n17499) );
  NAND2_X1 U12282 ( .A1(n17521), .A2(n11204), .ZN(n17494) );
  OR2_X1 U12283 ( .A1(n17276), .A2(n17275), .ZN(n17278) );
  AND2_X1 U12284 ( .A1(n12131), .A2(n12130), .ZN(n15098) );
  NAND2_X1 U12285 ( .A1(n17505), .A2(n17503), .ZN(n17508) );
  NAND2_X1 U12286 ( .A1(n17684), .A2(n17685), .ZN(n17517) );
  OR2_X1 U12287 ( .A1(n17689), .A2(n11650), .ZN(n16209) );
  NOR2_X1 U12288 ( .A1(n17689), .A2(n17690), .ZN(n17688) );
  AND2_X1 U12289 ( .A1(n12113), .A2(n12112), .ZN(n16229) );
  AND2_X1 U12290 ( .A1(n15883), .A2(n11252), .ZN(n16238) );
  NAND2_X1 U12291 ( .A1(n15883), .A2(n11615), .ZN(n16230) );
  NAND2_X1 U12292 ( .A1(n11707), .A2(n17752), .ZN(n17731) );
  OAI21_X1 U12293 ( .B1(n17531), .B2(n11454), .A(n11452), .ZN(n11707) );
  INV_X1 U12294 ( .A(n11453), .ZN(n11452) );
  OR2_X1 U12295 ( .A1(n16139), .A2(n11645), .ZN(n16101) );
  NAND2_X1 U12296 ( .A1(n17934), .A2(n14113), .ZN(n17749) );
  NAND2_X1 U12297 ( .A1(n17749), .A2(n17750), .ZN(n17748) );
  NAND2_X1 U12298 ( .A1(n17938), .A2(n17937), .ZN(n17940) );
  NAND2_X1 U12299 ( .A1(n17935), .A2(n17936), .ZN(n17934) );
  NAND2_X1 U12300 ( .A1(n16094), .A2(n16122), .ZN(n16121) );
  AND2_X1 U12301 ( .A1(n16094), .A2(n11228), .ZN(n15496) );
  NAND2_X1 U12302 ( .A1(n11239), .A2(n14107), .ZN(n11577) );
  AOI21_X1 U12303 ( .B1(n11430), .B2(n14106), .A(n11576), .ZN(n11429) );
  INV_X1 U12304 ( .A(n14100), .ZN(n11431) );
  NAND2_X1 U12305 ( .A1(n11574), .A2(n19317), .ZN(n14102) );
  AOI211_X1 U12306 ( .C1(n17759), .C2(n14208), .A(n14207), .B(n19237), .ZN(
        n17760) );
  OR2_X1 U12307 ( .A1(n16056), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11439) );
  AND2_X1 U12308 ( .A1(n16056), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11438) );
  OR2_X1 U12309 ( .A1(n14215), .A2(n15650), .ZN(n17759) );
  NOR2_X1 U12310 ( .A1(n14137), .A2(n15129), .ZN(n14138) );
  XNOR2_X1 U12311 ( .A(n14374), .B(n14372), .ZN(n15061) );
  NOR2_X1 U12312 ( .A1(n11171), .A2(n13840), .ZN(n13831) );
  OR2_X1 U12313 ( .A1(n19860), .A2(n19027), .ZN(n19899) );
  AND2_X1 U12314 ( .A1(n15439), .A2(n13838), .ZN(n13853) );
  OR2_X2 U12315 ( .A1(n13842), .A2(n17905), .ZN(n13924) );
  NAND2_X1 U12316 ( .A1(n11965), .A2(n11936), .ZN(n11346) );
  NAND2_X1 U12317 ( .A1(n11959), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11347) );
  INV_X1 U12318 ( .A(n14149), .ZN(n20112) );
  AND2_X1 U12319 ( .A1(n19982), .A2(n18023), .ZN(n19844) );
  AND2_X1 U12320 ( .A1(n19860), .A2(n19027), .ZN(n19962) );
  NOR2_X1 U12321 ( .A1(n21237), .A2(n21114), .ZN(n21238) );
  NOR2_X1 U12322 ( .A1(n21222), .A2(n21221), .ZN(n21237) );
  NOR2_X1 U12323 ( .A1(n21157), .A2(n21156), .ZN(n21166) );
  NOR2_X1 U12324 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n21048), .ZN(n21070) );
  NOR2_X1 U12325 ( .A1(n18766), .A2(n20974), .ZN(n20985) );
  NOR2_X1 U12326 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20971), .ZN(n20991) );
  NOR2_X1 U12327 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20943), .ZN(n20970) );
  NAND2_X1 U12328 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18407), .ZN(n18401) );
  NOR2_X1 U12329 ( .A1(n18166), .A2(n18150), .ZN(n18169) );
  NAND2_X1 U12330 ( .A1(n12611), .A2(n11223), .ZN(n21336) );
  INV_X1 U12331 ( .A(n12615), .ZN(n11538) );
  NOR2_X1 U12332 ( .A1(n20849), .A2(n12446), .ZN(n12609) );
  NOR2_X1 U12333 ( .A1(n20789), .A2(n17833), .ZN(n18940) );
  NOR2_X1 U12334 ( .A1(n21927), .A2(n20789), .ZN(n20790) );
  NAND2_X1 U12335 ( .A1(n18726), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n18694) );
  NOR2_X1 U12336 ( .A1(n18694), .A2(n20857), .ZN(n18717) );
  NAND2_X1 U12337 ( .A1(n18717), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18708) );
  NOR3_X1 U12338 ( .A1(n18653), .A2(n11471), .A3(n21203), .ZN(n18726) );
  NAND2_X1 U12339 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11471) );
  NOR3_X1 U12340 ( .A1(n18653), .A2(n21203), .A3(n21209), .ZN(n18651) );
  INV_X1 U12341 ( .A(n18656), .ZN(n18671) );
  NOR2_X1 U12342 ( .A1(n18653), .A2(n21203), .ZN(n18656) );
  NOR2_X1 U12343 ( .A1(n21771), .A2(n21690), .ZN(n18624) );
  AND2_X1 U12344 ( .A1(n18519), .A2(n11195), .ZN(n18642) );
  NAND2_X1 U12345 ( .A1(n18519), .A2(n11193), .ZN(n18615) );
  NAND2_X1 U12346 ( .A1(n21658), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18518) );
  INV_X1 U12347 ( .A(n18521), .ZN(n18519) );
  NAND2_X1 U12348 ( .A1(n18795), .A2(n18502), .ZN(n18766) );
  OR2_X1 U12349 ( .A1(n18891), .A2(n18501), .ZN(n18756) );
  AOI22_X1 U12350 ( .A1(n21903), .A2(n21895), .B1(n21901), .B2(n21898), .ZN(
        n21924) );
  AOI21_X2 U12351 ( .B1(n20786), .B2(n20846), .A(n18871), .ZN(n18840) );
  NOR2_X1 U12352 ( .A1(n18663), .A2(n18662), .ZN(n18670) );
  NOR2_X1 U12353 ( .A1(n18793), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18598) );
  NAND2_X1 U12354 ( .A1(n18515), .A2(n18596), .ZN(n18514) );
  NAND2_X1 U12355 ( .A1(n21657), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21817) );
  NOR2_X1 U12356 ( .A1(n12560), .A2(n12557), .ZN(n18539) );
  INV_X1 U12357 ( .A(n12558), .ZN(n12557) );
  NOR2_X1 U12358 ( .A1(n18552), .A2(n12553), .ZN(n18741) );
  AOI21_X1 U12359 ( .B1(n11178), .B2(n21589), .A(n11188), .ZN(n11555) );
  INV_X1 U12360 ( .A(n11545), .ZN(n11543) );
  NAND2_X1 U12361 ( .A1(n12735), .A2(n18791), .ZN(n21617) );
  INV_X1 U12362 ( .A(n12733), .ZN(n12731) );
  XNOR2_X1 U12363 ( .A(n12729), .B(n11586), .ZN(n18823) );
  INV_X1 U12364 ( .A(n12728), .ZN(n11586) );
  NOR2_X1 U12365 ( .A1(n12545), .A2(n18831), .ZN(n18820) );
  NAND2_X1 U12366 ( .A1(n18846), .A2(n12726), .ZN(n18829) );
  NAND2_X1 U12367 ( .A1(n18829), .A2(n18830), .ZN(n18828) );
  XNOR2_X1 U12368 ( .A(n12724), .B(n11585), .ZN(n18848) );
  NOR2_X1 U12369 ( .A1(n18856), .A2(n18855), .ZN(n18854) );
  NAND2_X1 U12370 ( .A1(n12721), .A2(n12722), .ZN(n18859) );
  NAND2_X1 U12371 ( .A1(n18859), .A2(n18860), .ZN(n18858) );
  XNOR2_X1 U12372 ( .A(n12718), .B(n12536), .ZN(n18868) );
  NAND2_X1 U12373 ( .A1(n11395), .A2(n11394), .ZN(n21528) );
  INV_X1 U12374 ( .A(n21503), .ZN(n11394) );
  OR2_X1 U12375 ( .A1(n12740), .A2(n11396), .ZN(n11395) );
  INV_X1 U12376 ( .A(n12746), .ZN(n11396) );
  NOR2_X1 U12377 ( .A1(n11382), .A2(n21279), .ZN(n12707) );
  NOR2_X1 U12378 ( .A1(n21865), .A2(n11393), .ZN(n21479) );
  AND2_X1 U12379 ( .A1(n21528), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11393) );
  INV_X1 U12380 ( .A(n12740), .ZN(n21499) );
  NOR2_X1 U12381 ( .A1(n12657), .A2(n12656), .ZN(n19592) );
  NOR2_X1 U12382 ( .A1(n12627), .A2(n12626), .ZN(n19550) );
  NOR2_X1 U12383 ( .A1(n12608), .A2(n12607), .ZN(n21335) );
  NOR3_X1 U12384 ( .A1(n16304), .A2(n16303), .A3(n16302), .ZN(n21925) );
  AND2_X1 U12385 ( .A1(n21918), .A2(n21916), .ZN(n11390) );
  INV_X1 U12386 ( .A(n21950), .ZN(n11387) );
  OAI21_X1 U12387 ( .B1(n15056), .B2(n15055), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n16354) );
  INV_X1 U12388 ( .A(n22265), .ZN(n20704) );
  OR2_X1 U12389 ( .A1(n15136), .A2(n22782), .ZN(n21953) );
  NAND2_X1 U12390 ( .A1(n16509), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n16492) );
  NOR2_X1 U12391 ( .A1(n16496), .A2(n20568), .ZN(n16509) );
  AND2_X1 U12392 ( .A1(n16542), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16535) );
  NAND2_X1 U12393 ( .A1(n16556), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n16543) );
  AND2_X1 U12394 ( .A1(n22197), .A2(n22190), .ZN(n22228) );
  NOR2_X1 U12395 ( .A1(n16543), .A2(n20563), .ZN(n16542) );
  INV_X1 U12396 ( .A(n22242), .ZN(n22204) );
  AND2_X1 U12397 ( .A1(n22190), .A2(n15806), .ZN(n22216) );
  NAND2_X1 U12398 ( .A1(n15812), .A2(n15804), .ZN(n22235) );
  NAND2_X1 U12399 ( .A1(n15812), .A2(n15811), .ZN(n22197) );
  INV_X1 U12400 ( .A(n22228), .ZN(n22161) );
  AND2_X1 U12401 ( .A1(n22238), .A2(n15800), .ZN(n22124) );
  AND2_X1 U12402 ( .A1(n16789), .A2(n16727), .ZN(n16778) );
  INV_X1 U12403 ( .A(n16725), .ZN(n16776) );
  NAND2_X1 U12404 ( .A1(n16789), .A2(n15183), .ZN(n16791) );
  INV_X1 U12405 ( .A(n15261), .ZN(n22377) );
  OR2_X1 U12406 ( .A1(n15122), .A2(n17862), .ZN(n22379) );
  NAND2_X1 U12407 ( .A1(n15261), .A2(n12891), .ZN(n22373) );
  OAI21_X1 U12408 ( .B1(n16474), .B2(n16475), .A(n16462), .ZN(n16810) );
  NAND2_X1 U12409 ( .A1(n16821), .A2(n13793), .ZN(n16812) );
  OR2_X1 U12410 ( .A1(n16485), .A2(n16484), .ZN(n16486) );
  XNOR2_X1 U12411 ( .A(n16443), .B(n16442), .ZN(n16940) );
  NAND2_X1 U12412 ( .A1(n16438), .A2(n16437), .ZN(n16443) );
  NAND2_X1 U12413 ( .A1(n16326), .A2(n16327), .ZN(n16793) );
  OR2_X1 U12414 ( .A1(n16830), .A2(n16829), .ZN(n16831) );
  NAND2_X1 U12415 ( .A1(n11664), .A2(n13761), .ZN(n16170) );
  NAND2_X1 U12416 ( .A1(n16201), .A2(n16202), .ZN(n11664) );
  AND2_X1 U12417 ( .A1(n15396), .A2(n22121), .ZN(n22016) );
  AND2_X1 U12418 ( .A1(n15395), .A2(n15383), .ZN(n22106) );
  AND2_X1 U12419 ( .A1(n15395), .A2(n15380), .ZN(n22118) );
  INV_X1 U12420 ( .A(n22497), .ZN(n22506) );
  INV_X1 U12421 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17889) );
  AND2_X1 U12422 ( .A1(n22417), .A2(n22396), .ZN(n22714) );
  AND2_X1 U12423 ( .A1(n22417), .A2(n15963), .ZN(n22720) );
  INV_X1 U12424 ( .A(n22428), .ZN(n22722) );
  NOR2_X2 U12425 ( .A1(n15621), .A2(n15733), .ZN(n22728) );
  OAI211_X1 U12426 ( .C1(n22733), .C2(n22452), .A(n22451), .B(n22465), .ZN(
        n22736) );
  NOR2_X1 U12427 ( .A1(n15846), .A2(n15733), .ZN(n22746) );
  OAI211_X1 U12428 ( .C1(n22514), .C2(n22769), .A(n22513), .B(n22512), .ZN(
        n22773) );
  NOR2_X1 U12429 ( .A1(n22493), .A2(n22486), .ZN(n22772) );
  NAND2_X1 U12430 ( .A1(n15913), .A2(n15963), .ZN(n22700) );
  NOR2_X1 U12431 ( .A1(n16371), .A2(n22452), .ZN(n22259) );
  INV_X2 U12432 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n22489) );
  INV_X1 U12433 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n22250) );
  INV_X1 U12434 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n22452) );
  INV_X1 U12435 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n22256) );
  INV_X1 U12436 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n22299) );
  NAND2_X1 U12437 ( .A1(n14272), .A2(n14271), .ZN(n17104) );
  OR2_X1 U12438 ( .A1(n14261), .A2(n14260), .ZN(n14258) );
  CLKBUF_X1 U12439 ( .A(n19124), .Z(n19208) );
  INV_X1 U12440 ( .A(n19147), .ZN(n19218) );
  INV_X1 U12441 ( .A(n19163), .ZN(n19210) );
  INV_X1 U12442 ( .A(n19199), .ZN(n19207) );
  AND2_X1 U12443 ( .A1(n15107), .A2(n12381), .ZN(n19140) );
  AND2_X1 U12444 ( .A1(n15107), .A2(n11993), .ZN(n19217) );
  INV_X1 U12445 ( .A(n19217), .ZN(n19165) );
  OR2_X1 U12446 ( .A1(n12345), .A2(n12344), .ZN(n16245) );
  NOR2_X1 U12447 ( .A1(n12317), .A2(n12316), .ZN(n16233) );
  OR2_X1 U12448 ( .A1(n12293), .A2(n12292), .ZN(n15882) );
  NOR2_X1 U12449 ( .A1(n12281), .A2(n12280), .ZN(n15957) );
  AND2_X1 U12450 ( .A1(n15536), .A2(n14381), .ZN(n11350) );
  INV_X1 U12451 ( .A(n17272), .ZN(n17274) );
  XNOR2_X1 U12452 ( .A(n11351), .B(n11595), .ZN(n17306) );
  OAI21_X1 U12453 ( .B1(n11600), .B2(n11599), .A(n17209), .ZN(n11351) );
  AND2_X1 U12454 ( .A1(n16355), .A2(n16354), .ZN(n20316) );
  AND2_X1 U12455 ( .A1(n16355), .A2(n16353), .ZN(n20317) );
  NAND2_X1 U12456 ( .A1(n14378), .A2(n14377), .ZN(n16070) );
  NAND2_X1 U12457 ( .A1(n11643), .A2(n12229), .ZN(n16058) );
  NAND2_X1 U12458 ( .A1(n20153), .A2(n19835), .ZN(n20154) );
  INV_X1 U12459 ( .A(n20154), .ZN(n20319) );
  BUF_X1 U12460 ( .A(n15296), .Z(n15303) );
  XNOR2_X1 U12461 ( .A(n11311), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17403) );
  NOR2_X1 U12462 ( .A1(n12388), .A2(n16319), .ZN(n11311) );
  XNOR2_X1 U12463 ( .A(n17488), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14179) );
  NAND2_X1 U12464 ( .A1(n17521), .A2(n11202), .ZN(n18011) );
  INV_X1 U12465 ( .A(n18002), .ZN(n18001) );
  INV_X1 U12466 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17932) );
  INV_X1 U12467 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17923) );
  NAND2_X1 U12468 ( .A1(n19353), .A2(n14141), .ZN(n17987) );
  INV_X1 U12469 ( .A(n18008), .ZN(n17983) );
  INV_X1 U12470 ( .A(n17987), .ZN(n18003) );
  XNOR2_X1 U12471 ( .A(n11415), .B(n11750), .ZN(n16325) );
  NAND2_X1 U12472 ( .A1(n17396), .A2(n17408), .ZN(n11415) );
  NAND2_X1 U12473 ( .A1(n11698), .A2(n11697), .ZN(n14298) );
  NAND2_X1 U12474 ( .A1(n17464), .A2(n11713), .ZN(n11712) );
  NAND2_X1 U12475 ( .A1(n17462), .A2(n14247), .ZN(n17451) );
  NOR2_X1 U12476 ( .A1(n14069), .A2(n14068), .ZN(n17470) );
  NOR2_X1 U12477 ( .A1(n14209), .A2(n19338), .ZN(n19253) );
  AND2_X1 U12478 ( .A1(n14102), .A2(n11573), .ZN(n19323) );
  NAND2_X1 U12479 ( .A1(n16088), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11573) );
  INV_X1 U12480 ( .A(n11574), .ZN(n16088) );
  INV_X1 U12481 ( .A(n19271), .ZN(n19332) );
  CLKBUF_X1 U12482 ( .A(n15439), .Z(n19330) );
  AND2_X1 U12483 ( .A1(n17759), .A2(n17756), .ZN(n19237) );
  INV_X1 U12484 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12216) );
  INV_X1 U12485 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19884) );
  INV_X1 U12486 ( .A(n19882), .ZN(n19900) );
  INV_X1 U12487 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17845) );
  OAI21_X1 U12488 ( .B1(n19023), .B2(n15712), .A(n14358), .ZN(n17771) );
  AND2_X1 U12489 ( .A1(n15641), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17803) );
  NOR2_X1 U12490 ( .A1(n19843), .A2(n20006), .ZN(n20414) );
  NOR2_X2 U12491 ( .A1(n20006), .A2(n16022), .ZN(n20415) );
  OAI21_X1 U12492 ( .B1(n19976), .B2(n19975), .A(n19974), .ZN(n20398) );
  INV_X1 U12493 ( .A(n20396), .ZN(n20293) );
  INV_X1 U12494 ( .A(n20382), .ZN(n20287) );
  OAI21_X1 U12495 ( .B1(n20364), .B2(n19915), .A(n19932), .ZN(n20367) );
  OAI21_X1 U12496 ( .B1(n19921), .B2(n19929), .A(n19920), .ZN(n20366) );
  NOR2_X1 U12497 ( .A1(n19900), .A2(n19899), .ZN(n20365) );
  INV_X1 U12498 ( .A(n20175), .ZN(n20353) );
  AND2_X1 U12499 ( .A1(n19882), .A2(n19936), .ZN(n20358) );
  AOI21_X1 U12500 ( .B1(n20330), .B2(n19932), .A(n19850), .ZN(n20333) );
  AND2_X1 U12501 ( .A1(n19844), .A2(n19924), .ZN(n20210) );
  AND2_X1 U12502 ( .A1(n19932), .A2(n20314), .ZN(n20434) );
  INV_X1 U12503 ( .A(n20403), .ZN(n20428) );
  INV_X1 U12504 ( .A(n20306), .ZN(n20309) );
  INV_X1 U12505 ( .A(n20198), .ZN(n20188) );
  AND2_X1 U12506 ( .A1(n16031), .A2(n16030), .ZN(n20194) );
  INV_X1 U12507 ( .A(n20146), .ZN(n20149) );
  INV_X1 U12508 ( .A(n20102), .ZN(n20105) );
  INV_X1 U12509 ( .A(n20056), .ZN(n20059) );
  AND2_X1 U12510 ( .A1(n19844), .A2(n19962), .ZN(n20430) );
  INV_X1 U12511 ( .A(n20015), .ZN(n20018) );
  AND2_X1 U12512 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n11917), .ZN(n19341) );
  AOI21_X1 U12513 ( .B1(n15712), .B2(n15711), .A(n15710), .ZN(n19345) );
  OAI21_X1 U12514 ( .B1(n22320), .B2(n22305), .A(n18099), .ZN(n22312) );
  INV_X1 U12515 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n22320) );
  OR2_X1 U12516 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n22307), .ZN(n18104) );
  INV_X2 U12517 ( .A(n18104), .ZN(n22306) );
  NAND2_X1 U12518 ( .A1(n21926), .A2(n21921), .ZN(n20789) );
  AND2_X1 U12519 ( .A1(n11457), .A2(n11268), .ZN(n21197) );
  NAND2_X1 U12520 ( .A1(n11457), .A2(n11458), .ZN(n21196) );
  NAND2_X1 U12521 ( .A1(n21126), .A2(n21125), .ZN(n11462) );
  NOR2_X1 U12522 ( .A1(n21126), .A2(n21114), .ZN(n21127) );
  NOR2_X1 U12523 ( .A1(n21127), .A2(n21128), .ZN(n21142) );
  NOR2_X1 U12524 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n21109), .ZN(n21130) );
  INV_X1 U12525 ( .A(n21152), .ZN(n21087) );
  INV_X1 U12526 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20857) );
  NAND4_X1 U12527 ( .A1(n21868), .A2(n20848), .A3(n21179), .A4(n21945), .ZN(
        n21272) );
  OAI211_X1 U12528 ( .C1(n20854), .C2(n21279), .A(n21928), .B(n20853), .ZN(
        n21268) );
  NAND4_X1 U12529 ( .A1(n20853), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n20850), 
        .A4(n20845), .ZN(n21267) );
  NOR2_X1 U12530 ( .A1(n21186), .A2(n18392), .ZN(n18397) );
  NOR2_X1 U12531 ( .A1(n21072), .A2(n18463), .ZN(n18485) );
  NAND2_X1 U12532 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18165), .ZN(n18463) );
  INV_X1 U12533 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18409) );
  AOI211_X1 U12534 ( .C1(n18319), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n12634), .B(n12633), .ZN(n12635) );
  NOR2_X1 U12535 ( .A1(n21376), .A2(n11329), .ZN(n21398) );
  NAND2_X1 U12536 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(P3_EAX_REG_27__SCAN_IN), 
        .ZN(n11329) );
  NOR2_X1 U12537 ( .A1(n21376), .A2(n21377), .ZN(n21404) );
  INV_X1 U12538 ( .A(n21408), .ZN(n21372) );
  NAND2_X1 U12539 ( .A1(n21372), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n21376) );
  NOR3_X1 U12540 ( .A1(n21420), .A2(n21370), .A3(n21369), .ZN(n21414) );
  INV_X1 U12541 ( .A(n21447), .ZN(n21389) );
  NAND2_X1 U12542 ( .A1(n21429), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n21420) );
  AND2_X1 U12543 ( .A1(n21335), .A2(n21389), .ZN(n21418) );
  OR2_X1 U12544 ( .A1(n21436), .A2(n11330), .ZN(n21431) );
  NOR2_X1 U12545 ( .A1(n21437), .A2(n21458), .ZN(n21435) );
  NOR2_X1 U12546 ( .A1(n12472), .A2(n12471), .ZN(n21326) );
  NOR3_X1 U12547 ( .A1(n11551), .A2(n12481), .A3(n11374), .ZN(n11373) );
  NOR2_X1 U12548 ( .A1(n11554), .A2(n11553), .ZN(n11552) );
  INV_X1 U12549 ( .A(n12483), .ZN(n11551) );
  OAI21_X1 U12550 ( .B1(n21282), .B2(n21281), .A(n21280), .ZN(n21456) );
  INV_X1 U12551 ( .A(n21450), .ZN(n21453) );
  INV_X1 U12552 ( .A(n21443), .ZN(n21454) );
  NOR2_X1 U12553 ( .A1(n18957), .A2(n18940), .ZN(n18949) );
  CLKBUF_X1 U12555 ( .A(n20826), .Z(n20842) );
  AND2_X1 U12557 ( .A1(n18731), .A2(n11549), .ZN(n18659) );
  NOR2_X1 U12558 ( .A1(n18640), .A2(n21783), .ZN(n11549) );
  NAND2_X1 U12559 ( .A1(n21519), .A2(n21709), .ZN(n21771) );
  NOR2_X1 U12560 ( .A1(n21817), .A2(n18640), .ZN(n21519) );
  INV_X1 U12561 ( .A(n18731), .ZN(n18639) );
  NAND2_X1 U12562 ( .A1(n18519), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18600) );
  NAND2_X1 U12563 ( .A1(n18503), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18521) );
  NOR2_X1 U12564 ( .A1(n18526), .A2(n18541), .ZN(n18728) );
  AND2_X1 U12565 ( .A1(n18535), .A2(n11550), .ZN(n18731) );
  INV_X1 U12566 ( .A(n21829), .ZN(n11550) );
  OAI22_X1 U12567 ( .A1(n21511), .A2(n18892), .B1(n21616), .B2(n18756), .ZN(
        n18535) );
  INV_X1 U12568 ( .A(n18535), .ZN(n18790) );
  INV_X1 U12569 ( .A(n11557), .ZN(n18807) );
  NAND2_X1 U12570 ( .A1(n11456), .A2(n11261), .ZN(n18824) );
  INV_X1 U12571 ( .A(n18851), .ZN(n11456) );
  INV_X1 U12572 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20922) );
  AND3_X1 U12573 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18835) );
  INV_X1 U12574 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20890) );
  NAND2_X1 U12575 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18851) );
  NAND2_X1 U12576 ( .A1(n19716), .A2(n18897), .ZN(n19549) );
  INV_X1 U12577 ( .A(n18885), .ZN(n18873) );
  NAND2_X1 U12578 ( .A1(n18871), .A2(n20850), .ZN(n18891) );
  NAND2_X1 U12579 ( .A1(n21279), .A2(n18871), .ZN(n18892) );
  NAND2_X1 U12580 ( .A1(n11605), .A2(n11604), .ZN(n21747) );
  NAND2_X1 U12581 ( .A1(n21731), .A2(n21898), .ZN(n11605) );
  NAND2_X1 U12582 ( .A1(n21730), .A2(n21819), .ZN(n11604) );
  NAND2_X1 U12583 ( .A1(n18662), .A2(n12571), .ZN(n21758) );
  OR3_X1 U12584 ( .A1(n12740), .A2(n11544), .A3(n21503), .ZN(n21788) );
  NAND2_X1 U12585 ( .A1(n11545), .A2(n21826), .ZN(n11544) );
  INV_X1 U12586 ( .A(n21528), .ZN(n21875) );
  NOR2_X1 U12587 ( .A1(n11372), .A2(n11256), .ZN(n18730) );
  INV_X1 U12588 ( .A(n12559), .ZN(n11372) );
  NOR2_X1 U12589 ( .A1(n21661), .A2(n18750), .ZN(n21657) );
  INV_X1 U12590 ( .A(n21885), .ZN(n21849) );
  OAI21_X1 U12591 ( .B1(n21665), .B2(n21613), .A(n21856), .ZN(n21890) );
  INV_X1 U12592 ( .A(n21794), .ZN(n21819) );
  INV_X1 U12593 ( .A(n21788), .ZN(n21843) );
  INV_X1 U12594 ( .A(n21773), .ZN(n21881) );
  INV_X1 U12595 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19403) );
  INV_X1 U12596 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19383) );
  INV_X1 U12597 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n21481) );
  NAND2_X1 U12598 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21485) );
  INV_X1 U12599 ( .A(n21892), .ZN(n16299) );
  INV_X1 U12600 ( .A(n21926), .ZN(n21948) );
  NAND2_X1 U12601 ( .A1(n21947), .A2(n11383), .ZN(n21936) );
  INV_X1 U12602 ( .A(n11384), .ZN(n11383) );
  INV_X1 U12603 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21937) );
  INV_X1 U12604 ( .A(n18990), .ZN(n18996) );
  CLKBUF_X1 U12605 ( .A(n19713), .Z(n19671) );
  OAI21_X1 U12606 ( .B1(n16943), .B2(n20696), .A(n13805), .ZN(P1_U2968) );
  AND2_X1 U12607 ( .A1(n14653), .A2(n14652), .ZN(n14654) );
  NOR2_X1 U12608 ( .A1(n11226), .A2(n11640), .ZN(n17545) );
  AND2_X1 U12609 ( .A1(n14296), .A2(n14295), .ZN(n14297) );
  OR2_X1 U12610 ( .A1(n15047), .A2(n15046), .ZN(n15087) );
  AOI21_X1 U12611 ( .B1(n11476), .B2(n21934), .A(n11472), .ZN(n21250) );
  NAND2_X1 U12612 ( .A1(n11474), .A2(n11473), .ZN(n11472) );
  OAI211_X1 U12613 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n21382), .A(n11327), .B(
        n11326), .ZN(P3_U2704) );
  NAND2_X1 U12614 ( .A1(n21419), .A2(BUF2_REG_31__SCAN_IN), .ZN(n11326) );
  NAND2_X1 U12615 ( .A1(n11328), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n11327) );
  OAI21_X1 U12616 ( .B1(n21742), .B2(n18765), .A(n11567), .ZN(P3_U2801) );
  AND2_X1 U12617 ( .A1(n11572), .A2(n11267), .ZN(n11567) );
  OR2_X1 U12618 ( .A1(n18723), .A2(n18722), .ZN(n11572) );
  AOI21_X1 U12619 ( .B1(n12754), .B2(n21856), .A(n12753), .ZN(n12755) );
  OR2_X1 U12620 ( .A1(n20711), .A2(n20764), .ZN(U212) );
  NOR2_X1 U12621 ( .A1(n12443), .A2(n12444), .ZN(n12498) );
  CLKBUF_X3 U12622 ( .A(n11969), .Z(n14616) );
  AND2_X1 U12623 ( .A1(n11714), .A2(n11711), .ZN(n11177) );
  NAND2_X1 U12624 ( .A1(n11582), .A2(n11580), .ZN(n17236) );
  INV_X1 U12625 ( .A(n12009), .ZN(n13915) );
  INV_X1 U12626 ( .A(n11721), .ZN(n11720) );
  NAND2_X1 U12627 ( .A1(n11582), .A2(n11755), .ZN(n17247) );
  OR2_X1 U12628 ( .A1(n18528), .A2(n12550), .ZN(n11178) );
  NAND2_X1 U12629 ( .A1(n11603), .A2(n11200), .ZN(n11179) );
  OR3_X1 U12630 ( .A1(n16258), .A2(n11245), .A3(n11630), .ZN(n11180) );
  AND2_X1 U12631 ( .A1(n11338), .A2(n11257), .ZN(n11181) );
  NAND2_X1 U12632 ( .A1(n11678), .A2(n11681), .ZN(n16592) );
  NAND2_X1 U12633 ( .A1(n14027), .A2(n11254), .ZN(n11182) );
  AND2_X1 U12634 ( .A1(n17475), .A2(n11298), .ZN(n11183) );
  AND2_X2 U12635 ( .A1(n14070), .A2(n11761), .ZN(n11937) );
  INV_X1 U12636 ( .A(n11937), .ZN(n11760) );
  AND2_X1 U12637 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11184) );
  INV_X1 U12638 ( .A(n11976), .ZN(n15643) );
  OR2_X1 U12639 ( .A1(n14240), .A2(n11731), .ZN(n11185) );
  AND2_X1 U12640 ( .A1(n21279), .A2(n18107), .ZN(n11186) );
  AND2_X1 U12641 ( .A1(n12229), .A2(n11241), .ZN(n11187) );
  INV_X1 U12642 ( .A(n11716), .ZN(n11713) );
  NAND2_X1 U12643 ( .A1(n11259), .A2(n14247), .ZN(n11716) );
  AND2_X1 U12644 ( .A1(n18793), .A2(n21600), .ZN(n11188) );
  AND2_X1 U12645 ( .A1(n11469), .A2(n11467), .ZN(n11189) );
  OR2_X1 U12646 ( .A1(n12740), .A2(n21503), .ZN(n11547) );
  AND2_X1 U12647 ( .A1(n11252), .A2(n16237), .ZN(n11190) );
  INV_X1 U12648 ( .A(n13250), .ZN(n13265) );
  AND2_X1 U12649 ( .A1(n11603), .A2(n14393), .ZN(n11191) );
  AND2_X1 U12650 ( .A1(n18793), .A2(n21844), .ZN(n11192) );
  AND2_X1 U12651 ( .A1(n11465), .A2(n11263), .ZN(n11193) );
  AND2_X1 U12652 ( .A1(n14003), .A2(n17752), .ZN(n11194) );
  INV_X1 U12653 ( .A(n17251), .ZN(n11582) );
  INV_X1 U12654 ( .A(n13920), .ZN(n11413) );
  AND2_X1 U12655 ( .A1(n11193), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11195) );
  NOR2_X1 U12656 ( .A1(n11272), .A2(n11408), .ZN(n11196) );
  AND2_X1 U12657 ( .A1(n11625), .A2(n16582), .ZN(n11197) );
  AND2_X1 U12658 ( .A1(n11264), .A2(n13038), .ZN(n11198) );
  AND2_X1 U12659 ( .A1(n16066), .A2(n11294), .ZN(n11199) );
  INV_X1 U12660 ( .A(n21114), .ZN(n11463) );
  AND2_X1 U12661 ( .A1(n11299), .A2(n14393), .ZN(n11200) );
  AND2_X1 U12662 ( .A1(n11480), .A2(n14754), .ZN(n11201) );
  INV_X1 U12663 ( .A(n14064), .ZN(n11421) );
  INV_X1 U12664 ( .A(n14260), .ZN(n11423) );
  AND2_X1 U12665 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11202) );
  AND2_X1 U12666 ( .A1(n11202), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11203) );
  AND2_X1 U12667 ( .A1(n11203), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11204) );
  INV_X1 U12668 ( .A(n12321), .ZN(n12352) );
  OR3_X1 U12669 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21492), .A3(
        n16298), .ZN(n11205) );
  INV_X1 U12670 ( .A(n18172), .ZN(n12489) );
  NAND2_X1 U12671 ( .A1(n11399), .A2(n12976), .ZN(n13071) );
  OR2_X1 U12672 ( .A1(n12421), .A2(n17443), .ZN(n11206) );
  OR2_X1 U12673 ( .A1(n14261), .A2(n11422), .ZN(n11207) );
  AND2_X1 U12674 ( .A1(n11447), .A2(n14234), .ZN(n11208) );
  NOR2_X1 U12675 ( .A1(n12587), .A2(n12586), .ZN(n21278) );
  INV_X1 U12676 ( .A(n21278), .ZN(n11381) );
  OR2_X1 U12677 ( .A1(n13105), .A2(n13050), .ZN(n11210) );
  NAND2_X1 U12678 ( .A1(n11709), .A2(n11710), .ZN(n17421) );
  AND2_X1 U12679 ( .A1(n16547), .A2(n11675), .ZN(n16524) );
  AND4_X1 U12680 ( .A1(n12494), .A2(n12493), .A3(n12492), .A4(n12491), .ZN(
        n11211) );
  NOR2_X1 U12681 ( .A1(n16712), .A2(n16713), .ZN(n16620) );
  NAND2_X1 U12682 ( .A1(n17123), .A2(n17227), .ZN(n17218) );
  NAND2_X1 U12683 ( .A1(n16225), .A2(n11687), .ZN(n16272) );
  AND2_X1 U12684 ( .A1(n17521), .A2(n11203), .ZN(n11212) );
  AND2_X1 U12685 ( .A1(n17123), .A2(n11610), .ZN(n11213) );
  OR2_X1 U12686 ( .A1(n11645), .A2(n16102), .ZN(n11214) );
  OR2_X1 U12687 ( .A1(n17232), .A2(n14553), .ZN(n11215) );
  AND2_X1 U12688 ( .A1(n11441), .A2(n11208), .ZN(n11216) );
  OR3_X1 U12689 ( .A1(n14177), .A2(n17470), .A3(n19304), .ZN(n11217) );
  INV_X1 U12690 ( .A(n14007), .ZN(n17717) );
  AND2_X1 U12691 ( .A1(n14063), .A2(n14062), .ZN(n11218) );
  AND2_X1 U12692 ( .A1(n16547), .A2(n16548), .ZN(n11219) );
  AND2_X1 U12693 ( .A1(n17475), .A2(n11433), .ZN(n11220) );
  INV_X1 U12694 ( .A(n11382), .ZN(n19632) );
  OR2_X1 U12695 ( .A1(n12598), .A2(n12597), .ZN(n11382) );
  NAND2_X1 U12696 ( .A1(n17940), .A2(n13998), .ZN(n17751) );
  OAI21_X1 U12697 ( .B1(n17966), .B2(n17967), .A(n14016), .ZN(n17702) );
  NAND2_X1 U12698 ( .A1(n11726), .A2(n11732), .ZN(n17684) );
  NAND2_X1 U12699 ( .A1(n11712), .A2(n11714), .ZN(n17439) );
  AND2_X1 U12700 ( .A1(n13793), .A2(n16963), .ZN(n11221) );
  OR3_X1 U12701 ( .A1(n14177), .A2(n17470), .A3(n18008), .ZN(n11222) );
  AND4_X1 U12702 ( .A1(n12613), .A2(n11539), .A3(n12612), .A4(n11538), .ZN(
        n11223) );
  AND2_X1 U12703 ( .A1(n11557), .A2(n11178), .ZN(n11224) );
  AND4_X1 U12704 ( .A1(n11764), .A2(n11765), .A3(n11936), .A4(n11766), .ZN(
        n11225) );
  AND2_X1 U12705 ( .A1(n17542), .A2(n19281), .ZN(n11226) );
  XNOR2_X1 U12706 ( .A(n17232), .B(n14550), .ZN(n17224) );
  OR3_X1 U12707 ( .A1(n14261), .A2(n14260), .A3(n11906), .ZN(n11227) );
  NOR2_X1 U12708 ( .A1(n15497), .A2(n11622), .ZN(n11228) );
  NAND2_X1 U12709 ( .A1(n17532), .A2(n17530), .ZN(n17531) );
  AND3_X1 U12710 ( .A1(n11940), .A2(n11941), .A3(n11939), .ZN(n11229) );
  AND2_X1 U12711 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11230) );
  NAND2_X1 U12712 ( .A1(n16225), .A2(n16269), .ZN(n16273) );
  OR2_X1 U12713 ( .A1(n18793), .A2(n18637), .ZN(n11231) );
  OR2_X1 U12714 ( .A1(n21758), .A2(n12572), .ZN(n11232) );
  INV_X1 U12715 ( .A(n11434), .ZN(n17452) );
  NAND2_X1 U12716 ( .A1(n17475), .A2(n14294), .ZN(n11434) );
  INV_X1 U12717 ( .A(n14106), .ZN(n14107) );
  AND2_X1 U12718 ( .A1(n12004), .A2(n11364), .ZN(n11233) );
  AND2_X1 U12719 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11234) );
  INV_X1 U12720 ( .A(n11321), .ZN(n16472) );
  NOR3_X1 U12721 ( .A1(n16492), .A2(n20573), .A3(n20570), .ZN(n11321) );
  NAND2_X1 U12722 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12541), .ZN(
        n11235) );
  NAND2_X1 U12723 ( .A1(n20681), .A2(n13778), .ZN(n11236) );
  INV_X1 U12724 ( .A(n11448), .ZN(n11447) );
  NAND2_X1 U12725 ( .A1(n11218), .A2(n11449), .ZN(n11448) );
  NAND2_X1 U12726 ( .A1(n14245), .A2(n14244), .ZN(n17462) );
  AND2_X1 U12727 ( .A1(n13770), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11237) );
  INV_X1 U12728 ( .A(n14316), .ZN(n11704) );
  OR2_X1 U12729 ( .A1(n16298), .A2(n12443), .ZN(n11238) );
  AND2_X1 U12730 ( .A1(n17245), .A2(n17136), .ZN(n17124) );
  AND2_X1 U12731 ( .A1(n16155), .A2(n16154), .ZN(n11239) );
  NOR2_X1 U12732 ( .A1(n11381), .A2(n21438), .ZN(n12689) );
  NAND2_X1 U12733 ( .A1(n11724), .A2(n11727), .ZN(n17464) );
  AND2_X1 U12734 ( .A1(n11671), .A2(n13788), .ZN(n11240) );
  AND2_X1 U12735 ( .A1(n11644), .A2(n16079), .ZN(n11241) );
  AND2_X1 U12736 ( .A1(n11559), .A2(n11235), .ZN(n11242) );
  AND2_X1 U12737 ( .A1(n11742), .A2(n14336), .ZN(n11243) );
  NAND2_X1 U12738 ( .A1(n11704), .A2(n14310), .ZN(n11244) );
  INV_X1 U12739 ( .A(n13786), .ZN(n11670) );
  OR2_X1 U12740 ( .A1(n16286), .A2(n20608), .ZN(n11245) );
  INV_X1 U12741 ( .A(n18766), .ZN(n11468) );
  NOR3_X1 U12742 ( .A1(n12740), .A2(n21503), .A3(n11543), .ZN(n11246) );
  NOR2_X1 U12743 ( .A1(n17689), .A2(n11649), .ZN(n16208) );
  NAND2_X1 U12744 ( .A1(n13903), .A2(n11412), .ZN(n13919) );
  OR2_X1 U12745 ( .A1(n13996), .A2(n11416), .ZN(n13999) );
  OR2_X1 U12746 ( .A1(n16046), .A2(n15862), .ZN(n16045) );
  AND2_X1 U12747 ( .A1(n17264), .A2(n17263), .ZN(n17255) );
  NAND2_X1 U12748 ( .A1(n15880), .A2(n11579), .ZN(n16039) );
  NOR2_X1 U12749 ( .A1(n16244), .A2(n11601), .ZN(n17253) );
  NOR2_X1 U12750 ( .A1(n17251), .A2(n11583), .ZN(n17240) );
  AND2_X1 U12751 ( .A1(n16232), .A2(n16241), .ZN(n16239) );
  NAND2_X1 U12752 ( .A1(n11468), .A2(n11469), .ZN(n18549) );
  AOI21_X1 U12753 ( .B1(n11734), .B2(n14016), .A(n11733), .ZN(n11732) );
  INV_X1 U12754 ( .A(n11732), .ZN(n11731) );
  AND2_X1 U12755 ( .A1(n14118), .A2(n17256), .ZN(n11247) );
  AND2_X1 U12756 ( .A1(n11247), .A2(n11618), .ZN(n11248) );
  AND2_X1 U12757 ( .A1(n18519), .A2(n11465), .ZN(n11249) );
  NAND2_X1 U12758 ( .A1(n11345), .A2(n11344), .ZN(n11342) );
  OR2_X1 U12759 ( .A1(n13996), .A2(n13995), .ZN(n11250) );
  OR3_X1 U12760 ( .A1(n21735), .A2(n21821), .A3(n21734), .ZN(n11251) );
  AND2_X1 U12761 ( .A1(n17124), .A2(n17125), .ZN(n17123) );
  AND2_X1 U12762 ( .A1(n11615), .A2(n11614), .ZN(n11252) );
  XNOR2_X1 U12763 ( .A(n14315), .B(n11414), .ZN(n14313) );
  OAI22_X1 U12764 ( .A1(n17251), .A2(n11348), .B1(n14531), .B2(n11354), .ZN(
        n17231) );
  NOR3_X1 U12765 ( .A1(n17556), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n17541), .ZN(n11253) );
  NAND2_X1 U12766 ( .A1(n17919), .A2(n17918), .ZN(n17917) );
  AND2_X1 U12767 ( .A1(n11427), .A2(n14028), .ZN(n11254) );
  AND2_X1 U12768 ( .A1(n14256), .A2(n17442), .ZN(n11255) );
  NAND2_X1 U12769 ( .A1(n13130), .A2(n13129), .ZN(n15861) );
  OR2_X1 U12770 ( .A1(n12560), .A2(n11192), .ZN(n11256) );
  AND2_X1 U12771 ( .A1(n11199), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11257) );
  OR2_X1 U12772 ( .A1(n14688), .A2(n14689), .ZN(n11258) );
  NAND2_X1 U12773 ( .A1(n14250), .A2(n17453), .ZN(n11259) );
  NOR2_X1 U12774 ( .A1(n17754), .A2(n11708), .ZN(n11260) );
  AND2_X1 U12775 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11261) );
  OR2_X1 U12776 ( .A1(n11845), .A2(n13908), .ZN(n11262) );
  AND2_X1 U12777 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11263) );
  INV_X1 U12778 ( .A(n17937), .ZN(n11454) );
  NAND2_X1 U12779 ( .A1(n16714), .A2(n11625), .ZN(n11629) );
  NAND2_X1 U12780 ( .A1(n18501), .A2(n12549), .ZN(n21762) );
  AND2_X1 U12781 ( .A1(n11409), .A2(n13132), .ZN(n11264) );
  AND3_X1 U12782 ( .A1(n11388), .A2(n11387), .A3(n11385), .ZN(n11265) );
  AND2_X1 U12783 ( .A1(n11675), .A2(n16525), .ZN(n11266) );
  AND2_X1 U12784 ( .A1(n11571), .A2(n11568), .ZN(n11267) );
  AND2_X1 U12785 ( .A1(n11458), .A2(n11463), .ZN(n11268) );
  AND2_X1 U12786 ( .A1(n11248), .A2(n11617), .ZN(n11269) );
  AND2_X1 U12787 ( .A1(n21125), .A2(n11464), .ZN(n11270) );
  AND2_X1 U12788 ( .A1(n11189), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11271) );
  AND2_X1 U12789 ( .A1(n11667), .A2(n16927), .ZN(n11272) );
  NOR2_X1 U12790 ( .A1(n16231), .A2(n16238), .ZN(n11273) );
  NAND2_X1 U12791 ( .A1(n11338), .A2(n16066), .ZN(n15498) );
  AND2_X1 U12792 ( .A1(n11338), .A2(n11199), .ZN(n15486) );
  NAND2_X1 U12793 ( .A1(n11181), .A2(n11350), .ZN(n15777) );
  NAND2_X1 U12794 ( .A1(n11181), .A2(n15536), .ZN(n15535) );
  NAND2_X1 U12795 ( .A1(n15880), .A2(n15882), .ZN(n15881) );
  INV_X1 U12796 ( .A(n11333), .ZN(n12705) );
  OR2_X1 U12797 ( .A1(n11382), .A2(n21335), .ZN(n11333) );
  INV_X1 U12798 ( .A(n11548), .ZN(n18871) );
  OR2_X1 U12799 ( .A1(n21924), .A2(n21948), .ZN(n11548) );
  INV_X1 U12800 ( .A(n13902), .ZN(n14324) );
  AND3_X1 U12801 ( .A1(n11995), .A2(n11722), .A3(n15153), .ZN(n14212) );
  AND2_X1 U12802 ( .A1(n16094), .A2(n11619), .ZN(n15531) );
  NOR2_X1 U12803 ( .A1(n16139), .A2(n16138), .ZN(n15233) );
  NOR2_X1 U12804 ( .A1(n11365), .A2(n14195), .ZN(n14202) );
  AND2_X1 U12805 ( .A1(n16096), .A2(n12078), .ZN(n16094) );
  OR3_X1 U12806 ( .A1(n16258), .A2(n11245), .A3(n11632), .ZN(n11274) );
  AND2_X1 U12807 ( .A1(n11843), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11275) );
  AND2_X1 U12808 ( .A1(n11636), .A2(n11635), .ZN(n11276) );
  AND2_X1 U12809 ( .A1(n11843), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11277) );
  AND2_X1 U12810 ( .A1(n11420), .A2(n11419), .ZN(n11278) );
  OR2_X1 U12811 ( .A1(n21458), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n11279) );
  XOR2_X1 U12812 ( .A(n22085), .B(n14752), .Z(n11280) );
  AND2_X1 U12813 ( .A1(n13203), .A2(n16269), .ZN(n11281) );
  AND2_X1 U12814 ( .A1(n11462), .A2(n11463), .ZN(n11282) );
  NOR2_X1 U12815 ( .A1(n14607), .A2(n11595), .ZN(n11283) );
  AND2_X1 U12816 ( .A1(n14011), .A2(n19246), .ZN(n17967) );
  INV_X1 U12817 ( .A(n17967), .ZN(n11735) );
  OR2_X1 U12818 ( .A1(n21180), .A2(n21168), .ZN(n11284) );
  AND2_X1 U12819 ( .A1(n22256), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11285) );
  OR2_X1 U12820 ( .A1(n14756), .A2(n14755), .ZN(n11286) );
  INV_X1 U12821 ( .A(n21143), .ZN(n11464) );
  AND2_X1 U12822 ( .A1(n12229), .A2(n11644), .ZN(n11287) );
  AND2_X1 U12823 ( .A1(n14727), .A2(n11536), .ZN(n11288) );
  AND2_X1 U12824 ( .A1(n11579), .A2(n11578), .ZN(n11289) );
  AND2_X1 U12825 ( .A1(n11460), .A2(n11463), .ZN(n11290) );
  NOR2_X2 U12826 ( .A1(n15113), .A2(n14120), .ZN(n11291) );
  AND2_X2 U12827 ( .A1(n13683), .A2(n22497), .ZN(n20689) );
  AND2_X1 U12828 ( .A1(n14780), .A2(n11491), .ZN(n11292) );
  INV_X1 U12829 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11312) );
  AND2_X1 U12830 ( .A1(n18728), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18503) );
  NOR2_X1 U12831 ( .A1(n18854), .A2(n12540), .ZN(n11293) );
  INV_X1 U12832 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11623) );
  AND2_X1 U12833 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11294) );
  AND4_X1 U12834 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n11295)
         );
  AND2_X1 U12835 ( .A1(n14568), .A2(n14588), .ZN(n11296) );
  INV_X1 U12836 ( .A(n14287), .ZN(n11657) );
  AND2_X1 U12837 ( .A1(n11468), .A2(n11189), .ZN(n11297) );
  INV_X1 U12838 ( .A(n17210), .ZN(n11595) );
  INV_X1 U12839 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11470) );
  AND2_X1 U12840 ( .A1(n14294), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11298) );
  OR2_X1 U12841 ( .A1(n14403), .A2(n14402), .ZN(n11299) );
  AND2_X1 U12842 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput_216), .ZN(n11300)
         );
  INV_X1 U12843 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11403) );
  INV_X1 U12844 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11585) );
  INV_X1 U12845 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11414) );
  NOR2_X1 U12846 ( .A1(n22335), .A2(n22333), .ZN(n18990) );
  OAI22_X2 U12847 ( .A1(n15555), .A2(n15596), .B1(n20759), .B2(n15595), .ZN(
        n22753) );
  OAI22_X2 U12848 ( .A1(n15574), .A2(n15596), .B1(n20755), .B2(n15595), .ZN(
        n22657) );
  INV_X1 U12849 ( .A(n22538), .ZN(n11301) );
  INV_X1 U12850 ( .A(n11301), .ZN(n11302) );
  AOI22_X2 U12851 ( .A1(n20264), .A2(BUF2_REG_31__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19979) );
  NOR3_X2 U12852 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21930), .A3(
        n19432), .ZN(n19775) );
  NOR3_X2 U12853 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21930), .A3(
        n19451), .ZN(n19800) );
  INV_X1 U12854 ( .A(n22546), .ZN(n11303) );
  INV_X1 U12855 ( .A(n11303), .ZN(n11304) );
  INV_X1 U12856 ( .A(n22665), .ZN(n11305) );
  INV_X1 U12857 ( .A(n11305), .ZN(n11306) );
  INV_X1 U12858 ( .A(n22771), .ZN(n11307) );
  INV_X1 U12859 ( .A(n11307), .ZN(n11308) );
  INV_X1 U12860 ( .A(n22635), .ZN(n11309) );
  INV_X1 U12861 ( .A(n11309), .ZN(n11310) );
  OAI22_X2 U12862 ( .A1(n15597), .A2(n15596), .B1(n20766), .B2(n15595), .ZN(
        n22576) );
  OAI21_X1 U12863 ( .B1(n16325), .B2(n19304), .A(n11243), .ZN(P2_U3016) );
  INV_X1 U12864 ( .A(n19304), .ZN(n19335) );
  NOR3_X2 U12865 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21930), .A3(
        n19412), .ZN(n19750) );
  AOI22_X2 U12866 ( .A1(n20264), .A2(BUF2_REG_26__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n20236) );
  NOR2_X2 U12867 ( .A1(n15306), .A2(n15057), .ZN(n20263) );
  OAI22_X2 U12868 ( .A1(n15543), .A2(n15596), .B1(n20745), .B2(n15595), .ZN(
        n22477) );
  INV_X2 U12869 ( .A(n11172), .ZN(n19193) );
  AND2_X4 U12870 ( .A1(n11312), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17051) );
  INV_X2 U12871 ( .A(n12895), .ZN(n15813) );
  NAND3_X1 U12872 ( .A1(n12854), .A2(n12860), .A3(n12851), .ZN(n11318) );
  NOR2_X2 U12873 ( .A1(n21500), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12521) );
  OR2_X2 U12874 ( .A1(n21492), .A2(n12444), .ZN(n21500) );
  INV_X2 U12875 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20877) );
  INV_X1 U12876 ( .A(n21398), .ZN(n21403) );
  NAND4_X1 U12877 ( .A1(n21334), .A2(P3_EAX_REG_11__SCAN_IN), .A3(
        P3_EAX_REG_14__SCAN_IN), .A4(n11295), .ZN(n11330) );
  NAND3_X1 U12878 ( .A1(n12688), .A2(n11334), .A3(n11333), .ZN(n11332) );
  AND2_X4 U12879 ( .A1(n14070), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11976) );
  AND2_X2 U12880 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14070) );
  XNOR2_X1 U12881 ( .A(n11335), .B(n13807), .ZN(n14368) );
  INV_X1 U12882 ( .A(n11594), .ZN(n17214) );
  NAND2_X1 U12883 ( .A1(n14352), .A2(n14351), .ZN(n14379) );
  NAND2_X1 U12884 ( .A1(n14352), .A2(n11336), .ZN(n14356) );
  NOR2_X1 U12885 ( .A1(n11337), .A2(n14355), .ZN(n11336) );
  INV_X1 U12886 ( .A(n14351), .ZN(n11337) );
  AOI21_X1 U12887 ( .B1(n11352), .B2(n13806), .A(n11752), .ZN(n16096) );
  XNOR2_X2 U12888 ( .A(n11352), .B(n13806), .ZN(n13822) );
  NAND2_X2 U12889 ( .A1(n11153), .A2(n11156), .ZN(n12003) );
  NAND2_X1 U12890 ( .A1(n11767), .A2(n11225), .ZN(n11353) );
  NAND3_X1 U12891 ( .A1(n11362), .A2(n12005), .A3(n11361), .ZN(n12051) );
  INV_X1 U12892 ( .A(n13963), .ZN(n13965) );
  NAND3_X1 U12893 ( .A1(n17532), .A2(n17530), .A3(n11367), .ZN(n11368) );
  NAND2_X2 U12894 ( .A1(n18004), .A2(n14236), .ZN(n17505) );
  NAND2_X1 U12895 ( .A1(n12559), .A2(n11371), .ZN(n18729) );
  NOR2_X2 U12896 ( .A1(n18553), .A2(n11376), .ZN(n18771) );
  NAND3_X1 U12897 ( .A1(n21491), .A2(n21460), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11377) );
  NAND2_X1 U12898 ( .A1(n11378), .A2(n12697), .ZN(n11379) );
  INV_X1 U12899 ( .A(n21473), .ZN(n11378) );
  OAI21_X1 U12900 ( .B1(n21927), .B2(n21928), .A(n21926), .ZN(n11384) );
  INV_X2 U12901 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21491) );
  NAND2_X1 U12902 ( .A1(n13092), .A2(n13063), .ZN(n15435) );
  NAND2_X2 U12903 ( .A1(n13007), .A2(n13060), .ZN(n13092) );
  NAND3_X1 U12904 ( .A1(n13601), .A2(n15382), .A3(n11398), .ZN(n11397) );
  NAND2_X1 U12905 ( .A1(n15121), .A2(n12889), .ZN(n11398) );
  AND2_X2 U12906 ( .A1(n13659), .A2(n12895), .ZN(n15121) );
  NAND2_X1 U12907 ( .A1(n15134), .A2(n16376), .ZN(n13601) );
  NOR2_X2 U12908 ( .A1(n12890), .A2(n13686), .ZN(n15134) );
  NAND2_X1 U12909 ( .A1(n11400), .A2(n12976), .ZN(n13061) );
  INV_X1 U12910 ( .A(n16876), .ZN(n11404) );
  NAND2_X1 U12911 ( .A1(n11672), .A2(n16903), .ZN(n11406) );
  NAND2_X1 U12912 ( .A1(n11221), .A2(n16821), .ZN(n16326) );
  NAND2_X1 U12913 ( .A1(n13039), .A2(n13038), .ZN(n13105) );
  INV_X1 U12914 ( .A(n13908), .ZN(n11411) );
  NAND2_X1 U12915 ( .A1(n13903), .A2(n11410), .ZN(n13991) );
  NAND3_X1 U12916 ( .A1(n14257), .A2(n14266), .A3(n11423), .ZN(n11422) );
  AND3_X4 U12917 ( .A1(n15673), .A2(n11428), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11969) );
  NOR2_X2 U12918 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11606) );
  NAND2_X2 U12919 ( .A1(n17748), .A2(n14115), .ZN(n17716) );
  NAND2_X1 U12920 ( .A1(n17529), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14111) );
  NAND2_X1 U12921 ( .A1(n11577), .A2(n11429), .ZN(n17529) );
  NAND2_X1 U12922 ( .A1(n14109), .A2(n16154), .ZN(n11430) );
  NAND2_X1 U12923 ( .A1(n18006), .A2(n18005), .ZN(n18004) );
  NAND2_X1 U12924 ( .A1(n13901), .A2(n14088), .ZN(n17915) );
  NAND2_X1 U12925 ( .A1(n11440), .A2(n16056), .ZN(n13917) );
  NAND2_X1 U12926 ( .A1(n11440), .A2(n11438), .ZN(n11437) );
  OR2_X1 U12927 ( .A1(n17505), .A2(n11451), .ZN(n11441) );
  XNOR2_X2 U12928 ( .A(n18708), .B(n18691), .ZN(n21114) );
  INV_X1 U12929 ( .A(n11460), .ZN(n21178) );
  NAND2_X1 U12930 ( .A1(n21126), .A2(n11270), .ZN(n11461) );
  OAI21_X1 U12931 ( .B1(n11463), .B2(n21143), .A(n11461), .ZN(n21155) );
  NAND2_X1 U12932 ( .A1(n11468), .A2(n11271), .ZN(n18526) );
  NAND2_X1 U12933 ( .A1(n11478), .A2(n11479), .ZN(n14762) );
  NAND2_X1 U12934 ( .A1(n14751), .A2(n11201), .ZN(n11478) );
  INV_X1 U12935 ( .A(n14770), .ZN(n11484) );
  OAI21_X1 U12936 ( .B1(n11484), .B2(n11486), .A(n11485), .ZN(n14785) );
  INV_X1 U12937 ( .A(n14773), .ZN(n11492) );
  NAND3_X1 U12938 ( .A1(n12614), .A2(n12616), .A3(n11541), .ZN(n11540) );
  INV_X1 U12939 ( .A(n11547), .ZN(n21471) );
  INV_X1 U12940 ( .A(n12741), .ZN(n11546) );
  NAND3_X1 U12941 ( .A1(n12478), .A2(n12479), .A3(n12480), .ZN(n11553) );
  XNOR2_X1 U12942 ( .A(n18528), .B(n12550), .ZN(n18808) );
  NAND2_X1 U12943 ( .A1(n11178), .A2(n18808), .ZN(n11556) );
  NOR2_X2 U12944 ( .A1(n12443), .A2(n12445), .ZN(n12476) );
  NAND2_X1 U12945 ( .A1(n12540), .A2(n11562), .ZN(n11559) );
  NAND2_X1 U12946 ( .A1(n11558), .A2(n11559), .ZN(n18843) );
  NAND2_X1 U12947 ( .A1(n11954), .A2(n11994), .ZN(n11967) );
  NAND3_X1 U12948 ( .A1(n11222), .A2(n14145), .A3(n11575), .ZN(P2_U2994) );
  OR2_X1 U12949 ( .A1(n14179), .A2(n17996), .ZN(n11575) );
  NAND3_X1 U12950 ( .A1(n12032), .A2(n12031), .A3(n12030), .ZN(n13810) );
  INV_X2 U12951 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21460) );
  INV_X1 U12952 ( .A(n11740), .ZN(n11591) );
  NAND2_X1 U12953 ( .A1(n11594), .A2(n11591), .ZN(n11600) );
  INV_X1 U12954 ( .A(n14607), .ZN(n11599) );
  NOR2_X2 U12955 ( .A1(n21747), .A2(n11251), .ZN(n21736) );
  AND2_X4 U12956 ( .A1(n11606), .A2(n11761), .ZN(n11968) );
  NOR2_X1 U12957 ( .A1(n14071), .A2(n11606), .ZN(n15667) );
  INV_X1 U12958 ( .A(n15701), .ZN(n15635) );
  NAND2_X1 U12959 ( .A1(n14164), .A2(n11156), .ZN(n11608) );
  NAND2_X1 U12960 ( .A1(n11986), .A2(n14154), .ZN(n12038) );
  NAND2_X1 U12961 ( .A1(n15883), .A2(n11190), .ZN(n16214) );
  INV_X1 U12962 ( .A(n16122), .ZN(n11622) );
  AND2_X4 U12963 ( .A1(n12762), .A2(n17051), .ZN(n12848) );
  AND2_X2 U12964 ( .A1(n11623), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12762) );
  NAND3_X1 U12965 ( .A1(n15385), .A2(n11166), .A3(n11624), .ZN(n15387) );
  INV_X1 U12966 ( .A(n11629), .ZN(n16595) );
  AND2_X4 U12967 ( .A1(n15677), .A2(n15673), .ZN(n11960) );
  AND2_X2 U12968 ( .A1(n11762), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15677) );
  NAND2_X1 U12969 ( .A1(n15213), .A2(n11187), .ZN(n16080) );
  CLKBUF_X1 U12970 ( .A(n15213), .Z(n11643) );
  NOR2_X1 U12971 ( .A1(n11209), .A2(n14301), .ZN(n14286) );
  OR3_X1 U12972 ( .A1(n11209), .A2(n11652), .A3(n14301), .ZN(n17288) );
  NAND2_X1 U12973 ( .A1(n16201), .A2(n11658), .ZN(n11660) );
  NAND2_X1 U12974 ( .A1(n16903), .A2(n11240), .ZN(n11669) );
  NAND2_X1 U12975 ( .A1(n11673), .A2(n11405), .ZN(n11671) );
  XNOR2_X2 U12976 ( .A(n12952), .B(n12954), .ZN(n13083) );
  NAND2_X2 U12977 ( .A1(n11674), .A2(n12913), .ZN(n12952) );
  NAND2_X1 U12978 ( .A1(n16547), .A2(n11266), .ZN(n16510) );
  INV_X1 U12979 ( .A(n16510), .ZN(n13473) );
  NAND2_X1 U12980 ( .A1(n11677), .A2(n11676), .ZN(n16224) );
  NOR2_X1 U12981 ( .A1(n16712), .A2(n11683), .ZN(n16607) );
  NAND2_X1 U12982 ( .A1(n16474), .A2(n11690), .ZN(n16463) );
  NAND2_X1 U12983 ( .A1(n16474), .A2(n16475), .ZN(n16462) );
  AND2_X4 U12984 ( .A1(n11792), .A2(n15673), .ZN(n14633) );
  OAI211_X1 U12986 ( .C1(n17425), .C2(n11696), .A(n11693), .B(n11244), .ZN(
        n11694) );
  NAND2_X1 U12987 ( .A1(n17425), .A2(n11695), .ZN(n11693) );
  AOI21_X1 U12988 ( .B1(n17425), .B2(n11703), .A(n11700), .ZN(n11697) );
  OR2_X1 U12989 ( .A1(n17425), .A2(n14310), .ZN(n11698) );
  INV_X1 U12990 ( .A(n11702), .ZN(n11700) );
  OR2_X2 U12991 ( .A1(n13897), .A2(n13898), .ZN(n11706) );
  NAND2_X1 U12992 ( .A1(n13867), .A2(n13866), .ZN(n13899) );
  NAND2_X1 U12993 ( .A1(n14245), .A2(n11177), .ZN(n11709) );
  NAND3_X1 U12994 ( .A1(n11721), .A2(n14353), .A3(n16031), .ZN(n11717) );
  NAND3_X1 U12995 ( .A1(n11720), .A2(n11719), .A3(n11343), .ZN(n11718) );
  NAND2_X2 U12996 ( .A1(n12003), .A2(n11996), .ZN(n15153) );
  NAND2_X1 U12997 ( .A1(n14154), .A2(n20262), .ZN(n11996) );
  NAND2_X1 U12998 ( .A1(n14007), .A2(n14006), .ZN(n17966) );
  NAND2_X1 U12999 ( .A1(n14007), .A2(n11725), .ZN(n11724) );
  AND2_X1 U13000 ( .A1(n14069), .A2(n14068), .ZN(n14177) );
  NAND2_X1 U13001 ( .A1(n15531), .A2(n15779), .ZN(n15953) );
  NAND2_X1 U13002 ( .A1(n12187), .A2(n12186), .ZN(n17085) );
  INV_X1 U13003 ( .A(n12885), .ZN(n12892) );
  NAND2_X1 U13004 ( .A1(n12884), .A2(n12843), .ZN(n12844) );
  AND2_X2 U13005 ( .A1(n15430), .A2(n15429), .ZN(n12936) );
  NAND2_X1 U13006 ( .A1(n14111), .A2(n14110), .ZN(n17935) );
  AND2_X2 U13007 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15429) );
  NAND2_X1 U13008 ( .A1(n16466), .A2(n16454), .ZN(n16437) );
  OR2_X1 U13009 ( .A1(n16466), .A2(n16400), .ZN(n16438) );
  NAND4_X4 U13010 ( .A1(n12882), .A2(n12881), .A3(n12880), .A4(n12879), .ZN(
        n12891) );
  NAND2_X1 U13011 ( .A1(n13857), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13860) );
  OR2_X1 U13012 ( .A1(n14179), .A2(n19332), .ZN(n14227) );
  AND2_X4 U13013 ( .A1(n14617), .A2(n11936), .ZN(n14485) );
  AND2_X4 U13014 ( .A1(n11786), .A2(n11936), .ZN(n14480) );
  AND2_X2 U13015 ( .A1(n15598), .A2(n15384), .ZN(n15330) );
  CLKBUF_X1 U13016 ( .A(n12038), .Z(n15634) );
  NAND2_X1 U13017 ( .A1(n15609), .A2(n12923), .ZN(n15842) );
  OR2_X1 U13018 ( .A1(n14353), .A2(n12009), .ZN(n12017) );
  NAND2_X1 U13019 ( .A1(n16378), .A2(n13665), .ZN(n13682) );
  NAND2_X1 U13020 ( .A1(n13083), .A2(n22256), .ZN(n12969) );
  OR3_X2 U13021 ( .A1(n13856), .A2(n11171), .A3(n15439), .ZN(n19970) );
  NAND2_X1 U13022 ( .A1(n15439), .A2(n13855), .ZN(n13845) );
  AOI21_X1 U13023 ( .B1(n11937), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n11756), .ZN(n11955) );
  AOI22_X1 U13024 ( .A1(n11968), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11803) );
  AND2_X1 U13025 ( .A1(n16347), .A2(n13696), .ZN(n22405) );
  INV_X1 U13026 ( .A(n13696), .ZN(n15614) );
  AOI21_X1 U13027 ( .B1(n12071), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n12070), .ZN(n12074) );
  INV_X1 U13028 ( .A(n12071), .ZN(n17084) );
  AND2_X4 U13029 ( .A1(n17051), .A2(n15430), .ZN(n12829) );
  INV_X1 U13030 ( .A(n13053), .ZN(n13589) );
  INV_X1 U13031 ( .A(n13589), .ZN(n13469) );
  NOR2_X1 U13032 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14357) );
  INV_X1 U13033 ( .A(n14357), .ZN(n20002) );
  INV_X1 U13034 ( .A(n12192), .ZN(n12350) );
  INV_X1 U13035 ( .A(n12191), .ZN(n12351) );
  INV_X1 U13036 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n14346) );
  NAND2_X1 U13037 ( .A1(n20621), .A2(n15557), .ZN(n16724) );
  NAND2_X2 U13038 ( .A1(n15449), .A2(n15448), .ZN(n20621) );
  NAND2_X1 U13039 ( .A1(n15395), .A2(n16366), .ZN(n22112) );
  AND2_X1 U13040 ( .A1(n14061), .A2(n17646), .ZN(n17485) );
  NAND2_X1 U13041 ( .A1(n14842), .A2(n14841), .ZN(n11738) );
  OR2_X1 U13042 ( .A1(n14706), .A2(n14705), .ZN(n11739) );
  AND2_X1 U13043 ( .A1(n14569), .A2(n11296), .ZN(n11740) );
  AND2_X1 U13044 ( .A1(n14227), .A2(n14226), .ZN(n11741) );
  OR2_X1 U13045 ( .A1(n16320), .A2(n19332), .ZN(n11742) );
  AND2_X1 U13046 ( .A1(n11768), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11743) );
  INV_X1 U13047 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12569) );
  INV_X1 U13048 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14777) );
  INV_X1 U13049 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14311) );
  AND2_X1 U13050 ( .A1(n12893), .A2(n12842), .ZN(n11745) );
  INV_X1 U13051 ( .A(n20426), .ZN(n20431) );
  INV_X1 U13052 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12570) );
  AND2_X1 U13053 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n22284), .ZN(n22288) );
  INV_X1 U13054 ( .A(n16637), .ZN(n13272) );
  AND2_X1 U13055 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11746) );
  INV_X1 U13056 ( .A(n14310), .ZN(n14269) );
  AND2_X1 U13057 ( .A1(n21688), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11747) );
  INV_X1 U13058 ( .A(n12040), .ZN(n12026) );
  INV_X1 U13059 ( .A(n15057), .ZN(n17998) );
  NAND3_X1 U13060 ( .A1(n19846), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19932), 
        .ZN(n15057) );
  AND2_X1 U13061 ( .A1(n13599), .A2(P1_EAX_REG_5__SCAN_IN), .ZN(n11748) );
  OR2_X1 U13062 ( .A1(n21481), .A2(n18888), .ZN(n21891) );
  INV_X1 U13063 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13204) );
  AND4_X1 U13064 ( .A1(n14239), .A2(n14238), .A3(n14237), .A4(n17471), .ZN(
        n11749) );
  INV_X1 U13065 ( .A(n17483), .ZN(n14063) );
  AND2_X1 U13066 ( .A1(n17393), .A2(n17394), .ZN(n11750) );
  INV_X1 U13067 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n18691) );
  NOR2_X1 U13068 ( .A1(n12425), .A2(n12392), .ZN(n11751) );
  NAND2_X1 U13069 ( .A1(n18652), .A2(n18887), .ZN(n18693) );
  AND2_X1 U13070 ( .A1(n12074), .A2(n12073), .ZN(n11752) );
  AND2_X1 U13071 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11753) );
  OAI21_X1 U13072 ( .B1(n15066), .B2(n15065), .A(n14366), .ZN(n14367) );
  INV_X1 U13073 ( .A(n16306), .ZN(n15712) );
  INV_X1 U13074 ( .A(n19347), .ZN(n19194) );
  INV_X2 U13075 ( .A(n19549), .ZN(n19715) );
  INV_X1 U13076 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n14726) );
  OR3_X1 U13077 ( .A1(n17556), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14332), .ZN(n11754) );
  NOR2_X1 U13078 ( .A1(n12256), .A2(n12255), .ZN(n15534) );
  INV_X1 U13079 ( .A(n15776), .ZN(n14381) );
  OR2_X1 U13080 ( .A1(n14434), .A2(n14433), .ZN(n11755) );
  NAND2_X1 U13081 ( .A1(n17253), .A2(n17254), .ZN(n17251) );
  AND4_X1 U13082 ( .A1(n12833), .A2(n12832), .A3(n12831), .A4(n12830), .ZN(
        n11757) );
  AND2_X2 U13083 ( .A1(n12765), .A2(n17059), .ZN(n12956) );
  AND2_X1 U13084 ( .A1(n12897), .A2(n12896), .ZN(n11758) );
  AND4_X1 U13085 ( .A1(n12837), .A2(n12836), .A3(n12835), .A4(n12834), .ZN(
        n11759) );
  XNOR2_X1 U13086 ( .A(n14662), .B(DATAI_28_), .ZN(n14663) );
  NOR2_X1 U13087 ( .A1(n14659), .A2(n14658), .ZN(n14665) );
  OAI22_X1 U13088 ( .A1(n15568), .A2(keyinput_140), .B1(n14673), .B2(DATAI_20_), .ZN(n14674) );
  INV_X1 U13089 ( .A(n14674), .ZN(n14675) );
  OAI21_X1 U13090 ( .B1(DATAI_2_), .B2(keyinput_158), .A(n14704), .ZN(n14705)
         );
  NOR2_X1 U13091 ( .A1(n11739), .A2(n14709), .ZN(n14710) );
  NOR2_X1 U13092 ( .A1(n14715), .A2(keyinput_164), .ZN(n14716) );
  OAI22_X1 U13093 ( .A1(n14914), .A2(keyinput_165), .B1(n14720), .B2(READY2), 
        .ZN(n14721) );
  INV_X1 U13094 ( .A(keyinput_167), .ZN(n14725) );
  NAND2_X1 U13095 ( .A1(n14726), .A2(n14725), .ZN(n14727) );
  OAI22_X1 U13096 ( .A1(n20574), .A2(n14743), .B1(P1_REIP_REG_31__SCAN_IN), 
        .B2(keyinput_180), .ZN(n14744) );
  INV_X1 U13097 ( .A(keyinput_184), .ZN(n14752) );
  NOR2_X1 U13098 ( .A1(n20565), .A2(keyinput_187), .ZN(n14755) );
  OAI22_X1 U13099 ( .A1(n20563), .A2(keyinput_188), .B1(n14757), .B2(
        P1_REIP_REG_23__SCAN_IN), .ZN(n14758) );
  OAI22_X1 U13100 ( .A1(n20561), .A2(keyinput_189), .B1(n14759), .B2(
        P1_REIP_REG_22__SCAN_IN), .ZN(n14760) );
  AOI21_X1 U13101 ( .B1(n14762), .B2(n14761), .A(n14760), .ZN(n14763) );
  INV_X1 U13102 ( .A(keyinput_201), .ZN(n14776) );
  NAND2_X1 U13103 ( .A1(n14777), .A2(n14776), .ZN(n14778) );
  AND2_X1 U13104 ( .A1(n14779), .A2(n14778), .ZN(n14780) );
  XNOR2_X1 U13105 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_209), .ZN(n14790)
         );
  NOR2_X1 U13106 ( .A1(n14791), .A2(n14790), .ZN(n14792) );
  AND2_X1 U13107 ( .A1(n14797), .A2(n14796), .ZN(n14798) );
  INV_X1 U13108 ( .A(n15168), .ZN(n12887) );
  OAI22_X1 U13109 ( .A1(n20616), .A2(n14655), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(keyinput_228), .ZN(n14656) );
  NAND2_X1 U13110 ( .A1(n12888), .A2(n12887), .ZN(n12889) );
  OAI22_X1 U13111 ( .A1(n16720), .A2(keyinput_230), .B1(n14817), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14818) );
  OR2_X1 U13112 ( .A1(n19904), .A2(n13854), .ZN(n13861) );
  OAI22_X1 U13113 ( .A1(n22210), .A2(keyinput_231), .B1(n14819), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n14820) );
  NOR2_X1 U13114 ( .A1(n12026), .A2(n11753), .ZN(n12027) );
  AND2_X1 U13115 ( .A1(n11807), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11811) );
  INV_X1 U13116 ( .A(n11994), .ZN(n11995) );
  OAI22_X1 U13117 ( .A1(n16290), .A2(n14823), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(keyinput_232), .ZN(n14824) );
  INV_X1 U13118 ( .A(n16291), .ZN(n13203) );
  INV_X1 U13119 ( .A(n13102), .ZN(n13038) );
  INV_X1 U13120 ( .A(n13903), .ZN(n11845) );
  INV_X1 U13121 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11763) );
  NAND2_X1 U13122 ( .A1(n13881), .A2(n13880), .ZN(n13898) );
  NAND2_X1 U13123 ( .A1(n14106), .A2(n14324), .ZN(n13992) );
  INV_X1 U13124 ( .A(n14824), .ZN(n14825) );
  AND4_X1 U13125 ( .A1(n15570), .A2(n15583), .A3(n12892), .A4(n12842), .ZN(
        n12886) );
  INV_X1 U13126 ( .A(n16513), .ZN(n13472) );
  INV_X1 U13127 ( .A(n13057), .ZN(n13058) );
  OR2_X1 U13128 ( .A1(n13124), .A2(n13123), .ZN(n13754) );
  INV_X1 U13129 ( .A(n17733), .ZN(n14003) );
  INV_X1 U13130 ( .A(n12183), .ZN(n12069) );
  AND2_X1 U13131 ( .A1(n11947), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11951) );
  INV_X1 U13132 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12552) );
  AND2_X1 U13133 ( .A1(n22487), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13626) );
  AOI22_X1 U13134 ( .A1(n12955), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12813) );
  INV_X1 U13135 ( .A(n16537), .ZN(n13426) );
  NOR2_X1 U13136 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13053) );
  NAND2_X1 U13137 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13094) );
  OR2_X1 U13138 ( .A1(n13786), .A2(n13771), .ZN(n13772) );
  OR2_X1 U13139 ( .A1(n13024), .A2(n13023), .ZN(n13721) );
  INV_X1 U13140 ( .A(n16038), .ZN(n14382) );
  INV_X1 U13141 ( .A(n17719), .ZN(n14006) );
  AND2_X1 U13142 ( .A1(n14265), .A2(n17434), .ZN(n14316) );
  AND2_X1 U13143 ( .A1(n19146), .A2(n14067), .ZN(n14234) );
  AND2_X1 U13144 ( .A1(n12196), .A2(n12195), .ZN(n12214) );
  NAND2_X1 U13145 ( .A1(n14347), .A2(n14346), .ZN(n14369) );
  INV_X1 U13146 ( .A(n14367), .ZN(n15062) );
  OAI22_X1 U13147 ( .A1(n22369), .A2(keyinput_246), .B1(n14843), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n14844) );
  OAI21_X1 U13148 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21491), .A(
        n12662), .ZN(n12663) );
  INV_X1 U13149 ( .A(n18632), .ZN(n18633) );
  NOR2_X1 U13150 ( .A1(n21438), .A2(n19592), .ZN(n12706) );
  NAND2_X1 U13151 ( .A1(n13156), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13171) );
  AND2_X1 U13152 ( .A1(n16402), .A2(n16401), .ZN(n16613) );
  INV_X1 U13153 ( .A(n13561), .ZN(n13593) );
  INV_X1 U13154 ( .A(n12899), .ZN(n12900) );
  INV_X1 U13155 ( .A(n13112), .ZN(n13113) );
  NAND2_X1 U13156 ( .A1(n13790), .A2(n11667), .ZN(n13791) );
  AND2_X1 U13157 ( .A1(n13786), .A2(n22025), .ZN(n16908) );
  BUF_X1 U13158 ( .A(n16903), .Z(n20669) );
  OAI211_X1 U13159 ( .C1(n13624), .C2(n12972), .A(n12971), .B(n12970), .ZN(
        n13080) );
  INV_X1 U13160 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n22409) );
  INV_X1 U13161 ( .A(n22253), .ZN(n15428) );
  INV_X1 U13162 ( .A(n15593), .ZN(n22388) );
  INV_X1 U13163 ( .A(n14005), .ZN(n11900) );
  INV_X1 U13164 ( .A(n16093), .ZN(n12078) );
  AND2_X1 U13165 ( .A1(n11779), .A2(n11936), .ZN(n11783) );
  AND2_X1 U13166 ( .A1(n14317), .A2(n14316), .ZN(n14318) );
  INV_X1 U13167 ( .A(n17465), .ZN(n14244) );
  AND2_X1 U13168 ( .A1(n14059), .A2(n17633), .ZN(n17483) );
  NAND2_X1 U13169 ( .A1(n15060), .A2(n14375), .ZN(n15059) );
  NAND2_X1 U13170 ( .A1(n15062), .A2(n15061), .ZN(n15060) );
  INV_X1 U13171 ( .A(n13947), .ZN(n16027) );
  NAND2_X1 U13172 ( .A1(n15175), .A2(keyinput_254), .ZN(n14855) );
  INV_X1 U13173 ( .A(n20959), .ZN(n18502) );
  INV_X1 U13174 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12536) );
  NOR2_X1 U13175 ( .A1(n18818), .A2(n12548), .ZN(n18528) );
  OAI21_X1 U13176 ( .B1(n21939), .B2(n17814), .A(n21505), .ZN(n19384) );
  AND2_X1 U13177 ( .A1(n13608), .A2(n13610), .ZN(n13623) );
  NOR2_X1 U13178 ( .A1(n13171), .A2(n22175), .ZN(n13188) );
  NOR2_X1 U13179 ( .A1(n15331), .A2(n17039), .ZN(n16366) );
  NAND2_X1 U13180 ( .A1(n13658), .A2(n13657), .ZN(n15348) );
  INV_X1 U13181 ( .A(n16578), .ZN(n16593) );
  OR2_X1 U13182 ( .A1(n13786), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n20681) );
  OR2_X1 U13183 ( .A1(n13052), .A2(n22489), .ZN(n13250) );
  AND2_X1 U13184 ( .A1(n16285), .A2(n16284), .ZN(n20608) );
  NAND2_X1 U13185 ( .A1(n13733), .A2(n13732), .ZN(n16013) );
  AND2_X1 U13186 ( .A1(n22122), .A2(n22111), .ZN(n22018) );
  NAND2_X1 U13187 ( .A1(n12988), .A2(n12987), .ZN(n12989) );
  AND2_X1 U13188 ( .A1(n16347), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22416) );
  INV_X1 U13189 ( .A(n15963), .ZN(n15615) );
  OR2_X1 U13190 ( .A1(n15961), .A2(n15539), .ZN(n15621) );
  INV_X1 U13191 ( .A(n22405), .ZN(n15733) );
  NOR3_X1 U13192 ( .A1(n17865), .A2(n22259), .A3(n15428), .ZN(n15551) );
  OR2_X1 U13193 ( .A1(n15961), .A2(n15506), .ZN(n22493) );
  AOI21_X1 U13194 ( .B1(n22487), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n22388), 
        .ZN(n22495) );
  NAND2_X1 U13195 ( .A1(n12387), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12388) );
  NOR2_X2 U13196 ( .A1(n17377), .A2(n17363), .ZN(n17365) );
  AND2_X1 U13197 ( .A1(n11843), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n14024) );
  OR2_X1 U13198 ( .A1(n15111), .A2(n12434), .ZN(n19199) );
  OAI21_X1 U13199 ( .B1(n14074), .B2(n11916), .A(n14137), .ZN(n15699) );
  OR2_X1 U13200 ( .A1(n14587), .A2(n14591), .ZN(n17203) );
  INV_X1 U13201 ( .A(n17771), .ZN(n15069) );
  NOR2_X1 U13202 ( .A1(n12123), .A2(n12411), .ZN(n12410) );
  INV_X1 U13203 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17523) );
  NOR2_X1 U13204 ( .A1(n17932), .A2(n12398), .ZN(n12401) );
  OR2_X1 U13205 ( .A1(n17577), .A2(n14275), .ZN(n17556) );
  AOI21_X1 U13206 ( .B1(n19329), .B2(n14225), .A(n14224), .ZN(n14226) );
  OR2_X1 U13207 ( .A1(n19103), .A2(n14037), .ZN(n17992) );
  NOR2_X1 U13208 ( .A1(n14087), .A2(n14324), .ZN(n14114) );
  INV_X2 U13209 ( .A(n14368), .ZN(n17172) );
  OR2_X1 U13210 ( .A1(n14215), .A2(n14085), .ZN(n14178) );
  AND2_X1 U13211 ( .A1(n15663), .A2(n15662), .ZN(n17773) );
  OR2_X1 U13212 ( .A1(n19982), .A2(n18023), .ZN(n20006) );
  OR2_X1 U13213 ( .A1(n19860), .A2(n18018), .ZN(n19843) );
  OR2_X1 U13214 ( .A1(n19982), .A2(n20200), .ZN(n19952) );
  NAND2_X1 U13215 ( .A1(n14856), .A2(n14855), .ZN(n14857) );
  AND2_X1 U13216 ( .A1(n19982), .A2(n20200), .ZN(n19882) );
  NAND2_X1 U13217 ( .A1(n19932), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20261) );
  OAI21_X1 U13218 ( .B1(n12674), .B2(n12673), .A(n12672), .ZN(n21897) );
  NOR2_X1 U13219 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20998), .ZN(n21014) );
  NAND2_X1 U13220 ( .A1(n20852), .A2(n20853), .ZN(n21269) );
  NAND2_X1 U13221 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18462), .ZN(n18370) );
  INV_X1 U13222 ( .A(n12485), .ZN(n12497) );
  INV_X1 U13223 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n20974) );
  XNOR2_X1 U13224 ( .A(n12537), .B(n12536), .ZN(n18865) );
  INV_X1 U13225 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12574) );
  AND2_X1 U13226 ( .A1(n18793), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12571) );
  INV_X1 U13227 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21661) );
  NAND2_X1 U13228 ( .A1(n16300), .A2(n17834), .ZN(n21826) );
  INV_X1 U13229 ( .A(n21865), .ZN(n21876) );
  NAND2_X1 U13230 ( .A1(n20846), .A2(n19384), .ZN(n19591) );
  INV_X1 U13231 ( .A(n12699), .ZN(n12702) );
  OR2_X1 U13232 ( .A1(n16370), .A2(n15135), .ZN(n16374) );
  NAND2_X1 U13233 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n13189), .ZN(
        n13230) );
  INV_X1 U13234 ( .A(n22235), .ZN(n22201) );
  INV_X1 U13235 ( .A(n22197), .ZN(n22222) );
  AND2_X1 U13236 ( .A1(n15812), .A2(n15801), .ZN(n22199) );
  INV_X1 U13237 ( .A(n16724), .ZN(n20617) );
  INV_X1 U13238 ( .A(n16789), .ZN(n16775) );
  NAND2_X1 U13239 ( .A1(n15348), .A2(n20704), .ZN(n13664) );
  INV_X1 U13240 ( .A(n22379), .ZN(n15257) );
  NAND2_X1 U13241 ( .A1(n13358), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13379) );
  AND2_X1 U13242 ( .A1(n20646), .A2(n20631), .ZN(n20676) );
  INV_X1 U13243 ( .A(n22112), .ZN(n22021) );
  INV_X1 U13244 ( .A(n22018), .ZN(n21982) );
  NOR2_X1 U13245 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n17824) );
  OAI211_X1 U13246 ( .C1(n22393), .C2(n22489), .A(n22465), .B(n22392), .ZN(
        n22702) );
  AND2_X1 U13247 ( .A1(n22417), .A2(n22380), .ZN(n22708) );
  AND2_X1 U13248 ( .A1(n22417), .A2(n22405), .ZN(n22721) );
  OAI21_X1 U13249 ( .B1(n15970), .B2(n16009), .A(n22512), .ZN(n16005) );
  NOR2_X1 U13250 ( .A1(n15621), .A2(n22470), .ZN(n15985) );
  NOR2_X2 U13251 ( .A1(n15621), .A2(n22486), .ZN(n22727) );
  NOR2_X2 U13252 ( .A1(n15621), .A2(n15615), .ZN(n22735) );
  INV_X1 U13253 ( .A(n22533), .ZN(n22740) );
  NOR2_X2 U13254 ( .A1(n15846), .A2(n22486), .ZN(n22747) );
  OAI21_X1 U13255 ( .B1(n15735), .B2(n15736), .A(n22495), .ZN(n15759) );
  INV_X1 U13256 ( .A(n22472), .ZN(n22754) );
  NOR2_X2 U13257 ( .A1(n22493), .A2(n22470), .ZN(n22762) );
  INV_X1 U13258 ( .A(n22485), .ZN(n22507) );
  AND2_X1 U13259 ( .A1(n22250), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17865) );
  INV_X1 U13260 ( .A(HOLD), .ZN(n22334) );
  OR2_X1 U13261 ( .A1(n14151), .A2(n14138), .ZN(n15641) );
  INV_X1 U13262 ( .A(n19124), .ZN(n19182) );
  NAND2_X1 U13263 ( .A1(n16065), .A2(n15111), .ZN(n15107) );
  NOR2_X1 U13264 ( .A1(n19163), .A2(n14346), .ZN(n19124) );
  NOR2_X1 U13265 ( .A1(n11354), .A2(n14591), .ZN(n17210) );
  OR2_X1 U13266 ( .A1(n14424), .A2(n14423), .ZN(n17254) );
  AND2_X1 U13267 ( .A1(n15069), .A2(n15068), .ZN(n19027) );
  NOR2_X1 U13268 ( .A1(n15303), .A2(n15112), .ZN(n15262) );
  INV_X1 U13269 ( .A(n15316), .ZN(n15296) );
  AOI21_X1 U13270 ( .B1(n14225), .B2(n17998), .A(n14144), .ZN(n14145) );
  NAND2_X1 U13271 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n12407), .ZN(
        n12406) );
  AND2_X1 U13272 ( .A1(n15533), .A2(n15532), .ZN(n19061) );
  AND2_X1 U13273 ( .A1(n17987), .A2(n14142), .ZN(n18002) );
  OAI211_X1 U13274 ( .C1(n14328), .C2(n14334), .A(n14333), .B(n11754), .ZN(
        n14335) );
  AND2_X1 U13275 ( .A1(n19253), .A2(n14293), .ZN(n17616) );
  INV_X1 U13276 ( .A(n18007), .ZN(n19265) );
  INV_X1 U13277 ( .A(n19285), .ZN(n19329) );
  OR2_X1 U13278 ( .A1(n14215), .A2(n14203), .ZN(n17756) );
  XNOR2_X1 U13279 ( .A(n15058), .B(n15059), .ZN(n19982) );
  NAND2_X1 U13280 ( .A1(n15060), .A2(n15064), .ZN(n20200) );
  OAI21_X1 U13281 ( .B1(n17792), .B2(n17796), .A(n17791), .ZN(n20433) );
  NOR2_X2 U13282 ( .A1(n19899), .A2(n20006), .ZN(n20432) );
  INV_X1 U13283 ( .A(n20404), .ZN(n20297) );
  OAI21_X1 U13284 ( .B1(n19976), .B2(n19973), .A(n19972), .ZN(n20399) );
  INV_X1 U13285 ( .A(n19899), .ZN(n19950) );
  INV_X1 U13286 ( .A(n19843), .ZN(n19936) );
  INV_X1 U13287 ( .A(n19952), .ZN(n19951) );
  OAI21_X1 U13288 ( .B1(n19907), .B2(n19911), .A(n19906), .ZN(n20359) );
  OAI21_X1 U13289 ( .B1(n19895), .B2(n19894), .A(n19893), .ZN(n20352) );
  AND2_X1 U13290 ( .A1(n19882), .A2(n19924), .ZN(n20351) );
  INV_X1 U13291 ( .A(n19869), .ZN(n20272) );
  AND2_X1 U13292 ( .A1(n19844), .A2(n19950), .ZN(n20339) );
  OAI21_X1 U13293 ( .B1(n19855), .B2(n19863), .A(n19854), .ZN(n20332) );
  INV_X1 U13294 ( .A(n20242), .ZN(n20245) );
  NOR2_X2 U13295 ( .A1(n16353), .A2(n15057), .ZN(n20264) );
  INV_X1 U13296 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n17901) );
  INV_X1 U13297 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n22307) );
  INV_X1 U13298 ( .A(n21919), .ZN(n18494) );
  NOR2_X1 U13299 ( .A1(n21238), .A2(n21239), .ZN(n21259) );
  NOR2_X1 U13300 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n21137), .ZN(n21162) );
  NOR2_X1 U13301 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n21084), .ZN(n21100) );
  NOR2_X1 U13302 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n21032), .ZN(n21044) );
  INV_X1 U13303 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21808) );
  NOR2_X1 U13304 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20916), .ZN(n20936) );
  INV_X1 U13305 ( .A(n21268), .ZN(n21253) );
  NOR2_X2 U13306 ( .A1(n21193), .A2(n21937), .ZN(n21254) );
  AND2_X1 U13307 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18377), .ZN(n18407) );
  NAND2_X1 U13308 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18485), .ZN(n18447) );
  NAND3_X1 U13309 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18489), .A3(n18111), .ZN(
        n18150) );
  NOR2_X1 U13310 ( .A1(n20842), .A2(n20790), .ZN(n20808) );
  NOR2_X1 U13311 ( .A1(n21893), .A2(n21281), .ZN(n20826) );
  INV_X1 U13312 ( .A(n18503), .ZN(n18504) );
  OAI21_X1 U13313 ( .B1(n20857), .B2(n18693), .A(n19549), .ZN(n18655) );
  AND2_X1 U13314 ( .A1(n12707), .A2(n21843), .ZN(n21895) );
  NOR2_X1 U13315 ( .A1(n21612), .A2(n21611), .ZN(n21665) );
  INV_X1 U13316 ( .A(n21821), .ZN(n21856) );
  NOR3_X1 U13317 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n22278), .ZN(n18897) );
  INV_X1 U13318 ( .A(n21938), .ZN(n21505) );
  INV_X1 U13319 ( .A(n19774), .ZN(n19782) );
  INV_X1 U13320 ( .A(n19732), .ZN(n19745) );
  INV_X1 U13321 ( .A(n19712), .ZN(n19703) );
  INV_X1 U13322 ( .A(n19458), .ZN(n19461) );
  INV_X1 U13323 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20846) );
  INV_X1 U13324 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n22284) );
  NOR2_X1 U13325 ( .A1(n16374), .A2(n22265), .ZN(n22782) );
  INV_X1 U13326 ( .A(n22199), .ZN(n22237) );
  INV_X1 U13327 ( .A(n22215), .ZN(n22238) );
  NAND2_X1 U13328 ( .A1(n20621), .A2(n12842), .ZN(n16723) );
  INV_X1 U13329 ( .A(n20504), .ZN(n20526) );
  AND2_X1 U13330 ( .A1(n15136), .A2(n15123), .ZN(n15261) );
  INV_X1 U13331 ( .A(n20676), .ZN(n20703) );
  INV_X1 U13332 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20645) );
  INV_X1 U13333 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20640) );
  INV_X1 U13334 ( .A(n20689), .ZN(n20697) );
  INV_X1 U13335 ( .A(n22106), .ZN(n22115) );
  INV_X1 U13336 ( .A(n22118), .ZN(n22043) );
  INV_X1 U13337 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17899) );
  AOI22_X1 U13338 ( .A1(n22391), .A2(n22389), .B1(n22393), .B2(n22459), .ZN(
        n22705) );
  INV_X1 U13339 ( .A(n22714), .ZN(n22712) );
  AOI22_X1 U13340 ( .A1(n22407), .A2(n22412), .B1(n22459), .B2(n22433), .ZN(
        n22718) );
  AOI22_X1 U13341 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22424), .B1(n22427), 
        .B2(n22423), .ZN(n22725) );
  INV_X1 U13342 ( .A(n22720), .ZN(n16012) );
  INV_X1 U13343 ( .A(n15542), .ZN(n15604) );
  AOI22_X1 U13344 ( .A1(n22434), .A2(n22439), .B1(n22503), .B2(n22433), .ZN(
        n22732) );
  INV_X1 U13345 ( .A(n15613), .ZN(n15731) );
  NAND2_X1 U13346 ( .A1(n15841), .A2(n22380), .ZN(n22744) );
  AOI22_X1 U13347 ( .A1(n22460), .A2(n22466), .B1(n22459), .B2(n22458), .ZN(
        n22751) );
  AND2_X1 U13348 ( .A1(n15563), .A2(n15562), .ZN(n22581) );
  AOI22_X1 U13349 ( .A1(n22475), .A2(n22481), .B1(n22503), .B2(n22474), .ZN(
        n22759) );
  INV_X1 U13350 ( .A(n22772), .ZN(n22766) );
  NAND2_X1 U13351 ( .A1(n15913), .A2(n22405), .ZN(n22776) );
  NAND2_X1 U13352 ( .A1(n17865), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n22265) );
  INV_X1 U13353 ( .A(n22271), .ZN(n17860) );
  INV_X1 U13354 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n22302) );
  OR2_X1 U13355 ( .A1(n15631), .A2(n19350), .ZN(n19353) );
  NAND2_X1 U13356 ( .A1(n15107), .A2(n11991), .ZN(n19147) );
  INV_X1 U13357 ( .A(n19140), .ZN(n19222) );
  INV_X1 U13358 ( .A(n17544), .ZN(n17193) );
  AND2_X2 U13359 ( .A1(n14650), .A2(n19341), .ZN(n17281) );
  OR2_X1 U13360 ( .A1(n14651), .A2(n19835), .ZN(n17272) );
  INV_X1 U13361 ( .A(n20313), .ZN(n20153) );
  INV_X1 U13362 ( .A(n16084), .ZN(n20257) );
  NAND2_X1 U13363 ( .A1(n18048), .A2(n15130), .ZN(n15420) );
  INV_X1 U13364 ( .A(n18048), .ZN(n18080) );
  OR2_X1 U13365 ( .A1(n15111), .A2(n11354), .ZN(n15316) );
  AND2_X1 U13366 ( .A1(n14343), .A2(n14342), .ZN(n14344) );
  OR2_X1 U13367 ( .A1(n19353), .A2(n14120), .ZN(n18008) );
  INV_X1 U13368 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17988) );
  INV_X1 U13369 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17958) );
  INV_X1 U13370 ( .A(n18010), .ZN(n17996) );
  NAND2_X1 U13371 ( .A1(n14176), .A2(n12005), .ZN(n19304) );
  INV_X1 U13372 ( .A(n17760), .ZN(n19338) );
  INV_X1 U13373 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17821) );
  AOI22_X1 U13374 ( .A1(n17797), .A2(n17796), .B1(n17795), .B2(n17794), .ZN(
        n20438) );
  INV_X1 U13375 ( .A(n20414), .ZN(n20425) );
  AOI211_X2 U13376 ( .C1(n16026), .C2(n19846), .A(n20259), .B(n16025), .ZN(
        n20419) );
  NAND2_X1 U13377 ( .A1(n19963), .A2(n19962), .ZN(n20404) );
  NAND2_X1 U13378 ( .A1(n19951), .A2(n19950), .ZN(n20396) );
  NAND2_X1 U13379 ( .A1(n19951), .A2(n19936), .ZN(n20393) );
  NAND2_X1 U13380 ( .A1(n19951), .A2(n19924), .ZN(n20382) );
  INV_X1 U13381 ( .A(n20373), .ZN(n20370) );
  INV_X1 U13382 ( .A(n20365), .ZN(n20363) );
  INV_X1 U13383 ( .A(n20358), .ZN(n20356) );
  AND2_X1 U13384 ( .A1(n19890), .A2(n19889), .ZN(n20175) );
  INV_X1 U13385 ( .A(n20351), .ZN(n20280) );
  INV_X1 U13386 ( .A(n20172), .ZN(n20349) );
  INV_X1 U13387 ( .A(n20339), .ZN(n20215) );
  INV_X1 U13388 ( .A(n20331), .ZN(n20343) );
  INV_X1 U13389 ( .A(n20210), .ZN(n20336) );
  AOI21_X1 U13390 ( .B1(n21282), .B2(n21894), .A(n20789), .ZN(n17836) );
  INV_X1 U13391 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n22278) );
  INV_X1 U13392 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21123) );
  INV_X1 U13393 ( .A(n21934), .ZN(n21179) );
  INV_X1 U13394 ( .A(n21254), .ZN(n21228) );
  AND2_X1 U13395 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18397), .ZN(n18391) );
  NOR2_X1 U13396 ( .A1(n21161), .A2(n18401), .ZN(n18406) );
  NOR2_X1 U13397 ( .A1(n21043), .A2(n18152), .ZN(n18165) );
  INV_X1 U13398 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18298) );
  AND2_X1 U13399 ( .A1(n18489), .A2(n21371), .ZN(n18491) );
  NOR2_X1 U13400 ( .A1(n21283), .A2(n21301), .ZN(n21305) );
  NOR2_X1 U13401 ( .A1(n12462), .A2(n12461), .ZN(n21317) );
  NAND2_X1 U13402 ( .A1(n21456), .A2(n21459), .ZN(n21450) );
  INV_X1 U13403 ( .A(n18940), .ZN(n18939) );
  INV_X1 U13404 ( .A(n18802), .ZN(n18765) );
  INV_X1 U13405 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21853) );
  OAI21_X2 U13406 ( .B1(n16302), .B2(n12684), .A(n21926), .ZN(n21821) );
  NAND2_X1 U13407 ( .A1(n21868), .A2(n21821), .ZN(n21773) );
  INV_X1 U13408 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17832) );
  INV_X1 U13409 ( .A(n19794), .ZN(n19806) );
  INV_X1 U13410 ( .A(n19771), .ZN(n19762) );
  INV_X1 U13411 ( .A(n19452), .ZN(n19468) );
  INV_X1 U13412 ( .A(n22281), .ZN(n17828) );
  NOR2_X1 U13413 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n15092), .ZN(n19713)
         );
  INV_X1 U13414 ( .A(n20500), .ZN(n20489) );
  OR4_X1 U13415 ( .A1(n15105), .A2(n15104), .A3(n15103), .A4(n15102), .ZN(
        P2_U2838) );
  NAND2_X1 U13416 ( .A1(n11217), .A2(n11741), .ZN(P2_U3026) );
  NAND2_X1 U13417 ( .A1(n12756), .A2(n12755), .ZN(P3_U2831) );
  INV_X1 U13418 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U13419 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U13420 ( .A1(n11968), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U13421 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11765) );
  AND2_X2 U13422 ( .A1(n11763), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15678) );
  AND3_X2 U13423 ( .A1(n11763), .A2(n11762), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U13424 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14630), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U13425 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U13426 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14630), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U13427 ( .A1(n11968), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U13428 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11769) );
  NAND4_X1 U13429 ( .A1(n11743), .A2(n11771), .A3(n11770), .A4(n11769), .ZN(
        n11772) );
  AOI22_X1 U13430 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U13431 ( .A1(n11169), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14636), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U13432 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U13433 ( .A1(n11968), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U13434 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U13435 ( .A1(n11968), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U13436 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U13437 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14630), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11780) );
  NAND4_X1 U13438 ( .A1(n11783), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(
        n11784) );
  NAND2_X4 U13439 ( .A1(n11785), .A2(n11784), .ZN(n14120) );
  CLKBUF_X3 U13440 ( .A(n11960), .Z(n14626) );
  AND2_X2 U13441 ( .A1(n14626), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14445) );
  AND2_X2 U13442 ( .A1(n14616), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14446) );
  AOI22_X1 U13443 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11790) );
  BUF_X4 U13444 ( .A(n11968), .Z(n14625) );
  AND2_X2 U13445 ( .A1(n14625), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14451) );
  AOI22_X1 U13446 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11789) );
  AND2_X2 U13447 ( .A1(n11975), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14414) );
  AND2_X2 U13448 ( .A1(n14627), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14456) );
  AOI22_X1 U13449 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11788) );
  INV_X1 U13450 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20248) );
  AOI22_X1 U13451 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n14480), .B1(
        n14460), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11787) );
  NAND4_X1 U13452 ( .A1(n11790), .A2(n11789), .A3(n11788), .A4(n11787), .ZN(
        n11798) );
  AOI22_X1 U13453 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14485), .B1(
        n11174), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11796) );
  AND2_X2 U13454 ( .A1(n14630), .A2(n11936), .ZN(n14486) );
  AOI22_X1 U13455 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11795) );
  AND2_X2 U13456 ( .A1(n15678), .A2(n14497), .ZN(n14488) );
  NOR2_X1 U13457 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U13459 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11794) );
  AND2_X2 U13460 ( .A1(n15677), .A2(n14497), .ZN(n14490) );
  AOI22_X1 U13462 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11793) );
  NAND4_X1 U13463 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n11793), .ZN(
        n11797) );
  NAND2_X1 U13464 ( .A1(n12005), .A2(n13865), .ZN(n11801) );
  MUX2_X1 U13465 ( .A(n12216), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11910) );
  NAND2_X1 U13466 ( .A1(n20000), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13912) );
  INV_X1 U13467 ( .A(n13912), .ZN(n11911) );
  NAND2_X1 U13468 ( .A1(n11910), .A2(n11911), .ZN(n11800) );
  NAND2_X1 U13469 ( .A1(n12216), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11799) );
  NAND2_X1 U13470 ( .A1(n11800), .A2(n11799), .ZN(n11839) );
  XNOR2_X1 U13471 ( .A(n15673), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11837) );
  XNOR2_X1 U13472 ( .A(n11839), .B(n11837), .ZN(n14119) );
  NAND2_X1 U13473 ( .A1(n12003), .A2(n14119), .ZN(n14129) );
  NAND2_X1 U13474 ( .A1(n11801), .A2(n14129), .ZN(n14077) );
  AOI22_X1 U13475 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14636), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U13476 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11804) );
  NAND2_X1 U13477 ( .A1(n11806), .A2(n11936), .ZN(n11813) );
  AOI22_X1 U13478 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U13479 ( .A1(n11968), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U13480 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U13481 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14636), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11808) );
  NAND4_X1 U13482 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(
        n11812) );
  INV_X1 U13483 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12028) );
  AND2_X1 U13484 ( .A1(n11720), .A2(n12028), .ZN(n13914) );
  INV_X1 U13485 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n11814) );
  NAND2_X1 U13486 ( .A1(n13914), .A2(n11814), .ZN(n11826) );
  AOI22_X1 U13487 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U13488 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11817) );
  AOI22_X1 U13489 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11816) );
  INV_X1 U13490 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20312) );
  AOI22_X1 U13491 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14480), .B1(
        n14460), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11815) );
  NAND4_X1 U13492 ( .A1(n11818), .A2(n11817), .A3(n11816), .A4(n11815), .ZN(
        n11825) );
  AOI22_X1 U13493 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14485), .B1(
        n11174), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U13494 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U13495 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U13496 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11820) );
  NAND4_X1 U13497 ( .A1(n11823), .A2(n11822), .A3(n11821), .A4(n11820), .ZN(
        n11824) );
  NAND2_X1 U13498 ( .A1(n13915), .A2(n14093), .ZN(n12219) );
  NAND2_X1 U13499 ( .A1(n11826), .A2(n12219), .ZN(n13905) );
  AOI22_X1 U13500 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n14445), .B1(
        n14414), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U13501 ( .A1(n14451), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U13502 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n14479), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U13503 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14480), .B1(
        n11174), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11827) );
  NAND4_X1 U13504 ( .A1(n11830), .A2(n11829), .A3(n11828), .A4(n11827), .ZN(
        n11836) );
  AOI22_X1 U13505 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n14460), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U13506 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U13507 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n14490), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U13508 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n14488), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11831) );
  NAND4_X1 U13509 ( .A1(n11834), .A2(n11833), .A3(n11832), .A4(n11831), .ZN(
        n11835) );
  INV_X1 U13510 ( .A(n11837), .ZN(n11838) );
  NAND2_X1 U13511 ( .A1(n11839), .A2(n11838), .ZN(n11841) );
  NAND2_X1 U13512 ( .A1(n19884), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11840) );
  XNOR2_X1 U13513 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11857) );
  INV_X1 U13514 ( .A(n11857), .ZN(n11842) );
  XNOR2_X1 U13515 ( .A(n11858), .B(n11842), .ZN(n11908) );
  MUX2_X1 U13516 ( .A(n13894), .B(n11908), .S(n12003), .Z(n14081) );
  INV_X1 U13517 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11844) );
  MUX2_X1 U13518 ( .A(n14081), .B(n11844), .S(n11843), .Z(n13903) );
  AOI22_X1 U13519 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U13520 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U13521 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U13522 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11846) );
  NAND4_X1 U13523 ( .A1(n11849), .A2(n11848), .A3(n11847), .A4(n11846), .ZN(
        n11855) );
  AOI22_X1 U13524 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n14485), .B1(
        n11174), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U13525 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U13526 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U13527 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11850) );
  NAND4_X1 U13528 ( .A1(n11853), .A2(n11852), .A3(n11851), .A4(n11850), .ZN(
        n11854) );
  NOR2_X1 U13529 ( .A1(n11936), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11856) );
  NOR2_X1 U13530 ( .A1(n17845), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11859) );
  NAND2_X1 U13531 ( .A1(n11913), .A2(n11859), .ZN(n11909) );
  MUX2_X1 U13532 ( .A(n14089), .B(n11909), .S(n12003), .Z(n14080) );
  INV_X1 U13533 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11860) );
  MUX2_X1 U13534 ( .A(n14080), .B(n11860), .S(n11843), .Z(n13920) );
  AOI22_X1 U13535 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U13536 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U13537 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11862) );
  INV_X1 U13538 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20108) );
  AOI22_X1 U13539 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n14480), .B1(
        n14460), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11861) );
  NAND4_X1 U13540 ( .A1(n11864), .A2(n11863), .A3(n11862), .A4(n11861), .ZN(
        n11870) );
  AOI22_X1 U13541 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n14485), .B1(
        n11174), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U13542 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U13543 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U13544 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11865) );
  NAND4_X1 U13545 ( .A1(n11868), .A2(n11867), .A3(n11866), .A4(n11865), .ZN(
        n11869) );
  NOR2_X1 U13546 ( .A1(n11870), .A2(n11869), .ZN(n13956) );
  MUX2_X1 U13547 ( .A(n13956), .B(P2_EBX_REG_5__SCAN_IN), .S(n11843), .Z(
        n13959) );
  INV_X1 U13548 ( .A(n13959), .ZN(n11871) );
  INV_X1 U13549 ( .A(n13991), .ZN(n11883) );
  AOI22_X1 U13550 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U13551 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U13552 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U13553 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n14485), .B1(
        n11174), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11872) );
  NAND4_X1 U13554 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n11881) );
  AOI22_X1 U13555 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U13556 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U13557 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14490), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U13558 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14488), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11876) );
  NAND4_X1 U13559 ( .A1(n11879), .A2(n11878), .A3(n11877), .A4(n11876), .ZN(
        n11880) );
  MUX2_X1 U13560 ( .A(n13983), .B(P2_EBX_REG_6__SCAN_IN), .S(n11843), .Z(
        n13990) );
  INV_X1 U13561 ( .A(n13990), .ZN(n11882) );
  NAND2_X1 U13562 ( .A1(n11883), .A2(n11882), .ZN(n13996) );
  NAND2_X1 U13563 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11887) );
  NAND2_X1 U13564 ( .A1(n14479), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11886) );
  NAND2_X1 U13565 ( .A1(n14456), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11885) );
  NAND2_X1 U13566 ( .A1(n14446), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11884) );
  AOI22_X1 U13567 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U13568 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11890) );
  NAND2_X1 U13569 ( .A1(n11819), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11889) );
  NAND2_X1 U13570 ( .A1(n14486), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11888) );
  NAND2_X1 U13571 ( .A1(n14445), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11895) );
  NAND2_X1 U13572 ( .A1(n14451), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11894) );
  NAND2_X1 U13573 ( .A1(n14480), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11893) );
  NAND2_X1 U13574 ( .A1(n14485), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11892) );
  AOI22_X1 U13575 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n14460), .B1(
        n11174), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11896) );
  NAND4_X1 U13576 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n13902) );
  MUX2_X1 U13577 ( .A(n14324), .B(P2_EBX_REG_7__SCAN_IN), .S(n11843), .Z(
        n13995) );
  NAND2_X1 U13578 ( .A1(n11843), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n14002) );
  NAND2_X1 U13579 ( .A1(n11843), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14004) );
  NAND2_X1 U13580 ( .A1(n11900), .A2(n14004), .ZN(n14009) );
  INV_X1 U13581 ( .A(n14009), .ZN(n11902) );
  NAND2_X1 U13582 ( .A1(n11843), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14017) );
  INV_X1 U13583 ( .A(n14017), .ZN(n11903) );
  NAND2_X1 U13584 ( .A1(n11843), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n14021) );
  INV_X1 U13585 ( .A(n14021), .ZN(n11904) );
  NAND2_X1 U13586 ( .A1(n11843), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14028) );
  NAND2_X1 U13587 ( .A1(n11843), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n14038) );
  AND2_X1 U13588 ( .A1(n11843), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14044) );
  NAND2_X1 U13589 ( .A1(n11843), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14047) );
  AND2_X1 U13590 ( .A1(n11843), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14054) );
  NAND2_X1 U13591 ( .A1(n11843), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14064) );
  AND2_X1 U13592 ( .A1(n11843), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14241) );
  NAND2_X1 U13593 ( .A1(n11843), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14248) );
  INV_X1 U13594 ( .A(n14248), .ZN(n11905) );
  NAND2_X1 U13595 ( .A1(n11843), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n14252) );
  AND2_X1 U13596 ( .A1(n11843), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n14260) );
  NAND2_X1 U13597 ( .A1(n11843), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14257) );
  INV_X1 U13598 ( .A(n14257), .ZN(n11906) );
  NAND2_X1 U13599 ( .A1(n11843), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14266) );
  AND2_X1 U13600 ( .A1(n11843), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14270) );
  NAND2_X1 U13601 ( .A1(n11843), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14320) );
  NAND2_X1 U13602 ( .A1(n14321), .A2(n14320), .ZN(n17074) );
  AND2_X1 U13603 ( .A1(n11843), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11907) );
  XNOR2_X1 U13604 ( .A(n17074), .B(n11907), .ZN(n14325) );
  INV_X1 U13605 ( .A(n14325), .ZN(n14327) );
  NAND2_X1 U13606 ( .A1(n11909), .A2(n11908), .ZN(n14131) );
  INV_X1 U13607 ( .A(n14119), .ZN(n14127) );
  OR2_X1 U13608 ( .A1(n14131), .A2(n14127), .ZN(n14074) );
  INV_X1 U13609 ( .A(n11910), .ZN(n14124) );
  XNOR2_X1 U13610 ( .A(n14124), .B(n11911), .ZN(n14121) );
  INV_X1 U13611 ( .A(n14121), .ZN(n11916) );
  NAND2_X1 U13612 ( .A1(n17845), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11912) );
  NAND2_X1 U13613 ( .A1(n11913), .A2(n11912), .ZN(n11915) );
  NAND2_X1 U13614 ( .A1(n17821), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11914) );
  INV_X2 U13615 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n12085) );
  NAND2_X1 U13616 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12085), .ZN(n15706) );
  INV_X1 U13617 ( .A(n15706), .ZN(n11917) );
  INV_X1 U13618 ( .A(n19341), .ZN(n19350) );
  OR2_X1 U13619 ( .A1(n15699), .A2(n19350), .ZN(n11987) );
  AOI22_X1 U13620 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11921) );
  AOI22_X1 U13621 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14630), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11920) );
  AOI22_X1 U13622 ( .A1(n11968), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U13623 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11918) );
  NAND4_X1 U13624 ( .A1(n11921), .A2(n11920), .A3(n11919), .A4(n11918), .ZN(
        n11922) );
  NAND2_X1 U13625 ( .A1(n11922), .A2(n11936), .ZN(n11930) );
  AOI22_X1 U13626 ( .A1(n11968), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U13627 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U13628 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14636), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11924) );
  NAND4_X1 U13629 ( .A1(n11927), .A2(n11926), .A3(n11925), .A4(n11924), .ZN(
        n11928) );
  NAND2_X1 U13630 ( .A1(n11928), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11929) );
  NAND2_X2 U13631 ( .A1(n11930), .A2(n11929), .ZN(n12006) );
  AOI22_X1 U13632 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14630), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U13633 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U13634 ( .A1(n11968), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11931) );
  NAND4_X1 U13635 ( .A1(n11934), .A2(n11933), .A3(n11932), .A4(n11931), .ZN(
        n11935) );
  AOI22_X1 U13636 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14636), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U13637 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U13638 ( .A1(n11968), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U13639 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U13640 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14630), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U13641 ( .A1(n11968), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U13642 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U13643 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11945) );
  NAND2_X1 U13644 ( .A1(n11946), .A2(n11945), .ZN(n11953) );
  AOI22_X1 U13645 ( .A1(n11968), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U13646 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14630), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U13647 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U13648 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11948) );
  NAND4_X1 U13649 ( .A1(n11951), .A2(n11950), .A3(n11949), .A4(n11948), .ZN(
        n11952) );
  NAND2_X1 U13650 ( .A1(n11997), .A2(n11983), .ZN(n11954) );
  AOI22_X1 U13651 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11969), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U13652 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14636), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U13653 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11956) );
  NAND4_X1 U13654 ( .A1(n11958), .A2(n11957), .A3(n11956), .A4(n11955), .ZN(
        n11959) );
  AOI22_X1 U13655 ( .A1(n11969), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U13656 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U13657 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14636), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U13658 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11968), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11961) );
  NAND4_X1 U13659 ( .A1(n11964), .A2(n11963), .A3(n11962), .A4(n11961), .ZN(
        n11965) );
  NAND2_X1 U13660 ( .A1(n12014), .A2(n16031), .ZN(n11966) );
  NAND2_X1 U13661 ( .A1(n11967), .A2(n11966), .ZN(n12016) );
  INV_X1 U13662 ( .A(n12016), .ZN(n11985) );
  AOI22_X1 U13663 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14627), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U13664 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14636), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U13665 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14616), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U13666 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11970) );
  NAND4_X1 U13667 ( .A1(n11973), .A2(n11972), .A3(n11971), .A4(n11970), .ZN(
        n11974) );
  AOI22_X1 U13668 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14636), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U13669 ( .A1(n11937), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11977) );
  AND2_X1 U13670 ( .A1(n11978), .A2(n11977), .ZN(n11981) );
  AOI22_X1 U13671 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14627), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U13672 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14616), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11979) );
  NAND3_X1 U13673 ( .A1(n11981), .A2(n11980), .A3(n11979), .ZN(n11982) );
  AND4_X1 U13674 ( .A1(n11983), .A2(n12006), .A3(n13915), .A4(n14146), .ZN(
        n11984) );
  INV_X1 U13675 ( .A(n12018), .ZN(n11986) );
  OR2_X1 U13676 ( .A1(n11987), .A2(n15634), .ZN(n16065) );
  NAND2_X1 U13677 ( .A1(n14353), .A2(n12009), .ZN(n12010) );
  INV_X1 U13678 ( .A(n12010), .ZN(n11988) );
  NOR2_X1 U13679 ( .A1(n15706), .A2(n15699), .ZN(n11989) );
  NAND2_X1 U13680 ( .A1(n12002), .A2(n11989), .ZN(n15111) );
  NAND2_X1 U13681 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19342) );
  INV_X1 U13682 ( .A(n19342), .ZN(n22317) );
  NOR2_X1 U13683 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n22317), .ZN(n12431) );
  INV_X1 U13684 ( .A(n12431), .ZN(n11992) );
  NAND2_X1 U13685 ( .A1(n11992), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11990) );
  NOR2_X1 U13686 ( .A1(n12003), .A2(n11990), .ZN(n11991) );
  NOR2_X1 U13687 ( .A1(n12003), .A2(n11992), .ZN(n11993) );
  NAND2_X1 U13688 ( .A1(n14212), .A2(n12004), .ZN(n12033) );
  INV_X1 U13689 ( .A(n11996), .ZN(n11998) );
  NAND2_X1 U13690 ( .A1(n15157), .A2(n15161), .ZN(n12039) );
  NAND3_X1 U13691 ( .A1(n12033), .A2(n12038), .A3(n12039), .ZN(n11999) );
  NAND2_X1 U13692 ( .A1(n11999), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12001) );
  NAND2_X1 U13693 ( .A1(n12002), .A2(n20262), .ZN(n12000) );
  NAND2_X2 U13694 ( .A1(n12001), .A2(n12000), .ZN(n12071) );
  INV_X2 U13695 ( .A(n17084), .ZN(n12175) );
  INV_X1 U13696 ( .A(n12003), .ZN(n12005) );
  AOI22_X1 U13697 ( .A1(n12066), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12007) );
  OAI21_X1 U13698 ( .B1(n12069), .B2(n19302), .A(n12007), .ZN(n12008) );
  AOI21_X1 U13699 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n12175), .A(
        n12008), .ZN(n15497) );
  INV_X1 U13700 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19224) );
  NAND2_X1 U13701 ( .A1(n12071), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12032) );
  NAND2_X1 U13702 ( .A1(n14156), .A2(n20112), .ZN(n14157) );
  NAND2_X1 U13703 ( .A1(n12014), .A2(n14149), .ZN(n14160) );
  NAND2_X1 U13704 ( .A1(n14190), .A2(n16031), .ZN(n12013) );
  NAND2_X1 U13705 ( .A1(n12013), .A2(n12012), .ZN(n12015) );
  NAND3_X1 U13706 ( .A1(n14195), .A2(n20262), .A3(n12014), .ZN(n15156) );
  NAND2_X1 U13707 ( .A1(n12015), .A2(n15156), .ZN(n12024) );
  NAND2_X1 U13708 ( .A1(n12017), .A2(n20207), .ZN(n12019) );
  OAI211_X1 U13709 ( .C1(n12016), .C2(n12019), .A(n12018), .B(n14154), .ZN(
        n14199) );
  INV_X1 U13710 ( .A(n12017), .ZN(n12020) );
  NAND2_X1 U13711 ( .A1(n12021), .A2(n12020), .ZN(n14085) );
  AND2_X1 U13712 ( .A1(n20207), .A2(n11354), .ZN(n12022) );
  NAND2_X1 U13713 ( .A1(n14085), .A2(n12022), .ZN(n14211) );
  NAND3_X1 U13714 ( .A1(n14211), .A2(n11156), .A3(n15707), .ZN(n12023) );
  NAND3_X1 U13715 ( .A1(n12024), .A2(n14199), .A3(n12023), .ZN(n12025) );
  INV_X1 U13717 ( .A(n12063), .ZN(n12031) );
  NAND2_X1 U13718 ( .A1(n17901), .A2(n12085), .ZN(n12040) );
  AOI21_X1 U13719 ( .B1(n12183), .B2(P2_REIP_REG_0__SCAN_IN), .A(n12029), .ZN(
        n12030) );
  NAND2_X1 U13720 ( .A1(n12063), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12037) );
  OAI21_X1 U13722 ( .B1(n12040), .B2(n20000), .A(n12051), .ZN(n12035) );
  AOI21_X1 U13723 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n15644), .A(n12035), 
        .ZN(n12036) );
  NAND2_X1 U13724 ( .A1(n12037), .A2(n12036), .ZN(n13809) );
  NAND2_X1 U13725 ( .A1(n12063), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12043) );
  INV_X1 U13726 ( .A(n15707), .ZN(n14164) );
  NAND2_X1 U13727 ( .A1(n14180), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12042) );
  NAND2_X1 U13728 ( .A1(n12026), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12041) );
  INV_X1 U13729 ( .A(n12183), .ZN(n12055) );
  INV_X1 U13730 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n17185) );
  NAND2_X1 U13731 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12044) );
  OAI211_X1 U13732 ( .C1(n12055), .C2(n17185), .A(n12045), .B(n12044), .ZN(
        n12046) );
  NAND2_X1 U13733 ( .A1(n13808), .A2(n13814), .ZN(n12047) );
  INV_X1 U13734 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n12054) );
  INV_X1 U13735 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12049) );
  INV_X1 U13736 ( .A(n12052), .ZN(n12053) );
  OAI21_X1 U13737 ( .B1(n12055), .B2(n12054), .A(n12053), .ZN(n12056) );
  AOI21_X1 U13738 ( .B1(n17901), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12057) );
  INV_X1 U13739 ( .A(n12059), .ZN(n12061) );
  NAND2_X1 U13740 ( .A1(n12061), .A2(n12060), .ZN(n12062) );
  NAND2_X1 U13741 ( .A1(n12063), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12065) );
  NAND2_X1 U13742 ( .A1(n12026), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12064) );
  NAND2_X1 U13743 ( .A1(n12065), .A2(n12064), .ZN(n12072) );
  INV_X1 U13744 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19326) );
  INV_X1 U13745 ( .A(n12051), .ZN(n12066) );
  NAND2_X1 U13746 ( .A1(n12066), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n12068) );
  NAND2_X1 U13747 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12067) );
  OAI211_X1 U13748 ( .C1(n12069), .C2(n19326), .A(n12068), .B(n12067), .ZN(
        n12070) );
  INV_X1 U13749 ( .A(n12072), .ZN(n12073) );
  INV_X1 U13750 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U13751 ( .A1(n12066), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12075) );
  OAI21_X1 U13752 ( .B1(n12069), .B2(n12076), .A(n12075), .ZN(n12077) );
  AOI21_X1 U13753 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n12175), .A(
        n12077), .ZN(n16093) );
  INV_X1 U13754 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16166) );
  AOI22_X1 U13755 ( .A1(n12066), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12080) );
  NAND2_X1 U13756 ( .A1(n12160), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12079) );
  OAI211_X1 U13757 ( .C1(n17084), .C2(n16166), .A(n12080), .B(n12079), .ZN(
        n16122) );
  NAND2_X1 U13758 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12084) );
  INV_X1 U13759 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12081) );
  INV_X1 U13760 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16143) );
  OAI22_X1 U13761 ( .A1(n12181), .A2(n12081), .B1(n12085), .B2(n16143), .ZN(
        n12082) );
  AOI21_X1 U13762 ( .B1(n12160), .B2(P2_REIP_REG_7__SCAN_IN), .A(n12082), .ZN(
        n12083) );
  NAND2_X1 U13763 ( .A1(n12084), .A2(n12083), .ZN(n15487) );
  NAND2_X1 U13764 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12090) );
  INV_X1 U13765 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12087) );
  INV_X1 U13766 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12086) );
  OAI22_X1 U13767 ( .A1(n12181), .A2(n12087), .B1(n12085), .B2(n12086), .ZN(
        n12088) );
  AOI21_X1 U13768 ( .B1(n12160), .B2(P2_REIP_REG_8__SCAN_IN), .A(n12088), .ZN(
        n12089) );
  NAND2_X1 U13769 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12094) );
  INV_X1 U13770 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12091) );
  OAI22_X1 U13771 ( .A1(n12181), .A2(n12091), .B1(n12085), .B2(n17958), .ZN(
        n12092) );
  AOI21_X1 U13772 ( .B1(n12160), .B2(P2_REIP_REG_9__SCAN_IN), .A(n12092), .ZN(
        n12093) );
  NAND2_X1 U13773 ( .A1(n12094), .A2(n12093), .ZN(n15779) );
  NAND2_X1 U13774 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12099) );
  INV_X1 U13775 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12096) );
  INV_X1 U13776 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12095) );
  OAI22_X1 U13777 ( .A1(n12181), .A2(n12096), .B1(n12085), .B2(n12095), .ZN(
        n12097) );
  AOI21_X1 U13778 ( .B1(n12160), .B2(P2_REIP_REG_10__SCAN_IN), .A(n12097), 
        .ZN(n12098) );
  NAND2_X1 U13779 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12104) );
  INV_X1 U13780 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12101) );
  INV_X1 U13781 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12100) );
  OAI22_X1 U13782 ( .A1(n12181), .A2(n12101), .B1(n12085), .B2(n12100), .ZN(
        n12102) );
  AOI21_X1 U13783 ( .B1(n12160), .B2(P2_REIP_REG_11__SCAN_IN), .A(n12102), 
        .ZN(n12103) );
  NAND2_X1 U13784 ( .A1(n12104), .A2(n12103), .ZN(n15884) );
  NAND2_X1 U13785 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12109) );
  INV_X1 U13786 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12106) );
  INV_X1 U13787 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12105) );
  OAI22_X1 U13788 ( .A1(n12181), .A2(n12106), .B1(n12085), .B2(n12105), .ZN(
        n12107) );
  AOI21_X1 U13789 ( .B1(n12160), .B2(P2_REIP_REG_12__SCAN_IN), .A(n12107), 
        .ZN(n12108) );
  NAND2_X1 U13790 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12113) );
  INV_X1 U13791 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12110) );
  OAI22_X1 U13792 ( .A1(n12181), .A2(n12110), .B1(n12085), .B2(n17988), .ZN(
        n12111) );
  AOI21_X1 U13793 ( .B1(n12160), .B2(P2_REIP_REG_13__SCAN_IN), .A(n12111), 
        .ZN(n12112) );
  NAND2_X1 U13794 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12118) );
  INV_X1 U13795 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12115) );
  INV_X1 U13796 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12114) );
  OAI22_X1 U13797 ( .A1(n12181), .A2(n12115), .B1(n12085), .B2(n12114), .ZN(
        n12116) );
  AOI21_X1 U13798 ( .B1(n12160), .B2(P2_REIP_REG_14__SCAN_IN), .A(n12116), 
        .ZN(n12117) );
  NAND2_X1 U13799 ( .A1(n12118), .A2(n12117), .ZN(n16237) );
  NAND2_X1 U13800 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12122) );
  INV_X1 U13801 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12119) );
  OAI22_X1 U13802 ( .A1(n12181), .A2(n12119), .B1(n12085), .B2(n17523), .ZN(
        n12120) );
  AOI21_X1 U13803 ( .B1(n12160), .B2(P2_REIP_REG_15__SCAN_IN), .A(n12120), 
        .ZN(n12121) );
  NAND2_X1 U13804 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12127) );
  INV_X1 U13805 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12124) );
  INV_X1 U13806 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12123) );
  OAI22_X1 U13807 ( .A1(n12181), .A2(n12124), .B1(n12085), .B2(n12123), .ZN(
        n12125) );
  AOI21_X1 U13808 ( .B1(n12160), .B2(P2_REIP_REG_16__SCAN_IN), .A(n12125), 
        .ZN(n12126) );
  NAND2_X1 U13809 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12131) );
  INV_X1 U13810 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12128) );
  INV_X1 U13811 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17511) );
  OAI22_X1 U13812 ( .A1(n12181), .A2(n12128), .B1(n12085), .B2(n17511), .ZN(
        n12129) );
  AOI21_X1 U13813 ( .B1(n12160), .B2(P2_REIP_REG_17__SCAN_IN), .A(n12129), 
        .ZN(n12130) );
  NAND2_X1 U13814 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12135) );
  INV_X1 U13815 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n12132) );
  INV_X1 U13816 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17495) );
  OAI22_X1 U13817 ( .A1(n12181), .A2(n12132), .B1(n12085), .B2(n17495), .ZN(
        n12133) );
  AOI21_X1 U13818 ( .B1(n12160), .B2(P2_REIP_REG_18__SCAN_IN), .A(n12133), 
        .ZN(n12134) );
  NAND2_X1 U13819 ( .A1(n12135), .A2(n12134), .ZN(n17263) );
  NAND2_X1 U13820 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12139) );
  INV_X1 U13821 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12136) );
  INV_X1 U13822 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17489) );
  OAI22_X1 U13823 ( .A1(n12181), .A2(n12136), .B1(n12085), .B2(n17489), .ZN(
        n12137) );
  AOI21_X1 U13824 ( .B1(n12160), .B2(P2_REIP_REG_19__SCAN_IN), .A(n12137), 
        .ZN(n12138) );
  NAND2_X1 U13825 ( .A1(n12139), .A2(n12138), .ZN(n17256) );
  NAND2_X1 U13826 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12143) );
  INV_X1 U13827 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n19149) );
  INV_X1 U13828 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12140) );
  OAI22_X1 U13829 ( .A1(n12181), .A2(n19149), .B1(n12085), .B2(n12140), .ZN(
        n12141) );
  AOI21_X1 U13830 ( .B1(n12160), .B2(P2_REIP_REG_20__SCAN_IN), .A(n12141), 
        .ZN(n12142) );
  NAND2_X1 U13831 ( .A1(n12143), .A2(n12142), .ZN(n14118) );
  NAND2_X1 U13832 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12147) );
  INV_X1 U13833 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12144) );
  INV_X1 U13834 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17477) );
  OAI22_X1 U13835 ( .A1(n12181), .A2(n12144), .B1(n12085), .B2(n17477), .ZN(
        n12145) );
  AOI21_X1 U13836 ( .B1(n12160), .B2(P2_REIP_REG_21__SCAN_IN), .A(n12145), 
        .ZN(n12146) );
  NAND2_X1 U13837 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12151) );
  INV_X1 U13838 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n12148) );
  INV_X1 U13839 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12418) );
  OAI22_X1 U13840 ( .A1(n12181), .A2(n12148), .B1(n12085), .B2(n12418), .ZN(
        n12149) );
  AOI21_X1 U13841 ( .B1(n12160), .B2(P2_REIP_REG_22__SCAN_IN), .A(n12149), 
        .ZN(n12150) );
  NAND2_X1 U13842 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12154) );
  INV_X1 U13843 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n17140) );
  INV_X1 U13844 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17454) );
  OAI22_X1 U13845 ( .A1(n12181), .A2(n17140), .B1(n12085), .B2(n17454), .ZN(
        n12152) );
  AOI21_X1 U13846 ( .B1(n12160), .B2(P2_REIP_REG_23__SCAN_IN), .A(n12152), 
        .ZN(n12153) );
  NAND2_X1 U13847 ( .A1(n12154), .A2(n12153), .ZN(n17136) );
  NAND2_X1 U13848 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12157) );
  INV_X1 U13849 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n17128) );
  INV_X1 U13850 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17443) );
  OAI22_X1 U13851 ( .A1(n12181), .A2(n17128), .B1(n12085), .B2(n17443), .ZN(
        n12155) );
  AOI21_X1 U13852 ( .B1(n12160), .B2(P2_REIP_REG_24__SCAN_IN), .A(n12155), 
        .ZN(n12156) );
  NAND2_X1 U13853 ( .A1(n12157), .A2(n12156), .ZN(n17125) );
  NAND2_X1 U13854 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12162) );
  INV_X1 U13855 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n12158) );
  INV_X1 U13856 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n19183) );
  OAI22_X1 U13857 ( .A1(n12181), .A2(n12158), .B1(n12085), .B2(n19183), .ZN(
        n12159) );
  AOI21_X1 U13858 ( .B1(n12160), .B2(P2_REIP_REG_25__SCAN_IN), .A(n12159), 
        .ZN(n12161) );
  NAND2_X1 U13859 ( .A1(n12162), .A2(n12161), .ZN(n17227) );
  NAND2_X1 U13860 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12167) );
  INV_X1 U13861 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12164) );
  INV_X1 U13862 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12163) );
  OAI22_X1 U13863 ( .A1(n12181), .A2(n12164), .B1(n12085), .B2(n12163), .ZN(
        n12165) );
  AOI21_X1 U13864 ( .B1(n12160), .B2(P2_REIP_REG_26__SCAN_IN), .A(n12165), 
        .ZN(n12166) );
  AND2_X1 U13865 ( .A1(n12167), .A2(n12166), .ZN(n17221) );
  NAND2_X1 U13866 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12170) );
  INV_X1 U13867 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n17112) );
  INV_X1 U13868 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17111) );
  OAI22_X1 U13869 ( .A1(n12181), .A2(n17112), .B1(n12085), .B2(n17111), .ZN(
        n12168) );
  AOI21_X1 U13870 ( .B1(n12160), .B2(P2_REIP_REG_27__SCAN_IN), .A(n12168), 
        .ZN(n12169) );
  NAND2_X1 U13871 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12174) );
  INV_X1 U13872 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12171) );
  INV_X1 U13873 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17099) );
  OAI22_X1 U13874 ( .A1(n12181), .A2(n12171), .B1(n12085), .B2(n17099), .ZN(
        n12172) );
  AOI21_X1 U13875 ( .B1(n12160), .B2(P2_REIP_REG_28__SCAN_IN), .A(n12172), 
        .ZN(n12173) );
  NAND2_X1 U13876 ( .A1(n12174), .A2(n12173), .ZN(n14284) );
  NAND2_X1 U13877 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12179) );
  INV_X1 U13878 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12176) );
  INV_X1 U13879 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17415) );
  OAI22_X1 U13880 ( .A1(n12181), .A2(n12176), .B1(n12085), .B2(n17415), .ZN(
        n12177) );
  AOI21_X1 U13881 ( .B1(n12183), .B2(P2_REIP_REG_29__SCAN_IN), .A(n12177), 
        .ZN(n12178) );
  NAND2_X1 U13882 ( .A1(n12179), .A2(n12178), .ZN(n17198) );
  NAND2_X1 U13883 ( .A1(n17199), .A2(n17198), .ZN(n12188) );
  INV_X1 U13884 ( .A(n12188), .ZN(n12187) );
  NAND2_X1 U13885 ( .A1(n12175), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12185) );
  INV_X1 U13886 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12180) );
  INV_X1 U13887 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16319) );
  OAI22_X1 U13888 ( .A1(n12181), .A2(n12180), .B1(n12085), .B2(n16319), .ZN(
        n12182) );
  AOI21_X1 U13889 ( .B1(n12183), .B2(P2_REIP_REG_30__SCAN_IN), .A(n12182), 
        .ZN(n12184) );
  AND2_X1 U13890 ( .A1(n12185), .A2(n12184), .ZN(n12189) );
  INV_X1 U13891 ( .A(n12189), .ZN(n12186) );
  NAND2_X1 U13892 ( .A1(n12188), .A2(n12189), .ZN(n12190) );
  INV_X2 U13893 ( .A(n12351), .ZN(n12368) );
  INV_X2 U13894 ( .A(n12350), .ZN(n12367) );
  AOI22_X1 U13895 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12194) );
  NAND2_X1 U13896 ( .A1(n12321), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12193) );
  NAND2_X1 U13897 ( .A1(n12194), .A2(n12193), .ZN(n17375) );
  AOI22_X1 U13898 ( .A1(n12191), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n12192), .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12196) );
  NAND2_X1 U13899 ( .A1(n12321), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12195) );
  NAND2_X1 U13900 ( .A1(n19835), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12197) );
  OAI211_X1 U13901 ( .C1(n20262), .C2(n19224), .A(n12197), .B(n14346), .ZN(
        n12198) );
  INV_X1 U13902 ( .A(n12198), .ZN(n12199) );
  NAND2_X1 U13903 ( .A1(n12200), .A2(n12199), .ZN(n15148) );
  AOI22_X1 U13904 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U13905 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U13906 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12202) );
  INV_X1 U13907 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20437) );
  AOI22_X1 U13908 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n14480), .B1(
        n14460), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12201) );
  NAND4_X1 U13909 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12211) );
  AOI22_X1 U13910 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n14485), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U13911 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U13912 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U13913 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12206) );
  NAND4_X1 U13914 ( .A1(n12209), .A2(n12208), .A3(n12207), .A4(n12206), .ZN(
        n12210) );
  OR2_X2 U13915 ( .A1(n12211), .A2(n12210), .ZN(n14094) );
  INV_X1 U13916 ( .A(n14094), .ZN(n13913) );
  AND2_X1 U13917 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12212) );
  NOR2_X1 U13918 ( .A1(n12192), .A2(n12212), .ZN(n12213) );
  INV_X1 U13919 ( .A(n12014), .ZN(n15160) );
  NAND2_X1 U13920 ( .A1(n12191), .A2(n15160), .ZN(n12222) );
  OAI211_X1 U13921 ( .C1(n12334), .C2(n13913), .A(n12213), .B(n12222), .ZN(
        n15147) );
  NAND2_X1 U13922 ( .A1(n15148), .A2(n15147), .ZN(n15149) );
  NAND2_X1 U13923 ( .A1(n12214), .A2(n15149), .ZN(n12221) );
  XNOR2_X1 U13924 ( .A(n15149), .B(n12214), .ZN(n15202) );
  INV_X1 U13925 ( .A(n12215), .ZN(n12220) );
  NAND2_X1 U13926 ( .A1(n12014), .A2(n12006), .ZN(n12217) );
  MUX2_X1 U13927 ( .A(n12217), .B(n12216), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12218) );
  OAI21_X1 U13928 ( .B1(n12220), .B2(n12219), .A(n12218), .ZN(n15201) );
  OR2_X2 U13929 ( .A1(n15202), .A2(n15201), .ZN(n15204) );
  NAND2_X1 U13930 ( .A1(n12221), .A2(n15204), .ZN(n12227) );
  OAI21_X1 U13931 ( .B1(n14346), .B2(n19884), .A(n12222), .ZN(n12223) );
  AOI21_X1 U13932 ( .B1(n12346), .B2(n13865), .A(n12223), .ZN(n12228) );
  INV_X1 U13933 ( .A(n12228), .ZN(n12224) );
  XNOR2_X1 U13934 ( .A(n12227), .B(n12224), .ZN(n15215) );
  AOI22_X1 U13935 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12226) );
  NAND2_X1 U13936 ( .A1(n12321), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12225) );
  AND2_X1 U13937 ( .A1(n12226), .A2(n12225), .ZN(n15214) );
  NAND2_X1 U13938 ( .A1(n12228), .A2(n12227), .ZN(n12229) );
  NAND2_X1 U13939 ( .A1(n12346), .A2(n13894), .ZN(n12233) );
  AOI22_X1 U13940 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12232) );
  NAND2_X1 U13941 ( .A1(n12367), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12231) );
  NAND2_X1 U13942 ( .A1(n12321), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12230) );
  INV_X1 U13943 ( .A(n14089), .ZN(n12236) );
  AOI22_X1 U13944 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12235) );
  NAND2_X1 U13945 ( .A1(n12321), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12234) );
  OAI211_X1 U13946 ( .C1(n12236), .C2(n12334), .A(n12235), .B(n12234), .ZN(
        n16079) );
  INV_X1 U13947 ( .A(n16080), .ZN(n12239) );
  AOI22_X1 U13948 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12238) );
  NAND2_X1 U13949 ( .A1(n12321), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12237) );
  OAI211_X1 U13950 ( .C1(n13956), .C2(n12334), .A(n12238), .B(n12237), .ZN(
        n16123) );
  NAND2_X1 U13951 ( .A1(n12239), .A2(n16123), .ZN(n16124) );
  INV_X1 U13952 ( .A(n13983), .ZN(n12240) );
  NAND2_X1 U13953 ( .A1(n12346), .A2(n12240), .ZN(n12241) );
  NAND2_X1 U13954 ( .A1(n16124), .A2(n12241), .ZN(n15189) );
  AOI22_X1 U13955 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n12192), .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12243) );
  NAND2_X1 U13956 ( .A1(n12321), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12242) );
  NAND2_X1 U13957 ( .A1(n12243), .A2(n12242), .ZN(n15188) );
  NAND2_X1 U13958 ( .A1(n15189), .A2(n15188), .ZN(n15191) );
  NAND2_X1 U13959 ( .A1(n12346), .A2(n14067), .ZN(n12244) );
  AOI22_X1 U13960 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12246) );
  NAND2_X1 U13961 ( .A1(n12321), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U13962 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n14479), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U13963 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n14445), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U13964 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U13965 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n14485), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12247) );
  NAND4_X1 U13966 ( .A1(n12250), .A2(n12249), .A3(n12248), .A4(n12247), .ZN(
        n12256) );
  AOI22_X1 U13967 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n11174), .B1(
        n14460), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U13968 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U13969 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n14490), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U13970 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n14488), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12251) );
  NAND4_X1 U13971 ( .A1(n12254), .A2(n12253), .A3(n12252), .A4(n12251), .ZN(
        n12255) );
  AOI22_X1 U13972 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U13973 ( .A1(n12321), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12257) );
  OAI211_X1 U13974 ( .C1(n15534), .C2(n12334), .A(n12258), .B(n12257), .ZN(
        n15234) );
  AOI22_X1 U13975 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12262) );
  AOI22_X1 U13976 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U13977 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U13978 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12259) );
  NAND4_X1 U13979 ( .A1(n12262), .A2(n12261), .A3(n12260), .A4(n12259), .ZN(
        n12268) );
  AOI22_X1 U13980 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U13981 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U13982 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U13983 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12263) );
  NAND4_X1 U13984 ( .A1(n12266), .A2(n12265), .A3(n12264), .A4(n12263), .ZN(
        n12267) );
  NOR2_X1 U13985 ( .A1(n12268), .A2(n12267), .ZN(n15776) );
  NOR2_X1 U13986 ( .A1(n12334), .A2(n15776), .ZN(n12271) );
  INV_X1 U13987 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17742) );
  INV_X1 U13988 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n12269) );
  OAI22_X1 U13989 ( .A1(n12351), .A2(n17742), .B1(n12350), .B2(n12269), .ZN(
        n12270) );
  AOI211_X1 U13990 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n12321), .A(n12271), .B(
        n12270), .ZN(n16102) );
  AOI22_X1 U13991 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U13992 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U13993 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U13994 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12272) );
  NAND4_X1 U13995 ( .A1(n12275), .A2(n12274), .A3(n12273), .A4(n12272), .ZN(
        n12281) );
  AOI22_X1 U13996 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U13997 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U13998 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U13999 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12276) );
  NAND4_X1 U14000 ( .A1(n12279), .A2(n12278), .A3(n12277), .A4(n12276), .ZN(
        n12280) );
  AOI22_X1 U14001 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n12283) );
  NAND2_X1 U14002 ( .A1(n12321), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12282) );
  OAI211_X1 U14003 ( .C1(n15957), .C2(n12334), .A(n12283), .B(n12282), .ZN(
        n15425) );
  AOI22_X1 U14004 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U14005 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U14006 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U14007 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12284) );
  NAND4_X1 U14008 ( .A1(n12287), .A2(n12286), .A3(n12285), .A4(n12284), .ZN(
        n12293) );
  AOI22_X1 U14009 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U14010 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U14011 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U14012 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12288) );
  NAND4_X1 U14013 ( .A1(n12291), .A2(n12290), .A3(n12289), .A4(n12288), .ZN(
        n12292) );
  INV_X1 U14014 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n16116) );
  AOI22_X1 U14015 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12294) );
  OAI21_X1 U14016 ( .B1(n12352), .B2(n16116), .A(n12294), .ZN(n12295) );
  AOI21_X1 U14017 ( .B1(n12346), .B2(n15882), .A(n12295), .ZN(n15493) );
  AOI22_X1 U14018 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n14445), .B1(
        n14414), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U14019 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n14446), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U14020 ( .A1(n14479), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U14021 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11174), .B1(
        n14460), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12296) );
  NAND4_X1 U14022 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12305) );
  AOI22_X1 U14023 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n14485), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U14024 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U14025 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14490), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U14026 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14488), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12300) );
  NAND4_X1 U14027 ( .A1(n12303), .A2(n12302), .A3(n12301), .A4(n12300), .ZN(
        n12304) );
  NOR2_X1 U14028 ( .A1(n12305), .A2(n12304), .ZN(n16038) );
  AOI22_X1 U14029 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n12307) );
  NAND2_X1 U14030 ( .A1(n12321), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12306) );
  OAI211_X1 U14031 ( .C1(n16038), .C2(n12334), .A(n12307), .B(n12306), .ZN(
        n15503) );
  AOI22_X1 U14032 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U14033 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U14034 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U14035 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12308) );
  NAND4_X1 U14036 ( .A1(n12311), .A2(n12310), .A3(n12309), .A4(n12308), .ZN(
        n12317) );
  AOI22_X1 U14037 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U14038 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U14039 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U14040 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12312) );
  NAND4_X1 U14041 ( .A1(n12315), .A2(n12314), .A3(n12313), .A4(n12312), .ZN(
        n12316) );
  NOR2_X1 U14042 ( .A1(n12334), .A2(n16233), .ZN(n12320) );
  INV_X1 U14043 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17696) );
  INV_X1 U14044 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n12318) );
  OAI22_X1 U14045 ( .A1(n12351), .A2(n17696), .B1(n12350), .B2(n12318), .ZN(
        n12319) );
  AOI211_X1 U14046 ( .C1(n12321), .C2(P2_REIP_REG_13__SCAN_IN), .A(n12320), 
        .B(n12319), .ZN(n17690) );
  AOI22_X1 U14047 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U14048 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U14049 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U14050 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11174), .B1(
        n14460), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12322) );
  NAND4_X1 U14051 ( .A1(n12325), .A2(n12324), .A3(n12323), .A4(n12322), .ZN(
        n12331) );
  AOI22_X1 U14052 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n14485), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U14053 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U14054 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14490), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U14055 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14488), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12326) );
  NAND4_X1 U14056 ( .A1(n12329), .A2(n12328), .A3(n12327), .A4(n12326), .ZN(
        n12330) );
  OR2_X1 U14057 ( .A1(n12331), .A2(n12330), .ZN(n16241) );
  INV_X1 U14058 ( .A(n16241), .ZN(n12335) );
  AOI22_X1 U14059 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n12333) );
  NAND2_X1 U14060 ( .A1(n12321), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12332) );
  OAI211_X1 U14061 ( .C1(n12335), .C2(n12334), .A(n12333), .B(n12332), .ZN(
        n15790) );
  AOI22_X1 U14062 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U14063 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U14064 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U14065 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12336) );
  NAND4_X1 U14066 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12345) );
  AOI22_X1 U14067 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U14068 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U14069 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U14070 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12340) );
  NAND4_X1 U14071 ( .A1(n12343), .A2(n12342), .A3(n12341), .A4(n12340), .ZN(
        n12344) );
  NAND2_X1 U14072 ( .A1(n12346), .A2(n16245), .ZN(n12349) );
  AOI22_X1 U14073 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n12348) );
  NAND2_X1 U14074 ( .A1(n12321), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12347) );
  INV_X1 U14075 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n18087) );
  INV_X1 U14076 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n19268) );
  INV_X1 U14077 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n15401) );
  OAI222_X1 U14078 ( .A1(n12352), .A2(n18087), .B1(n12351), .B2(n19268), .C1(
        n12350), .C2(n15401), .ZN(n19116) );
  AOI22_X1 U14079 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12354) );
  NAND2_X1 U14080 ( .A1(n12321), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12353) );
  NOR2_X2 U14081 ( .A1(n15099), .A2(n15100), .ZN(n17374) );
  NAND2_X1 U14082 ( .A1(n17375), .A2(n17374), .ZN(n17377) );
  AOI22_X1 U14083 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12356) );
  NAND2_X1 U14084 ( .A1(n12321), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U14085 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12358) );
  NAND2_X1 U14086 ( .A1(n12321), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12357) );
  NAND2_X1 U14087 ( .A1(n12358), .A2(n12357), .ZN(n14216) );
  AND2_X2 U14088 ( .A1(n17365), .A2(n14216), .ZN(n17156) );
  AOI22_X1 U14089 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12360) );
  NAND2_X1 U14090 ( .A1(n12321), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12359) );
  NAND2_X1 U14091 ( .A1(n12360), .A2(n12359), .ZN(n17157) );
  AOI22_X1 U14092 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n12362) );
  NAND2_X1 U14093 ( .A1(n12321), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12361) );
  AND2_X1 U14094 ( .A1(n12362), .A2(n12361), .ZN(n17340) );
  AOI22_X1 U14095 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12364) );
  NAND2_X1 U14096 ( .A1(n12321), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12363) );
  AND2_X1 U14097 ( .A1(n12364), .A2(n12363), .ZN(n17137) );
  AOI22_X1 U14098 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n12366) );
  NAND2_X1 U14099 ( .A1(n12321), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12365) );
  NOR2_X2 U14100 ( .A1(n17139), .A2(n17127), .ZN(n17319) );
  AOI22_X1 U14101 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n12370) );
  NAND2_X1 U14102 ( .A1(n12321), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12369) );
  NAND2_X1 U14103 ( .A1(n12370), .A2(n12369), .ZN(n17318) );
  NAND2_X1 U14104 ( .A1(n17319), .A2(n17318), .ZN(n17307) );
  AOI22_X1 U14105 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n12372) );
  NAND2_X1 U14106 ( .A1(n12321), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12371) );
  AND2_X1 U14107 ( .A1(n12372), .A2(n12371), .ZN(n17308) );
  AOI22_X1 U14108 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12374) );
  NAND2_X1 U14109 ( .A1(n12321), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12373) );
  AND2_X1 U14110 ( .A1(n12374), .A2(n12373), .ZN(n14301) );
  AOI22_X1 U14111 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n12376) );
  NAND2_X1 U14112 ( .A1(n12321), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12375) );
  NAND2_X1 U14113 ( .A1(n12376), .A2(n12375), .ZN(n14287) );
  AOI22_X1 U14114 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n12378) );
  NAND2_X1 U14115 ( .A1(n12321), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12377) );
  NAND2_X1 U14116 ( .A1(n12378), .A2(n12377), .ZN(n17285) );
  AOI22_X1 U14117 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n12367), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n12380) );
  NAND2_X1 U14118 ( .A1(n12321), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12379) );
  AND2_X1 U14119 ( .A1(n12380), .A2(n12379), .ZN(n17087) );
  INV_X1 U14120 ( .A(n16359), .ZN(n12382) );
  INV_X1 U14121 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n22323) );
  NAND2_X1 U14122 ( .A1(n22307), .A2(n22323), .ZN(n22305) );
  NAND2_X1 U14123 ( .A1(n22312), .A2(n12431), .ZN(n15709) );
  AND2_X1 U14124 ( .A1(n11156), .A2(n20262), .ZN(n14155) );
  INV_X1 U14125 ( .A(n14155), .ZN(n15708) );
  NOR2_X1 U14126 ( .A1(n15709), .A2(n15708), .ZN(n12381) );
  AOI222_X1 U14127 ( .A1(n14327), .A2(n19218), .B1(n19217), .B2(n16323), .C1(
        n12382), .C2(n19140), .ZN(n12438) );
  NOR2_X1 U14128 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17842) );
  INV_X1 U14129 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n22273) );
  NAND3_X1 U14130 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n17842), .A3(n22273), 
        .ZN(n19347) );
  NAND2_X1 U14131 ( .A1(n12085), .A2(n14346), .ZN(n18021) );
  INV_X1 U14132 ( .A(n17842), .ZN(n12383) );
  OR2_X2 U14133 ( .A1(n18021), .A2(n12383), .ZN(n19325) );
  NOR4_X1 U14134 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n17901), .A4(n14346), .ZN(n17807) );
  INV_X1 U14135 ( .A(n17807), .ZN(n12384) );
  NAND3_X1 U14136 ( .A1(n19347), .A2(n19325), .A3(n12384), .ZN(n12385) );
  NOR2_X2 U14137 ( .A1(n15107), .A2(n12385), .ZN(n19163) );
  XNOR2_X1 U14138 ( .A(n12388), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16316) );
  INV_X1 U14139 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17083) );
  NOR2_X1 U14140 ( .A1(n16316), .A2(n19193), .ZN(n17080) );
  INV_X1 U14141 ( .A(n12387), .ZN(n12429) );
  NAND2_X1 U14142 ( .A1(n12429), .A2(n17415), .ZN(n12389) );
  AND2_X1 U14143 ( .A1(n12389), .A2(n12388), .ZN(n17417) );
  INV_X1 U14144 ( .A(n17417), .ZN(n19213) );
  NOR2_X1 U14145 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n12390), .ZN(
        n12391) );
  NOR2_X1 U14146 ( .A1(n12426), .A2(n12391), .ZN(n17105) );
  AND2_X1 U14147 ( .A1(n11206), .A2(n19183), .ZN(n12392) );
  OAI21_X1 U14148 ( .B1(n12419), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n12421), .ZN(n12393) );
  INV_X1 U14149 ( .A(n12393), .ZN(n17456) );
  NAND2_X1 U14150 ( .A1(n17477), .A2(n12415), .ZN(n12394) );
  AND2_X1 U14151 ( .A1(n12394), .A2(n12417), .ZN(n17479) );
  AOI21_X1 U14152 ( .B1(n12413), .B2(n17489), .A(n12416), .ZN(n19135) );
  OAI21_X1 U14153 ( .B1(n12410), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n12395), .ZN(n15095) );
  INV_X1 U14154 ( .A(n15095), .ZN(n17509) );
  AOI21_X1 U14155 ( .B1(n12408), .B2(n17523), .A(n12396), .ZN(n17526) );
  AOI21_X1 U14156 ( .B1(n17988), .B2(n12406), .A(n12409), .ZN(n19095) );
  AOI21_X1 U14157 ( .B1(n12100), .B2(n12404), .A(n12407), .ZN(n17964) );
  AOI21_X1 U14158 ( .B1(n17958), .B2(n12402), .A(n12405), .ZN(n17951) );
  AOI21_X1 U14159 ( .B1(n16143), .B2(n12400), .A(n12403), .ZN(n17933) );
  AOI21_X1 U14160 ( .B1(n17932), .B2(n12398), .A(n12401), .ZN(n17924) );
  AOI21_X1 U14161 ( .B1(n17923), .B2(n12397), .A(n12399), .ZN(n17912) );
  OAI22_X1 U14162 ( .A1(n17901), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19030) );
  INV_X1 U14163 ( .A(n19030), .ZN(n17181) );
  INV_X1 U14164 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15206) );
  AOI22_X1 U14165 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15206), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17901), .ZN(n17180) );
  NOR2_X1 U14166 ( .A1(n17181), .A2(n17180), .ZN(n17179) );
  OAI21_X1 U14167 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12397), .ZN(n17174) );
  NAND2_X1 U14168 ( .A1(n17179), .A2(n17174), .ZN(n16052) );
  NOR2_X1 U14169 ( .A1(n17912), .A2(n16052), .ZN(n19031) );
  OAI21_X1 U14170 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12399), .A(
        n12398), .ZN(n19032) );
  NAND2_X1 U14171 ( .A1(n19031), .A2(n19032), .ZN(n16127) );
  NOR2_X1 U14172 ( .A1(n17924), .A2(n16127), .ZN(n19049) );
  OAI21_X1 U14173 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12401), .A(
        n12400), .ZN(n19050) );
  NAND2_X1 U14174 ( .A1(n19049), .A2(n19050), .ZN(n16140) );
  NOR2_X1 U14175 ( .A1(n17933), .A2(n16140), .ZN(n19058) );
  OAI21_X1 U14176 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12403), .A(
        n12402), .ZN(n19059) );
  NAND2_X1 U14177 ( .A1(n19058), .A2(n19059), .ZN(n16103) );
  NOR2_X1 U14178 ( .A1(n17951), .A2(n16103), .ZN(n19070) );
  OAI21_X1 U14179 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12405), .A(
        n12404), .ZN(n19071) );
  NAND2_X1 U14180 ( .A1(n19070), .A2(n19071), .ZN(n16111) );
  NOR2_X1 U14181 ( .A1(n17964), .A2(n16111), .ZN(n19082) );
  OAI21_X1 U14182 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12407), .A(
        n12406), .ZN(n19083) );
  NAND2_X1 U14183 ( .A1(n19082), .A2(n19083), .ZN(n19096) );
  NOR2_X1 U14184 ( .A1(n19095), .A2(n19096), .ZN(n19094) );
  OAI21_X1 U14185 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12409), .A(
        n12408), .ZN(n19105) );
  NAND2_X1 U14186 ( .A1(n19094), .A2(n19105), .ZN(n16211) );
  NOR2_X1 U14187 ( .A1(n17526), .A2(n16211), .ZN(n19110) );
  AOI21_X1 U14188 ( .B1(n12123), .B2(n12411), .A(n12410), .ZN(n19112) );
  INV_X1 U14189 ( .A(n19112), .ZN(n12412) );
  NAND2_X1 U14190 ( .A1(n19110), .A2(n12412), .ZN(n15093) );
  NOR2_X1 U14191 ( .A1(n17509), .A2(n15093), .ZN(n19125) );
  OAI21_X1 U14192 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12414), .A(
        n12413), .ZN(n19126) );
  NAND2_X1 U14193 ( .A1(n19125), .A2(n19126), .ZN(n19133) );
  NOR2_X1 U14194 ( .A1(n19135), .A2(n19133), .ZN(n19156) );
  OAI21_X1 U14195 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12416), .A(
        n12415), .ZN(n19159) );
  NAND2_X1 U14196 ( .A1(n19156), .A2(n19159), .ZN(n17151) );
  NOR2_X1 U14197 ( .A1(n17479), .A2(n17151), .ZN(n19170) );
  AND2_X1 U14198 ( .A1(n12418), .A2(n12417), .ZN(n12420) );
  OR2_X1 U14199 ( .A1(n12420), .A2(n12419), .ZN(n19169) );
  NAND2_X1 U14200 ( .A1(n19170), .A2(n19169), .ZN(n17144) );
  NOR2_X1 U14201 ( .A1(n17456), .A2(n17144), .ZN(n17119) );
  NAND2_X1 U14202 ( .A1(n12421), .A2(n17443), .ZN(n12422) );
  AND2_X1 U14203 ( .A1(n11206), .A2(n12422), .ZN(n17445) );
  INV_X1 U14204 ( .A(n17445), .ZN(n12423) );
  NAND2_X1 U14205 ( .A1(n17119), .A2(n12423), .ZN(n19177) );
  NOR2_X1 U14206 ( .A1(n11751), .A2(n19177), .ZN(n19192) );
  OAI21_X1 U14207 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n12425), .A(
        n12424), .ZN(n19191) );
  NAND2_X1 U14208 ( .A1(n19192), .A2(n19191), .ZN(n17106) );
  NOR2_X1 U14209 ( .A1(n17105), .A2(n17106), .ZN(n17093) );
  INV_X1 U14210 ( .A(n12426), .ZN(n12427) );
  NAND2_X1 U14211 ( .A1(n12427), .A2(n17099), .ZN(n12428) );
  NAND2_X1 U14212 ( .A1(n12429), .A2(n12428), .ZN(n17095) );
  NAND2_X1 U14213 ( .A1(n17093), .A2(n17095), .ZN(n12430) );
  NAND2_X1 U14214 ( .A1(n11173), .A2(n12430), .ZN(n19215) );
  AOI21_X1 U14215 ( .B1(n19213), .B2(n19215), .A(n19347), .ZN(n19214) );
  AOI22_X1 U14216 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19208), .B1(
        n17080), .B2(n19214), .ZN(n12437) );
  NOR3_X1 U14217 ( .A1(n17417), .A2(n19347), .A3(n12430), .ZN(n17079) );
  NOR2_X1 U14218 ( .A1(n11173), .A2(n19347), .ZN(n19092) );
  OAI21_X1 U14219 ( .B1(n17079), .B2(n19092), .A(n16316), .ZN(n12436) );
  INV_X1 U14220 ( .A(n15709), .ZN(n12432) );
  OAI22_X1 U14221 ( .A1(n12432), .A2(n11354), .B1(P2_EBX_REG_31__SCAN_IN), 
        .B2(n12431), .ZN(n12433) );
  INV_X1 U14222 ( .A(n12433), .ZN(n12434) );
  AOI22_X1 U14223 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19207), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19163), .ZN(n12435) );
  NAND4_X1 U14224 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        P2_U2825) );
  AOI22_X1 U14225 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12442) );
  INV_X2 U14226 ( .A(n11238), .ZN(n18466) );
  AOI22_X1 U14227 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18329), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12441) );
  NOR2_X2 U14228 ( .A1(n21460), .A2(n21500), .ZN(n12486) );
  BUF_X4 U14229 ( .A(n12486), .Z(n18468) );
  AOI22_X1 U14230 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U14231 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12439) );
  NAND4_X1 U14232 ( .A1(n12442), .A2(n12441), .A3(n12440), .A4(n12439), .ZN(
        n12452) );
  NOR2_X2 U14233 ( .A1(n20849), .A2(n16298), .ZN(n18475) );
  AOI22_X1 U14234 ( .A1(n18475), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18474), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U14235 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12449) );
  NOR2_X2 U14236 ( .A1(n20849), .A2(n12444), .ZN(n12576) );
  INV_X2 U14237 ( .A(n11205), .ZN(n18449) );
  AOI22_X1 U14238 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18449), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12448) );
  NOR2_X2 U14239 ( .A1(n12445), .A2(n21485), .ZN(n12475) );
  AOI22_X1 U14240 ( .A1(n12475), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12447) );
  NAND4_X1 U14241 ( .A1(n12450), .A2(n12449), .A3(n12448), .A4(n12447), .ZN(
        n12451) );
  AOI22_X1 U14242 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U14243 ( .A1(n18475), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U14244 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U14245 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12453) );
  NAND4_X1 U14246 ( .A1(n12456), .A2(n12455), .A3(n12454), .A4(n12453), .ZN(
        n12462) );
  AOI22_X1 U14247 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U14248 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18449), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U14249 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U14250 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12457) );
  NAND4_X1 U14251 ( .A1(n12460), .A2(n12459), .A3(n12458), .A4(n12457), .ZN(
        n12461) );
  AOI22_X1 U14252 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18416), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U14253 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18449), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U14254 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U14255 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12463) );
  NAND4_X1 U14256 ( .A1(n12466), .A2(n12465), .A3(n12464), .A4(n12463), .ZN(
        n12472) );
  AOI22_X1 U14257 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U14258 ( .A1(n18475), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18474), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U14259 ( .A1(n18476), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12468) );
  AOI22_X1 U14260 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12467) );
  NAND4_X1 U14261 ( .A1(n12470), .A2(n12469), .A3(n12468), .A4(n12467), .ZN(
        n12471) );
  INV_X2 U14262 ( .A(n11238), .ZN(n18439) );
  AOI22_X1 U14263 ( .A1(n12592), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U14264 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18449), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12482) );
  INV_X1 U14265 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18309) );
  AOI22_X1 U14266 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12474) );
  OAI21_X1 U14267 ( .B1(n12523), .B2(n18309), .A(n12474), .ZN(n12481) );
  AOI22_X1 U14268 ( .A1(n12609), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12475), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12480) );
  AOI22_X1 U14269 ( .A1(n18475), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12576), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U14270 ( .A1(n12490), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12489), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U14271 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12524), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12477) );
  INV_X1 U14272 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18488) );
  AOI22_X1 U14273 ( .A1(n12473), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n11167), .ZN(n12484) );
  OAI21_X1 U14274 ( .B1(n18488), .B2(n12523), .A(n12484), .ZN(n12485) );
  AOI22_X1 U14275 ( .A1(n12592), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n12475), .ZN(n12487) );
  INV_X1 U14276 ( .A(n12487), .ZN(n12488) );
  AOI22_X1 U14277 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12476), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12495) );
  AOI22_X1 U14278 ( .A1(n12609), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12489), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U14279 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n12524), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U14280 ( .A1(n18475), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12576), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U14281 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12490), .B1(
        n18449), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U14282 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18449), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12508) );
  AOI22_X1 U14283 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12507) );
  INV_X1 U14284 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18321) );
  AOI22_X1 U14285 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12499) );
  OAI21_X1 U14286 ( .B1(n12523), .B2(n18321), .A(n12499), .ZN(n12505) );
  AOI22_X1 U14287 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12503) );
  AOI22_X1 U14288 ( .A1(n18475), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U14289 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U14290 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18416), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12500) );
  NAND4_X1 U14291 ( .A1(n12503), .A2(n12502), .A3(n12501), .A4(n12500), .ZN(
        n12504) );
  AOI211_X1 U14292 ( .C1(n18454), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n12505), .B(n12504), .ZN(n12506) );
  NAND3_X1 U14293 ( .A1(n12508), .A2(n12507), .A3(n12506), .ZN(n12708) );
  NAND2_X1 U14294 ( .A1(n12519), .A2(n12708), .ZN(n12542) );
  AOI22_X1 U14295 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U14296 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12517) );
  AOI22_X1 U14297 ( .A1(n18469), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12509) );
  OAI21_X1 U14298 ( .B1(n12523), .B2(n18409), .A(n12509), .ZN(n12515) );
  AOI22_X1 U14299 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12513) );
  AOI22_X1 U14300 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12512) );
  CLKBUF_X3 U14301 ( .A(n12592), .Z(n18319) );
  AOI22_X1 U14302 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12511) );
  AOI22_X1 U14303 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18449), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12510) );
  NAND4_X1 U14304 ( .A1(n12513), .A2(n12512), .A3(n12511), .A4(n12510), .ZN(
        n12514) );
  AOI211_X1 U14305 ( .C1(n18468), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n12515), .B(n12514), .ZN(n12516) );
  NAND3_X1 U14306 ( .A1(n12518), .A2(n12517), .A3(n12516), .ZN(n12709) );
  INV_X1 U14307 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21600) );
  INV_X1 U14308 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21589) );
  INV_X1 U14309 ( .A(n12708), .ZN(n21322) );
  XNOR2_X1 U14310 ( .A(n21322), .B(n12519), .ZN(n12541) );
  INV_X1 U14311 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21564) );
  INV_X1 U14312 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21543) );
  NOR2_X1 U14313 ( .A1(n12520), .A2(n21543), .ZN(n12534) );
  XNOR2_X1 U14314 ( .A(n21451), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18880) );
  AOI22_X1 U14315 ( .A1(n12609), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12489), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12533) );
  AOI22_X1 U14316 ( .A1(n12592), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12576), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12532) );
  INV_X1 U14317 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18287) );
  AOI22_X1 U14318 ( .A1(n12486), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12522) );
  OAI21_X1 U14319 ( .B1(n12523), .B2(n18287), .A(n12522), .ZN(n12530) );
  AOI22_X1 U14320 ( .A1(n12473), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18449), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12528) );
  AOI22_X1 U14321 ( .A1(n12498), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12524), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12527) );
  AOI22_X1 U14322 ( .A1(n18475), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12526) );
  AOI22_X1 U14323 ( .A1(n12490), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12475), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12525) );
  NAND4_X1 U14324 ( .A1(n12528), .A2(n12527), .A3(n12526), .A4(n12525), .ZN(
        n12529) );
  AOI211_X1 U14325 ( .C1(n18454), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n12530), .B(n12529), .ZN(n12531) );
  NAND3_X1 U14326 ( .A1(n12533), .A2(n12532), .A3(n12531), .ZN(n21452) );
  NAND2_X1 U14327 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n11152), .ZN(
        n18886) );
  NOR2_X1 U14328 ( .A1(n18880), .A2(n18886), .ZN(n18879) );
  NOR2_X1 U14329 ( .A1(n12534), .A2(n18879), .ZN(n18866) );
  OR2_X1 U14330 ( .A1(n21330), .A2(n12520), .ZN(n12535) );
  NOR2_X1 U14331 ( .A1(n18866), .A2(n18865), .ZN(n18864) );
  NOR2_X1 U14332 ( .A1(n12536), .A2(n12537), .ZN(n12538) );
  XNOR2_X1 U14333 ( .A(n21326), .B(n12717), .ZN(n18855) );
  NOR2_X1 U14334 ( .A1(n12539), .A2(n21564), .ZN(n12540) );
  XNOR2_X1 U14335 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12541), .ZN(
        n18844) );
  XNOR2_X1 U14336 ( .A(n21317), .B(n12542), .ZN(n12544) );
  NOR2_X1 U14337 ( .A1(n12543), .A2(n12544), .ZN(n12545) );
  INV_X1 U14338 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18833) );
  NOR2_X1 U14339 ( .A1(n18833), .A2(n18832), .ZN(n18831) );
  INV_X1 U14340 ( .A(n12709), .ZN(n21313) );
  XNOR2_X1 U14341 ( .A(n21313), .B(n12546), .ZN(n12547) );
  XNOR2_X1 U14342 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12547), .ZN(
        n18819) );
  NOR2_X1 U14343 ( .A1(n18820), .A2(n18819), .ZN(n18818) );
  OAI21_X1 U14344 ( .B1(n12549), .B2(n18501), .A(n21762), .ZN(n12550) );
  NOR2_X1 U14345 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18773) );
  INV_X1 U14346 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21852) );
  AND2_X1 U14347 ( .A1(n18773), .A2(n21852), .ZN(n12551) );
  NAND2_X1 U14348 ( .A1(n21853), .A2(n12552), .ZN(n12553) );
  NOR2_X1 U14349 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12554) );
  INV_X1 U14350 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21889) );
  INV_X1 U14351 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21862) );
  NOR2_X1 U14352 ( .A1(n21889), .A2(n21862), .ZN(n21621) );
  NAND2_X1 U14353 ( .A1(n21621), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n21635) );
  NOR2_X1 U14354 ( .A1(n21635), .A2(n21853), .ZN(n21629) );
  NAND2_X1 U14355 ( .A1(n21629), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n21645) );
  NOR2_X1 U14356 ( .A1(n21661), .A2(n21645), .ZN(n21664) );
  NAND2_X1 U14357 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21664), .ZN(
        n21829) );
  INV_X1 U14358 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21770) );
  INV_X1 U14359 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21844) );
  INV_X1 U14360 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21837) );
  NOR2_X1 U14361 ( .A1(n21844), .A2(n21837), .ZN(n21816) );
  NAND2_X1 U14362 ( .A1(n21816), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n21510) );
  INV_X1 U14363 ( .A(n21510), .ZN(n12742) );
  NAND2_X1 U14364 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18592) );
  INV_X1 U14365 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18586) );
  NOR2_X1 U14366 ( .A1(n18592), .A2(n18586), .ZN(n21688) );
  NAND2_X1 U14367 ( .A1(n12742), .A2(n21688), .ZN(n18640) );
  NOR2_X1 U14368 ( .A1(n21770), .A2(n18640), .ZN(n12745) );
  INV_X1 U14369 ( .A(n12745), .ZN(n12555) );
  OAI21_X1 U14370 ( .B1(n18539), .B2(n12555), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12562) );
  INV_X1 U14371 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21800) );
  NAND2_X1 U14372 ( .A1(n18598), .A2(n21800), .ZN(n12556) );
  NOR2_X1 U14373 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12556), .ZN(
        n18585) );
  NAND2_X1 U14374 ( .A1(n18585), .A2(n18586), .ZN(n18576) );
  NOR2_X1 U14375 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18576), .ZN(
        n18618) );
  OR2_X1 U14376 ( .A1(n18618), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12561) );
  NAND3_X1 U14377 ( .A1(n12562), .A2(n12561), .A3(n18596), .ZN(n18638) );
  NOR2_X2 U14378 ( .A1(n18638), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18637) );
  INV_X1 U14379 ( .A(n18637), .ZN(n12564) );
  INV_X1 U14380 ( .A(n21816), .ZN(n18511) );
  NAND2_X1 U14381 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21783) );
  NAND2_X1 U14382 ( .A1(n12564), .A2(n12563), .ZN(n18632) );
  INV_X1 U14383 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21711) );
  INV_X1 U14384 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21695) );
  NOR2_X1 U14385 ( .A1(n21711), .A2(n21695), .ZN(n21705) );
  INV_X1 U14386 ( .A(n21705), .ZN(n12567) );
  AOI21_X1 U14387 ( .B1(n21711), .B2(n21695), .A(n18793), .ZN(n12565) );
  INV_X1 U14388 ( .A(n12565), .ZN(n12566) );
  OAI211_X1 U14389 ( .C1(n18632), .C2(n12567), .A(n12566), .B(n11231), .ZN(
        n12568) );
  INV_X1 U14390 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21759) );
  NOR2_X1 U14391 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18793), .ZN(
        n18661) );
  NAND2_X1 U14392 ( .A1(n18663), .A2(n18661), .ZN(n18720) );
  NAND2_X1 U14393 ( .A1(n12570), .A2(n12569), .ZN(n12573) );
  NAND2_X1 U14394 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12572) );
  OAI21_X1 U14395 ( .B1(n18720), .B2(n12573), .A(n11232), .ZN(n12575) );
  XNOR2_X1 U14396 ( .A(n12575), .B(n12574), .ZN(n18700) );
  AOI22_X1 U14397 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U14398 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U14399 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U14400 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12578) );
  NAND4_X1 U14401 ( .A1(n12581), .A2(n12580), .A3(n12579), .A4(n12578), .ZN(
        n12587) );
  AOI22_X1 U14402 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U14403 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U14404 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12583) );
  INV_X2 U14405 ( .A(n18172), .ZN(n18363) );
  AOI22_X1 U14406 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12582) );
  NAND4_X1 U14407 ( .A1(n12585), .A2(n12584), .A3(n12583), .A4(n12582), .ZN(
        n12586) );
  AOI22_X1 U14408 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U14409 ( .A1(n18439), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18474), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12590) );
  INV_X2 U14410 ( .A(n11205), .ZN(n18477) );
  AOI22_X1 U14411 ( .A1(n18477), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U14412 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12588) );
  NAND4_X1 U14413 ( .A1(n12591), .A2(n12590), .A3(n12589), .A4(n12588), .ZN(
        n12598) );
  AOI22_X1 U14414 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U14415 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U14416 ( .A1(n18476), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U14417 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18416), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12593) );
  NAND4_X1 U14418 ( .A1(n12596), .A2(n12595), .A3(n12594), .A4(n12593), .ZN(
        n12597) );
  AOI22_X1 U14419 ( .A1(n18477), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U14420 ( .A1(n18476), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12601) );
  AOI22_X1 U14421 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U14422 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12599) );
  NAND4_X1 U14423 ( .A1(n12602), .A2(n12601), .A3(n12600), .A4(n12599), .ZN(
        n12608) );
  AOI22_X1 U14424 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U14425 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U14426 ( .A1(n18439), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18416), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U14427 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12603) );
  NAND4_X1 U14428 ( .A1(n12606), .A2(n12605), .A3(n12604), .A4(n12603), .ZN(
        n12607) );
  AOI22_X1 U14429 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18329), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U14430 ( .A1(n18476), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U14431 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12610) );
  OAI21_X1 U14432 ( .B1(n18172), .B2(n18409), .A(n12610), .ZN(n12615) );
  AOI22_X1 U14433 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U14434 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18474), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U14435 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12612) );
  AOI22_X1 U14436 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12611) );
  AOI22_X1 U14437 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18449), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U14438 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18416), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U14439 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U14440 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12618) );
  NAND4_X1 U14441 ( .A1(n12621), .A2(n12620), .A3(n12619), .A4(n12618), .ZN(
        n12627) );
  AOI22_X1 U14442 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12625) );
  AOI22_X1 U14443 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U14444 ( .A1(n12475), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12623) );
  AOI22_X1 U14445 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12622) );
  NAND4_X1 U14446 ( .A1(n12625), .A2(n12624), .A3(n12623), .A4(n12622), .ZN(
        n12626) );
  NAND2_X1 U14447 ( .A1(n19632), .A2(n19550), .ZN(n12685) );
  AOI22_X1 U14448 ( .A1(n18477), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12637) );
  AOI22_X1 U14449 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12636) );
  AOI22_X1 U14450 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12628) );
  OAI21_X1 U14451 ( .B1(n18172), .B2(n18298), .A(n12628), .ZN(n12634) );
  AOI22_X1 U14452 ( .A1(n18439), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18329), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U14453 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U14454 ( .A1(n18475), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U14455 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12629) );
  NAND4_X1 U14456 ( .A1(n12632), .A2(n12631), .A3(n12630), .A4(n12629), .ZN(
        n12633) );
  NOR2_X1 U14457 ( .A1(n21438), .A2(n21459), .ZN(n21284) );
  AOI22_X1 U14458 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18329), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U14459 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18319), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U14460 ( .A1(n12475), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12638) );
  OAI21_X1 U14461 ( .B1(n18172), .B2(n18488), .A(n12638), .ZN(n12644) );
  AOI22_X1 U14462 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12642) );
  AOI22_X1 U14463 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18416), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12641) );
  AOI22_X1 U14464 ( .A1(n18469), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U14465 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12639) );
  NAND4_X1 U14466 ( .A1(n12642), .A2(n12641), .A3(n12640), .A4(n12639), .ZN(
        n12643) );
  NOR3_X1 U14467 ( .A1(n21278), .A2(n21284), .A3(n20850), .ZN(n12695) );
  INV_X1 U14468 ( .A(n12695), .ZN(n12660) );
  NAND2_X1 U14469 ( .A1(n20850), .A2(n21278), .ZN(n12701) );
  NAND2_X1 U14470 ( .A1(n12701), .A2(n19632), .ZN(n12690) );
  AOI22_X1 U14471 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18416), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U14472 ( .A1(n18477), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U14473 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U14474 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12648) );
  NAND4_X1 U14475 ( .A1(n12651), .A2(n12650), .A3(n12649), .A4(n12648), .ZN(
        n12657) );
  AOI22_X1 U14476 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U14477 ( .A1(n18363), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U14478 ( .A1(n18439), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18474), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U14479 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12652) );
  NAND4_X1 U14480 ( .A1(n12655), .A2(n12654), .A3(n12653), .A4(n12652), .ZN(
        n12656) );
  NAND2_X1 U14481 ( .A1(n21335), .A2(n21336), .ZN(n12697) );
  OAI211_X1 U14482 ( .C1(n21459), .C2(n19550), .A(n12706), .B(n12697), .ZN(
        n12658) );
  INV_X1 U14483 ( .A(n21336), .ZN(n19470) );
  NAND4_X1 U14484 ( .A1(n19592), .A2(n19550), .A3(n12689), .A4(n12692), .ZN(
        n12741) );
  OR2_X1 U14485 ( .A1(n12741), .A2(n19632), .ZN(n12700) );
  OAI21_X1 U14486 ( .B1(n12690), .B2(n12658), .A(n12700), .ZN(n12659) );
  OAI211_X1 U14487 ( .C1(n12687), .C2(n12685), .A(n12660), .B(n12659), .ZN(
        n16302) );
  AOI21_X1 U14488 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n21460), .A(
        n12671), .ZN(n12676) );
  OAI22_X1 U14489 ( .A1(n21491), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n19383), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12669) );
  AOI22_X1 U14490 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19403), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n21492), .ZN(n12675) );
  NAND2_X1 U14491 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12663), .ZN(
        n12665) );
  OAI22_X1 U14492 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17832), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12663), .ZN(n12667) );
  AOI21_X1 U14493 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12665), .A(
        n12667), .ZN(n12664) );
  NOR2_X1 U14494 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17832), .ZN(
        n12666) );
  AOI22_X1 U14495 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12667), .B1(
        n12666), .B2(n12665), .ZN(n12679) );
  NAND2_X1 U14496 ( .A1(n12670), .A2(n12669), .ZN(n12668) );
  OAI211_X1 U14497 ( .C1(n12670), .C2(n12669), .A(n12679), .B(n12668), .ZN(
        n12674) );
  NAND2_X1 U14498 ( .A1(n12672), .A2(n12674), .ZN(n12677) );
  XNOR2_X1 U14499 ( .A(n12671), .B(n12675), .ZN(n12673) );
  AOI21_X1 U14500 ( .B1(n12676), .B2(n12677), .A(n21897), .ZN(n21903) );
  NAND2_X1 U14501 ( .A1(n12707), .A2(n21903), .ZN(n12683) );
  AND2_X1 U14502 ( .A1(n12676), .A2(n12675), .ZN(n12678) );
  XOR2_X1 U14503 ( .A(n21279), .B(n19632), .Z(n12680) );
  INV_X2 U14504 ( .A(n22288), .ZN(n22333) );
  NAND2_X1 U14505 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22284), .ZN(n22330) );
  INV_X1 U14506 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n22335) );
  AOI21_X1 U14507 ( .B1(n22333), .B2(n22330), .A(n18990), .ZN(n20851) );
  NAND2_X1 U14508 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n22332) );
  OAI21_X1 U14509 ( .B1(n12680), .B2(n20851), .A(n22332), .ZN(n21920) );
  OAI21_X1 U14510 ( .B1(n21897), .B2(n21920), .A(n11333), .ZN(n12681) );
  OAI21_X1 U14511 ( .B1(n21901), .B2(n11333), .A(n12681), .ZN(n12682) );
  OAI21_X1 U14512 ( .B1(n19470), .B2(n12683), .A(n12682), .ZN(n12684) );
  NAND2_X1 U14513 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21481), .ZN(n21929) );
  INV_X1 U14514 ( .A(n12685), .ZN(n12686) );
  NAND2_X1 U14515 ( .A1(n12686), .A2(n12697), .ZN(n12688) );
  NOR2_X1 U14516 ( .A1(n19550), .A2(n21336), .ZN(n21473) );
  INV_X1 U14517 ( .A(n12689), .ZN(n12703) );
  NOR2_X1 U14518 ( .A1(n21438), .A2(n12692), .ZN(n12693) );
  INV_X1 U14519 ( .A(n12690), .ZN(n12691) );
  OAI22_X1 U14520 ( .A1(n19550), .A2(n12693), .B1(n12692), .B2(n12691), .ZN(
        n12694) );
  AOI211_X1 U14521 ( .C1(n19592), .C2(n12703), .A(n12695), .B(n12694), .ZN(
        n12696) );
  NAND2_X1 U14522 ( .A1(n12698), .A2(n12696), .ZN(n21503) );
  NAND2_X1 U14523 ( .A1(n19632), .A2(n19592), .ZN(n12704) );
  NOR2_X1 U14524 ( .A1(n12697), .A2(n12704), .ZN(n18107) );
  NAND3_X1 U14525 ( .A1(n21335), .A2(n12706), .A3(n12698), .ZN(n12699) );
  NAND2_X1 U14526 ( .A1(n12700), .A2(n12699), .ZN(n21919) );
  INV_X1 U14527 ( .A(n12704), .ZN(n21472) );
  NOR2_X1 U14528 ( .A1(n21279), .A2(n12706), .ZN(n21470) );
  AND3_X1 U14529 ( .A1(n12706), .A2(n12705), .A3(n21473), .ZN(n16300) );
  XNOR2_X1 U14530 ( .A(n21279), .B(n21278), .ZN(n17834) );
  NAND2_X1 U14531 ( .A1(n18700), .A2(n21885), .ZN(n12756) );
  NAND2_X1 U14532 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12744) );
  INV_X1 U14533 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21690) );
  INV_X1 U14534 ( .A(n21783), .ZN(n21709) );
  INV_X1 U14535 ( .A(n21645), .ZN(n21642) );
  NOR2_X1 U14536 ( .A1(n21326), .A2(n12714), .ZN(n12725) );
  NAND2_X1 U14537 ( .A1(n12725), .A2(n12708), .ZN(n12712) );
  NOR2_X1 U14538 ( .A1(n21317), .A2(n12712), .ZN(n12711) );
  NAND2_X1 U14539 ( .A1(n12711), .A2(n12709), .ZN(n12710) );
  NOR2_X1 U14540 ( .A1(n21751), .A2(n12710), .ZN(n12734) );
  XNOR2_X1 U14541 ( .A(n18501), .B(n12710), .ZN(n18810) );
  XNOR2_X1 U14542 ( .A(n21313), .B(n12711), .ZN(n12728) );
  XOR2_X1 U14543 ( .A(n21317), .B(n12712), .Z(n12713) );
  NAND2_X1 U14544 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12713), .ZN(
        n12727) );
  XNOR2_X1 U14545 ( .A(n18833), .B(n12713), .ZN(n18830) );
  XNOR2_X1 U14546 ( .A(n21326), .B(n12716), .ZN(n12715) );
  NAND2_X1 U14547 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12715), .ZN(
        n12723) );
  XNOR2_X1 U14548 ( .A(n21564), .B(n12715), .ZN(n18860) );
  NAND2_X1 U14549 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12718), .ZN(
        n12722) );
  AOI21_X1 U14550 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12520), .A(
        n11152), .ZN(n12720) );
  INV_X1 U14551 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21615) );
  NOR2_X1 U14552 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12520), .ZN(
        n12719) );
  NAND2_X1 U14553 ( .A1(n18868), .A2(n18867), .ZN(n12721) );
  NAND2_X1 U14554 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12724), .ZN(
        n12726) );
  XNOR2_X1 U14555 ( .A(n21322), .B(n12725), .ZN(n18847) );
  NAND2_X1 U14556 ( .A1(n18848), .A2(n18847), .ZN(n18846) );
  NAND2_X1 U14557 ( .A1(n12728), .A2(n12729), .ZN(n12730) );
  NAND2_X1 U14558 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18823), .ZN(
        n18822) );
  NAND2_X1 U14559 ( .A1(n12734), .A2(n12731), .ZN(n12735) );
  NAND2_X1 U14560 ( .A1(n18810), .A2(n18811), .ZN(n18809) );
  NAND2_X1 U14561 ( .A1(n12734), .A2(n12733), .ZN(n12732) );
  OAI211_X1 U14562 ( .C1(n12734), .C2(n12733), .A(n18809), .B(n12732), .ZN(
        n18792) );
  NAND2_X1 U14563 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18792), .ZN(
        n18791) );
  NAND2_X1 U14564 ( .A1(n21642), .A2(n21617), .ZN(n18750) );
  NAND2_X1 U14565 ( .A1(n21705), .A2(n18624), .ZN(n21707) );
  NAND3_X1 U14566 ( .A1(n21753), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12736) );
  XOR2_X1 U14567 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12736), .Z(
        n18704) );
  NAND2_X1 U14568 ( .A1(n21895), .A2(n21751), .ZN(n21794) );
  NAND2_X1 U14569 ( .A1(n21762), .A2(n11224), .ZN(n18754) );
  INV_X1 U14570 ( .A(n18754), .ZN(n18742) );
  NOR2_X2 U14571 ( .A1(n18742), .A2(n21600), .ZN(n18757) );
  NAND2_X1 U14572 ( .A1(n18757), .A2(n21642), .ZN(n18751) );
  NOR2_X2 U14573 ( .A1(n18751), .A2(n21661), .ZN(n21658) );
  NOR2_X2 U14574 ( .A1(n18640), .A2(n18518), .ZN(n21515) );
  NAND2_X1 U14575 ( .A1(n21709), .A2(n21515), .ZN(n21772) );
  NOR2_X2 U14576 ( .A1(n21772), .A2(n21690), .ZN(n18631) );
  NOR2_X2 U14577 ( .A1(n12744), .A2(n21719), .ZN(n21754) );
  NAND3_X1 U14578 ( .A1(n21754), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12737) );
  XNOR2_X1 U14579 ( .A(n12737), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n18701) );
  NOR3_X1 U14580 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n12569), .A3(
        n12570), .ZN(n12743) );
  NAND3_X1 U14581 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n21705), .ZN(n21718) );
  NOR2_X1 U14582 ( .A1(n21770), .A2(n21718), .ZN(n21722) );
  INV_X1 U14583 ( .A(n12744), .ZN(n21733) );
  AOI21_X1 U14584 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21555) );
  INV_X1 U14585 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12738) );
  NAND3_X1 U14586 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21580) );
  NOR2_X1 U14587 ( .A1(n12738), .A2(n21580), .ZN(n21601) );
  NAND3_X1 U14588 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n21601), .ZN(n21611) );
  NOR2_X1 U14589 ( .A1(n21555), .A2(n21611), .ZN(n21663) );
  INV_X1 U14590 ( .A(n21663), .ZN(n12739) );
  NOR3_X1 U14591 ( .A1(n21829), .A2(n18511), .A3(n12739), .ZN(n21827) );
  NAND2_X1 U14592 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21827), .ZN(
        n21516) );
  INV_X1 U14593 ( .A(n11246), .ZN(n21828) );
  NAND2_X1 U14594 ( .A1(n21499), .A2(n21892), .ZN(n21865) );
  NAND2_X1 U14595 ( .A1(n21876), .A2(n21615), .ZN(n21535) );
  NAND2_X1 U14596 ( .A1(n21828), .A2(n21535), .ZN(n21554) );
  NAND2_X1 U14597 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21553) );
  INV_X1 U14598 ( .A(n21553), .ZN(n21552) );
  AND2_X1 U14599 ( .A1(n21552), .A2(n21601), .ZN(n21877) );
  NAND3_X1 U14600 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n21877), .ZN(n21864) );
  NOR2_X1 U14601 ( .A1(n21829), .A2(n21864), .ZN(n21820) );
  NAND2_X1 U14602 ( .A1(n12742), .A2(n21820), .ZN(n21522) );
  OAI22_X1 U14603 ( .A1(n21826), .A2(n21516), .B1(n21554), .B2(n21522), .ZN(
        n21687) );
  AND4_X1 U14604 ( .A1(n21688), .A2(n21722), .A3(n21733), .A4(n21687), .ZN(
        n21738) );
  AOI22_X1 U14605 ( .A1(n21819), .A2(n18701), .B1(n12743), .B2(n21738), .ZN(
        n12751) );
  NOR2_X1 U14606 ( .A1(n12744), .A2(n12570), .ZN(n18706) );
  INV_X1 U14607 ( .A(n21718), .ZN(n12749) );
  AND2_X1 U14608 ( .A1(n21827), .A2(n12745), .ZN(n21691) );
  AOI21_X1 U14609 ( .B1(n12749), .B2(n21691), .A(n21826), .ZN(n21717) );
  NAND2_X1 U14610 ( .A1(n21820), .A2(n12745), .ZN(n12748) );
  INV_X1 U14611 ( .A(n12748), .ZN(n12747) );
  AOI21_X1 U14612 ( .B1(n12747), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n21875), .ZN(n21681) );
  AOI21_X1 U14613 ( .B1(n21865), .B2(n12748), .A(n21681), .ZN(n21775) );
  OAI221_X1 U14614 ( .B1(n11246), .B2(n12749), .C1(n11246), .C2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n21775), .ZN(n21735) );
  NOR2_X1 U14615 ( .A1(n21717), .A2(n21735), .ZN(n21752) );
  OAI211_X1 U14616 ( .C1(n21843), .C2(n18706), .A(n21752), .B(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21746) );
  NAND3_X1 U14617 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21788), .A3(
        n21746), .ZN(n12750) );
  OAI211_X1 U14618 ( .C1(n18704), .C2(n21792), .A(n12751), .B(n12750), .ZN(
        n12754) );
  NOR2_X1 U14619 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21939) );
  INV_X1 U14620 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n21262) );
  NOR2_X1 U14621 ( .A1(n21868), .A2(n21262), .ZN(n18699) );
  INV_X1 U14622 ( .A(n18699), .ZN(n12752) );
  OAI21_X1 U14623 ( .B1(n21773), .B2(n12574), .A(n12752), .ZN(n12753) );
  AND2_X4 U14624 ( .A1(n12757), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17054) );
  AOI22_X1 U14625 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12848), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12761) );
  AND2_X2 U14626 ( .A1(n17051), .A2(n12763), .ZN(n12994) );
  AND2_X2 U14627 ( .A1(n12763), .A2(n12765), .ZN(n12924) );
  AND2_X4 U14628 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17059) );
  AND2_X2 U14629 ( .A1(n17054), .A2(n17059), .ZN(n13241) );
  AOI22_X1 U14630 ( .A1(n13241), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12956), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12759) );
  NOR2_X4 U14631 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15430) );
  AOI22_X1 U14632 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12758) );
  NAND4_X1 U14633 ( .A1(n12761), .A2(n12760), .A3(n12759), .A4(n12758), .ZN(
        n12771) );
  AND2_X4 U14634 ( .A1(n17054), .A2(n12762), .ZN(n13018) );
  AND2_X2 U14635 ( .A1(n17054), .A2(n15430), .ZN(n12955) );
  AOI22_X1 U14636 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12955), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12769) );
  AND2_X2 U14637 ( .A1(n12762), .A2(n12765), .ZN(n12808) );
  AND2_X2 U14638 ( .A1(n12763), .A2(n15429), .ZN(n12818) );
  AOI22_X1 U14639 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12936), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12766) );
  NAND4_X1 U14640 ( .A1(n12769), .A2(n12768), .A3(n12767), .A4(n12766), .ZN(
        n12770) );
  OR2_X2 U14641 ( .A1(n12771), .A2(n12770), .ZN(n12885) );
  AOI22_X1 U14642 ( .A1(n12809), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12775) );
  AOI22_X1 U14643 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12848), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U14644 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12817), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U14645 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12955), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12772) );
  AOI22_X1 U14646 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12924), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12780) );
  BUF_X4 U14647 ( .A(n13241), .Z(n13566) );
  AOI22_X1 U14648 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U14649 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12956), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12777) );
  AOI22_X1 U14650 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12936), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12776) );
  AND2_X1 U14651 ( .A1(n12777), .A2(n12776), .ZN(n12778) );
  AND2_X2 U14653 ( .A1(n12885), .A2(n15583), .ZN(n12899) );
  NAND2_X1 U14654 ( .A1(n12955), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12785) );
  NAND2_X1 U14655 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12784) );
  NAND2_X1 U14656 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12783) );
  NAND3_X1 U14657 ( .A1(n12785), .A2(n12784), .A3(n12783), .ZN(n12786) );
  AOI21_X2 U14658 ( .B1(n12829), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n12786), .ZN(n12802) );
  NAND2_X1 U14659 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12790) );
  NAND2_X1 U14660 ( .A1(n12817), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12789) );
  NAND2_X1 U14661 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12788) );
  NAND2_X1 U14662 ( .A1(n12818), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12787) );
  NAND2_X1 U14663 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12794) );
  NAND2_X1 U14664 ( .A1(n12924), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12793) );
  NAND2_X1 U14665 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12792) );
  NAND2_X1 U14666 ( .A1(n12936), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12791) );
  NAND2_X1 U14667 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12798) );
  NAND2_X1 U14668 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12797) );
  NAND2_X1 U14669 ( .A1(n12956), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12796) );
  NAND2_X1 U14670 ( .A1(n17061), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12795) );
  AOI22_X1 U14671 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12924), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U14672 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12848), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12806) );
  AOI22_X1 U14673 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12817), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U14674 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12936), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12804) );
  NAND4_X1 U14675 ( .A1(n12807), .A2(n12806), .A3(n12805), .A4(n12804), .ZN(
        n12815) );
  AOI22_X1 U14676 ( .A1(n12809), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U14677 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12956), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U14678 ( .A1(n13241), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11175), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12810) );
  NAND4_X1 U14679 ( .A1(n12813), .A2(n12812), .A3(n12811), .A4(n12810), .ZN(
        n12814) );
  OR2_X2 U14680 ( .A1(n12815), .A2(n12814), .ZN(n12842) );
  INV_X1 U14681 ( .A(n12843), .ZN(n12816) );
  INV_X1 U14682 ( .A(n12902), .ZN(n12846) );
  AOI22_X1 U14683 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12955), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12822) );
  AOI22_X1 U14684 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12848), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U14685 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12817), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U14686 ( .A1(n12809), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12819) );
  NAND4_X1 U14687 ( .A1(n12822), .A2(n12821), .A3(n12820), .A4(n12819), .ZN(
        n12828) );
  AOI22_X1 U14688 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12936), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12826) );
  AOI22_X1 U14689 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12924), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12825) );
  AOI22_X1 U14690 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12956), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12824) );
  BUF_X4 U14691 ( .A(n13241), .Z(n13387) );
  NAND4_X1 U14692 ( .A1(n12826), .A2(n12825), .A3(n12824), .A4(n12823), .ZN(
        n12827) );
  INV_X2 U14693 ( .A(n15583), .ZN(n13052) );
  NAND2_X1 U14694 ( .A1(n13052), .A2(n12885), .ZN(n12838) );
  AOI22_X1 U14695 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12955), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U14696 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13260), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U14697 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12817), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12831) );
  AOI22_X1 U14698 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12818), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12830) );
  AOI22_X1 U14699 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12936), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U14700 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12924), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U14701 ( .A1(n13387), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12956), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U14702 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12834) );
  NAND2_X2 U14703 ( .A1(n11757), .A2(n11759), .ZN(n12883) );
  NAND2_X1 U14704 ( .A1(n12838), .A2(n15598), .ZN(n12841) );
  INV_X1 U14705 ( .A(n12894), .ZN(n12839) );
  AND2_X2 U14706 ( .A1(n12839), .A2(n12885), .ZN(n12847) );
  NAND2_X1 U14707 ( .A1(n12847), .A2(n12883), .ZN(n12840) );
  NAND2_X2 U14708 ( .A1(n13052), .A2(n12842), .ZN(n12884) );
  OAI211_X2 U14709 ( .C1(n12846), .C2(n15564), .A(n12845), .B(n12844), .ZN(
        n12890) );
  NAND2_X1 U14710 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12851) );
  NAND2_X1 U14711 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12850) );
  NAND2_X1 U14712 ( .A1(n12955), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12849) );
  NAND2_X1 U14713 ( .A1(n12817), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12854) );
  NAND2_X1 U14714 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12853) );
  NAND2_X1 U14715 ( .A1(n12818), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12852) );
  NAND2_X1 U14716 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12858) );
  NAND2_X1 U14717 ( .A1(n12924), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12857) );
  NAND2_X1 U14718 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12856) );
  NAND2_X1 U14719 ( .A1(n12936), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12855) );
  NAND2_X1 U14720 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12861) );
  NAND2_X1 U14721 ( .A1(n12956), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12860) );
  NAND2_X1 U14722 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12859) );
  NAND2_X1 U14723 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12866) );
  NAND2_X1 U14724 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12865) );
  NAND2_X1 U14725 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12864) );
  NAND2_X1 U14726 ( .A1(n12817), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12863) );
  NAND2_X1 U14727 ( .A1(n12924), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12870) );
  NAND2_X1 U14728 ( .A1(n13387), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12869) );
  NAND2_X1 U14729 ( .A1(n12956), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12868) );
  NAND2_X1 U14730 ( .A1(n17061), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12867) );
  AND4_X2 U14731 ( .A1(n12870), .A2(n12869), .A3(n12868), .A4(n12867), .ZN(
        n12881) );
  NAND2_X1 U14732 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12874) );
  NAND2_X1 U14733 ( .A1(n12994), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12873) );
  NAND2_X1 U14734 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12872) );
  NAND2_X1 U14735 ( .A1(n12936), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12871) );
  NAND2_X1 U14736 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12878) );
  NAND2_X1 U14737 ( .A1(n12955), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12877) );
  NAND2_X1 U14738 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12876) );
  NAND2_X1 U14739 ( .A1(n12818), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12875) );
  NOR2_X4 U14740 ( .A1(n12895), .A2(n12891), .ZN(n16376) );
  NAND3_X1 U14741 ( .A1(n17062), .A2(n16726), .A3(n16376), .ZN(n13660) );
  XNOR2_X1 U14742 ( .A(n22299), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n15168) );
  NAND2_X1 U14743 ( .A1(n12914), .A2(n15813), .ZN(n12905) );
  INV_X1 U14744 ( .A(n17062), .ZN(n15319) );
  NAND2_X1 U14745 ( .A1(n12892), .A2(n13052), .ZN(n12893) );
  NAND2_X1 U14746 ( .A1(n11745), .A2(n15570), .ZN(n12898) );
  NAND2_X1 U14747 ( .A1(n12898), .A2(n21956), .ZN(n12897) );
  INV_X1 U14748 ( .A(n16376), .ZN(n12915) );
  OAI21_X1 U14749 ( .B1(n15813), .B2(n12883), .A(n12915), .ZN(n12896) );
  INV_X1 U14750 ( .A(n12898), .ZN(n12901) );
  NAND2_X1 U14751 ( .A1(n15323), .A2(n17039), .ZN(n12903) );
  NAND4_X1 U14752 ( .A1(n12905), .A2(n12904), .A3(n11758), .A4(n12903), .ZN(
        n12906) );
  NAND2_X1 U14753 ( .A1(n12906), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12907) );
  NAND2_X1 U14754 ( .A1(n12982), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12910) );
  NAND2_X1 U14755 ( .A1(n17824), .A2(n22256), .ZN(n13687) );
  XNOR2_X1 U14756 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22445) );
  OR2_X1 U14757 ( .A1(n17865), .A2(n22476), .ZN(n12977) );
  OAI21_X1 U14758 ( .B1(n13687), .B2(n22445), .A(n12977), .ZN(n12908) );
  INV_X1 U14759 ( .A(n12908), .ZN(n12909) );
  NAND2_X1 U14760 ( .A1(n12910), .A2(n12909), .ZN(n12912) );
  MUX2_X1 U14761 ( .A(n13687), .B(n17865), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n12913) );
  NAND3_X1 U14762 ( .A1(n12900), .A2(n12915), .A3(n15384), .ZN(n12916) );
  NAND2_X1 U14763 ( .A1(n12914), .A2(n12916), .ZN(n12922) );
  NAND3_X1 U14764 ( .A1(n15323), .A2(n17039), .A3(n12891), .ZN(n12921) );
  NAND2_X1 U14765 ( .A1(n17062), .A2(n15583), .ZN(n12918) );
  NAND2_X1 U14766 ( .A1(n12917), .A2(n12918), .ZN(n15389) );
  NAND2_X1 U14767 ( .A1(n17824), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12919) );
  NOR2_X1 U14768 ( .A1(n15389), .A2(n12919), .ZN(n12920) );
  NAND4_X1 U14769 ( .A1(n12922), .A2(n11758), .A3(n12921), .A4(n12920), .ZN(
        n12953) );
  OR2_X2 U14770 ( .A1(n15609), .A2(n12923), .ZN(n12981) );
  INV_X1 U14771 ( .A(n12992), .ZN(n12973) );
  AOI22_X1 U14772 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13018), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12928) );
  AOI22_X1 U14773 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12927) );
  AOI22_X1 U14774 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12926) );
  AOI22_X1 U14775 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12925) );
  NAND4_X1 U14776 ( .A1(n12928), .A2(n12927), .A3(n12926), .A4(n12925), .ZN(
        n12934) );
  AOI22_X1 U14777 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13260), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12932) );
  AOI22_X1 U14778 ( .A1(n12809), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U14779 ( .A1(n13523), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12956), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12930) );
  AOI22_X1 U14780 ( .A1(n13387), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12929) );
  NAND4_X1 U14781 ( .A1(n12932), .A2(n12931), .A3(n12930), .A4(n12929), .ZN(
        n12933) );
  NAND2_X1 U14782 ( .A1(n12973), .A2(n13709), .ZN(n12935) );
  AOI22_X1 U14783 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U14784 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12939) );
  AOI22_X1 U14785 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U14786 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12937) );
  NAND4_X1 U14787 ( .A1(n12940), .A2(n12939), .A3(n12938), .A4(n12937), .ZN(
        n12946) );
  AOI22_X1 U14788 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12944) );
  AOI22_X1 U14789 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U14790 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12956), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U14791 ( .A1(n13387), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12941) );
  NAND4_X1 U14792 ( .A1(n12944), .A2(n12943), .A3(n12942), .A4(n12941), .ZN(
        n12945) );
  NAND2_X1 U14793 ( .A1(n13642), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12949) );
  INV_X1 U14794 ( .A(n12993), .ZN(n12947) );
  NAND2_X1 U14795 ( .A1(n12947), .A2(n13709), .ZN(n12948) );
  OAI211_X1 U14796 ( .C1(n12992), .C2(n13766), .A(n12949), .B(n12948), .ZN(
        n12950) );
  NAND2_X1 U14797 ( .A1(n13697), .A2(n12950), .ZN(n12951) );
  INV_X1 U14798 ( .A(n12953), .ZN(n12954) );
  AOI22_X1 U14799 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n13569), .B1(
        n12829), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12960) );
  BUF_X1 U14800 ( .A(n12808), .Z(n13549) );
  AOI22_X1 U14801 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n13549), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U14802 ( .A1(n13018), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12958) );
  AOI22_X1 U14803 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n13550), .B1(
        n12956), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12957) );
  NAND4_X1 U14804 ( .A1(n12960), .A2(n12959), .A3(n12958), .A4(n12957), .ZN(
        n12966) );
  AOI22_X1 U14805 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13566), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U14806 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n12809), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U14807 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12962) );
  AOI22_X1 U14808 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12961) );
  NAND4_X1 U14809 ( .A1(n12964), .A2(n12963), .A3(n12962), .A4(n12961), .ZN(
        n12965) );
  XNOR2_X1 U14810 ( .A(n13698), .B(n13766), .ZN(n12967) );
  NAND2_X1 U14811 ( .A1(n12967), .A2(n12973), .ZN(n12968) );
  INV_X1 U14812 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12972) );
  AOI21_X1 U14813 ( .B1(n15570), .B2(n13766), .A(n22256), .ZN(n12971) );
  NAND2_X1 U14814 ( .A1(n15813), .A2(n13708), .ZN(n12970) );
  NAND2_X1 U14815 ( .A1(n13081), .A2(n13080), .ZN(n12974) );
  NAND2_X1 U14816 ( .A1(n12973), .A2(n13766), .ZN(n13763) );
  NAND2_X1 U14817 ( .A1(n12974), .A2(n13763), .ZN(n13072) );
  INV_X1 U14818 ( .A(n13072), .ZN(n12975) );
  INV_X1 U14819 ( .A(n13061), .ZN(n13007) );
  INV_X1 U14820 ( .A(n12977), .ZN(n12979) );
  OAI21_X1 U14821 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n12979), .A(
        n12978), .ZN(n12980) );
  NAND2_X1 U14822 ( .A1(n12981), .A2(n12980), .ZN(n12990) );
  NAND2_X1 U14823 ( .A1(n12982), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12988) );
  NAND2_X1 U14824 ( .A1(n12983), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15611) );
  INV_X1 U14825 ( .A(n12983), .ZN(n12984) );
  NAND2_X1 U14826 ( .A1(n12984), .A2(n22408), .ZN(n12985) );
  NAND2_X1 U14827 ( .A1(n15611), .A2(n12985), .ZN(n15973) );
  OAI22_X1 U14828 ( .A1(n15973), .A2(n13687), .B1(n17865), .B2(n22408), .ZN(
        n12986) );
  INV_X1 U14829 ( .A(n12986), .ZN(n12987) );
  NAND2_X2 U14830 ( .A1(n12990), .A2(n12989), .ZN(n15875) );
  OR2_X2 U14831 ( .A1(n12990), .A2(n12989), .ZN(n12991) );
  OR2_X2 U14832 ( .A1(n16674), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U14833 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13018), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U14834 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U14835 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U14836 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12995) );
  NAND4_X1 U14837 ( .A1(n12998), .A2(n12997), .A3(n12996), .A4(n12995), .ZN(
        n13004) );
  AOI22_X1 U14838 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U14839 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13566), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U14840 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13000) );
  AOI22_X1 U14841 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12999) );
  NAND4_X1 U14842 ( .A1(n13002), .A2(n13001), .A3(n13000), .A4(n12999), .ZN(
        n13003) );
  AOI22_X1 U14843 ( .A1(n13640), .A2(n13707), .B1(n13642), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13005) );
  NAND2_X2 U14844 ( .A1(n13006), .A2(n13005), .ZN(n13060) );
  NAND2_X1 U14845 ( .A1(n12982), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13013) );
  INV_X1 U14846 ( .A(n15611), .ZN(n13008) );
  NAND2_X1 U14847 ( .A1(n13008), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15936) );
  NAND2_X1 U14848 ( .A1(n15611), .A2(n22409), .ZN(n13009) );
  INV_X1 U14849 ( .A(n13687), .ZN(n13011) );
  NOR2_X1 U14850 ( .A1(n17865), .A2(n22409), .ZN(n13010) );
  AOI21_X1 U14851 ( .B1(n22446), .B2(n13011), .A(n13010), .ZN(n13012) );
  XNOR2_X2 U14852 ( .A(n15875), .B(n15874), .ZN(n22384) );
  AOI22_X1 U14853 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13017) );
  AOI22_X1 U14854 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13016) );
  AOI22_X1 U14855 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13015) );
  AOI22_X1 U14856 ( .A1(n12809), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13014) );
  NAND4_X1 U14857 ( .A1(n13017), .A2(n13016), .A3(n13015), .A4(n13014), .ZN(
        n13024) );
  AOI22_X1 U14858 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13022) );
  AOI22_X1 U14859 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U14860 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13020) );
  AOI22_X1 U14861 ( .A1(n13387), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13019) );
  NAND4_X1 U14862 ( .A1(n13022), .A2(n13021), .A3(n13020), .A4(n13019), .ZN(
        n13023) );
  AOI22_X1 U14863 ( .A1(n13640), .A2(n13721), .B1(n13642), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13025) );
  INV_X1 U14864 ( .A(n13103), .ZN(n13039) );
  AOI22_X1 U14865 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13031) );
  AOI22_X1 U14866 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13030) );
  AOI22_X1 U14867 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13029) );
  AOI22_X1 U14868 ( .A1(n13387), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13028) );
  NAND4_X1 U14869 ( .A1(n13031), .A2(n13030), .A3(n13029), .A4(n13028), .ZN(
        n13037) );
  AOI22_X1 U14870 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13260), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13035) );
  AOI22_X1 U14871 ( .A1(n12809), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13034) );
  AOI22_X1 U14872 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13033) );
  AOI22_X1 U14873 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13032) );
  NAND4_X1 U14874 ( .A1(n13035), .A2(n13034), .A3(n13033), .A4(n13032), .ZN(
        n13036) );
  AOI22_X1 U14875 ( .A1(n13640), .A2(n13734), .B1(n13642), .B2(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13102) );
  AOI22_X1 U14876 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U14877 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U14878 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13041) );
  AOI22_X1 U14879 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13040) );
  NAND4_X1 U14880 ( .A1(n13043), .A2(n13042), .A3(n13041), .A4(n13040), .ZN(
        n13049) );
  AOI22_X1 U14881 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13047) );
  AOI22_X1 U14882 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U14883 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U14884 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13044) );
  NAND4_X1 U14885 ( .A1(n13047), .A2(n13046), .A3(n13045), .A4(n13044), .ZN(
        n13048) );
  AOI22_X1 U14886 ( .A1(n13640), .A2(n13737), .B1(n13642), .B2(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13050) );
  NAND2_X1 U14887 ( .A1(n13105), .A2(n13050), .ZN(n13051) );
  NAND2_X1 U14888 ( .A1(n11210), .A2(n13051), .ZN(n13740) );
  INV_X1 U14889 ( .A(n13106), .ZN(n13056) );
  INV_X1 U14890 ( .A(n13125), .ZN(n13055) );
  OAI21_X1 U14891 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n13056), .A(
        n13055), .ZN(n15890) );
  AOI22_X1 U14892 ( .A1(n13469), .A2(n15890), .B1(n13598), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13057) );
  INV_X1 U14893 ( .A(n13060), .ZN(n13062) );
  NAND2_X1 U14894 ( .A1(n13062), .A2(n13061), .ZN(n13063) );
  INV_X1 U14895 ( .A(n12884), .ZN(n13064) );
  INV_X1 U14896 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13067) );
  XNOR2_X1 U14897 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16677) );
  AOI21_X1 U14898 ( .B1(n13053), .B2(n16677), .A(n13598), .ZN(n13066) );
  OAI21_X1 U14899 ( .B1(n13065), .B2(n13067), .A(n13066), .ZN(n13068) );
  AOI21_X1 U14900 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13100), .A(
        n13068), .ZN(n13069) );
  OAI21_X2 U14901 ( .B1(n15435), .B2(n13250), .A(n13069), .ZN(n13070) );
  NAND2_X1 U14902 ( .A1(n13598), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13091) );
  NAND2_X1 U14903 ( .A1(n13070), .A2(n13091), .ZN(n15514) );
  INV_X1 U14904 ( .A(n15514), .ZN(n13090) );
  NAND2_X1 U14905 ( .A1(n13073), .A2(n13072), .ZN(n13074) );
  NAND2_X1 U14906 ( .A1(n16347), .A2(n13265), .ZN(n13079) );
  INV_X1 U14907 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n13076) );
  INV_X1 U14908 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13075) );
  OAI22_X1 U14909 ( .A1(n13065), .A2(n13076), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13075), .ZN(n13077) );
  AOI21_X1 U14910 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13100), .A(
        n13077), .ZN(n13078) );
  NAND2_X1 U14911 ( .A1(n13696), .A2(n15583), .ZN(n13082) );
  NAND2_X1 U14912 ( .A1(n13082), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15178) );
  INV_X1 U14913 ( .A(n13100), .ZN(n13110) );
  INV_X1 U14914 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15353) );
  NAND2_X1 U14915 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13085) );
  NAND2_X1 U14916 ( .A1(n13599), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n13084) );
  OAI211_X1 U14917 ( .C1(n13110), .C2(n15353), .A(n13085), .B(n13084), .ZN(
        n13086) );
  AOI21_X1 U14918 ( .B1(n13083), .B2(n13265), .A(n13086), .ZN(n13087) );
  OR2_X1 U14919 ( .A1(n15178), .A2(n13087), .ZN(n15179) );
  INV_X1 U14920 ( .A(n13087), .ZN(n15180) );
  OR2_X1 U14921 ( .A1(n15180), .A2(n13589), .ZN(n13088) );
  NAND2_X1 U14922 ( .A1(n15179), .A2(n13088), .ZN(n15442) );
  NAND2_X1 U14923 ( .A1(n15444), .A2(n15442), .ZN(n15513) );
  INV_X1 U14924 ( .A(n15513), .ZN(n13089) );
  NAND2_X1 U14925 ( .A1(n13090), .A2(n13089), .ZN(n15511) );
  INV_X1 U14926 ( .A(n15539), .ZN(n15506) );
  INV_X1 U14927 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n13098) );
  INV_X1 U14928 ( .A(n13094), .ZN(n13096) );
  INV_X1 U14929 ( .A(n13107), .ZN(n13095) );
  OAI21_X1 U14930 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13096), .A(
        n13095), .ZN(n15827) );
  AOI22_X1 U14931 ( .A1(n13469), .A2(n15827), .B1(n13598), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13097) );
  OAI21_X1 U14932 ( .B1(n13065), .B2(n13098), .A(n13097), .ZN(n13099) );
  AOI21_X1 U14933 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13100), .A(
        n13099), .ZN(n13101) );
  NAND2_X1 U14934 ( .A1(n15607), .A2(n15606), .ZN(n15605) );
  NAND2_X1 U14935 ( .A1(n13103), .A2(n13102), .ZN(n13104) );
  NAND2_X1 U14936 ( .A1(n13105), .A2(n13104), .ZN(n13727) );
  INV_X1 U14937 ( .A(n13727), .ZN(n13114) );
  OAI21_X1 U14938 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13107), .A(
        n13106), .ZN(n15866) );
  INV_X1 U14939 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n22268) );
  OAI21_X1 U14940 ( .B1(n22268), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n22489), .ZN(n13109) );
  NAND2_X1 U14941 ( .A1(n13599), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n13108) );
  OAI211_X1 U14942 ( .C1(n13110), .C2(n17889), .A(n13109), .B(n13108), .ZN(
        n13111) );
  OAI21_X1 U14943 ( .B1(n13589), .B2(n15866), .A(n13111), .ZN(n13112) );
  AOI21_X1 U14944 ( .B1(n13114), .B2(n13265), .A(n13113), .ZN(n15767) );
  NOR2_X2 U14945 ( .A1(n15605), .A2(n15767), .ZN(n15766) );
  AOI22_X1 U14946 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13118) );
  AOI22_X1 U14947 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13117) );
  AOI22_X1 U14948 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U14949 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13115) );
  NAND4_X1 U14950 ( .A1(n13118), .A2(n13117), .A3(n13116), .A4(n13115), .ZN(
        n13124) );
  AOI22_X1 U14951 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U14952 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13121) );
  AOI22_X1 U14953 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U14954 ( .A1(n13387), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13119) );
  NAND4_X1 U14955 ( .A1(n13122), .A2(n13121), .A3(n13120), .A4(n13119), .ZN(
        n13123) );
  AOI22_X1 U14956 ( .A1(n13640), .A2(n13754), .B1(n13642), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13131) );
  NAND2_X1 U14957 ( .A1(n13744), .A2(n13265), .ZN(n13130) );
  INV_X1 U14958 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13127) );
  OAI21_X1 U14959 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13125), .A(
        n13136), .ZN(n22141) );
  AOI22_X1 U14960 ( .A1(n13469), .A2(n22141), .B1(n13598), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13126) );
  OAI21_X1 U14961 ( .B1(n13065), .B2(n13127), .A(n13126), .ZN(n13128) );
  INV_X1 U14962 ( .A(n13128), .ZN(n13129) );
  NAND2_X1 U14963 ( .A1(n15836), .A2(n15861), .ZN(n15862) );
  INV_X1 U14964 ( .A(n13131), .ZN(n13132) );
  INV_X1 U14965 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13134) );
  NAND2_X1 U14966 ( .A1(n13640), .A2(n13766), .ZN(n13133) );
  OAI21_X1 U14967 ( .B1(n13134), .B2(n13624), .A(n13133), .ZN(n13135) );
  INV_X1 U14968 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13140) );
  INV_X1 U14969 ( .A(n13136), .ZN(n13138) );
  INV_X1 U14970 ( .A(n13156), .ZN(n13137) );
  OAI21_X1 U14971 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13138), .A(
        n13137), .ZN(n22148) );
  AOI22_X1 U14972 ( .A1(n13469), .A2(n22148), .B1(n13598), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13139) );
  OAI21_X1 U14973 ( .B1(n13065), .B2(n13140), .A(n13139), .ZN(n13141) );
  AOI21_X1 U14974 ( .B1(n13752), .B2(n13265), .A(n13141), .ZN(n16046) );
  INV_X1 U14975 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n16199) );
  XNOR2_X1 U14976 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n13156), .ZN(
        n22166) );
  AOI22_X1 U14977 ( .A1(n13469), .A2(n22166), .B1(n13598), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13142) );
  OAI21_X1 U14978 ( .B1(n13065), .B2(n16199), .A(n13142), .ZN(n13155) );
  AOI22_X1 U14979 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13575), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13146) );
  AOI22_X1 U14980 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13145) );
  AOI22_X1 U14981 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n13578), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13144) );
  AOI22_X1 U14982 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n11168), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13143) );
  NAND4_X1 U14983 ( .A1(n13146), .A2(n13145), .A3(n13144), .A4(n13143), .ZN(
        n13152) );
  AOI22_X1 U14984 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n13549), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13150) );
  AOI22_X1 U14985 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13149) );
  AOI22_X1 U14986 ( .A1(n13387), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13148) );
  AOI22_X1 U14987 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13147) );
  NAND4_X1 U14988 ( .A1(n13150), .A2(n13149), .A3(n13148), .A4(n13147), .ZN(
        n13151) );
  NOR2_X1 U14989 ( .A1(n13152), .A2(n13151), .ZN(n13153) );
  NOR2_X1 U14990 ( .A1(n13250), .A2(n13153), .ZN(n13154) );
  NOR2_X1 U14991 ( .A1(n13155), .A2(n13154), .ZN(n16190) );
  XNOR2_X1 U14992 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n13171), .ZN(
        n16263) );
  INV_X1 U14993 ( .A(n16263), .ZN(n22178) );
  AOI22_X1 U14994 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13160) );
  AOI22_X1 U14995 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13159) );
  AOI22_X1 U14996 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13158) );
  AOI22_X1 U14997 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13157) );
  NAND4_X1 U14998 ( .A1(n13160), .A2(n13159), .A3(n13158), .A4(n13157), .ZN(
        n13166) );
  AOI22_X1 U14999 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13543), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13164) );
  AOI22_X1 U15000 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13549), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13163) );
  AOI22_X1 U15001 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13162) );
  AOI22_X1 U15002 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13161) );
  NAND4_X1 U15003 ( .A1(n13164), .A2(n13163), .A3(n13162), .A4(n13161), .ZN(
        n13165) );
  OAI21_X1 U15004 ( .B1(n13166), .B2(n13165), .A(n13265), .ZN(n13169) );
  NAND2_X1 U15005 ( .A1(n13599), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13168) );
  NAND2_X1 U15006 ( .A1(n13598), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13167) );
  NAND3_X1 U15007 ( .A1(n13169), .A2(n13168), .A3(n13167), .ZN(n13170) );
  XNOR2_X1 U15008 ( .A(n13188), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n20650) );
  NAND2_X1 U15009 ( .A1(n20650), .A2(n13469), .ZN(n13187) );
  INV_X1 U15010 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n16271) );
  INV_X1 U15011 ( .A(n13598), .ZN(n13248) );
  INV_X1 U15012 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13172) );
  OAI22_X1 U15013 ( .A1(n13065), .A2(n16271), .B1(n13248), .B2(n13172), .ZN(
        n13185) );
  AOI22_X1 U15014 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13549), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13176) );
  AOI22_X1 U15015 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U15016 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13174) );
  AOI22_X1 U15017 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13173) );
  NAND4_X1 U15018 ( .A1(n13176), .A2(n13175), .A3(n13174), .A4(n13173), .ZN(
        n13182) );
  AOI22_X1 U15019 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13543), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U15020 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13179) );
  AOI22_X1 U15021 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13178) );
  AOI22_X1 U15022 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13177) );
  NAND4_X1 U15023 ( .A1(n13180), .A2(n13179), .A3(n13178), .A4(n13177), .ZN(
        n13181) );
  NOR2_X1 U15024 ( .A1(n13182), .A2(n13181), .ZN(n13183) );
  NOR2_X1 U15025 ( .A1(n13250), .A2(n13183), .ZN(n13184) );
  NOR2_X1 U15026 ( .A1(n13185), .A2(n13184), .ZN(n13186) );
  NAND2_X1 U15027 ( .A1(n13187), .A2(n13186), .ZN(n16269) );
  INV_X1 U15028 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n16279) );
  OAI21_X1 U15029 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13189), .A(
        n13230), .ZN(n22209) );
  AOI22_X1 U15030 ( .A1(n13469), .A2(n22209), .B1(n13598), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13190) );
  OAI21_X1 U15031 ( .B1(n13065), .B2(n16279), .A(n13190), .ZN(n13191) );
  INV_X1 U15032 ( .A(n13191), .ZN(n16274) );
  AOI22_X1 U15033 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13543), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13195) );
  AOI22_X1 U15034 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13194) );
  AOI22_X1 U15035 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13193) );
  AOI22_X1 U15036 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13192) );
  NAND4_X1 U15037 ( .A1(n13195), .A2(n13194), .A3(n13193), .A4(n13192), .ZN(
        n13201) );
  AOI22_X1 U15038 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U15039 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13198) );
  AOI22_X1 U15040 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13197) );
  AOI22_X1 U15041 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13196) );
  NAND4_X1 U15042 ( .A1(n13199), .A2(n13198), .A3(n13197), .A4(n13196), .ZN(
        n13200) );
  OR2_X1 U15043 ( .A1(n13201), .A2(n13200), .ZN(n13202) );
  NAND2_X1 U15044 ( .A1(n13265), .A2(n13202), .ZN(n16291) );
  XNOR2_X1 U15045 ( .A(n13236), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16912) );
  NAND2_X1 U15046 ( .A1(n16912), .A2(n13469), .ZN(n13219) );
  INV_X1 U15047 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n16790) );
  INV_X1 U15048 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16665) );
  OAI22_X1 U15049 ( .A1(n13065), .A2(n16790), .B1(n13248), .B2(n16665), .ZN(
        n13217) );
  AOI22_X1 U15050 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13208) );
  AOI22_X1 U15051 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13207) );
  AOI22_X1 U15052 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13549), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13206) );
  AOI22_X1 U15053 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13205) );
  NAND4_X1 U15054 ( .A1(n13208), .A2(n13207), .A3(n13206), .A4(n13205), .ZN(
        n13214) );
  AOI22_X1 U15055 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13566), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13212) );
  AOI22_X1 U15056 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13211) );
  AOI22_X1 U15057 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13210) );
  AOI22_X1 U15058 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13209) );
  NAND4_X1 U15059 ( .A1(n13212), .A2(n13211), .A3(n13210), .A4(n13209), .ZN(
        n13213) );
  NOR2_X1 U15060 ( .A1(n13214), .A2(n13213), .ZN(n13215) );
  NOR2_X1 U15061 ( .A1(n13250), .A2(n13215), .ZN(n13216) );
  NOR2_X1 U15062 ( .A1(n13217), .A2(n13216), .ZN(n13218) );
  NAND2_X1 U15063 ( .A1(n13219), .A2(n13218), .ZN(n16660) );
  AOI22_X1 U15064 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13223) );
  AOI22_X1 U15065 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13222) );
  AOI22_X1 U15066 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13221) );
  AOI22_X1 U15067 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13220) );
  NAND4_X1 U15068 ( .A1(n13223), .A2(n13222), .A3(n13221), .A4(n13220), .ZN(
        n13229) );
  AOI22_X1 U15069 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U15070 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13226) );
  AOI22_X1 U15071 ( .A1(n13387), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13225) );
  AOI22_X1 U15072 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13224) );
  NAND4_X1 U15073 ( .A1(n13227), .A2(n13226), .A3(n13225), .A4(n13224), .ZN(
        n13228) );
  NOR2_X1 U15074 ( .A1(n13229), .A2(n13228), .ZN(n13234) );
  NAND2_X1 U15075 ( .A1(n13599), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n13233) );
  XNOR2_X1 U15076 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n13230), .ZN(
        n22217) );
  OAI22_X1 U15077 ( .A1(n22217), .A2(n13589), .B1(n13248), .B2(n13204), .ZN(
        n13231) );
  INV_X1 U15078 ( .A(n13231), .ZN(n13232) );
  OAI211_X1 U15079 ( .C1(n13234), .C2(n13250), .A(n13233), .B(n13232), .ZN(
        n16293) );
  NAND2_X1 U15080 ( .A1(n16660), .A2(n16293), .ZN(n13235) );
  XOR2_X1 U15081 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n13254), .Z(
        n20675) );
  AOI22_X1 U15082 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13240) );
  AOI22_X1 U15083 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13549), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13239) );
  AOI22_X1 U15084 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13238) );
  AOI22_X1 U15085 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13237) );
  NAND4_X1 U15086 ( .A1(n13240), .A2(n13239), .A3(n13238), .A4(n13237), .ZN(
        n13247) );
  AOI22_X1 U15087 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13245) );
  AOI22_X1 U15088 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U15089 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U15090 ( .A1(n13543), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13242) );
  NAND4_X1 U15091 ( .A1(n13245), .A2(n13244), .A3(n13243), .A4(n13242), .ZN(
        n13246) );
  NOR2_X1 U15092 ( .A1(n13247), .A2(n13246), .ZN(n13249) );
  INV_X1 U15093 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16653) );
  OAI22_X1 U15094 ( .A1(n13250), .A2(n13249), .B1(n13248), .B2(n16653), .ZN(
        n13252) );
  INV_X1 U15095 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n16786) );
  NOR2_X1 U15096 ( .A1(n13065), .A2(n16786), .ZN(n13251) );
  NOR2_X1 U15097 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  OAI21_X1 U15098 ( .B1(n20675), .B2(n13589), .A(n13253), .ZN(n16648) );
  NAND2_X1 U15099 ( .A1(n16647), .A2(n16648), .ZN(n16636) );
  INV_X1 U15100 ( .A(n16636), .ZN(n13273) );
  INV_X1 U15101 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n13255) );
  XNOR2_X1 U15102 ( .A(n13274), .B(n13255), .ZN(n16900) );
  AOI22_X1 U15103 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13259) );
  AOI22_X1 U15104 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13258) );
  AOI22_X1 U15105 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13257) );
  AOI22_X1 U15106 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13256) );
  NAND4_X1 U15107 ( .A1(n13259), .A2(n13258), .A3(n13257), .A4(n13256), .ZN(
        n13267) );
  AOI22_X1 U15108 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13260), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13264) );
  AOI22_X1 U15109 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13263) );
  AOI22_X1 U15110 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13262) );
  AOI22_X1 U15111 ( .A1(n13543), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13261) );
  NAND4_X1 U15112 ( .A1(n13264), .A2(n13263), .A3(n13262), .A4(n13261), .ZN(
        n13266) );
  OAI21_X1 U15113 ( .B1(n13267), .B2(n13266), .A(n13265), .ZN(n13270) );
  NAND2_X1 U15114 ( .A1(n13599), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13269) );
  NAND2_X1 U15115 ( .A1(n13598), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13268) );
  NAND3_X1 U15116 ( .A1(n13270), .A2(n13269), .A3(n13268), .ZN(n13271) );
  AOI21_X1 U15117 ( .B1(n16900), .B2(n13469), .A(n13271), .ZN(n16637) );
  OR2_X1 U15118 ( .A1(n13275), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13276) );
  NAND2_X1 U15119 ( .A1(n13276), .A2(n13322), .ZN(n22245) );
  AOI22_X1 U15120 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13569), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13280) );
  AOI22_X1 U15121 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n13518), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13279) );
  AOI22_X1 U15122 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13278) );
  AOI22_X1 U15123 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n13550), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13277) );
  NAND4_X1 U15124 ( .A1(n13280), .A2(n13279), .A3(n13278), .A4(n13277), .ZN(
        n13286) );
  AOI22_X1 U15125 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13566), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13284) );
  AOI22_X1 U15126 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n13549), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13283) );
  AOI22_X1 U15127 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U15128 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13281) );
  NAND4_X1 U15129 ( .A1(n13284), .A2(n13283), .A3(n13282), .A4(n13281), .ZN(
        n13285) );
  OAI21_X1 U15130 ( .B1(n13286), .B2(n13285), .A(n13561), .ZN(n13289) );
  NAND2_X1 U15131 ( .A1(n13599), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n13288) );
  NAND2_X1 U15132 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13287) );
  NAND4_X1 U15133 ( .A1(n13289), .A2(n13589), .A3(n13288), .A4(n13287), .ZN(
        n13290) );
  AOI22_X1 U15134 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13574), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13294) );
  AOI22_X1 U15135 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13293) );
  AOI22_X1 U15136 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13292) );
  AOI22_X1 U15137 ( .A1(n13543), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13291) );
  NAND4_X1 U15138 ( .A1(n13294), .A2(n13293), .A3(n13292), .A4(n13291), .ZN(
        n13300) );
  AOI22_X1 U15139 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13298) );
  AOI22_X1 U15140 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13297) );
  AOI22_X1 U15141 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13296) );
  AOI22_X1 U15142 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13295) );
  NAND4_X1 U15143 ( .A1(n13298), .A2(n13297), .A3(n13296), .A4(n13295), .ZN(
        n13299) );
  OR2_X1 U15144 ( .A1(n13300), .A2(n13299), .ZN(n13301) );
  NAND2_X1 U15145 ( .A1(n13561), .A2(n13301), .ZN(n13307) );
  INV_X1 U15146 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13304) );
  INV_X1 U15147 ( .A(n13322), .ZN(n13302) );
  XNOR2_X1 U15148 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n13302), .ZN(
        n16890) );
  AOI22_X1 U15149 ( .A1(n13469), .A2(n16890), .B1(n13598), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13303) );
  OAI21_X1 U15150 ( .B1(n13065), .B2(n13304), .A(n13303), .ZN(n13305) );
  INV_X1 U15151 ( .A(n13305), .ZN(n13306) );
  NAND2_X1 U15152 ( .A1(n13307), .A2(n13306), .ZN(n16619) );
  AOI22_X1 U15153 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13311) );
  AOI22_X1 U15154 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13518), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13310) );
  AOI22_X1 U15155 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13309) );
  AOI22_X1 U15156 ( .A1(n13543), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13308) );
  NAND4_X1 U15157 ( .A1(n13311), .A2(n13310), .A3(n13309), .A4(n13308), .ZN(
        n13317) );
  AOI22_X1 U15158 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13315) );
  AOI22_X1 U15159 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13314) );
  AOI22_X1 U15160 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13313) );
  AOI22_X1 U15161 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13312) );
  NAND4_X1 U15162 ( .A1(n13315), .A2(n13314), .A3(n13313), .A4(n13312), .ZN(
        n13316) );
  NOR2_X1 U15163 ( .A1(n13317), .A2(n13316), .ZN(n13320) );
  OAI21_X1 U15164 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n22268), .A(
        n22489), .ZN(n13319) );
  NAND2_X1 U15165 ( .A1(n13599), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n13318) );
  OAI211_X1 U15166 ( .C1(n13593), .C2(n13320), .A(n13319), .B(n13318), .ZN(
        n13325) );
  OAI21_X1 U15167 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n13323), .A(
        n13357), .ZN(n16879) );
  OR2_X1 U15168 ( .A1(n13589), .A2(n16879), .ZN(n13324) );
  AOI22_X1 U15169 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13329) );
  AOI22_X1 U15170 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13328) );
  AOI22_X1 U15171 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13327) );
  AOI22_X1 U15172 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13326) );
  NAND4_X1 U15173 ( .A1(n13329), .A2(n13328), .A3(n13327), .A4(n13326), .ZN(
        n13335) );
  AOI22_X1 U15174 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13543), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13333) );
  AOI22_X1 U15175 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U15176 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13331) );
  AOI22_X1 U15177 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13330) );
  NAND4_X1 U15178 ( .A1(n13333), .A2(n13332), .A3(n13331), .A4(n13330), .ZN(
        n13334) );
  NOR2_X1 U15179 ( .A1(n13335), .A2(n13334), .ZN(n13339) );
  INV_X1 U15180 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15241) );
  NAND2_X1 U15181 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13336) );
  OAI211_X1 U15182 ( .C1(n13065), .C2(n15241), .A(n13589), .B(n13336), .ZN(
        n13337) );
  INV_X1 U15183 ( .A(n13337), .ZN(n13338) );
  OAI21_X1 U15184 ( .B1(n13593), .B2(n13339), .A(n13338), .ZN(n13341) );
  XNOR2_X1 U15185 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n13357), .ZN(
        n16869) );
  NAND2_X1 U15186 ( .A1(n13053), .A2(n16869), .ZN(n13340) );
  NAND2_X1 U15187 ( .A1(n13341), .A2(n13340), .ZN(n16594) );
  AOI22_X1 U15188 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13345) );
  AOI22_X1 U15189 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13344) );
  AOI22_X1 U15190 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13343) );
  AOI22_X1 U15191 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13342) );
  NAND4_X1 U15192 ( .A1(n13345), .A2(n13344), .A3(n13343), .A4(n13342), .ZN(
        n13351) );
  AOI22_X1 U15193 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13349) );
  AOI22_X1 U15194 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U15195 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13347) );
  AOI22_X1 U15196 ( .A1(n13543), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13346) );
  NAND4_X1 U15197 ( .A1(n13349), .A2(n13348), .A3(n13347), .A4(n13346), .ZN(
        n13350) );
  NOR2_X1 U15198 ( .A1(n13351), .A2(n13350), .ZN(n13355) );
  INV_X1 U15199 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n15483) );
  NAND2_X1 U15200 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13352) );
  OAI211_X1 U15201 ( .C1(n13065), .C2(n15483), .A(n13589), .B(n13352), .ZN(
        n13353) );
  INV_X1 U15202 ( .A(n13353), .ZN(n13354) );
  OAI21_X1 U15203 ( .B1(n13593), .B2(n13355), .A(n13354), .ZN(n13360) );
  OAI21_X1 U15204 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n13358), .A(
        n13379), .ZN(n20693) );
  OR2_X1 U15205 ( .A1(n13589), .A2(n20693), .ZN(n13359) );
  NAND2_X1 U15206 ( .A1(n13360), .A2(n13359), .ZN(n16580) );
  NAND2_X1 U15207 ( .A1(n16578), .A2(n13361), .ZN(n16566) );
  AOI22_X1 U15208 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13365) );
  AOI22_X1 U15209 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13364) );
  AOI22_X1 U15210 ( .A1(n13568), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13363) );
  AOI22_X1 U15211 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13362) );
  NAND4_X1 U15212 ( .A1(n13365), .A2(n13364), .A3(n13363), .A4(n13362), .ZN(
        n13371) );
  AOI22_X1 U15213 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13543), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13369) );
  AOI22_X1 U15214 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13368) );
  AOI22_X1 U15215 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13367) );
  AOI22_X1 U15216 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13366) );
  NAND4_X1 U15217 ( .A1(n13369), .A2(n13368), .A3(n13367), .A4(n13366), .ZN(
        n13370) );
  NOR2_X1 U15218 ( .A1(n13371), .A2(n13370), .ZN(n13375) );
  INV_X1 U15219 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15175) );
  NAND2_X1 U15220 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13372) );
  OAI211_X1 U15221 ( .C1(n13065), .C2(n15175), .A(n13589), .B(n13372), .ZN(
        n13373) );
  INV_X1 U15222 ( .A(n13373), .ZN(n13374) );
  OAI21_X1 U15223 ( .B1(n13593), .B2(n13375), .A(n13374), .ZN(n13377) );
  XNOR2_X1 U15224 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n13379), .ZN(
        n16861) );
  NAND2_X1 U15225 ( .A1(n13053), .A2(n16861), .ZN(n13376) );
  NAND2_X1 U15226 ( .A1(n13377), .A2(n13376), .ZN(n16568) );
  INV_X1 U15227 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n13378) );
  OR2_X1 U15228 ( .A1(n13380), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13381) );
  NAND2_X1 U15229 ( .A1(n13381), .A2(n13444), .ZN(n20702) );
  AOI22_X1 U15230 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13386) );
  AOI22_X1 U15231 ( .A1(n12829), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13569), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13385) );
  AOI22_X1 U15232 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13549), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13384) );
  AOI22_X1 U15233 ( .A1(n12803), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13383) );
  NAND4_X1 U15234 ( .A1(n13386), .A2(n13385), .A3(n13384), .A4(n13383), .ZN(
        n13393) );
  AOI22_X1 U15235 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13391) );
  AOI22_X1 U15236 ( .A1(n13568), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13390) );
  AOI22_X1 U15237 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13389) );
  AOI22_X1 U15238 ( .A1(n13387), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13388) );
  NAND4_X1 U15239 ( .A1(n13391), .A2(n13390), .A3(n13389), .A4(n13388), .ZN(
        n13392) );
  NOR2_X1 U15240 ( .A1(n13393), .A2(n13392), .ZN(n13396) );
  OAI21_X1 U15241 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n22268), .A(
        n22489), .ZN(n13395) );
  NAND2_X1 U15242 ( .A1(n13599), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n13394) );
  OAI211_X1 U15243 ( .C1(n13593), .C2(n13396), .A(n13395), .B(n13394), .ZN(
        n13397) );
  OAI21_X1 U15244 ( .B1(n20702), .B2(n13589), .A(n13397), .ZN(n13398) );
  INV_X1 U15245 ( .A(n13398), .ZN(n16548) );
  AOI22_X1 U15246 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13566), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U15247 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12829), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13401) );
  AOI22_X1 U15248 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n12818), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13400) );
  AOI22_X1 U15249 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13399) );
  NAND4_X1 U15250 ( .A1(n13402), .A2(n13401), .A3(n13400), .A4(n13399), .ZN(
        n13408) );
  AOI22_X1 U15251 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13406) );
  AOI22_X1 U15252 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n13518), .B1(
        n13549), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13405) );
  AOI22_X1 U15253 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13404) );
  AOI22_X1 U15254 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n13569), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13403) );
  NAND4_X1 U15255 ( .A1(n13406), .A2(n13405), .A3(n13404), .A4(n13403), .ZN(
        n13407) );
  NOR2_X1 U15256 ( .A1(n13408), .A2(n13407), .ZN(n13428) );
  AOI22_X1 U15257 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13412) );
  AOI22_X1 U15258 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13411) );
  AOI22_X1 U15259 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13410) );
  AOI22_X1 U15260 ( .A1(n13543), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13409) );
  NAND4_X1 U15261 ( .A1(n13412), .A2(n13411), .A3(n13410), .A4(n13409), .ZN(
        n13419) );
  AOI22_X1 U15262 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12829), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U15263 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13416) );
  AOI22_X1 U15264 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U15265 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13414) );
  NAND4_X1 U15266 ( .A1(n13417), .A2(n13416), .A3(n13415), .A4(n13414), .ZN(
        n13418) );
  NOR2_X1 U15267 ( .A1(n13419), .A2(n13418), .ZN(n13427) );
  XOR2_X1 U15268 ( .A(n13428), .B(n13427), .Z(n13420) );
  NAND2_X1 U15269 ( .A1(n13420), .A2(n13561), .ZN(n13425) );
  INV_X1 U15270 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n15250) );
  NAND2_X1 U15271 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13421) );
  OAI211_X1 U15272 ( .C1(n13065), .C2(n15250), .A(n13589), .B(n13421), .ZN(
        n13422) );
  INV_X1 U15273 ( .A(n13422), .ZN(n13424) );
  XNOR2_X1 U15274 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n13444), .ZN(
        n16855) );
  AOI21_X1 U15275 ( .B1(n13425), .B2(n13424), .A(n13423), .ZN(n16537) );
  NOR2_X1 U15276 ( .A1(n13428), .A2(n13427), .ZN(n13463) );
  AOI22_X1 U15277 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13432) );
  AOI22_X1 U15278 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13431) );
  AOI22_X1 U15279 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U15280 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13429) );
  NAND4_X1 U15281 ( .A1(n13432), .A2(n13431), .A3(n13430), .A4(n13429), .ZN(
        n13438) );
  AOI22_X1 U15282 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13436) );
  AOI22_X1 U15283 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U15284 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13434) );
  AOI22_X1 U15285 ( .A1(n13543), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13433) );
  NAND4_X1 U15286 ( .A1(n13436), .A2(n13435), .A3(n13434), .A4(n13433), .ZN(
        n13437) );
  OR2_X1 U15287 ( .A1(n13438), .A2(n13437), .ZN(n13462) );
  INV_X1 U15288 ( .A(n13462), .ZN(n13439) );
  XNOR2_X1 U15289 ( .A(n13463), .B(n13439), .ZN(n13440) );
  NAND2_X1 U15290 ( .A1(n13440), .A2(n13561), .ZN(n13451) );
  INV_X1 U15291 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13442) );
  NAND2_X1 U15292 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13441) );
  OAI211_X1 U15293 ( .C1(n13065), .C2(n13442), .A(n13589), .B(n13441), .ZN(
        n13443) );
  INV_X1 U15294 ( .A(n13443), .ZN(n13450) );
  INV_X1 U15295 ( .A(n13446), .ZN(n13447) );
  INV_X1 U15296 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16526) );
  NAND2_X1 U15297 ( .A1(n13447), .A2(n16526), .ZN(n13448) );
  NAND2_X1 U15298 ( .A1(n13491), .A2(n13448), .ZN(n16845) );
  NOR2_X1 U15299 ( .A1(n16845), .A2(n13589), .ZN(n13449) );
  AOI21_X1 U15300 ( .B1(n13451), .B2(n13450), .A(n13449), .ZN(n16525) );
  AOI22_X1 U15301 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12808), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13455) );
  AOI22_X1 U15302 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13413), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13454) );
  AOI22_X1 U15303 ( .A1(n13543), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13453) );
  AOI22_X1 U15304 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13452) );
  NAND4_X1 U15305 ( .A1(n13455), .A2(n13454), .A3(n13453), .A4(n13452), .ZN(
        n13461) );
  AOI22_X1 U15306 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13459) );
  AOI22_X1 U15307 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13458) );
  AOI22_X1 U15308 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U15309 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13456) );
  NAND4_X1 U15310 ( .A1(n13459), .A2(n13458), .A3(n13457), .A4(n13456), .ZN(
        n13460) );
  NOR2_X1 U15311 ( .A1(n13461), .A2(n13460), .ZN(n13475) );
  NAND2_X1 U15312 ( .A1(n13463), .A2(n13462), .ZN(n13474) );
  XOR2_X1 U15313 ( .A(n13475), .B(n13474), .Z(n13467) );
  INV_X1 U15314 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13465) );
  NAND2_X1 U15315 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13464) );
  OAI211_X1 U15316 ( .C1(n13065), .C2(n13465), .A(n13589), .B(n13464), .ZN(
        n13466) );
  AOI21_X1 U15317 ( .B1(n13467), .B2(n13561), .A(n13466), .ZN(n13468) );
  INV_X1 U15318 ( .A(n13468), .ZN(n13471) );
  XNOR2_X1 U15319 ( .A(n13491), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16835) );
  NAND2_X1 U15320 ( .A1(n16835), .A2(n13469), .ZN(n13470) );
  NAND2_X1 U15321 ( .A1(n13471), .A2(n13470), .ZN(n16513) );
  NAND2_X1 U15322 ( .A1(n13473), .A2(n13472), .ZN(n16497) );
  NOR2_X1 U15323 ( .A1(n13475), .A2(n13474), .ZN(n13508) );
  AOI22_X1 U15324 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13479) );
  AOI22_X1 U15325 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13478) );
  AOI22_X1 U15326 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13477) );
  AOI22_X1 U15327 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13476) );
  NAND4_X1 U15328 ( .A1(n13479), .A2(n13478), .A3(n13477), .A4(n13476), .ZN(
        n13485) );
  AOI22_X1 U15329 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13483) );
  AOI22_X1 U15330 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13482) );
  AOI22_X1 U15331 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13481) );
  AOI22_X1 U15332 ( .A1(n13543), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13480) );
  NAND4_X1 U15333 ( .A1(n13483), .A2(n13482), .A3(n13481), .A4(n13480), .ZN(
        n13484) );
  OR2_X1 U15334 ( .A1(n13485), .A2(n13484), .ZN(n13507) );
  INV_X1 U15335 ( .A(n13507), .ZN(n13486) );
  XNOR2_X1 U15336 ( .A(n13508), .B(n13486), .ZN(n13490) );
  INV_X1 U15337 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13488) );
  NAND2_X1 U15338 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13487) );
  OAI211_X1 U15339 ( .C1(n13065), .C2(n13488), .A(n13589), .B(n13487), .ZN(
        n13489) );
  AOI21_X1 U15340 ( .B1(n13490), .B2(n13561), .A(n13489), .ZN(n13496) );
  INV_X1 U15341 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16833) );
  INV_X1 U15342 ( .A(n13492), .ZN(n13493) );
  INV_X1 U15343 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16500) );
  NAND2_X1 U15344 ( .A1(n13493), .A2(n16500), .ZN(n13494) );
  NAND2_X1 U15345 ( .A1(n13535), .A2(n13494), .ZN(n16823) );
  NOR2_X1 U15346 ( .A1(n16823), .A2(n13589), .ZN(n13495) );
  AOI22_X1 U15347 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13500) );
  AOI22_X1 U15348 ( .A1(n12848), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12829), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13499) );
  AOI22_X1 U15349 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13549), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13498) );
  AOI22_X1 U15350 ( .A1(n13543), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13497) );
  NAND4_X1 U15351 ( .A1(n13500), .A2(n13499), .A3(n13498), .A4(n13497), .ZN(
        n13506) );
  AOI22_X1 U15352 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13504) );
  AOI22_X1 U15353 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13503) );
  AOI22_X1 U15354 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13502) );
  AOI22_X1 U15355 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13501) );
  NAND4_X1 U15356 ( .A1(n13504), .A2(n13503), .A3(n13502), .A4(n13501), .ZN(
        n13505) );
  NOR2_X1 U15357 ( .A1(n13506), .A2(n13505), .ZN(n13517) );
  NAND2_X1 U15358 ( .A1(n13508), .A2(n13507), .ZN(n13516) );
  XOR2_X1 U15359 ( .A(n13517), .B(n13516), .Z(n13509) );
  NAND2_X1 U15360 ( .A1(n13509), .A2(n13561), .ZN(n13515) );
  INV_X1 U15361 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13511) );
  NAND2_X1 U15362 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13510) );
  OAI211_X1 U15363 ( .C1(n13065), .C2(n13511), .A(n13589), .B(n13510), .ZN(
        n13512) );
  INV_X1 U15364 ( .A(n13512), .ZN(n13514) );
  XNOR2_X1 U15365 ( .A(n13535), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16817) );
  NOR2_X1 U15366 ( .A1(n13517), .A2(n13516), .ZN(n13558) );
  AOI22_X1 U15367 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13550), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13522) );
  AOI22_X1 U15368 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13521) );
  AOI22_X1 U15369 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13520) );
  AOI22_X1 U15370 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13519) );
  NAND4_X1 U15371 ( .A1(n13522), .A2(n13521), .A3(n13520), .A4(n13519), .ZN(
        n13529) );
  AOI22_X1 U15372 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13527) );
  AOI22_X1 U15373 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13526) );
  AOI22_X1 U15374 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13525) );
  AOI22_X1 U15375 ( .A1(n13543), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13524) );
  NAND4_X1 U15376 ( .A1(n13527), .A2(n13526), .A3(n13525), .A4(n13524), .ZN(
        n13528) );
  OR2_X1 U15377 ( .A1(n13529), .A2(n13528), .ZN(n13557) );
  INV_X1 U15378 ( .A(n13557), .ZN(n13530) );
  XNOR2_X1 U15379 ( .A(n13558), .B(n13530), .ZN(n13531) );
  NAND2_X1 U15380 ( .A1(n13531), .A2(n13561), .ZN(n13542) );
  INV_X1 U15381 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13533) );
  NAND2_X1 U15382 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13532) );
  OAI211_X1 U15383 ( .C1(n13065), .C2(n13533), .A(n13589), .B(n13532), .ZN(
        n13534) );
  INV_X1 U15384 ( .A(n13534), .ZN(n13541) );
  INV_X1 U15385 ( .A(n13535), .ZN(n13536) );
  INV_X1 U15386 ( .A(n13537), .ZN(n13538) );
  INV_X1 U15387 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16476) );
  NAND2_X1 U15388 ( .A1(n13538), .A2(n16476), .ZN(n13539) );
  NAND2_X1 U15389 ( .A1(n13595), .A2(n13539), .ZN(n16801) );
  NOR2_X1 U15390 ( .A1(n16801), .A2(n13589), .ZN(n13540) );
  AOI21_X1 U15391 ( .B1(n13542), .B2(n13541), .A(n13540), .ZN(n16475) );
  AOI22_X1 U15392 ( .A1(n13574), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13543), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13547) );
  AOI22_X1 U15393 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13546) );
  AOI22_X1 U15394 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13545) );
  AOI22_X1 U15395 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17061), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13544) );
  NAND4_X1 U15396 ( .A1(n13547), .A2(n13546), .A3(n13545), .A4(n13544), .ZN(
        n13556) );
  AOI22_X1 U15397 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13567), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13554) );
  AOI22_X1 U15398 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13548), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13553) );
  AOI22_X1 U15399 ( .A1(n13549), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13552) );
  AOI22_X1 U15400 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13551) );
  NAND4_X1 U15401 ( .A1(n13554), .A2(n13553), .A3(n13552), .A4(n13551), .ZN(
        n13555) );
  NOR2_X1 U15402 ( .A1(n13556), .A2(n13555), .ZN(n13586) );
  NAND2_X1 U15403 ( .A1(n13558), .A2(n13557), .ZN(n13585) );
  XOR2_X1 U15404 ( .A(n13586), .B(n13585), .Z(n13562) );
  INV_X1 U15405 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n22369) );
  OAI21_X1 U15406 ( .B1(n22268), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n22489), .ZN(n13559) );
  OAI21_X1 U15407 ( .B1(n13065), .B2(n22369), .A(n13559), .ZN(n13560) );
  AOI21_X1 U15408 ( .B1(n13562), .B2(n13561), .A(n13560), .ZN(n13563) );
  INV_X1 U15409 ( .A(n13563), .ZN(n13565) );
  XNOR2_X1 U15410 ( .A(n13595), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16798) );
  NAND2_X1 U15411 ( .A1(n16798), .A2(n13469), .ZN(n13564) );
  NAND2_X1 U15412 ( .A1(n13565), .A2(n13564), .ZN(n16465) );
  AOI22_X1 U15413 ( .A1(n13567), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13566), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13573) );
  AOI22_X1 U15414 ( .A1(n13569), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13568), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13572) );
  AOI22_X1 U15415 ( .A1(n13413), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13523), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13571) );
  AOI22_X1 U15416 ( .A1(n13550), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11175), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13570) );
  NAND4_X1 U15417 ( .A1(n13573), .A2(n13572), .A3(n13571), .A4(n13570), .ZN(
        n13584) );
  AOI22_X1 U15418 ( .A1(n13575), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13574), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13582) );
  AOI22_X1 U15419 ( .A1(n13548), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13549), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13581) );
  AOI22_X1 U15420 ( .A1(n13518), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13580) );
  AOI22_X1 U15421 ( .A1(n13578), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13577), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13579) );
  NAND4_X1 U15422 ( .A1(n13582), .A2(n13581), .A3(n13580), .A4(n13579), .ZN(
        n13583) );
  NOR2_X1 U15423 ( .A1(n13584), .A2(n13583), .ZN(n13588) );
  NOR2_X1 U15424 ( .A1(n13586), .A2(n13585), .ZN(n13587) );
  XOR2_X1 U15425 ( .A(n13588), .B(n13587), .Z(n13594) );
  INV_X1 U15426 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n22375) );
  NAND2_X1 U15427 ( .A1(n22489), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13590) );
  OAI211_X1 U15428 ( .C1(n13065), .C2(n22375), .A(n13590), .B(n13589), .ZN(
        n13591) );
  INV_X1 U15429 ( .A(n13591), .ZN(n13592) );
  OAI21_X1 U15430 ( .B1(n13594), .B2(n13593), .A(n13592), .ZN(n13597) );
  INV_X1 U15431 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16796) );
  XNOR2_X1 U15432 ( .A(n13691), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16457) );
  NAND2_X1 U15433 ( .A1(n16457), .A2(n13469), .ZN(n13596) );
  NAND2_X1 U15434 ( .A1(n13597), .A2(n13596), .ZN(n16331) );
  AOI22_X1 U15435 ( .A1(n13599), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13598), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13600) );
  XNOR2_X1 U15436 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13609) );
  NAND2_X1 U15437 ( .A1(n13626), .A2(n13609), .ZN(n13603) );
  NAND2_X1 U15438 ( .A1(n22476), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13602) );
  NAND2_X1 U15439 ( .A1(n13603), .A2(n13602), .ZN(n13618) );
  XNOR2_X1 U15440 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13617) );
  NAND2_X1 U15441 ( .A1(n13618), .A2(n13617), .ZN(n13620) );
  NAND2_X1 U15442 ( .A1(n22408), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13604) );
  NAND2_X1 U15443 ( .A1(n13620), .A2(n13604), .ZN(n13614) );
  XNOR2_X1 U15444 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13612) );
  NAND2_X1 U15445 ( .A1(n13614), .A2(n13612), .ZN(n13606) );
  NAND2_X1 U15446 ( .A1(n22409), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13605) );
  NAND2_X1 U15447 ( .A1(n13606), .A2(n13605), .ZN(n13611) );
  AND2_X1 U15448 ( .A1(n17899), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13607) );
  NAND2_X1 U15449 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17889), .ZN(
        n13610) );
  XNOR2_X1 U15450 ( .A(n13609), .B(n13626), .ZN(n13634) );
  OR2_X1 U15451 ( .A1(n13611), .A2(n13610), .ZN(n13616) );
  INV_X1 U15452 ( .A(n13612), .ZN(n13613) );
  XNOR2_X1 U15453 ( .A(n13614), .B(n13613), .ZN(n13615) );
  NAND2_X1 U15454 ( .A1(n13616), .A2(n13615), .ZN(n13650) );
  OR2_X1 U15455 ( .A1(n13618), .A2(n13617), .ZN(n13619) );
  NAND2_X1 U15456 ( .A1(n13620), .A2(n13619), .ZN(n13641) );
  OR2_X1 U15457 ( .A1(n13650), .A2(n13641), .ZN(n13621) );
  NOR2_X1 U15458 ( .A1(n13634), .A2(n13621), .ZN(n13622) );
  NOR2_X1 U15459 ( .A1(n13623), .A2(n13622), .ZN(n16369) );
  NAND2_X1 U15460 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n22248) );
  NAND2_X1 U15461 ( .A1(n16369), .A2(n22248), .ZN(n15360) );
  OR2_X1 U15462 ( .A1(n13601), .A2(n15360), .ZN(n13658) );
  NAND2_X1 U15463 ( .A1(n13651), .A2(n13623), .ZN(n13654) );
  NAND2_X1 U15464 ( .A1(n13624), .A2(n13650), .ZN(n13649) );
  AND2_X1 U15465 ( .A1(n15353), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13625) );
  NOR2_X1 U15466 ( .A1(n13626), .A2(n13625), .ZN(n13629) );
  INV_X1 U15467 ( .A(n13629), .ZN(n13627) );
  AOI21_X1 U15468 ( .B1(n12847), .B2(n12895), .A(n13627), .ZN(n13631) );
  AND2_X1 U15469 ( .A1(n12888), .A2(n12885), .ZN(n13628) );
  AOI21_X1 U15470 ( .B1(n13629), .B2(n13640), .A(n13651), .ZN(n13630) );
  AOI21_X1 U15471 ( .B1(n13631), .B2(n13645), .A(n13630), .ZN(n13638) );
  AOI22_X1 U15472 ( .A1(n13642), .A2(n13634), .B1(n16726), .B2(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n13632) );
  NAND3_X1 U15473 ( .A1(n12888), .A2(n13634), .A3(n13632), .ZN(n13637) );
  INV_X1 U15474 ( .A(n13640), .ZN(n13633) );
  OAI21_X1 U15475 ( .B1(n13633), .B2(n12888), .A(n13632), .ZN(n13636) );
  OAI21_X1 U15476 ( .B1(n13640), .B2(n13762), .A(n13634), .ZN(n13635) );
  AOI22_X1 U15477 ( .A1(n13638), .A2(n13637), .B1(n13636), .B2(n13635), .ZN(
        n13647) );
  INV_X1 U15478 ( .A(n13641), .ZN(n13639) );
  NAND2_X1 U15479 ( .A1(n13640), .A2(n13639), .ZN(n13644) );
  NAND2_X1 U15480 ( .A1(n13642), .A2(n13641), .ZN(n13643) );
  AND3_X1 U15481 ( .A1(n13645), .A2(n13644), .A3(n13643), .ZN(n13646) );
  OAI22_X1 U15482 ( .A1(n13647), .A2(n13646), .B1(n13645), .B2(n13644), .ZN(
        n13648) );
  AOI22_X1 U15483 ( .A1(n13651), .A2(n13650), .B1(n13649), .B2(n13648), .ZN(
        n13652) );
  INV_X1 U15484 ( .A(n13652), .ZN(n13653) );
  INV_X1 U15485 ( .A(n16371), .ZN(n16365) );
  INV_X1 U15486 ( .A(n15330), .ZN(n15324) );
  OR2_X1 U15487 ( .A1(n15324), .A2(n12915), .ZN(n13656) );
  NOR2_X1 U15488 ( .A1(n17039), .A2(n13656), .ZN(n15373) );
  NAND2_X1 U15489 ( .A1(n16365), .A2(n15373), .ZN(n13657) );
  INV_X1 U15490 ( .A(n13659), .ZN(n15328) );
  OR2_X1 U15491 ( .A1(n15328), .A2(n16439), .ZN(n15378) );
  INV_X1 U15492 ( .A(n22248), .ZN(n22296) );
  NOR2_X1 U15493 ( .A1(n15378), .A2(n22296), .ZN(n13662) );
  INV_X1 U15494 ( .A(n12842), .ZN(n15557) );
  NAND4_X1 U15495 ( .A1(n15557), .A2(n15570), .A3(n20704), .A4(n13052), .ZN(
        n15446) );
  NOR2_X1 U15496 ( .A1(n13660), .A2(n15446), .ZN(n13661) );
  AOI21_X1 U15497 ( .B1(n15370), .B2(n13662), .A(n13661), .ZN(n13663) );
  AND2_X1 U15498 ( .A1(n16789), .A2(n15557), .ZN(n13665) );
  NOR4_X1 U15499 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13669) );
  NOR4_X1 U15500 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13668) );
  NOR4_X1 U15501 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13667) );
  NOR4_X1 U15502 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13666) );
  AND4_X1 U15503 ( .A1(n13669), .A2(n13668), .A3(n13667), .A4(n13666), .ZN(
        n13674) );
  NOR4_X1 U15504 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n13672) );
  NOR4_X1 U15505 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13671) );
  NOR4_X1 U15506 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13670) );
  INV_X1 U15507 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20528) );
  AND4_X1 U15508 ( .A1(n13672), .A2(n13671), .A3(n13670), .A4(n20528), .ZN(
        n13673) );
  NAND2_X1 U15509 ( .A1(n13674), .A2(n13673), .ZN(n13675) );
  AND2_X2 U15510 ( .A1(n13675), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n16731)
         );
  INV_X1 U15511 ( .A(n16731), .ZN(n16277) );
  NOR3_X1 U15512 ( .A1(n16775), .A2(n12884), .A3(n16277), .ZN(n13676) );
  AOI22_X1 U15513 ( .A1(n16779), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n16775), .ZN(n13677) );
  INV_X1 U15514 ( .A(n13677), .ZN(n13680) );
  NOR2_X1 U15515 ( .A1(n12884), .A2(n16731), .ZN(n13678) );
  NAND2_X1 U15516 ( .A1(n16789), .A2(n13678), .ZN(n16725) );
  INV_X1 U15517 ( .A(DATAI_31_), .ZN(n15556) );
  NOR2_X1 U15518 ( .A1(n16725), .A2(n15556), .ZN(n13679) );
  NOR2_X1 U15519 ( .A1(n13680), .A2(n13679), .ZN(n13681) );
  NAND2_X1 U15520 ( .A1(n13682), .A2(n13681), .ZN(P1_U2873) );
  NAND3_X1 U15521 ( .A1(n22256), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n22252) );
  INV_X1 U15522 ( .A(n22252), .ZN(n13683) );
  NAND2_X1 U15523 ( .A1(n12847), .A2(n15583), .ZN(n13684) );
  AND2_X1 U15524 ( .A1(n11745), .A2(n13684), .ZN(n15320) );
  NAND2_X1 U15525 ( .A1(n17039), .A2(n15813), .ZN(n13685) );
  NAND3_X1 U15526 ( .A1(n15320), .A2(n15330), .A3(n13685), .ZN(n15341) );
  OR2_X1 U15527 ( .A1(n15341), .A2(n13686), .ZN(n15375) );
  INV_X1 U15528 ( .A(n15375), .ZN(n17879) );
  NAND2_X1 U15529 ( .A1(n22506), .A2(n13687), .ZN(n21954) );
  NAND2_X1 U15530 ( .A1(n21954), .A2(n22256), .ZN(n13688) );
  NAND2_X1 U15531 ( .A1(n22256), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13690) );
  NAND2_X1 U15532 ( .A1(n22268), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13689) );
  NAND2_X1 U15533 ( .A1(n13690), .A2(n13689), .ZN(n20631) );
  INV_X1 U15534 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16333) );
  XNOR2_X1 U15535 ( .A(n13692), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15805) );
  NAND2_X1 U15536 ( .A1(n22497), .A2(n22250), .ZN(n20706) );
  OR2_X2 U15537 ( .A1(n20706), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n22093) );
  INV_X1 U15538 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20574) );
  NOR2_X1 U15539 ( .A1(n22093), .A2(n20574), .ZN(n16938) );
  AOI21_X1 U15540 ( .B1(n20694), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16938), .ZN(n13693) );
  OAI21_X1 U15541 ( .B1(n20703), .B2(n15805), .A(n13693), .ZN(n13694) );
  AOI21_X1 U15542 ( .B1(n16378), .B2(n20689), .A(n13694), .ZN(n13805) );
  AND2_X1 U15543 ( .A1(n15813), .A2(n15384), .ZN(n13712) );
  AOI21_X1 U15544 ( .B1(n13698), .B2(n21956), .A(n13712), .ZN(n13695) );
  OR2_X1 U15545 ( .A1(n13697), .A2(n13762), .ZN(n13702) );
  XNOR2_X1 U15546 ( .A(n13698), .B(n13709), .ZN(n13699) );
  NAND2_X1 U15547 ( .A1(n13699), .A2(n21956), .ZN(n13700) );
  AND3_X1 U15548 ( .A1(n13700), .A2(n15330), .A3(n12885), .ZN(n13701) );
  NAND2_X1 U15549 ( .A1(n13702), .A2(n13701), .ZN(n13703) );
  NAND2_X1 U15550 ( .A1(n15359), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13706) );
  INV_X1 U15551 ( .A(n13703), .ZN(n13704) );
  OR2_X1 U15552 ( .A1(n20628), .A2(n13704), .ZN(n13705) );
  NAND2_X1 U15553 ( .A1(n13706), .A2(n13705), .ZN(n13716) );
  INV_X1 U15554 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15456) );
  XNOR2_X1 U15555 ( .A(n13716), .B(n15456), .ZN(n15455) );
  OR2_X1 U15556 ( .A1(n15435), .A2(n13762), .ZN(n13715) );
  INV_X1 U15557 ( .A(n13707), .ZN(n13711) );
  NAND2_X1 U15558 ( .A1(n13709), .A2(n13708), .ZN(n13710) );
  NAND2_X1 U15559 ( .A1(n13710), .A2(n13711), .ZN(n13720) );
  OAI21_X1 U15560 ( .B1(n13711), .B2(n13710), .A(n13720), .ZN(n13713) );
  AOI21_X1 U15561 ( .B1(n13713), .B2(n21956), .A(n13712), .ZN(n13714) );
  NAND2_X1 U15562 ( .A1(n13715), .A2(n13714), .ZN(n15454) );
  NAND2_X1 U15563 ( .A1(n15455), .A2(n15454), .ZN(n13718) );
  NAND2_X1 U15564 ( .A1(n13716), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13717) );
  INV_X1 U15565 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13719) );
  OR2_X1 U15566 ( .A1(n15962), .A2(n13762), .ZN(n13723) );
  NAND2_X1 U15567 ( .A1(n13720), .A2(n13721), .ZN(n13736) );
  OAI211_X1 U15568 ( .C1(n13721), .C2(n13720), .A(n13736), .B(n21956), .ZN(
        n13722) );
  NAND2_X1 U15569 ( .A1(n13723), .A2(n13722), .ZN(n15819) );
  NAND2_X1 U15570 ( .A1(n15818), .A2(n15819), .ZN(n13726) );
  NAND2_X1 U15571 ( .A1(n13724), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13725) );
  NAND2_X1 U15572 ( .A1(n13726), .A2(n13725), .ZN(n15785) );
  OR2_X1 U15573 ( .A1(n13727), .A2(n13762), .ZN(n13730) );
  XNOR2_X1 U15574 ( .A(n13736), .B(n13734), .ZN(n13728) );
  NAND2_X1 U15575 ( .A1(n13728), .A2(n21956), .ZN(n13729) );
  NAND2_X1 U15576 ( .A1(n13730), .A2(n13729), .ZN(n13731) );
  INV_X1 U15577 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21986) );
  XNOR2_X1 U15578 ( .A(n13731), .B(n21986), .ZN(n15784) );
  NAND2_X1 U15579 ( .A1(n15785), .A2(n15784), .ZN(n13733) );
  NAND2_X1 U15580 ( .A1(n13731), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13732) );
  INV_X1 U15581 ( .A(n13734), .ZN(n13735) );
  NOR2_X1 U15582 ( .A1(n13736), .A2(n13735), .ZN(n13738) );
  NAND2_X1 U15583 ( .A1(n13738), .A2(n13737), .ZN(n13753) );
  OAI211_X1 U15584 ( .C1(n13738), .C2(n13737), .A(n13753), .B(n21956), .ZN(
        n13739) );
  OAI21_X1 U15585 ( .B1(n13740), .B2(n13762), .A(n13739), .ZN(n13741) );
  INV_X1 U15586 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16923) );
  XNOR2_X1 U15587 ( .A(n13741), .B(n16923), .ZN(n16014) );
  NAND2_X1 U15588 ( .A1(n16013), .A2(n16014), .ZN(n13743) );
  NAND2_X1 U15589 ( .A1(n13741), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13742) );
  NAND2_X1 U15590 ( .A1(n13743), .A2(n13742), .ZN(n15981) );
  NAND3_X1 U15591 ( .A1(n13765), .A2(n13751), .A3(n13744), .ZN(n13747) );
  XNOR2_X1 U15592 ( .A(n13753), .B(n13754), .ZN(n13745) );
  NAND2_X1 U15593 ( .A1(n13745), .A2(n21956), .ZN(n13746) );
  NAND2_X1 U15594 ( .A1(n13747), .A2(n13746), .ZN(n13748) );
  INV_X1 U15595 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n22006) );
  XNOR2_X1 U15596 ( .A(n13748), .B(n22006), .ZN(n15980) );
  NAND2_X1 U15597 ( .A1(n15981), .A2(n15980), .ZN(n13750) );
  NAND2_X1 U15598 ( .A1(n13748), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13749) );
  NAND2_X1 U15599 ( .A1(n13750), .A2(n13749), .ZN(n16201) );
  NAND2_X1 U15600 ( .A1(n13752), .A2(n13751), .ZN(n13758) );
  INV_X1 U15601 ( .A(n13753), .ZN(n13755) );
  NAND2_X1 U15602 ( .A1(n13755), .A2(n13754), .ZN(n13768) );
  XNOR2_X1 U15603 ( .A(n13768), .B(n13766), .ZN(n13756) );
  NAND2_X1 U15604 ( .A1(n13756), .A2(n21956), .ZN(n13757) );
  NAND2_X1 U15605 ( .A1(n13758), .A2(n13757), .ZN(n13760) );
  INV_X1 U15606 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13759) );
  XNOR2_X1 U15607 ( .A(n13760), .B(n13759), .ZN(n16202) );
  NAND2_X1 U15608 ( .A1(n13760), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13761) );
  NOR2_X1 U15609 ( .A1(n13763), .A2(n13762), .ZN(n13764) );
  NAND2_X1 U15610 ( .A1(n21956), .A2(n13766), .ZN(n13767) );
  OR2_X1 U15611 ( .A1(n13768), .A2(n13767), .ZN(n13769) );
  NAND2_X1 U15612 ( .A1(n13786), .A2(n13769), .ZN(n13770) );
  INV_X1 U15613 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16179) );
  XNOR2_X1 U15614 ( .A(n13770), .B(n16179), .ZN(n16169) );
  XNOR2_X1 U15615 ( .A(n13786), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16249) );
  INV_X1 U15616 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13771) );
  INV_X1 U15617 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13773) );
  NAND2_X1 U15618 ( .A1(n13786), .A2(n13773), .ZN(n13774) );
  NAND2_X1 U15619 ( .A1(n20670), .A2(n13774), .ZN(n16909) );
  NAND2_X1 U15620 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13775) );
  AND2_X1 U15621 ( .A1(n13786), .A2(n13775), .ZN(n16905) );
  INV_X1 U15622 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n22025) );
  INV_X1 U15623 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16386) );
  AND2_X1 U15624 ( .A1(n13786), .A2(n16386), .ZN(n13776) );
  NOR2_X1 U15625 ( .A1(n20671), .A2(n13776), .ZN(n13777) );
  NAND2_X1 U15626 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n22060) );
  INV_X1 U15627 ( .A(n22060), .ZN(n22049) );
  NAND2_X1 U15628 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n22049), .ZN(
        n13778) );
  NOR2_X1 U15629 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13779) );
  OR2_X1 U15630 ( .A1(n13786), .A2(n13779), .ZN(n16904) );
  OR2_X1 U15631 ( .A1(n13786), .A2(n22025), .ZN(n16906) );
  NAND2_X1 U15632 ( .A1(n16904), .A2(n16906), .ZN(n20668) );
  INV_X1 U15633 ( .A(n20670), .ZN(n13781) );
  NOR2_X1 U15634 ( .A1(n13786), .A2(n16386), .ZN(n13780) );
  NOR3_X2 U15635 ( .A1(n20668), .A2(n13781), .A3(n13780), .ZN(n16895) );
  INV_X1 U15636 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17030) );
  OR2_X1 U15637 ( .A1(n13786), .A2(n17030), .ZN(n13782) );
  NOR2_X1 U15638 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13783) );
  NOR2_X1 U15639 ( .A1(n13786), .A2(n13783), .ZN(n13784) );
  INV_X1 U15640 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16859) );
  INV_X1 U15641 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16857) );
  NAND2_X1 U15642 ( .A1(n16859), .A2(n16857), .ZN(n13785) );
  NAND3_X1 U15643 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16919) );
  INV_X1 U15644 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n22048) );
  NOR2_X1 U15645 ( .A1(n16919), .A2(n22048), .ZN(n13788) );
  NAND2_X2 U15646 ( .A1(n16991), .A2(n16827), .ZN(n16850) );
  INV_X1 U15647 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16838) );
  INV_X1 U15648 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16842) );
  INV_X1 U15649 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13789) );
  NAND3_X1 U15650 ( .A1(n16838), .A2(n16842), .A3(n13789), .ZN(n16803) );
  OR2_X2 U15651 ( .A1(n16850), .A2(n16803), .ZN(n13792) );
  NAND3_X1 U15652 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16926) );
  NOR2_X1 U15653 ( .A1(n16827), .A2(n16926), .ZN(n13790) );
  NAND2_X1 U15654 ( .A1(n13792), .A2(n11670), .ZN(n13793) );
  NOR2_X1 U15655 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16963) );
  NAND2_X1 U15656 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16965) );
  INV_X1 U15657 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16927) );
  INV_X1 U15658 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16934) );
  XNOR2_X1 U15659 ( .A(n11667), .B(n16934), .ZN(n13799) );
  INV_X1 U15660 ( .A(n13799), .ZN(n13794) );
  INV_X1 U15661 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16933) );
  NAND2_X1 U15662 ( .A1(n13786), .A2(n16933), .ZN(n13796) );
  NAND2_X1 U15663 ( .A1(n13794), .A2(n13796), .ZN(n13802) );
  NOR2_X1 U15664 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13795) );
  OR2_X1 U15665 ( .A1(n11667), .A2(n13795), .ZN(n13798) );
  NAND2_X1 U15666 ( .A1(n13798), .A2(n13796), .ZN(n13797) );
  NAND2_X1 U15667 ( .A1(n13797), .A2(n16934), .ZN(n13801) );
  NAND3_X1 U15668 ( .A1(n13803), .A2(n13799), .A3(n13798), .ZN(n13800) );
  INV_X1 U15669 ( .A(n20696), .ZN(n13804) );
  BUF_X4 U15670 ( .A(n13822), .Z(n15439) );
  INV_X1 U15671 ( .A(n13809), .ZN(n13812) );
  INV_X1 U15672 ( .A(n13810), .ZN(n13811) );
  NAND2_X1 U15673 ( .A1(n13812), .A2(n13811), .ZN(n13813) );
  INV_X1 U15674 ( .A(n19023), .ZN(n19230) );
  OR2_X1 U15675 ( .A1(n14368), .A2(n19230), .ZN(n13840) );
  NOR2_X1 U15676 ( .A1(n15439), .A2(n13840), .ZN(n13820) );
  INV_X1 U15677 ( .A(n13814), .ZN(n13817) );
  INV_X1 U15678 ( .A(n13818), .ZN(n13819) );
  NAND2_X1 U15679 ( .A1(n16027), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13828) );
  INV_X2 U15680 ( .A(n17172), .ZN(n17905) );
  AND2_X1 U15681 ( .A1(n19230), .A2(n13823), .ZN(n13838) );
  INV_X1 U15682 ( .A(n13838), .ZN(n13824) );
  OR3_X2 U15683 ( .A1(n15439), .A2(n17905), .A3(n13824), .ZN(n19999) );
  INV_X1 U15684 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13821) );
  OR2_X1 U15685 ( .A1(n19999), .A2(n13821), .ZN(n13827) );
  OR2_X1 U15686 ( .A1(n13823), .A2(n19023), .ZN(n13858) );
  OR3_X2 U15687 ( .A1(n15439), .A2(n17905), .A3(n13858), .ZN(n19983) );
  INV_X1 U15688 ( .A(n19983), .ZN(n19989) );
  NAND2_X1 U15689 ( .A1(n19989), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13826) );
  INV_X1 U15690 ( .A(n13940), .ZN(n19956) );
  NAND2_X1 U15691 ( .A1(n19956), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13825) );
  NAND4_X1 U15692 ( .A1(n13828), .A2(n13827), .A3(n13826), .A4(n13825), .ZN(
        n13837) );
  AND2_X1 U15693 ( .A1(n14368), .A2(n19023), .ZN(n13855) );
  OR2_X2 U15694 ( .A1(n13845), .A2(n11171), .ZN(n15078) );
  INV_X1 U15695 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13835) );
  NAND2_X1 U15696 ( .A1(n13855), .A2(n11171), .ZN(n13829) );
  INV_X1 U15697 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13830) );
  OR2_X1 U15698 ( .A1(n19942), .A2(n13830), .ZN(n13834) );
  INV_X1 U15699 ( .A(n13822), .ZN(n13832) );
  OAI211_X1 U15700 ( .C1(n15078), .C2(n13835), .A(n13834), .B(n13833), .ZN(
        n13836) );
  NOR2_X1 U15701 ( .A1(n13837), .A2(n13836), .ZN(n13864) );
  INV_X1 U15702 ( .A(n19864), .ZN(n19858) );
  INV_X1 U15703 ( .A(n13858), .ZN(n13839) );
  INV_X1 U15704 ( .A(n13924), .ZN(n19874) );
  AOI22_X1 U15705 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19858), .B1(
        n19874), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13852) );
  INV_X1 U15706 ( .A(n13840), .ZN(n13841) );
  NAND2_X1 U15707 ( .A1(n13841), .A2(n15439), .ZN(n13843) );
  INV_X1 U15708 ( .A(n19886), .ZN(n19892) );
  INV_X1 U15709 ( .A(n13931), .ZN(n19831) );
  AOI22_X1 U15710 ( .A1(n19892), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n19831), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13851) );
  OR2_X2 U15711 ( .A1(n13843), .A2(n11171), .ZN(n19917) );
  INV_X1 U15712 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13844) );
  INV_X1 U15713 ( .A(n13845), .ZN(n13846) );
  NAND2_X2 U15714 ( .A1(n13846), .A2(n11171), .ZN(n19851) );
  INV_X1 U15715 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13847) );
  NOR2_X1 U15716 ( .A1(n19851), .A2(n13847), .ZN(n13848) );
  NOR2_X1 U15717 ( .A1(n13849), .A2(n13848), .ZN(n13850) );
  AND3_X1 U15718 ( .A1(n13852), .A2(n13851), .A3(n13850), .ZN(n13863) );
  INV_X1 U15719 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13854) );
  INV_X1 U15720 ( .A(n13855), .ZN(n13856) );
  INV_X1 U15721 ( .A(n19970), .ZN(n13857) );
  INV_X1 U15722 ( .A(n19930), .ZN(n19925) );
  NAND2_X1 U15723 ( .A1(n19925), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13859) );
  NAND3_X1 U15724 ( .A1(n13864), .A2(n13863), .A3(n13862), .ZN(n13867) );
  AND2_X1 U15725 ( .A1(n20262), .A2(n14094), .ZN(n16307) );
  NAND2_X1 U15726 ( .A1(n16307), .A2(n14093), .ZN(n14090) );
  INV_X1 U15727 ( .A(n13865), .ZN(n14091) );
  NAND2_X1 U15728 ( .A1(n14090), .A2(n14091), .ZN(n13866) );
  INV_X1 U15729 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13869) );
  INV_X1 U15730 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13868) );
  OAI22_X1 U15731 ( .A1(n13869), .A2(n13940), .B1(n19930), .B2(n13868), .ZN(
        n13873) );
  INV_X1 U15732 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13871) );
  INV_X1 U15733 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13870) );
  OAI22_X1 U15734 ( .A1(n13871), .A2(n19983), .B1(n19999), .B2(n13870), .ZN(
        n13872) );
  NOR2_X1 U15735 ( .A1(n13873), .A2(n13872), .ZN(n13881) );
  INV_X1 U15736 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13875) );
  INV_X1 U15737 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13874) );
  OAI22_X1 U15738 ( .A1(n13875), .A2(n15078), .B1(n19904), .B2(n13874), .ZN(
        n13879) );
  INV_X1 U15739 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13877) );
  INV_X1 U15740 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13876) );
  OAI22_X1 U15741 ( .A1(n13877), .A2(n13924), .B1(n19864), .B2(n13876), .ZN(
        n13878) );
  NOR2_X1 U15742 ( .A1(n13879), .A2(n13878), .ZN(n13880) );
  INV_X1 U15743 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13883) );
  INV_X1 U15744 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13882) );
  OAI22_X1 U15745 ( .A1(n13883), .A2(n19886), .B1(n13931), .B2(n13882), .ZN(
        n13887) );
  INV_X1 U15746 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13885) );
  INV_X1 U15747 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13884) );
  OAI22_X1 U15748 ( .A1(n13885), .A2(n19917), .B1(n19851), .B2(n13884), .ZN(
        n13886) );
  NOR2_X1 U15749 ( .A1(n13887), .A2(n13886), .ZN(n13893) );
  INV_X1 U15750 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13888) );
  INV_X1 U15751 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17800) );
  OAI22_X1 U15752 ( .A1(n19970), .A2(n13888), .B1(n13945), .B2(n17800), .ZN(
        n13891) );
  INV_X1 U15753 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13889) );
  INV_X1 U15754 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16034) );
  OAI22_X1 U15755 ( .A1(n19942), .A2(n13889), .B1(n13947), .B2(n16034), .ZN(
        n13890) );
  NOR2_X1 U15756 ( .A1(n13891), .A2(n13890), .ZN(n13892) );
  NAND2_X1 U15757 ( .A1(n13893), .A2(n13892), .ZN(n13897) );
  INV_X1 U15758 ( .A(n13894), .ZN(n13895) );
  NAND2_X1 U15759 ( .A1(n13895), .A2(n20262), .ZN(n13896) );
  NAND2_X1 U15760 ( .A1(n13900), .A2(n13899), .ZN(n13901) );
  XNOR2_X1 U15761 ( .A(n13908), .B(n11845), .ZN(n16056) );
  INV_X1 U15762 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19339) );
  INV_X1 U15763 ( .A(n13904), .ZN(n13906) );
  INV_X1 U15764 ( .A(n13905), .ZN(n13910) );
  NAND2_X1 U15765 ( .A1(n13906), .A2(n13910), .ZN(n13907) );
  NAND2_X1 U15766 ( .A1(n13908), .A2(n13907), .ZN(n17169) );
  INV_X1 U15767 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15222) );
  NAND3_X1 U15768 ( .A1(n11843), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n13909) );
  NAND2_X1 U15769 ( .A1(n13910), .A2(n13909), .ZN(n17182) );
  NAND2_X1 U15770 ( .A1(n11761), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13911) );
  NAND2_X1 U15771 ( .A1(n13912), .A2(n13911), .ZN(n14123) );
  MUX2_X1 U15772 ( .A(n13913), .B(n14123), .S(n12003), .Z(n14079) );
  AOI21_X1 U15773 ( .B1(n14079), .B2(n13915), .A(n13914), .ZN(n19019) );
  NAND2_X1 U15774 ( .A1(n19019), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16311) );
  NOR2_X1 U15775 ( .A1(n17182), .A2(n16311), .ZN(n13916) );
  XNOR2_X1 U15776 ( .A(n17182), .B(n16311), .ZN(n15140) );
  NOR2_X1 U15777 ( .A1(n15206), .A2(n15140), .ZN(n15139) );
  NOR2_X1 U15778 ( .A1(n13916), .A2(n15139), .ZN(n15217) );
  XNOR2_X1 U15779 ( .A(n17169), .B(n15222), .ZN(n15216) );
  OR2_X1 U15780 ( .A1(n15217), .A2(n15216), .ZN(n15219) );
  OAI21_X1 U15781 ( .B1(n17169), .B2(n15222), .A(n15219), .ZN(n17918) );
  NAND2_X1 U15782 ( .A1(n13917), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13918) );
  NAND2_X1 U15783 ( .A1(n17917), .A2(n13918), .ZN(n16090) );
  NAND2_X1 U15784 ( .A1(n11262), .A2(n11413), .ZN(n13921) );
  NAND2_X1 U15785 ( .A1(n13919), .A2(n13921), .ZN(n19034) );
  XNOR2_X1 U15786 ( .A(n19034), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16089) );
  NAND2_X1 U15787 ( .A1(n16090), .A2(n16089), .ZN(n16092) );
  INV_X1 U15788 ( .A(n19034), .ZN(n13922) );
  NAND2_X1 U15789 ( .A1(n13922), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13923) );
  NAND2_X1 U15790 ( .A1(n16092), .A2(n13923), .ZN(n16152) );
  INV_X1 U15791 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13926) );
  INV_X1 U15792 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13925) );
  OAI22_X1 U15793 ( .A1(n13926), .A2(n19864), .B1(n13924), .B2(n13925), .ZN(
        n13930) );
  INV_X1 U15794 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13928) );
  INV_X1 U15795 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13927) );
  OAI22_X1 U15796 ( .A1(n13928), .A2(n19904), .B1(n19851), .B2(n13927), .ZN(
        n13929) );
  NOR2_X1 U15797 ( .A1(n13930), .A2(n13929), .ZN(n13955) );
  INV_X1 U15798 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13933) );
  INV_X1 U15799 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13932) );
  OAI22_X1 U15800 ( .A1(n13933), .A2(n19886), .B1(n13931), .B2(n13932), .ZN(
        n13937) );
  INV_X1 U15801 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13935) );
  INV_X1 U15802 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13934) );
  OAI22_X1 U15803 ( .A1(n13935), .A2(n19917), .B1(n15078), .B2(n13934), .ZN(
        n13936) );
  NOR2_X1 U15804 ( .A1(n13937), .A2(n13936), .ZN(n13954) );
  INV_X1 U15805 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13939) );
  INV_X1 U15806 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13938) );
  OAI22_X1 U15807 ( .A1(n13939), .A2(n19999), .B1(n19930), .B2(n13938), .ZN(
        n13944) );
  INV_X1 U15808 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13942) );
  INV_X1 U15809 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13941) );
  OAI22_X1 U15810 ( .A1(n13942), .A2(n13940), .B1(n19983), .B2(n13941), .ZN(
        n13943) );
  NOR2_X1 U15811 ( .A1(n13944), .A2(n13943), .ZN(n13953) );
  INV_X1 U15812 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13946) );
  OAI22_X1 U15813 ( .A1(n19970), .A2(n13946), .B1(n13945), .B2(n20108), .ZN(
        n13951) );
  INV_X1 U15814 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13949) );
  INV_X1 U15815 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13948) );
  OAI22_X1 U15816 ( .A1(n19942), .A2(n13949), .B1(n13947), .B2(n13948), .ZN(
        n13950) );
  NOR2_X1 U15817 ( .A1(n13951), .A2(n13950), .ZN(n13952) );
  NAND4_X1 U15818 ( .A1(n13955), .A2(n13954), .A3(n13953), .A4(n13952), .ZN(
        n13958) );
  NAND2_X1 U15819 ( .A1(n13956), .A2(n14120), .ZN(n13957) );
  NAND2_X1 U15820 ( .A1(n14104), .A2(n14324), .ZN(n13960) );
  XNOR2_X1 U15821 ( .A(n13919), .B(n13959), .ZN(n16131) );
  NAND2_X1 U15822 ( .A1(n13960), .A2(n16131), .ZN(n13961) );
  XNOR2_X1 U15823 ( .A(n13961), .B(n16166), .ZN(n16151) );
  NAND2_X1 U15824 ( .A1(n16152), .A2(n16151), .ZN(n16150) );
  NAND2_X1 U15825 ( .A1(n13961), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13962) );
  NAND2_X1 U15826 ( .A1(n16150), .A2(n13962), .ZN(n17532) );
  NAND2_X1 U15827 ( .A1(n13965), .A2(n13964), .ZN(n13988) );
  INV_X1 U15828 ( .A(n13988), .ZN(n13986) );
  INV_X1 U15829 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14457) );
  INV_X1 U15830 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13966) );
  OAI22_X1 U15831 ( .A1(n14457), .A2(n19851), .B1(n13931), .B2(n13966), .ZN(
        n13969) );
  INV_X1 U15832 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14455) );
  INV_X1 U15833 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13967) );
  OAI22_X1 U15834 ( .A1(n14455), .A2(n19917), .B1(n19904), .B2(n13967), .ZN(
        n13968) );
  NOR2_X1 U15835 ( .A1(n13969), .A2(n13968), .ZN(n13982) );
  INV_X1 U15836 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14450) );
  INV_X1 U15837 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14447) );
  OAI22_X1 U15838 ( .A1(n14450), .A2(n19864), .B1(n15078), .B2(n14447), .ZN(
        n13971) );
  INV_X1 U15839 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n20036) );
  INV_X1 U15840 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14452) );
  OAI22_X1 U15841 ( .A1(n20036), .A2(n19886), .B1(n13924), .B2(n14452), .ZN(
        n13970) );
  NOR2_X1 U15842 ( .A1(n13971), .A2(n13970), .ZN(n13981) );
  INV_X1 U15843 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14469) );
  INV_X1 U15844 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13972) );
  OAI22_X1 U15845 ( .A1(n14469), .A2(n19983), .B1(n19930), .B2(n13972), .ZN(
        n13976) );
  INV_X1 U15846 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13974) );
  INV_X1 U15847 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13973) );
  OAI22_X1 U15848 ( .A1(n13974), .A2(n13940), .B1(n19999), .B2(n13973), .ZN(
        n13975) );
  NOR2_X1 U15849 ( .A1(n13976), .A2(n13975), .ZN(n13980) );
  INV_X1 U15850 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14472) );
  INV_X1 U15851 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20062) );
  OAI22_X1 U15852 ( .A1(n19970), .A2(n14472), .B1(n13945), .B2(n20062), .ZN(
        n13978) );
  INV_X1 U15853 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14467) );
  INV_X1 U15854 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14462) );
  OAI22_X1 U15855 ( .A1(n19942), .A2(n14467), .B1(n13947), .B2(n14462), .ZN(
        n13977) );
  NOR2_X1 U15856 ( .A1(n13978), .A2(n13977), .ZN(n13979) );
  NAND4_X1 U15857 ( .A1(n13982), .A2(n13981), .A3(n13980), .A4(n13979), .ZN(
        n13985) );
  NAND2_X1 U15858 ( .A1(n13983), .A2(n14120), .ZN(n13984) );
  NAND2_X1 U15859 ( .A1(n13986), .A2(n14108), .ZN(n14087) );
  INV_X1 U15860 ( .A(n14108), .ZN(n13987) );
  NAND2_X1 U15861 ( .A1(n13988), .A2(n13987), .ZN(n13989) );
  XNOR2_X1 U15862 ( .A(n13991), .B(n13990), .ZN(n19045) );
  NAND2_X1 U15863 ( .A1(n13992), .A2(n19045), .ZN(n13993) );
  INV_X1 U15864 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n19299) );
  XNOR2_X1 U15865 ( .A(n13993), .B(n19299), .ZN(n17530) );
  NAND2_X1 U15866 ( .A1(n13993), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13994) );
  XNOR2_X1 U15867 ( .A(n13996), .B(n13995), .ZN(n16144) );
  XNOR2_X1 U15868 ( .A(n16144), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17937) );
  INV_X1 U15869 ( .A(n16144), .ZN(n13997) );
  NAND2_X1 U15870 ( .A1(n13997), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13998) );
  NAND2_X1 U15871 ( .A1(n11250), .A2(n11275), .ZN(n14000) );
  NAND2_X1 U15872 ( .A1(n13999), .A2(n14000), .ZN(n19056) );
  OR2_X1 U15873 ( .A1(n19056), .A2(n14324), .ZN(n14001) );
  NOR2_X1 U15874 ( .A1(n14001), .A2(n17761), .ZN(n17754) );
  NAND2_X1 U15875 ( .A1(n14001), .A2(n17761), .ZN(n17752) );
  XNOR2_X1 U15876 ( .A(n13999), .B(n14002), .ZN(n16106) );
  AOI21_X1 U15877 ( .B1(n16106), .B2(n14067), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17733) );
  XNOR2_X1 U15878 ( .A(n14005), .B(n14004), .ZN(n19066) );
  NAND2_X1 U15879 ( .A1(n19066), .A2(n14067), .ZN(n14014) );
  INV_X1 U15880 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14013) );
  AND2_X1 U15881 ( .A1(n14014), .A2(n14013), .ZN(n17719) );
  NAND2_X1 U15882 ( .A1(n14009), .A2(n14008), .ZN(n14010) );
  NAND2_X1 U15883 ( .A1(n14018), .A2(n14010), .ZN(n16120) );
  NOR2_X1 U15884 ( .A1(n16120), .A2(n14324), .ZN(n14012) );
  INV_X1 U15885 ( .A(n14012), .ZN(n14011) );
  NAND2_X1 U15886 ( .A1(n14012), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17968) );
  OR2_X1 U15887 ( .A1(n14014), .A2(n14013), .ZN(n17718) );
  AND2_X1 U15888 ( .A1(n14067), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14015) );
  NAND2_X1 U15889 ( .A1(n16106), .A2(n14015), .ZN(n17730) );
  AND2_X1 U15890 ( .A1(n17718), .A2(n17730), .ZN(n17965) );
  AND2_X1 U15891 ( .A1(n17968), .A2(n17965), .ZN(n14016) );
  XNOR2_X1 U15892 ( .A(n14018), .B(n14017), .ZN(n19078) );
  AND2_X1 U15893 ( .A1(n14067), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14019) );
  AND2_X1 U15894 ( .A1(n19078), .A2(n14019), .ZN(n17703) );
  NAND2_X1 U15895 ( .A1(n19078), .A2(n14067), .ZN(n14020) );
  INV_X1 U15896 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17695) );
  NAND2_X1 U15897 ( .A1(n14020), .A2(n17695), .ZN(n17704) );
  XNOR2_X1 U15898 ( .A(n14022), .B(n14021), .ZN(n19093) );
  AND2_X1 U15899 ( .A1(n14067), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14023) );
  NAND2_X1 U15900 ( .A1(n19093), .A2(n14023), .ZN(n17685) );
  NAND2_X1 U15901 ( .A1(n14032), .A2(n14024), .ZN(n14025) );
  NAND2_X1 U15902 ( .A1(n11182), .A2(n14025), .ZN(n16222) );
  INV_X1 U15903 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17662) );
  OAI21_X1 U15904 ( .B1(n16222), .B2(n14324), .A(n17662), .ZN(n17516) );
  NAND2_X1 U15905 ( .A1(n19093), .A2(n14067), .ZN(n14026) );
  NAND2_X1 U15906 ( .A1(n14026), .A2(n17696), .ZN(n17686) );
  INV_X1 U15907 ( .A(n14027), .ZN(n14030) );
  INV_X1 U15908 ( .A(n14028), .ZN(n14029) );
  NAND2_X1 U15909 ( .A1(n14030), .A2(n14029), .ZN(n14031) );
  NAND2_X1 U15910 ( .A1(n14032), .A2(n14031), .ZN(n19103) );
  OR2_X1 U15911 ( .A1(n19103), .A2(n14324), .ZN(n14034) );
  INV_X1 U15912 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14033) );
  NAND2_X1 U15913 ( .A1(n14034), .A2(n14033), .ZN(n17993) );
  AND3_X1 U15914 ( .A1(n17516), .A2(n17686), .A3(n17993), .ZN(n14231) );
  INV_X1 U15915 ( .A(n16222), .ZN(n14036) );
  AND2_X1 U15916 ( .A1(n14067), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14035) );
  NAND2_X1 U15917 ( .A1(n14036), .A2(n14035), .ZN(n17515) );
  NAND2_X1 U15918 ( .A1(n14067), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14037) );
  AND2_X1 U15919 ( .A1(n17515), .A2(n17992), .ZN(n14235) );
  INV_X1 U15920 ( .A(n14038), .ZN(n14039) );
  NAND2_X1 U15921 ( .A1(n11182), .A2(n14039), .ZN(n14040) );
  NAND2_X1 U15922 ( .A1(n14045), .A2(n14040), .ZN(n19113) );
  OR2_X1 U15923 ( .A1(n19113), .A2(n14324), .ZN(n14041) );
  XNOR2_X1 U15924 ( .A(n14041), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n18005) );
  INV_X1 U15925 ( .A(n14041), .ZN(n14042) );
  NAND2_X1 U15926 ( .A1(n14042), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14236) );
  INV_X1 U15927 ( .A(n14043), .ZN(n14049) );
  NAND2_X1 U15928 ( .A1(n14045), .A2(n14044), .ZN(n14046) );
  AND2_X1 U15929 ( .A1(n14049), .A2(n14046), .ZN(n15096) );
  NAND2_X1 U15930 ( .A1(n15096), .A2(n14067), .ZN(n14051) );
  INV_X1 U15931 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17663) );
  NAND2_X1 U15932 ( .A1(n14051), .A2(n17663), .ZN(n17503) );
  INV_X1 U15933 ( .A(n14047), .ZN(n14048) );
  NAND2_X1 U15934 ( .A1(n14049), .A2(n14048), .ZN(n14050) );
  NAND2_X1 U15935 ( .A1(n14055), .A2(n14050), .ZN(n19121) );
  NOR2_X1 U15936 ( .A1(n19121), .A2(n14324), .ZN(n14060) );
  NAND2_X1 U15937 ( .A1(n14060), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17498) );
  INV_X1 U15938 ( .A(n14051), .ZN(n14052) );
  NAND2_X1 U15939 ( .A1(n14052), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17504) );
  AND2_X1 U15940 ( .A1(n17498), .A2(n17504), .ZN(n14057) );
  INV_X1 U15941 ( .A(n14053), .ZN(n14065) );
  NAND2_X1 U15942 ( .A1(n14055), .A2(n14054), .ZN(n14056) );
  NAND2_X1 U15943 ( .A1(n14065), .A2(n14056), .ZN(n19137) );
  NOR2_X1 U15944 ( .A1(n19137), .A2(n14324), .ZN(n14058) );
  NAND2_X1 U15945 ( .A1(n14058), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17484) );
  AND2_X1 U15946 ( .A1(n14057), .A2(n17484), .ZN(n14238) );
  INV_X1 U15947 ( .A(n14058), .ZN(n14059) );
  INV_X1 U15948 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17633) );
  INV_X1 U15949 ( .A(n14060), .ZN(n14061) );
  INV_X1 U15950 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17646) );
  NAND2_X1 U15951 ( .A1(n14065), .A2(n11421), .ZN(n14066) );
  AND2_X1 U15952 ( .A1(n14228), .A2(n14066), .ZN(n19146) );
  INV_X1 U15953 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14068) );
  NAND2_X1 U15954 ( .A1(n14071), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14072) );
  NAND2_X1 U15955 ( .A1(n14072), .A2(n17821), .ZN(n15632) );
  INV_X1 U15956 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n14073) );
  OAI21_X1 U15957 ( .B1(n14414), .B2(n15632), .A(n14073), .ZN(n18015) );
  NOR2_X1 U15958 ( .A1(n14074), .A2(n14123), .ZN(n14075) );
  NOR2_X1 U15959 ( .A1(n15699), .A2(n14075), .ZN(n14076) );
  MUX2_X1 U15960 ( .A(n18015), .B(n14076), .S(n12085), .Z(n17843) );
  NAND2_X1 U15961 ( .A1(n17843), .A2(n12005), .ZN(n14084) );
  INV_X1 U15962 ( .A(n14077), .ZN(n14078) );
  OAI21_X1 U15963 ( .B1(n14079), .B2(n14124), .A(n14078), .ZN(n14082) );
  NAND3_X1 U15964 ( .A1(n14082), .A2(n14081), .A3(n14080), .ZN(n14083) );
  AND2_X1 U15965 ( .A1(n14083), .A2(n14137), .ZN(n15636) );
  NAND2_X1 U15966 ( .A1(n15636), .A2(n14155), .ZN(n14166) );
  NAND2_X1 U15967 ( .A1(n14084), .A2(n14166), .ZN(n14086) );
  INV_X1 U15968 ( .A(n14085), .ZN(n15637) );
  NAND2_X1 U15969 ( .A1(n14086), .A2(n15637), .ZN(n15631) );
  XNOR2_X1 U15970 ( .A(n14087), .B(n14067), .ZN(n14112) );
  NAND2_X1 U15971 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n14112), .ZN(
        n14113) );
  NAND2_X1 U15972 ( .A1(n14104), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16153) );
  XOR2_X1 U15973 ( .A(n14091), .B(n14090), .Z(n14092) );
  OR2_X1 U15974 ( .A1(n15222), .A2(n14092), .ZN(n14098) );
  XNOR2_X1 U15975 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n14092), .ZN(
        n15227) );
  XOR2_X1 U15976 ( .A(n14094), .B(n14093), .Z(n14095) );
  NOR2_X1 U15977 ( .A1(n16307), .A2(n19224), .ZN(n16309) );
  NAND2_X1 U15978 ( .A1(n14095), .A2(n16309), .ZN(n14097) );
  XOR2_X1 U15979 ( .A(n14095), .B(n16309), .Z(n15142) );
  NAND2_X1 U15980 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15142), .ZN(
        n14096) );
  NAND2_X1 U15981 ( .A1(n14097), .A2(n14096), .ZN(n15226) );
  NAND2_X1 U15982 ( .A1(n15227), .A2(n15226), .ZN(n15225) );
  NAND2_X1 U15983 ( .A1(n14098), .A2(n15225), .ZN(n17914) );
  NOR2_X1 U15984 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17914), .ZN(
        n14099) );
  NAND2_X1 U15985 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17914), .ZN(
        n17913) );
  OR2_X1 U15986 ( .A1(n14100), .A2(n14101), .ZN(n14103) );
  NAND2_X1 U15987 ( .A1(n14103), .A2(n14102), .ZN(n14105) );
  NAND2_X1 U15988 ( .A1(n16153), .A2(n14105), .ZN(n14109) );
  INV_X1 U15989 ( .A(n14105), .ZN(n16155) );
  NAND3_X1 U15990 ( .A1(n14106), .A2(n14109), .A3(n16154), .ZN(n14110) );
  INV_X1 U15991 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19294) );
  XNOR2_X1 U15992 ( .A(n19294), .B(n14112), .ZN(n17936) );
  INV_X1 U15993 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17761) );
  XNOR2_X1 U15994 ( .A(n17761), .B(n14114), .ZN(n17750) );
  NAND2_X1 U15995 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n14114), .ZN(
        n14115) );
  NAND3_X1 U15996 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17693) );
  NOR3_X1 U15997 ( .A1(n17696), .A2(n17695), .A3(n17693), .ZN(n19254) );
  AND2_X1 U15998 ( .A1(n19254), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14116) );
  NOR2_X1 U15999 ( .A1(n19353), .A2(n11354), .ZN(n14117) );
  OAI21_X1 U16000 ( .B1(n17258), .B2(n14118), .A(n17154), .ZN(n19152) );
  INV_X1 U16001 ( .A(n19152), .ZN(n14225) );
  NAND2_X1 U16002 ( .A1(n20262), .A2(n14123), .ZN(n14122) );
  AOI22_X1 U16003 ( .A1(n14122), .A2(n14121), .B1(n20262), .B2(n14119), .ZN(
        n14126) );
  OAI21_X1 U16004 ( .B1(n14124), .B2(n14123), .A(n12005), .ZN(n14125) );
  OAI21_X1 U16005 ( .B1(n14126), .B2(n11156), .A(n14125), .ZN(n14135) );
  NAND2_X1 U16006 ( .A1(n11354), .A2(n15129), .ZN(n14128) );
  NAND2_X1 U16007 ( .A1(n14128), .A2(n14127), .ZN(n14130) );
  AOI21_X1 U16008 ( .B1(n14130), .B2(n14129), .A(n14131), .ZN(n14134) );
  INV_X1 U16009 ( .A(n14131), .ZN(n14132) );
  OAI21_X1 U16010 ( .B1(n14132), .B2(n12003), .A(n14137), .ZN(n14133) );
  AOI21_X1 U16011 ( .B1(n14135), .B2(n14134), .A(n14133), .ZN(n14136) );
  MUX2_X1 U16012 ( .A(n17821), .B(n14136), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n14151) );
  NOR2_X1 U16013 ( .A1(n12085), .A2(n19916), .ZN(n15131) );
  OAI21_X1 U16014 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n17901), .ZN(n19010) );
  NOR2_X1 U16015 ( .A1(n15131), .A2(n19010), .ZN(n15070) );
  INV_X1 U16016 ( .A(n15070), .ZN(n14139) );
  AND2_X1 U16017 ( .A1(n20002), .A2(n18021), .ZN(n19014) );
  OR2_X1 U16018 ( .A1(n19014), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14141) );
  OAI21_X1 U16019 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n12085), .A(n15712), 
        .ZN(n14142) );
  INV_X1 U16020 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19150) );
  NOR2_X1 U16021 ( .A1(n19325), .A2(n19150), .ZN(n14221) );
  AOI21_X1 U16022 ( .B1(n18003), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14221), .ZN(n14143) );
  OAI21_X1 U16023 ( .B1(n18001), .B2(n19159), .A(n14143), .ZN(n14144) );
  AND2_X1 U16024 ( .A1(n15641), .A2(n11354), .ZN(n14148) );
  NAND2_X1 U16025 ( .A1(n14148), .A2(n22312), .ZN(n15126) );
  OAI21_X1 U16026 ( .B1(n15699), .B2(n11354), .A(n15126), .ZN(n14147) );
  NAND3_X1 U16027 ( .A1(n14147), .A2(n11342), .A3(n19342), .ZN(n14174) );
  INV_X1 U16028 ( .A(n14148), .ZN(n14150) );
  OAI211_X1 U16029 ( .C1(n11156), .C2(n14151), .A(n14150), .B(n14149), .ZN(
        n14172) );
  NAND2_X1 U16030 ( .A1(n14149), .A2(n20262), .ZN(n14182) );
  INV_X1 U16031 ( .A(n14152), .ZN(n14153) );
  AOI21_X1 U16032 ( .B1(n14154), .B2(n14182), .A(n14153), .ZN(n14158) );
  OAI21_X1 U16033 ( .B1(n14156), .B2(n19835), .A(n14155), .ZN(n14191) );
  OAI211_X1 U16034 ( .C1(n14158), .C2(n11342), .A(n14191), .B(n14157), .ZN(
        n14159) );
  INV_X1 U16035 ( .A(n14159), .ZN(n14163) );
  NAND2_X1 U16036 ( .A1(n14160), .A2(n20207), .ZN(n14161) );
  NAND2_X1 U16037 ( .A1(n15634), .A2(n14161), .ZN(n14162) );
  NOR2_X1 U16038 ( .A1(n15699), .A2(n22317), .ZN(n14169) );
  NAND3_X1 U16039 ( .A1(n14169), .A2(n14164), .A3(n22312), .ZN(n14165) );
  AND2_X1 U16040 ( .A1(n14184), .A2(n14165), .ZN(n15658) );
  NAND2_X1 U16041 ( .A1(n17843), .A2(n11354), .ZN(n14167) );
  NAND2_X1 U16042 ( .A1(n14167), .A2(n14166), .ZN(n14168) );
  NAND2_X1 U16043 ( .A1(n14168), .A2(n15637), .ZN(n14171) );
  NAND3_X1 U16044 ( .A1(n14169), .A2(n14164), .A3(n11354), .ZN(n14170) );
  NAND2_X1 U16045 ( .A1(n14174), .A2(n14173), .ZN(n14175) );
  INV_X1 U16046 ( .A(n14178), .ZN(n14176) );
  AOI21_X1 U16047 ( .B1(n14180), .B2(n14120), .A(n15644), .ZN(n14181) );
  INV_X1 U16048 ( .A(n14182), .ZN(n14183) );
  NOR2_X1 U16049 ( .A1(n15206), .A2(n19224), .ZN(n16157) );
  NOR2_X1 U16050 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n16157), .ZN(
        n14207) );
  INV_X1 U16051 ( .A(n14207), .ZN(n14185) );
  NAND2_X1 U16052 ( .A1(n14215), .A2(n19325), .ZN(n19225) );
  OAI21_X1 U16053 ( .B1(n17759), .B2(n14185), .A(n19225), .ZN(n16160) );
  INV_X1 U16054 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19317) );
  NOR3_X1 U16055 ( .A1(n19339), .A2(n16166), .A3(n19317), .ZN(n19296) );
  NAND4_X1 U16056 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n19296), .ZN(n14209) );
  INV_X1 U16057 ( .A(n14209), .ZN(n14186) );
  NOR2_X1 U16058 ( .A1(n17759), .A2(n14186), .ZN(n14187) );
  OR2_X1 U16059 ( .A1(n16160), .A2(n14187), .ZN(n14279) );
  NAND2_X1 U16060 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19254), .ZN(
        n17655) );
  INV_X1 U16061 ( .A(n17655), .ZN(n14188) );
  NOR2_X1 U16062 ( .A1(n17759), .A2(n14188), .ZN(n14189) );
  NOR2_X1 U16063 ( .A1(n14279), .A2(n14189), .ZN(n17659) );
  NAND2_X1 U16064 ( .A1(n14190), .A2(n11354), .ZN(n15675) );
  NAND2_X1 U16065 ( .A1(n15675), .A2(n14191), .ZN(n14192) );
  NAND2_X1 U16066 ( .A1(n14192), .A2(n16031), .ZN(n14201) );
  INV_X1 U16067 ( .A(n12004), .ZN(n14193) );
  NAND2_X1 U16068 ( .A1(n14193), .A2(n20112), .ZN(n14194) );
  INV_X1 U16069 ( .A(n15153), .ZN(n19009) );
  AOI22_X1 U16070 ( .A1(n14194), .A2(n19009), .B1(n11156), .B2(n11342), .ZN(
        n14198) );
  AND2_X1 U16071 ( .A1(n14195), .A2(n12004), .ZN(n14196) );
  OAI21_X1 U16072 ( .B1(n15157), .B2(n14196), .A(n15156), .ZN(n14197) );
  AND2_X1 U16073 ( .A1(n14198), .A2(n14197), .ZN(n14200) );
  NAND3_X1 U16074 ( .A1(n14201), .A2(n14200), .A3(n14199), .ZN(n15681) );
  NOR2_X1 U16075 ( .A1(n15681), .A2(n14202), .ZN(n14203) );
  NOR3_X1 U16076 ( .A1(n19268), .A2(n17662), .A3(n17663), .ZN(n14273) );
  NAND2_X1 U16077 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n16157), .ZN(
        n14208) );
  OR2_X1 U16078 ( .A1(n14209), .A2(n14208), .ZN(n17654) );
  INV_X1 U16079 ( .A(n17756), .ZN(n17656) );
  OAI21_X1 U16080 ( .B1(n17654), .B2(n17655), .A(n17656), .ZN(n14204) );
  OAI21_X1 U16081 ( .B1(n19237), .B2(n14273), .A(n14204), .ZN(n14205) );
  INV_X1 U16082 ( .A(n14205), .ZN(n14206) );
  AND2_X1 U16083 ( .A1(n17659), .A2(n14206), .ZN(n17647) );
  INV_X1 U16084 ( .A(n14273), .ZN(n14218) );
  NAND3_X1 U16085 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19254), .A3(
        n19253), .ZN(n17675) );
  NOR2_X1 U16086 ( .A1(n14218), .A2(n17675), .ZN(n14210) );
  NAND2_X1 U16087 ( .A1(n17646), .A2(n14210), .ZN(n17644) );
  AND2_X1 U16088 ( .A1(n17647), .A2(n17644), .ZN(n17634) );
  INV_X1 U16089 ( .A(n14211), .ZN(n14213) );
  AND2_X1 U16090 ( .A1(n14213), .A2(n14212), .ZN(n15648) );
  AOI21_X1 U16091 ( .B1(n11354), .B2(n15635), .A(n15648), .ZN(n14214) );
  NOR2_X1 U16092 ( .A1(n17365), .A2(n14216), .ZN(n14217) );
  OR2_X1 U16093 ( .A1(n17156), .A2(n14217), .ZN(n19151) );
  INV_X1 U16094 ( .A(n19151), .ZN(n14222) );
  XNOR2_X1 U16095 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14219) );
  OR3_X1 U16096 ( .A1(n17646), .A2(n14218), .A3(n17675), .ZN(n17636) );
  NOR2_X1 U16097 ( .A1(n14219), .A2(n17636), .ZN(n14220) );
  AOI211_X1 U16098 ( .C1(n19281), .C2(n14222), .A(n14221), .B(n14220), .ZN(
        n14223) );
  OAI21_X1 U16099 ( .B1(n17634), .B2(n14068), .A(n14223), .ZN(n14224) );
  NAND2_X1 U16100 ( .A1(n14228), .A2(n11277), .ZN(n14229) );
  NAND2_X1 U16101 ( .A1(n14242), .A2(n14229), .ZN(n17166) );
  OR2_X1 U16102 ( .A1(n17166), .A2(n14324), .ZN(n14230) );
  INV_X1 U16103 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17621) );
  NAND2_X1 U16104 ( .A1(n14230), .A2(n17621), .ZN(n17472) );
  NAND4_X1 U16105 ( .A1(n14062), .A2(n18005), .A3(n14231), .A4(n17503), .ZN(
        n14232) );
  NOR2_X1 U16106 ( .A1(n14232), .A2(n17483), .ZN(n14233) );
  OAI211_X1 U16107 ( .C1(n14234), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n17472), .B(n14233), .ZN(n14240) );
  NAND2_X1 U16108 ( .A1(n14234), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14239) );
  AND3_X1 U16109 ( .A1(n14236), .A2(n14235), .A3(n17685), .ZN(n14237) );
  OR3_X1 U16110 ( .A1(n17166), .A2(n14324), .A3(n17621), .ZN(n17471) );
  INV_X1 U16111 ( .A(n17464), .ZN(n14245) );
  NAND2_X1 U16112 ( .A1(n14242), .A2(n14241), .ZN(n14243) );
  NAND2_X1 U16113 ( .A1(n14249), .A2(n14243), .ZN(n19161) );
  OR2_X1 U16114 ( .A1(n19161), .A2(n14324), .ZN(n14246) );
  INV_X1 U16115 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17615) );
  XNOR2_X1 U16116 ( .A(n14246), .B(n17615), .ZN(n17465) );
  NAND2_X1 U16117 ( .A1(n14246), .A2(n17615), .ZN(n14247) );
  XNOR2_X1 U16118 ( .A(n14249), .B(n14248), .ZN(n17149) );
  NAND2_X1 U16119 ( .A1(n17149), .A2(n14067), .ZN(n14250) );
  INV_X1 U16120 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17453) );
  OR2_X1 U16121 ( .A1(n14250), .A2(n17453), .ZN(n17449) );
  INV_X1 U16122 ( .A(n14251), .ZN(n14254) );
  INV_X1 U16123 ( .A(n14252), .ZN(n14253) );
  NAND2_X1 U16124 ( .A1(n14254), .A2(n14253), .ZN(n14255) );
  NAND2_X1 U16125 ( .A1(n14261), .A2(n14255), .ZN(n17122) );
  INV_X1 U16126 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17442) );
  NOR2_X1 U16127 ( .A1(n14256), .A2(n17442), .ZN(n17440) );
  XNOR2_X1 U16128 ( .A(n14258), .B(n14257), .ZN(n19203) );
  NAND2_X1 U16129 ( .A1(n19203), .A2(n14067), .ZN(n14259) );
  XNOR2_X1 U16130 ( .A(n14259), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17423) );
  XNOR2_X1 U16131 ( .A(n14261), .B(n11423), .ZN(n19187) );
  NAND2_X1 U16132 ( .A1(n19187), .A2(n14067), .ZN(n14262) );
  INV_X1 U16133 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17567) );
  NAND2_X1 U16134 ( .A1(n14262), .A2(n17567), .ZN(n17435) );
  NAND2_X1 U16135 ( .A1(n17423), .A2(n17435), .ZN(n14263) );
  INV_X1 U16136 ( .A(n14314), .ZN(n17425) );
  NAND3_X1 U16137 ( .A1(n19203), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14067), .ZN(n14265) );
  INV_X1 U16138 ( .A(n19187), .ZN(n14264) );
  INV_X1 U16139 ( .A(n14266), .ZN(n14267) );
  NAND2_X1 U16140 ( .A1(n11227), .A2(n14267), .ZN(n14268) );
  NAND2_X1 U16141 ( .A1(n11207), .A2(n14268), .ZN(n17118) );
  NOR2_X1 U16142 ( .A1(n17118), .A2(n14324), .ZN(n14310) );
  NAND2_X1 U16143 ( .A1(n11207), .A2(n14270), .ZN(n14271) );
  NAND4_X1 U16144 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14273), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17619) );
  NOR3_X1 U16145 ( .A1(n17621), .A2(n17655), .A3(n17619), .ZN(n14293) );
  NAND2_X1 U16146 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17596) );
  INV_X1 U16147 ( .A(n17596), .ZN(n14294) );
  AND2_X1 U16148 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n14294), .ZN(
        n14274) );
  NAND2_X1 U16149 ( .A1(n17616), .A2(n14274), .ZN(n17577) );
  INV_X1 U16150 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17566) );
  NOR2_X1 U16151 ( .A1(n17567), .A2(n17566), .ZN(n17565) );
  INV_X1 U16152 ( .A(n17565), .ZN(n14275) );
  INV_X1 U16153 ( .A(n17556), .ZN(n14285) );
  NAND2_X1 U16154 ( .A1(n14285), .A2(n14311), .ZN(n14304) );
  NOR2_X1 U16155 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17596), .ZN(
        n14276) );
  NAND2_X1 U16156 ( .A1(n17616), .A2(n14276), .ZN(n17590) );
  INV_X1 U16157 ( .A(n17654), .ZN(n14277) );
  NOR2_X1 U16158 ( .A1(n17756), .A2(n14277), .ZN(n14278) );
  NOR2_X1 U16159 ( .A1(n14279), .A2(n14278), .ZN(n17743) );
  INV_X1 U16160 ( .A(n19237), .ZN(n16161) );
  INV_X1 U16161 ( .A(n14293), .ZN(n14280) );
  NAND2_X1 U16162 ( .A1(n16161), .A2(n14280), .ZN(n14281) );
  NAND2_X1 U16163 ( .A1(n17743), .A2(n14281), .ZN(n17626) );
  NOR2_X1 U16164 ( .A1(n19237), .A2(n14294), .ZN(n14282) );
  NOR2_X1 U16165 ( .A1(n17626), .A2(n14282), .ZN(n17584) );
  NAND2_X1 U16166 ( .A1(n17590), .A2(n17584), .ZN(n17579) );
  NOR2_X1 U16167 ( .A1(n19237), .A2(n17565), .ZN(n14283) );
  NOR2_X1 U16168 ( .A1(n17579), .A2(n14283), .ZN(n14329) );
  NAND2_X1 U16169 ( .A1(n14304), .A2(n14329), .ZN(n17549) );
  XNOR2_X1 U16170 ( .A(n11213), .B(n14284), .ZN(n17206) );
  NAND3_X1 U16171 ( .A1(n14285), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n11414), .ZN(n14291) );
  NOR2_X1 U16172 ( .A1(n14286), .A2(n14287), .ZN(n14288) );
  OR2_X2 U16173 ( .A1(n17286), .A2(n14288), .ZN(n17296) );
  INV_X1 U16174 ( .A(n17296), .ZN(n14289) );
  INV_X1 U16175 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n18095) );
  NOR2_X1 U16176 ( .A1(n19325), .A2(n18095), .ZN(n16341) );
  AOI21_X1 U16177 ( .B1(n14289), .B2(n19281), .A(n16341), .ZN(n14290) );
  OAI211_X1 U16178 ( .C1(n17206), .C2(n19285), .A(n14291), .B(n14290), .ZN(
        n14292) );
  AOI21_X1 U16179 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17549), .A(
        n14292), .ZN(n14296) );
  AND2_X2 U16180 ( .A1(n17716), .A2(n14293), .ZN(n17475) );
  XNOR2_X1 U16181 ( .A(n17411), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16344) );
  NAND2_X1 U16182 ( .A1(n16344), .A2(n19271), .ZN(n14295) );
  OAI21_X1 U16183 ( .B1(n16346), .B2(n19304), .A(n14297), .ZN(P2_U3018) );
  XNOR2_X1 U16184 ( .A(n14298), .B(n14311), .ZN(n14337) );
  NAND2_X1 U16185 ( .A1(n14337), .A2(n19335), .ZN(n14309) );
  AND2_X1 U16186 ( .A1(n17219), .A2(n14299), .ZN(n14300) );
  OR2_X1 U16187 ( .A1(n14300), .A2(n11213), .ZN(n17211) );
  INV_X1 U16188 ( .A(n17211), .ZN(n17115) );
  AND2_X1 U16189 ( .A1(n11209), .A2(n14301), .ZN(n14302) );
  OR2_X1 U16190 ( .A1(n14302), .A2(n14286), .ZN(n17303) );
  INV_X2 U16191 ( .A(n19325), .ZN(n19282) );
  NAND2_X1 U16192 ( .A1(n19282), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n14338) );
  OAI21_X1 U16193 ( .B1(n17303), .B2(n19327), .A(n14338), .ZN(n14303) );
  AOI21_X1 U16194 ( .B1(n17115), .B2(n19329), .A(n14303), .ZN(n14305) );
  OAI211_X1 U16195 ( .C1(n14329), .C2(n14311), .A(n14305), .B(n14304), .ZN(
        n14307) );
  OAI21_X1 U16196 ( .B1(n11220), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17411), .ZN(n14341) );
  NOR2_X1 U16197 ( .A1(n14341), .A2(n19332), .ZN(n14306) );
  NOR2_X1 U16198 ( .A1(n14307), .A2(n14306), .ZN(n14308) );
  NAND2_X1 U16199 ( .A1(n14309), .A2(n14308), .ZN(P2_U3019) );
  NAND2_X1 U16200 ( .A1(n14269), .A2(n14311), .ZN(n14312) );
  NAND2_X1 U16201 ( .A1(n14314), .A2(n11744), .ZN(n14319) );
  OAI21_X1 U16202 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n14315), .ZN(n14317) );
  XNOR2_X1 U16203 ( .A(n14321), .B(n14320), .ZN(n14323) );
  INV_X1 U16204 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14322) );
  OAI21_X1 U16205 ( .B1(n14323), .B2(n14324), .A(n14322), .ZN(n17407) );
  NAND2_X1 U16206 ( .A1(n17409), .A2(n17407), .ZN(n17396) );
  INV_X1 U16207 ( .A(n14323), .ZN(n19219) );
  NAND3_X1 U16208 ( .A1(n19219), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14067), .ZN(n17408) );
  INV_X1 U16209 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14328) );
  OAI21_X1 U16210 ( .B1(n14325), .B2(n14324), .A(n14328), .ZN(n17393) );
  AND2_X1 U16211 ( .A1(n14067), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14326) );
  NAND2_X1 U16212 ( .A1(n14327), .A2(n14326), .ZN(n17394) );
  NAND3_X1 U16213 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14332) );
  NOR2_X1 U16214 ( .A1(n14328), .A2(n14332), .ZN(n17540) );
  OAI21_X1 U16215 ( .B1(n19237), .B2(n17540), .A(n14329), .ZN(n17539) );
  INV_X1 U16216 ( .A(n17539), .ZN(n14334) );
  NAND2_X1 U16217 ( .A1(n16323), .A2(n19329), .ZN(n14330) );
  NAND2_X1 U16218 ( .A1(n19282), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n16317) );
  OAI211_X1 U16219 ( .C1(n16359), .C2(n19327), .A(n14330), .B(n16317), .ZN(
        n14331) );
  INV_X1 U16220 ( .A(n14331), .ZN(n14333) );
  INV_X1 U16221 ( .A(n14335), .ZN(n14336) );
  NAND2_X1 U16222 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17548) );
  NOR2_X1 U16223 ( .A1(n17411), .A2(n17548), .ZN(n17413) );
  NAND2_X1 U16224 ( .A1(n11220), .A2(n17540), .ZN(n17401) );
  OAI21_X1 U16225 ( .B1(n17413), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n17401), .ZN(n16320) );
  NAND2_X1 U16226 ( .A1(n14337), .A2(n17983), .ZN(n14345) );
  OAI21_X1 U16227 ( .B1(n17987), .B2(n17111), .A(n14338), .ZN(n14340) );
  NOR2_X1 U16228 ( .A1(n17211), .A2(n15057), .ZN(n14339) );
  AOI211_X1 U16229 ( .C1(n18002), .C2(n17105), .A(n14340), .B(n14339), .ZN(
        n14343) );
  OR2_X1 U16230 ( .A1(n14341), .A2(n17996), .ZN(n14342) );
  NAND2_X1 U16231 ( .A1(n14345), .A2(n14344), .ZN(P2_U2987) );
  NAND2_X1 U16232 ( .A1(n15439), .A2(n16306), .ZN(n14352) );
  NAND2_X1 U16233 ( .A1(n11997), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14347) );
  NAND2_X1 U16234 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19980) );
  INV_X1 U16235 ( .A(n19980), .ZN(n19872) );
  INV_X1 U16236 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18034) );
  NAND2_X1 U16237 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18034), .ZN(
        n19964) );
  INV_X1 U16238 ( .A(n19964), .ZN(n14348) );
  NAND2_X1 U16239 ( .A1(n19872), .A2(n14348), .ZN(n19929) );
  NOR3_X1 U16240 ( .A1(n12216), .A2(n19884), .A3(n18034), .ZN(n19839) );
  INV_X1 U16241 ( .A(n19839), .ZN(n19845) );
  INV_X1 U16242 ( .A(n20325), .ZN(n14349) );
  NAND2_X1 U16243 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14349), .ZN(
        n14350) );
  NAND2_X1 U16244 ( .A1(n19929), .A2(n14350), .ZN(n19967) );
  INV_X1 U16245 ( .A(n20002), .ZN(n19846) );
  AOI21_X1 U16246 ( .B1(n14369), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n15080), .ZN(n14351) );
  INV_X1 U16247 ( .A(n14588), .ZN(n14354) );
  NOR2_X1 U16248 ( .A1(n14354), .A2(n17800), .ZN(n14355) );
  NAND2_X1 U16249 ( .A1(n14356), .A2(n16068), .ZN(n15058) );
  INV_X1 U16250 ( .A(n15058), .ZN(n14376) );
  AOI22_X1 U16251 ( .A1(n14369), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n14357), .B2(n20000), .ZN(n14358) );
  NAND2_X1 U16252 ( .A1(n14588), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14359) );
  NAND2_X1 U16253 ( .A1(n15069), .A2(n14359), .ZN(n14366) );
  INV_X1 U16254 ( .A(n14359), .ZN(n14360) );
  NAND2_X1 U16255 ( .A1(n17771), .A2(n14360), .ZN(n14361) );
  NAND2_X1 U16256 ( .A1(n14362), .A2(n16306), .ZN(n14365) );
  NAND2_X1 U16257 ( .A1(n12216), .A2(n20000), .ZN(n19965) );
  AND2_X1 U16258 ( .A1(n19980), .A2(n19965), .ZN(n15071) );
  NAND2_X1 U16259 ( .A1(n14357), .A2(n15071), .ZN(n19939) );
  INV_X1 U16260 ( .A(n19939), .ZN(n14363) );
  AOI21_X1 U16261 ( .B1(n14369), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n14363), .ZN(n14364) );
  NAND2_X1 U16262 ( .A1(n14368), .A2(n16306), .ZN(n14371) );
  XNOR2_X1 U16263 ( .A(n19980), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15072) );
  AOI22_X1 U16264 ( .A1(n14369), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n14357), .B2(n15072), .ZN(n14370) );
  NAND2_X1 U16265 ( .A1(n14588), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14372) );
  INV_X1 U16266 ( .A(n14372), .ZN(n14373) );
  NAND2_X1 U16267 ( .A1(n14374), .A2(n14373), .ZN(n14375) );
  NAND2_X1 U16268 ( .A1(n14376), .A2(n15059), .ZN(n14378) );
  NAND2_X1 U16269 ( .A1(n11997), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14377) );
  NAND2_X1 U16270 ( .A1(n16239), .A2(n16245), .ZN(n16244) );
  AOI22_X1 U16271 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14386) );
  AOI22_X1 U16272 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14385) );
  AOI22_X1 U16273 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14384) );
  AOI22_X1 U16274 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14383) );
  NAND4_X1 U16275 ( .A1(n14386), .A2(n14385), .A3(n14384), .A4(n14383), .ZN(
        n14392) );
  AOI22_X1 U16276 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14390) );
  AOI22_X1 U16277 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14389) );
  AOI22_X1 U16278 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14388) );
  AOI22_X1 U16279 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14387) );
  NAND4_X1 U16280 ( .A1(n14390), .A2(n14389), .A3(n14388), .A4(n14387), .ZN(
        n14391) );
  NOR2_X1 U16281 ( .A1(n14392), .A2(n14391), .ZN(n17273) );
  INV_X1 U16282 ( .A(n17273), .ZN(n14393) );
  AOI22_X1 U16283 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U16284 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14396) );
  AOI22_X1 U16285 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14395) );
  AOI22_X1 U16286 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14394) );
  NAND4_X1 U16287 ( .A1(n14397), .A2(n14396), .A3(n14395), .A4(n14394), .ZN(
        n14403) );
  AOI22_X1 U16288 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14401) );
  AOI22_X1 U16289 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14400) );
  AOI22_X1 U16290 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14399) );
  AOI22_X1 U16291 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14398) );
  NAND4_X1 U16292 ( .A1(n14401), .A2(n14400), .A3(n14399), .A4(n14398), .ZN(
        n14402) );
  AOI22_X1 U16293 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U16294 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U16295 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14405) );
  AOI22_X1 U16296 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14404) );
  NAND4_X1 U16297 ( .A1(n14407), .A2(n14406), .A3(n14405), .A4(n14404), .ZN(
        n14413) );
  AOI22_X1 U16298 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14411) );
  AOI22_X1 U16299 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14410) );
  AOI22_X1 U16300 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14409) );
  AOI22_X1 U16301 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14408) );
  NAND4_X1 U16302 ( .A1(n14411), .A2(n14410), .A3(n14409), .A4(n14408), .ZN(
        n14412) );
  NOR2_X1 U16303 ( .A1(n14413), .A2(n14412), .ZN(n17261) );
  AOI22_X1 U16304 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14418) );
  AOI22_X1 U16305 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U16306 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14416) );
  AOI22_X1 U16307 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14415) );
  NAND4_X1 U16308 ( .A1(n14418), .A2(n14417), .A3(n14416), .A4(n14415), .ZN(
        n14424) );
  AOI22_X1 U16309 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14422) );
  AOI22_X1 U16310 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14421) );
  AOI22_X1 U16311 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14420) );
  AOI22_X1 U16312 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14419) );
  NAND4_X1 U16313 ( .A1(n14422), .A2(n14421), .A3(n14420), .A4(n14419), .ZN(
        n14423) );
  AOI22_X1 U16314 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14428) );
  AOI22_X1 U16315 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14427) );
  AOI22_X1 U16316 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14426) );
  AOI22_X1 U16317 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14425) );
  NAND4_X1 U16318 ( .A1(n14428), .A2(n14427), .A3(n14426), .A4(n14425), .ZN(
        n14434) );
  AOI22_X1 U16319 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14432) );
  AOI22_X1 U16320 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14431) );
  AOI22_X1 U16321 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14430) );
  AOI22_X1 U16322 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14429) );
  NAND4_X1 U16323 ( .A1(n14432), .A2(n14431), .A3(n14430), .A4(n14429), .ZN(
        n14433) );
  AOI22_X1 U16324 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U16325 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14437) );
  AOI22_X1 U16326 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14436) );
  AOI22_X1 U16327 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14435) );
  NAND4_X1 U16328 ( .A1(n14438), .A2(n14437), .A3(n14436), .A4(n14435), .ZN(
        n14444) );
  AOI22_X1 U16329 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14442) );
  AOI22_X1 U16330 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14441) );
  AOI22_X1 U16331 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14440) );
  AOI22_X1 U16332 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14439) );
  NAND4_X1 U16333 ( .A1(n14442), .A2(n14441), .A3(n14440), .A4(n14439), .ZN(
        n14443) );
  NOR2_X1 U16334 ( .A1(n14444), .A2(n14443), .ZN(n17248) );
  INV_X1 U16335 ( .A(n14445), .ZN(n14449) );
  INV_X1 U16336 ( .A(n14446), .ZN(n14448) );
  OAI22_X1 U16337 ( .A1(n14450), .A2(n14449), .B1(n14448), .B2(n14447), .ZN(
        n14466) );
  INV_X1 U16338 ( .A(n14479), .ZN(n14454) );
  INV_X1 U16339 ( .A(n14451), .ZN(n14453) );
  OAI22_X1 U16340 ( .A1(n14455), .A2(n14454), .B1(n14453), .B2(n14452), .ZN(
        n14465) );
  INV_X1 U16341 ( .A(n14414), .ZN(n14459) );
  INV_X1 U16342 ( .A(n14456), .ZN(n14458) );
  OAI22_X1 U16343 ( .A1(n14459), .A2(n20062), .B1(n14458), .B2(n14457), .ZN(
        n14464) );
  INV_X1 U16344 ( .A(n14460), .ZN(n14461) );
  INV_X1 U16345 ( .A(n14480), .ZN(n15654) );
  OAI22_X1 U16346 ( .A1(n14462), .A2(n14461), .B1(n15654), .B2(n20036), .ZN(
        n14463) );
  NOR4_X1 U16347 ( .A1(n14466), .A2(n14465), .A3(n14464), .A4(n14463), .ZN(
        n14478) );
  AOI22_X1 U16348 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14477) );
  AOI22_X1 U16349 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14476) );
  INV_X1 U16350 ( .A(n14489), .ZN(n14468) );
  NOR2_X1 U16351 ( .A1(n14468), .A2(n14467), .ZN(n14474) );
  INV_X1 U16352 ( .A(n14488), .ZN(n14471) );
  INV_X1 U16353 ( .A(n14487), .ZN(n14470) );
  OAI22_X1 U16354 ( .A1(n14472), .A2(n14471), .B1(n14470), .B2(n14469), .ZN(
        n14473) );
  AOI211_X1 U16355 ( .C1(n14490), .C2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n14474), .B(n14473), .ZN(n14475) );
  NAND4_X1 U16356 ( .A1(n14478), .A2(n14477), .A3(n14476), .A4(n14475), .ZN(
        n17241) );
  AOI22_X1 U16357 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n14445), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14484) );
  AOI22_X1 U16358 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n14479), .B1(
        n14451), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14483) );
  AOI22_X1 U16359 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14456), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14482) );
  AOI22_X1 U16360 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n14460), .B1(
        n14480), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14481) );
  NAND4_X1 U16361 ( .A1(n14484), .A2(n14483), .A3(n14482), .A4(n14481), .ZN(
        n14496) );
  AOI22_X1 U16362 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11174), .B1(
        n14485), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14494) );
  AOI22_X1 U16363 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n14486), .B1(
        n11819), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14493) );
  AOI22_X1 U16364 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n14488), .B1(
        n14487), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14492) );
  AOI22_X1 U16365 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n14490), .B1(
        n14489), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14491) );
  NAND4_X1 U16366 ( .A1(n14494), .A2(n14493), .A3(n14492), .A4(n14491), .ZN(
        n14495) );
  NOR2_X1 U16367 ( .A1(n14496), .A2(n14495), .ZN(n14513) );
  AOI22_X1 U16368 ( .A1(n14626), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14504) );
  AND2_X1 U16369 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14498) );
  OR2_X1 U16370 ( .A1(n14498), .A2(n14497), .ZN(n14639) );
  INV_X1 U16371 ( .A(n14639), .ZN(n14594) );
  NAND2_X1 U16372 ( .A1(n11786), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14500) );
  NAND2_X1 U16373 ( .A1(n14636), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14499) );
  AND3_X1 U16374 ( .A1(n14594), .A2(n14500), .A3(n14499), .ZN(n14503) );
  AOI22_X1 U16375 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14627), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14502) );
  AOI22_X1 U16376 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14617), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14501) );
  NAND4_X1 U16377 ( .A1(n14504), .A2(n14503), .A3(n14502), .A4(n14501), .ZN(
        n14512) );
  AOI22_X1 U16378 ( .A1(n14626), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14510) );
  AOI22_X1 U16379 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14627), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14509) );
  AOI22_X1 U16380 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14617), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14508) );
  NAND2_X1 U16381 ( .A1(n11786), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n14506) );
  NAND2_X1 U16382 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14505) );
  AND3_X1 U16383 ( .A1(n14506), .A2(n14505), .A3(n14639), .ZN(n14507) );
  NAND4_X1 U16384 ( .A1(n14510), .A2(n14509), .A3(n14508), .A4(n14507), .ZN(
        n14511) );
  NAND2_X1 U16385 ( .A1(n14512), .A2(n14511), .ZN(n14514) );
  XNOR2_X1 U16386 ( .A(n14513), .B(n14514), .ZN(n17237) );
  INV_X1 U16387 ( .A(n14513), .ZN(n14516) );
  INV_X1 U16388 ( .A(n14514), .ZN(n14515) );
  NAND2_X1 U16389 ( .A1(n14516), .A2(n14515), .ZN(n14531) );
  AOI22_X1 U16390 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14616), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14522) );
  NAND2_X1 U16391 ( .A1(n11786), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14518) );
  NAND2_X1 U16392 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n14517) );
  AND3_X1 U16393 ( .A1(n14594), .A2(n14518), .A3(n14517), .ZN(n14521) );
  AOI22_X1 U16394 ( .A1(n14626), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14627), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14520) );
  AOI22_X1 U16395 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14617), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14519) );
  NAND4_X1 U16396 ( .A1(n14522), .A2(n14521), .A3(n14520), .A4(n14519), .ZN(
        n14530) );
  AOI22_X1 U16397 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14528) );
  AOI22_X1 U16398 ( .A1(n14626), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14627), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14527) );
  AOI22_X1 U16399 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11786), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14526) );
  INV_X1 U16400 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n20303) );
  NAND2_X1 U16401 ( .A1(n14617), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14524) );
  NAND2_X1 U16402 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14523) );
  AND3_X1 U16403 ( .A1(n14524), .A2(n14523), .A3(n14639), .ZN(n14525) );
  NAND4_X1 U16404 ( .A1(n14528), .A2(n14527), .A3(n14526), .A4(n14525), .ZN(
        n14529) );
  NAND2_X1 U16405 ( .A1(n14530), .A2(n14529), .ZN(n14533) );
  NOR2_X1 U16406 ( .A1(n14531), .A2(n14533), .ZN(n14549) );
  INV_X1 U16407 ( .A(n14531), .ZN(n14532) );
  NAND2_X1 U16408 ( .A1(n14588), .A2(n14532), .ZN(n14534) );
  AOI22_X1 U16409 ( .A1(n14549), .A2(n11354), .B1(n14534), .B2(n14533), .ZN(
        n17233) );
  AOI22_X1 U16410 ( .A1(n14626), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14540) );
  NAND2_X1 U16411 ( .A1(n11786), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14536) );
  NAND2_X1 U16412 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14535) );
  AND3_X1 U16413 ( .A1(n14594), .A2(n14536), .A3(n14535), .ZN(n14539) );
  AOI22_X1 U16414 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14538) );
  AOI22_X1 U16415 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14617), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14537) );
  NAND4_X1 U16416 ( .A1(n14540), .A2(n14539), .A3(n14538), .A4(n14537), .ZN(
        n14548) );
  AOI22_X1 U16417 ( .A1(n14626), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14546) );
  AOI22_X1 U16418 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14627), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14545) );
  AOI22_X1 U16419 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14617), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14544) );
  NAND2_X1 U16420 ( .A1(n11786), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14542) );
  NAND2_X1 U16421 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14541) );
  AND3_X1 U16422 ( .A1(n14542), .A2(n14541), .A3(n14639), .ZN(n14543) );
  NAND4_X1 U16423 ( .A1(n14546), .A2(n14545), .A3(n14544), .A4(n14543), .ZN(
        n14547) );
  AND2_X1 U16424 ( .A1(n14548), .A2(n14547), .ZN(n14551) );
  NAND2_X1 U16425 ( .A1(n14549), .A2(n14551), .ZN(n14572) );
  OAI211_X1 U16426 ( .C1(n14549), .C2(n14551), .A(n14588), .B(n14572), .ZN(
        n14553) );
  INV_X1 U16427 ( .A(n14553), .ZN(n14550) );
  INV_X1 U16428 ( .A(n14551), .ZN(n14552) );
  NOR2_X1 U16429 ( .A1(n11354), .A2(n14552), .ZN(n17226) );
  AOI22_X1 U16430 ( .A1(n14626), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14559) );
  NAND2_X1 U16431 ( .A1(n11786), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14555) );
  NAND2_X1 U16432 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14554) );
  AND3_X1 U16433 ( .A1(n14594), .A2(n14555), .A3(n14554), .ZN(n14558) );
  AOI22_X1 U16434 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14557) );
  AOI22_X1 U16435 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14617), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14556) );
  NAND4_X1 U16436 ( .A1(n14559), .A2(n14558), .A3(n14557), .A4(n14556), .ZN(
        n14567) );
  AOI22_X1 U16437 ( .A1(n14626), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14565) );
  AOI22_X1 U16438 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14627), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14564) );
  AOI22_X1 U16439 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14617), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14563) );
  NAND2_X1 U16440 ( .A1(n11786), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n14561) );
  NAND2_X1 U16441 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14560) );
  AND3_X1 U16442 ( .A1(n14561), .A2(n14560), .A3(n14639), .ZN(n14562) );
  NAND4_X1 U16443 ( .A1(n14565), .A2(n14564), .A3(n14563), .A4(n14562), .ZN(
        n14566) );
  AND2_X1 U16444 ( .A1(n14567), .A2(n14566), .ZN(n14570) );
  XNOR2_X1 U16445 ( .A(n14572), .B(n14570), .ZN(n14568) );
  NAND2_X1 U16446 ( .A1(n14120), .A2(n14570), .ZN(n17215) );
  INV_X1 U16447 ( .A(n14570), .ZN(n14571) );
  OR2_X1 U16448 ( .A1(n14572), .A2(n14571), .ZN(n14587) );
  INV_X1 U16449 ( .A(n14587), .ZN(n14590) );
  AOI22_X1 U16450 ( .A1(n14626), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14578) );
  AOI22_X1 U16451 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14627), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14577) );
  AOI22_X1 U16452 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14617), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14576) );
  NAND2_X1 U16453 ( .A1(n11786), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n14574) );
  NAND2_X1 U16454 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14573) );
  AND3_X1 U16455 ( .A1(n14574), .A2(n14573), .A3(n14639), .ZN(n14575) );
  NAND4_X1 U16456 ( .A1(n14578), .A2(n14577), .A3(n14576), .A4(n14575), .ZN(
        n14586) );
  AOI22_X1 U16457 ( .A1(n14626), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14584) );
  NAND2_X1 U16458 ( .A1(n11786), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14580) );
  NAND2_X1 U16459 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n14579) );
  AND3_X1 U16460 ( .A1(n14594), .A2(n14580), .A3(n14579), .ZN(n14583) );
  AOI22_X1 U16461 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14582) );
  AOI22_X1 U16462 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14617), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14581) );
  NAND4_X1 U16463 ( .A1(n14584), .A2(n14583), .A3(n14582), .A4(n14581), .ZN(
        n14585) );
  NAND2_X1 U16464 ( .A1(n14586), .A2(n14585), .ZN(n14591) );
  INV_X1 U16465 ( .A(n14591), .ZN(n14589) );
  OAI211_X1 U16466 ( .C1(n14590), .C2(n14589), .A(n14588), .B(n17203), .ZN(
        n14607) );
  AOI22_X1 U16467 ( .A1(n14626), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14598) );
  NAND2_X1 U16468 ( .A1(n11786), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14593) );
  NAND2_X1 U16469 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14592) );
  AND3_X1 U16470 ( .A1(n14594), .A2(n14593), .A3(n14592), .ZN(n14597) );
  AOI22_X1 U16471 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14627), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14596) );
  AOI22_X1 U16472 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14617), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14595) );
  NAND4_X1 U16473 ( .A1(n14598), .A2(n14597), .A3(n14596), .A4(n14595), .ZN(
        n14606) );
  AOI22_X1 U16474 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14604) );
  AOI22_X1 U16475 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14603) );
  AOI22_X1 U16476 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14617), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14602) );
  NAND2_X1 U16477 ( .A1(n11786), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n14600) );
  NAND2_X1 U16478 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14599) );
  AND3_X1 U16479 ( .A1(n14600), .A2(n14599), .A3(n14639), .ZN(n14601) );
  NAND4_X1 U16480 ( .A1(n14604), .A2(n14603), .A3(n14602), .A4(n14601), .ZN(
        n14605) );
  AND2_X1 U16481 ( .A1(n14606), .A2(n14605), .ZN(n17204) );
  INV_X1 U16482 ( .A(n17203), .ZN(n14608) );
  NAND3_X1 U16483 ( .A1(n14608), .A2(n17204), .A3(n11354), .ZN(n17195) );
  AOI22_X1 U16484 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14616), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14610) );
  AOI22_X1 U16485 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14609) );
  NAND2_X1 U16486 ( .A1(n14610), .A2(n14609), .ZN(n14624) );
  AOI22_X1 U16487 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11786), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14612) );
  AOI21_X1 U16488 ( .B1(n14630), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n14639), .ZN(n14611) );
  OAI211_X1 U16489 ( .C1(n11760), .C2(n20036), .A(n14612), .B(n14611), .ZN(
        n14623) );
  AOI22_X1 U16490 ( .A1(n14613), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14615) );
  AOI22_X1 U16491 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14614) );
  NAND2_X1 U16492 ( .A1(n14615), .A2(n14614), .ZN(n14622) );
  AOI22_X1 U16493 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11786), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14620) );
  NAND2_X1 U16494 ( .A1(n14617), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n14619) );
  NAND2_X1 U16495 ( .A1(n14630), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n14618) );
  NAND4_X1 U16496 ( .A1(n14620), .A2(n14639), .A3(n14619), .A4(n14618), .ZN(
        n14621) );
  OAI22_X1 U16497 ( .A1(n14624), .A2(n14623), .B1(n14622), .B2(n14621), .ZN(
        n17194) );
  AOI21_X1 U16498 ( .B1(n17197), .B2(n17195), .A(n17194), .ZN(n14647) );
  AOI22_X1 U16499 ( .A1(n14626), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14629) );
  AOI22_X1 U16500 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14627), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14628) );
  NAND2_X1 U16501 ( .A1(n14629), .A2(n14628), .ZN(n14644) );
  INV_X1 U16502 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n19898) );
  AOI21_X1 U16503 ( .B1(n14630), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n14639), .ZN(n14632) );
  AOI22_X1 U16504 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14631) );
  OAI211_X1 U16505 ( .C1(n11760), .C2(n19898), .A(n14632), .B(n14631), .ZN(
        n14643) );
  AOI22_X1 U16506 ( .A1(n11170), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14625), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14635) );
  AOI22_X1 U16507 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14633), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14634) );
  NAND2_X1 U16508 ( .A1(n14635), .A2(n14634), .ZN(n14642) );
  AOI22_X1 U16509 ( .A1(n14616), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11976), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14640) );
  NAND2_X1 U16510 ( .A1(n14617), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14638) );
  NAND2_X1 U16511 ( .A1(n14636), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14637) );
  NAND4_X1 U16512 ( .A1(n14640), .A2(n14639), .A3(n14638), .A4(n14637), .ZN(
        n14641) );
  OAI22_X1 U16513 ( .A1(n14644), .A2(n14643), .B1(n14642), .B2(n14641), .ZN(
        n14645) );
  INV_X1 U16514 ( .A(n14645), .ZN(n14646) );
  XNOR2_X1 U16515 ( .A(n14647), .B(n14646), .ZN(n16363) );
  INV_X1 U16516 ( .A(n15641), .ZN(n14648) );
  NAND2_X1 U16517 ( .A1(n14648), .A2(n15648), .ZN(n15659) );
  INV_X1 U16518 ( .A(n14202), .ZN(n14649) );
  NAND2_X1 U16519 ( .A1(n15659), .A2(n14649), .ZN(n14650) );
  NAND2_X1 U16520 ( .A1(n16323), .A2(n17281), .ZN(n14653) );
  NAND2_X1 U16521 ( .A1(n14651), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14652) );
  OAI21_X1 U16522 ( .B1(n16363), .B2(n17272), .A(n14654), .ZN(P2_U2857) );
  INV_X1 U16523 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n20616) );
  INV_X1 U16524 ( .A(keyinput_228), .ZN(n14655) );
  INV_X1 U16525 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n22234) );
  INV_X1 U16526 ( .A(keyinput_227), .ZN(n14814) );
  INV_X1 U16527 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n16700) );
  INV_X1 U16528 ( .A(keyinput_220), .ZN(n14806) );
  INV_X1 U16529 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20559) );
  INV_X1 U16530 ( .A(keyinput_190), .ZN(n14765) );
  INV_X1 U16531 ( .A(keyinput_173), .ZN(n14735) );
  INV_X1 U16532 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17878) );
  INV_X1 U16533 ( .A(keyinput_172), .ZN(n14734) );
  INV_X1 U16534 ( .A(keyinput_171), .ZN(n14733) );
  INV_X1 U16535 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21963) );
  INV_X1 U16536 ( .A(keyinput_170), .ZN(n14731) );
  INV_X1 U16537 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20710) );
  INV_X1 U16538 ( .A(keyinput_169), .ZN(n14729) );
  INV_X1 U16539 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22779) );
  INV_X1 U16540 ( .A(DATAI_15_), .ZN(n14682) );
  INV_X1 U16541 ( .A(keyinput_145), .ZN(n14681) );
  INV_X1 U16542 ( .A(DATAI_25_), .ZN(n15588) );
  INV_X1 U16543 ( .A(keyinput_135), .ZN(n14667) );
  INV_X1 U16544 ( .A(DATAI_26_), .ZN(n15597) );
  INV_X1 U16545 ( .A(keyinput_134), .ZN(n14666) );
  INV_X1 U16546 ( .A(DATAI_29_), .ZN(n15575) );
  XNOR2_X1 U16547 ( .A(keyinput_131), .B(n15575), .ZN(n14659) );
  AOI22_X1 U16548 ( .A1(DATAI_31_), .A2(keyinput_129), .B1(
        P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_128), .ZN(n14660) );
  AOI22_X1 U16549 ( .A1(DATAI_24_), .A2(keyinput_136), .B1(DATAI_23_), .B2(
        keyinput_137), .ZN(n14668) );
  OAI221_X1 U16550 ( .B1(DATAI_24_), .B2(keyinput_136), .C1(DATAI_23_), .C2(
        keyinput_137), .A(n14668), .ZN(n14671) );
  INV_X1 U16551 ( .A(DATAI_22_), .ZN(n15579) );
  OAI22_X1 U16552 ( .A1(n15579), .A2(keyinput_138), .B1(keyinput_139), .B2(
        DATAI_21_), .ZN(n14669) );
  AOI221_X1 U16553 ( .B1(n15579), .B2(keyinput_138), .C1(DATAI_21_), .C2(
        keyinput_139), .A(n14669), .ZN(n14670) );
  OAI21_X1 U16554 ( .B1(n14672), .B2(n14671), .A(n14670), .ZN(n14676) );
  INV_X1 U16555 ( .A(DATAI_20_), .ZN(n15568) );
  INV_X1 U16556 ( .A(keyinput_140), .ZN(n14673) );
  INV_X1 U16557 ( .A(DATAI_19_), .ZN(n15561) );
  OAI22_X1 U16558 ( .A1(n15561), .A2(keyinput_141), .B1(DATAI_18_), .B2(
        keyinput_142), .ZN(n14677) );
  AOI221_X1 U16559 ( .B1(n15561), .B2(keyinput_141), .C1(keyinput_142), .C2(
        DATAI_18_), .A(n14677), .ZN(n14680) );
  INV_X1 U16560 ( .A(DATAI_17_), .ZN(n15587) );
  INV_X1 U16561 ( .A(DATAI_16_), .ZN(n15543) );
  AOI22_X1 U16562 ( .A1(n15587), .A2(keyinput_143), .B1(n15543), .B2(
        keyinput_144), .ZN(n14678) );
  OAI221_X1 U16563 ( .B1(n15587), .B2(keyinput_143), .C1(n15543), .C2(
        keyinput_144), .A(n14678), .ZN(n14679) );
  INV_X1 U16564 ( .A(DATAI_12_), .ZN(n14684) );
  INV_X1 U16565 ( .A(DATAI_11_), .ZN(n16278) );
  AOI22_X1 U16566 ( .A1(n14684), .A2(keyinput_148), .B1(n16278), .B2(
        keyinput_149), .ZN(n14683) );
  OAI221_X1 U16567 ( .B1(n14684), .B2(keyinput_148), .C1(n16278), .C2(
        keyinput_149), .A(n14683), .ZN(n14689) );
  INV_X1 U16568 ( .A(DATAI_14_), .ZN(n14687) );
  INV_X1 U16569 ( .A(DATAI_13_), .ZN(n14686) );
  AOI22_X1 U16570 ( .A1(n14687), .A2(keyinput_146), .B1(n14686), .B2(
        keyinput_147), .ZN(n14685) );
  OAI221_X1 U16571 ( .B1(n14687), .B2(keyinput_146), .C1(n14686), .C2(
        keyinput_147), .A(n14685), .ZN(n14688) );
  XNOR2_X1 U16572 ( .A(DATAI_10_), .B(keyinput_150), .ZN(n14697) );
  INV_X1 U16573 ( .A(DATAI_9_), .ZN(n14692) );
  INV_X1 U16574 ( .A(DATAI_8_), .ZN(n14691) );
  OAI22_X1 U16575 ( .A1(n14692), .A2(keyinput_151), .B1(n14691), .B2(
        keyinput_152), .ZN(n14690) );
  AOI221_X1 U16576 ( .B1(n14692), .B2(keyinput_151), .C1(keyinput_152), .C2(
        n14691), .A(n14690), .ZN(n14695) );
  OAI22_X1 U16577 ( .A1(DATAI_6_), .A2(keyinput_154), .B1(keyinput_153), .B2(
        DATAI_7_), .ZN(n14693) );
  AOI221_X1 U16578 ( .B1(DATAI_6_), .B2(keyinput_154), .C1(DATAI_7_), .C2(
        keyinput_153), .A(n14693), .ZN(n14694) );
  AND2_X1 U16579 ( .A1(n14695), .A2(n14694), .ZN(n14696) );
  OAI21_X1 U16580 ( .B1(n14698), .B2(n14697), .A(n14696), .ZN(n14701) );
  OAI22_X1 U16581 ( .A1(DATAI_4_), .A2(keyinput_156), .B1(DATAI_5_), .B2(
        keyinput_155), .ZN(n14699) );
  AOI221_X1 U16582 ( .B1(DATAI_4_), .B2(keyinput_156), .C1(keyinput_155), .C2(
        DATAI_5_), .A(n14699), .ZN(n14700) );
  NAND2_X1 U16583 ( .A1(n14701), .A2(n14700), .ZN(n14711) );
  INV_X1 U16584 ( .A(DATAI_1_), .ZN(n14703) );
  AOI22_X1 U16585 ( .A1(DATAI_0_), .A2(keyinput_160), .B1(n14703), .B2(
        keyinput_159), .ZN(n14702) );
  OAI221_X1 U16586 ( .B1(DATAI_0_), .B2(keyinput_160), .C1(n14703), .C2(
        keyinput_159), .A(n14702), .ZN(n14706) );
  NAND2_X1 U16587 ( .A1(DATAI_2_), .A2(keyinput_158), .ZN(n14704) );
  INV_X1 U16588 ( .A(DATAI_3_), .ZN(n14708) );
  AOI22_X1 U16589 ( .A1(n22334), .A2(keyinput_161), .B1(keyinput_157), .B2(
        n14708), .ZN(n14707) );
  OAI221_X1 U16590 ( .B1(n22334), .B2(keyinput_161), .C1(n14708), .C2(
        keyinput_157), .A(n14707), .ZN(n14709) );
  NAND2_X1 U16591 ( .A1(n14711), .A2(n14710), .ZN(n14714) );
  INV_X1 U16592 ( .A(NA), .ZN(n22336) );
  OAI22_X1 U16593 ( .A1(n22336), .A2(keyinput_162), .B1(keyinput_163), .B2(
        BS16), .ZN(n14712) );
  AOI221_X1 U16594 ( .B1(n22336), .B2(keyinput_162), .C1(BS16), .C2(
        keyinput_163), .A(n14712), .ZN(n14713) );
  NAND2_X1 U16595 ( .A1(n14714), .A2(n14713), .ZN(n14719) );
  INV_X1 U16596 ( .A(READY1), .ZN(n14715) );
  AND2_X1 U16597 ( .A1(n14715), .A2(keyinput_164), .ZN(n14717) );
  NOR2_X1 U16598 ( .A1(n14717), .A2(n14716), .ZN(n14718) );
  NAND2_X1 U16599 ( .A1(n14719), .A2(n14718), .ZN(n14723) );
  INV_X1 U16600 ( .A(READY2), .ZN(n14914) );
  INV_X1 U16601 ( .A(keyinput_165), .ZN(n14720) );
  INV_X1 U16602 ( .A(n14721), .ZN(n14722) );
  OAI22_X1 U16603 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(keyinput_166), .B1(
        keyinput_168), .B2(P1_CODEFETCH_REG_SCAN_IN), .ZN(n14724) );
  AOI221_X1 U16604 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_166), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(keyinput_168), .A(n14724), .ZN(n14728)
         );
  AOI221_X1 U16605 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(n14731), .C1(n20710), .C2(
        keyinput_170), .A(n14730), .ZN(n14732) );
  INV_X1 U16606 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20779) );
  INV_X1 U16607 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n22246) );
  AOI22_X1 U16608 ( .A1(n20779), .A2(keyinput_175), .B1(n22246), .B2(
        keyinput_174), .ZN(n14736) );
  OAI221_X1 U16609 ( .B1(n20779), .B2(keyinput_175), .C1(n22246), .C2(
        keyinput_174), .A(n14736), .ZN(n14740) );
  INV_X1 U16610 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20599) );
  INV_X1 U16611 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20602) );
  OAI22_X1 U16612 ( .A1(n20599), .A2(keyinput_177), .B1(n20602), .B2(
        keyinput_176), .ZN(n14737) );
  AOI221_X1 U16613 ( .B1(n20599), .B2(keyinput_177), .C1(keyinput_176), .C2(
        n20602), .A(n14737), .ZN(n14739) );
  XNOR2_X1 U16614 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_178), .ZN(
        n14738) );
  INV_X1 U16615 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20579) );
  INV_X1 U16616 ( .A(keyinput_179), .ZN(n14741) );
  OAI22_X1 U16617 ( .A1(n20579), .A2(n14741), .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_179), .ZN(n14742) );
  INV_X1 U16618 ( .A(n14742), .ZN(n14745) );
  INV_X1 U16619 ( .A(keyinput_180), .ZN(n14743) );
  INV_X1 U16620 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20576) );
  INV_X1 U16621 ( .A(keyinput_181), .ZN(n14747) );
  OAI22_X1 U16622 ( .A1(n20576), .A2(n14747), .B1(P1_REIP_REG_30__SCAN_IN), 
        .B2(keyinput_181), .ZN(n14750) );
  OAI22_X1 U16623 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(keyinput_183), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_182), .ZN(n14748) );
  AOI221_X1 U16624 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_183), .C1(
        keyinput_182), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14748), .ZN(n14749)
         );
  INV_X1 U16625 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n22085) );
  INV_X1 U16626 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20568) );
  OAI22_X1 U16627 ( .A1(n20568), .A2(keyinput_185), .B1(keyinput_186), .B2(
        P1_REIP_REG_25__SCAN_IN), .ZN(n14753) );
  AOI221_X1 U16628 ( .B1(n20568), .B2(keyinput_185), .C1(
        P1_REIP_REG_25__SCAN_IN), .C2(keyinput_186), .A(n14753), .ZN(n14754)
         );
  INV_X1 U16629 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20565) );
  AND2_X1 U16630 ( .A1(n20565), .A2(keyinput_187), .ZN(n14756) );
  INV_X1 U16631 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20563) );
  INV_X1 U16632 ( .A(keyinput_188), .ZN(n14757) );
  INV_X1 U16633 ( .A(n14758), .ZN(n14761) );
  INV_X1 U16634 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20561) );
  INV_X1 U16635 ( .A(keyinput_189), .ZN(n14759) );
  INV_X1 U16636 ( .A(n14763), .ZN(n14764) );
  OAI221_X1 U16637 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_190), .C1(
        n20559), .C2(n14765), .A(n14764), .ZN(n14770) );
  INV_X1 U16638 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n22067) );
  OAI22_X1 U16639 ( .A1(n22067), .A2(keyinput_192), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_191), .ZN(n14766) );
  AOI221_X1 U16640 ( .B1(n22067), .B2(keyinput_192), .C1(keyinput_191), .C2(
        P1_REIP_REG_20__SCAN_IN), .A(n14766), .ZN(n14769) );
  INV_X1 U16641 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20551) );
  AOI22_X1 U16642 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(keyinput_193), .B1(
        n20551), .B2(keyinput_194), .ZN(n14767) );
  OAI221_X1 U16643 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(keyinput_193), .C1(
        n20551), .C2(keyinput_194), .A(n14767), .ZN(n14768) );
  INV_X1 U16644 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n22227) );
  INV_X1 U16645 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20549) );
  AOI22_X1 U16646 ( .A1(n22227), .A2(keyinput_195), .B1(keyinput_196), .B2(
        n20549), .ZN(n14771) );
  OAI221_X1 U16647 ( .B1(n22227), .B2(keyinput_195), .C1(n20549), .C2(
        keyinput_196), .A(n14771), .ZN(n14774) );
  INV_X1 U16648 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21966) );
  OAI22_X1 U16649 ( .A1(n21966), .A2(keyinput_198), .B1(keyinput_197), .B2(
        P1_REIP_REG_14__SCAN_IN), .ZN(n14772) );
  AOI221_X1 U16650 ( .B1(n21966), .B2(keyinput_198), .C1(
        P1_REIP_REG_14__SCAN_IN), .C2(keyinput_197), .A(n14772), .ZN(n14773)
         );
  OAI22_X1 U16651 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(keyinput_200), .B1(
        keyinput_199), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n14775) );
  AOI221_X1 U16652 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(keyinput_200), .C1(
        P1_REIP_REG_12__SCAN_IN), .C2(keyinput_199), .A(n14775), .ZN(n14779)
         );
  INV_X1 U16653 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n22164) );
  AOI22_X1 U16654 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(keyinput_202), .B1(n22164), .B2(keyinput_203), .ZN(n14781) );
  OAI221_X1 U16655 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(keyinput_202), .C1(
        n22164), .C2(keyinput_203), .A(n14781), .ZN(n14784) );
  INV_X1 U16656 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20536) );
  INV_X1 U16657 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n22158) );
  OAI22_X1 U16658 ( .A1(n20536), .A2(keyinput_205), .B1(n22158), .B2(
        keyinput_204), .ZN(n14782) );
  AOI221_X1 U16659 ( .B1(n20536), .B2(keyinput_205), .C1(keyinput_204), .C2(
        n22158), .A(n14782), .ZN(n14783) );
  OAI21_X1 U16660 ( .B1(n14785), .B2(n14784), .A(n14783), .ZN(n14788) );
  INV_X1 U16661 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20535) );
  OAI22_X1 U16662 ( .A1(n20535), .A2(keyinput_206), .B1(keyinput_207), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n14786) );
  AOI221_X1 U16663 ( .B1(n20535), .B2(keyinput_206), .C1(
        P1_REIP_REG_4__SCAN_IN), .C2(keyinput_207), .A(n14786), .ZN(n14787) );
  NAND2_X1 U16664 ( .A1(n14788), .A2(n14787), .ZN(n14793) );
  AOI22_X1 U16665 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(keyinput_208), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(keyinput_210), .ZN(n14789) );
  OAI221_X1 U16666 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(keyinput_208), .C1(
        P1_REIP_REG_1__SCAN_IN), .C2(keyinput_210), .A(n14789), .ZN(n14791) );
  NAND2_X1 U16667 ( .A1(n14793), .A2(n14792), .ZN(n14799) );
  INV_X1 U16668 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n16686) );
  INV_X1 U16669 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14795) );
  OAI22_X1 U16670 ( .A1(n16686), .A2(keyinput_212), .B1(n14795), .B2(
        keyinput_211), .ZN(n14794) );
  AOI221_X1 U16671 ( .B1(n16686), .B2(keyinput_212), .C1(keyinput_211), .C2(
        n14795), .A(n14794), .ZN(n14797) );
  XNOR2_X1 U16672 ( .A(P1_EBX_REG_30__SCAN_IN), .B(keyinput_213), .ZN(n14796)
         );
  INV_X1 U16673 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n16691) );
  INV_X1 U16674 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n16692) );
  OAI22_X1 U16675 ( .A1(n16691), .A2(keyinput_214), .B1(n16692), .B2(
        keyinput_215), .ZN(n14800) );
  AOI221_X1 U16676 ( .B1(n16691), .B2(keyinput_214), .C1(keyinput_215), .C2(
        n16692), .A(n14800), .ZN(n14802) );
  NOR2_X1 U16677 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput_216), .ZN(n14801)
         );
  INV_X1 U16678 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n16518) );
  AOI22_X1 U16679 ( .A1(P1_EBX_REG_26__SCAN_IN), .A2(keyinput_217), .B1(n16518), .B2(keyinput_218), .ZN(n14803) );
  OAI221_X1 U16680 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(keyinput_217), .C1(
        n16518), .C2(keyinput_218), .A(n14803), .ZN(n14804) );
  AOI221_X1 U16681 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(keyinput_220), .C1(
        n16700), .C2(n14806), .A(n14805), .ZN(n14813) );
  INV_X1 U16682 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n16702) );
  AOI22_X1 U16683 ( .A1(P1_EBX_REG_22__SCAN_IN), .A2(keyinput_221), .B1(n16702), .B2(keyinput_222), .ZN(n14807) );
  OAI221_X1 U16684 ( .B1(P1_EBX_REG_22__SCAN_IN), .B2(keyinput_221), .C1(
        n16702), .C2(keyinput_222), .A(n14807), .ZN(n14812) );
  INV_X1 U16685 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n16711) );
  OAI22_X1 U16686 ( .A1(n16711), .A2(keyinput_226), .B1(keyinput_225), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n14808) );
  AOI221_X1 U16687 ( .B1(n16711), .B2(keyinput_226), .C1(
        P1_EBX_REG_18__SCAN_IN), .C2(keyinput_225), .A(n14808), .ZN(n14811) );
  OAI22_X1 U16688 ( .A1(P1_EBX_REG_20__SCAN_IN), .A2(keyinput_223), .B1(
        P1_EBX_REG_19__SCAN_IN), .B2(keyinput_224), .ZN(n14809) );
  AOI221_X1 U16689 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(keyinput_223), .C1(
        keyinput_224), .C2(P1_EBX_REG_19__SCAN_IN), .A(n14809), .ZN(n14810) );
  INV_X1 U16690 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n20620) );
  INV_X1 U16691 ( .A(keyinput_229), .ZN(n14815) );
  OAI22_X1 U16692 ( .A1(n20620), .A2(n14815), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(keyinput_229), .ZN(n14816) );
  INV_X1 U16693 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n16720) );
  INV_X1 U16694 ( .A(keyinput_230), .ZN(n14817) );
  INV_X1 U16695 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n22210) );
  INV_X1 U16696 ( .A(keyinput_231), .ZN(n14819) );
  INV_X1 U16697 ( .A(n14820), .ZN(n14821) );
  OAI21_X1 U16698 ( .B1(n14822), .B2(n14818), .A(n14821), .ZN(n14826) );
  INV_X1 U16699 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n16290) );
  INV_X1 U16700 ( .A(keyinput_232), .ZN(n14823) );
  NAND2_X1 U16701 ( .A1(n14826), .A2(n14825), .ZN(n14832) );
  INV_X1 U16702 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n20611) );
  OAI22_X1 U16703 ( .A1(n20611), .A2(keyinput_233), .B1(P1_EBX_REG_9__SCAN_IN), 
        .B2(keyinput_234), .ZN(n14827) );
  AOI221_X1 U16704 ( .B1(n20611), .B2(keyinput_233), .C1(keyinput_234), .C2(
        P1_EBX_REG_9__SCAN_IN), .A(n14827), .ZN(n14831) );
  XOR2_X1 U16705 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_236), .Z(n14830) );
  INV_X1 U16706 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n16197) );
  INV_X1 U16707 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n22138) );
  AOI22_X1 U16708 ( .A1(n16197), .A2(keyinput_235), .B1(keyinput_237), .B2(
        n22138), .ZN(n14828) );
  OAI221_X1 U16709 ( .B1(n16197), .B2(keyinput_235), .C1(n22138), .C2(
        keyinput_237), .A(n14828), .ZN(n14829) );
  AOI211_X1 U16710 ( .C1(n14832), .C2(n14831), .A(n14830), .B(n14829), .ZN(
        n14839) );
  INV_X1 U16711 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n20607) );
  INV_X1 U16712 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n22129) );
  AOI22_X1 U16713 ( .A1(n20607), .A2(keyinput_240), .B1(keyinput_242), .B2(
        n22129), .ZN(n14833) );
  OAI221_X1 U16714 ( .B1(n20607), .B2(keyinput_240), .C1(n22129), .C2(
        keyinput_242), .A(n14833), .ZN(n14836) );
  INV_X1 U16715 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n15459) );
  AOI22_X1 U16716 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(keyinput_238), .B1(n15459), 
        .B2(keyinput_241), .ZN(n14834) );
  OAI221_X1 U16717 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(keyinput_238), .C1(n15459), .C2(keyinput_241), .A(n14834), .ZN(n14835) );
  AOI211_X1 U16718 ( .C1(keyinput_239), .C2(P1_EBX_REG_4__SCAN_IN), .A(n14836), 
        .B(n14835), .ZN(n14837) );
  OAI21_X1 U16719 ( .B1(keyinput_239), .B2(P1_EBX_REG_4__SCAN_IN), .A(n14837), 
        .ZN(n14838) );
  NOR2_X1 U16720 ( .A1(n14839), .A2(n14838), .ZN(n14846) );
  OAI22_X1 U16721 ( .A1(P1_EAX_REG_31__SCAN_IN), .A2(keyinput_244), .B1(
        P1_EBX_REG_0__SCAN_IN), .B2(keyinput_243), .ZN(n14840) );
  AOI221_X1 U16722 ( .B1(P1_EAX_REG_31__SCAN_IN), .B2(keyinput_244), .C1(
        keyinput_243), .C2(P1_EBX_REG_0__SCAN_IN), .A(n14840), .ZN(n14842) );
  XNOR2_X1 U16723 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_245), .ZN(n14841)
         );
  INV_X1 U16724 ( .A(keyinput_246), .ZN(n14843) );
  INV_X1 U16725 ( .A(n14844), .ZN(n14845) );
  OAI21_X1 U16726 ( .B1(n14846), .B2(n11738), .A(n14845), .ZN(n14859) );
  OAI22_X1 U16727 ( .A1(n13533), .A2(keyinput_247), .B1(P1_EAX_REG_26__SCAN_IN), .B2(keyinput_249), .ZN(n14847) );
  AOI221_X1 U16728 ( .B1(n13533), .B2(keyinput_247), .C1(keyinput_249), .C2(
        P1_EAX_REG_26__SCAN_IN), .A(n14847), .ZN(n14850) );
  OAI22_X1 U16729 ( .A1(n13465), .A2(keyinput_250), .B1(n13442), .B2(
        keyinput_251), .ZN(n14848) );
  AOI221_X1 U16730 ( .B1(n13465), .B2(keyinput_250), .C1(keyinput_251), .C2(
        n13442), .A(n14848), .ZN(n14849) );
  OAI211_X1 U16731 ( .C1(P1_EAX_REG_27__SCAN_IN), .C2(keyinput_248), .A(n14850), .B(n14849), .ZN(n14851) );
  AOI21_X1 U16732 ( .B1(P1_EAX_REG_27__SCAN_IN), .B2(keyinput_248), .A(n14851), 
        .ZN(n14858) );
  OAI22_X1 U16733 ( .A1(n15175), .A2(keyinput_254), .B1(keyinput_253), .B2(
        P1_EAX_REG_22__SCAN_IN), .ZN(n14854) );
  AOI22_X1 U16734 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(keyinput_253), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(keyinput_252), .ZN(n14852) );
  OAI21_X1 U16735 ( .B1(keyinput_252), .B2(P1_EAX_REG_23__SCAN_IN), .A(n14852), 
        .ZN(n14853) );
  NOR2_X1 U16736 ( .A1(n14854), .A2(n14853), .ZN(n14856) );
  AOI21_X1 U16737 ( .B1(n14859), .B2(n14858), .A(n14857), .ZN(n15047) );
  XNOR2_X1 U16738 ( .A(keyinput_55), .B(P1_REIP_REG_28__SCAN_IN), .ZN(n14861)
         );
  XNOR2_X1 U16739 ( .A(keyinput_54), .B(P1_REIP_REG_29__SCAN_IN), .ZN(n14860)
         );
  NAND2_X1 U16740 ( .A1(n14861), .A2(n14860), .ZN(n14937) );
  INV_X1 U16741 ( .A(n14937), .ZN(n14943) );
  XNOR2_X1 U16742 ( .A(keyinput_53), .B(P1_REIP_REG_30__SCAN_IN), .ZN(n14942)
         );
  XOR2_X1 U16743 ( .A(keyinput_56), .B(P1_REIP_REG_27__SCAN_IN), .Z(n14941) );
  XOR2_X1 U16744 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_0), .Z(n14865)
         );
  XOR2_X1 U16745 ( .A(keyinput_1), .B(DATAI_31_), .Z(n14864) );
  XNOR2_X1 U16746 ( .A(keyinput_3), .B(DATAI_29_), .ZN(n14863) );
  XOR2_X1 U16747 ( .A(keyinput_2), .B(DATAI_30_), .Z(n14862) );
  AOI211_X1 U16748 ( .C1(n14865), .C2(n14864), .A(n14863), .B(n14862), .ZN(
        n14868) );
  XOR2_X1 U16749 ( .A(keyinput_5), .B(DATAI_27_), .Z(n14867) );
  XNOR2_X1 U16750 ( .A(keyinput_4), .B(DATAI_28_), .ZN(n14866) );
  NOR3_X1 U16751 ( .A1(n14868), .A2(n14867), .A3(n14866), .ZN(n14871) );
  XNOR2_X1 U16752 ( .A(keyinput_6), .B(DATAI_26_), .ZN(n14870) );
  XNOR2_X1 U16753 ( .A(keyinput_7), .B(DATAI_25_), .ZN(n14869) );
  OAI21_X1 U16754 ( .B1(n14871), .B2(n14870), .A(n14869), .ZN(n14874) );
  XNOR2_X1 U16755 ( .A(keyinput_9), .B(DATAI_23_), .ZN(n14873) );
  XNOR2_X1 U16756 ( .A(keyinput_8), .B(DATAI_24_), .ZN(n14872) );
  NAND3_X1 U16757 ( .A1(n14874), .A2(n14873), .A3(n14872), .ZN(n14877) );
  XOR2_X1 U16758 ( .A(keyinput_11), .B(DATAI_21_), .Z(n14876) );
  XNOR2_X1 U16759 ( .A(keyinput_10), .B(DATAI_22_), .ZN(n14875) );
  NAND3_X1 U16760 ( .A1(n14877), .A2(n14876), .A3(n14875), .ZN(n14881) );
  XOR2_X1 U16761 ( .A(keyinput_12), .B(DATAI_20_), .Z(n14880) );
  XOR2_X1 U16762 ( .A(keyinput_13), .B(DATAI_19_), .Z(n14879) );
  XOR2_X1 U16763 ( .A(keyinput_14), .B(DATAI_18_), .Z(n14878) );
  AOI211_X1 U16764 ( .C1(n14881), .C2(n14880), .A(n14879), .B(n14878), .ZN(
        n14884) );
  XOR2_X1 U16765 ( .A(keyinput_15), .B(DATAI_17_), .Z(n14883) );
  XNOR2_X1 U16766 ( .A(DATAI_16_), .B(keyinput_16), .ZN(n14882) );
  NOR3_X1 U16767 ( .A1(n14884), .A2(n14883), .A3(n14882), .ZN(n14891) );
  XNOR2_X1 U16768 ( .A(keyinput_17), .B(DATAI_15_), .ZN(n14890) );
  XOR2_X1 U16769 ( .A(keyinput_18), .B(DATAI_14_), .Z(n14888) );
  XNOR2_X1 U16770 ( .A(keyinput_19), .B(DATAI_13_), .ZN(n14887) );
  XNOR2_X1 U16771 ( .A(DATAI_11_), .B(keyinput_21), .ZN(n14886) );
  XNOR2_X1 U16772 ( .A(keyinput_20), .B(DATAI_12_), .ZN(n14885) );
  NOR4_X1 U16773 ( .A1(n14888), .A2(n14887), .A3(n14886), .A4(n14885), .ZN(
        n14889) );
  OAI21_X1 U16774 ( .B1(n14891), .B2(n14890), .A(n14889), .ZN(n14898) );
  XOR2_X1 U16775 ( .A(keyinput_22), .B(DATAI_10_), .Z(n14897) );
  XOR2_X1 U16776 ( .A(DATAI_9_), .B(keyinput_23), .Z(n14895) );
  XOR2_X1 U16777 ( .A(keyinput_26), .B(DATAI_6_), .Z(n14894) );
  XNOR2_X1 U16778 ( .A(keyinput_25), .B(DATAI_7_), .ZN(n14893) );
  XNOR2_X1 U16779 ( .A(keyinput_24), .B(DATAI_8_), .ZN(n14892) );
  NAND4_X1 U16780 ( .A1(n14895), .A2(n14894), .A3(n14893), .A4(n14892), .ZN(
        n14896) );
  AOI21_X1 U16781 ( .B1(n14898), .B2(n14897), .A(n14896), .ZN(n14901) );
  XNOR2_X1 U16782 ( .A(keyinput_28), .B(DATAI_4_), .ZN(n14900) );
  XNOR2_X1 U16783 ( .A(keyinput_27), .B(DATAI_5_), .ZN(n14899) );
  NOR3_X1 U16784 ( .A1(n14901), .A2(n14900), .A3(n14899), .ZN(n14913) );
  XNOR2_X1 U16785 ( .A(keyinput_32), .B(DATAI_0_), .ZN(n14903) );
  XNOR2_X1 U16786 ( .A(DATAI_3_), .B(keyinput_29), .ZN(n14902) );
  NOR2_X1 U16787 ( .A1(n14903), .A2(n14902), .ZN(n14909) );
  INV_X1 U16788 ( .A(keyinput_31), .ZN(n14904) );
  XNOR2_X1 U16789 ( .A(n14904), .B(DATAI_1_), .ZN(n14908) );
  INV_X1 U16790 ( .A(keyinput_30), .ZN(n14905) );
  XNOR2_X1 U16791 ( .A(n14905), .B(DATAI_2_), .ZN(n14907) );
  XNOR2_X1 U16792 ( .A(keyinput_33), .B(HOLD), .ZN(n14906) );
  NAND4_X1 U16793 ( .A1(n14909), .A2(n14908), .A3(n14907), .A4(n14906), .ZN(
        n14912) );
  XOR2_X1 U16794 ( .A(NA), .B(keyinput_34), .Z(n14911) );
  XOR2_X1 U16795 ( .A(BS16), .B(keyinput_35), .Z(n14910) );
  OAI211_X1 U16796 ( .C1(n14913), .C2(n14912), .A(n14911), .B(n14910), .ZN(
        n14917) );
  XNOR2_X1 U16797 ( .A(keyinput_36), .B(READY1), .ZN(n14916) );
  XNOR2_X1 U16798 ( .A(n14914), .B(keyinput_37), .ZN(n14915) );
  AOI21_X1 U16799 ( .B1(n14917), .B2(n14916), .A(n14915), .ZN(n14921) );
  INV_X1 U16800 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n20707) );
  XNOR2_X1 U16801 ( .A(n20707), .B(keyinput_40), .ZN(n14920) );
  XNOR2_X1 U16802 ( .A(P1_ADS_N_REG_SCAN_IN), .B(keyinput_39), .ZN(n14919) );
  XNOR2_X1 U16803 ( .A(keyinput_38), .B(P1_READREQUEST_REG_SCAN_IN), .ZN(
        n14918) );
  NOR4_X1 U16804 ( .A1(n14921), .A2(n14920), .A3(n14919), .A4(n14918), .ZN(
        n14924) );
  XNOR2_X1 U16805 ( .A(keyinput_41), .B(P1_M_IO_N_REG_SCAN_IN), .ZN(n14923) );
  XOR2_X1 U16806 ( .A(keyinput_42), .B(P1_D_C_N_REG_SCAN_IN), .Z(n14922) );
  OAI21_X1 U16807 ( .B1(n14924), .B2(n14923), .A(n14922), .ZN(n14927) );
  XOR2_X1 U16808 ( .A(keyinput_43), .B(P1_REQUESTPENDING_REG_SCAN_IN), .Z(
        n14926) );
  XNOR2_X1 U16809 ( .A(keyinput_44), .B(P1_STATEBS16_REG_SCAN_IN), .ZN(n14925)
         );
  AOI21_X1 U16810 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n14931) );
  XNOR2_X1 U16811 ( .A(n17878), .B(keyinput_45), .ZN(n14930) );
  XOR2_X1 U16812 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_47), .Z(n14929) );
  XNOR2_X1 U16813 ( .A(keyinput_46), .B(P1_FLUSH_REG_SCAN_IN), .ZN(n14928) );
  OAI211_X1 U16814 ( .C1(n14931), .C2(n14930), .A(n14929), .B(n14928), .ZN(
        n14935) );
  XOR2_X1 U16815 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_49), .Z(
        n14934) );
  XOR2_X1 U16816 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_50), .Z(
        n14933) );
  XOR2_X1 U16817 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_48), .Z(
        n14932) );
  NAND4_X1 U16818 ( .A1(n14935), .A2(n14934), .A3(n14933), .A4(n14932), .ZN(
        n14939) );
  XNOR2_X1 U16819 ( .A(keyinput_51), .B(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(
        n14938) );
  XNOR2_X1 U16820 ( .A(keyinput_52), .B(P1_REIP_REG_31__SCAN_IN), .ZN(n14936)
         );
  AOI211_X1 U16821 ( .C1(n14939), .C2(n14938), .A(n14937), .B(n14936), .ZN(
        n14940) );
  AOI211_X1 U16822 ( .C1(n14943), .C2(n14942), .A(n14941), .B(n14940), .ZN(
        n14946) );
  XNOR2_X1 U16823 ( .A(keyinput_57), .B(P1_REIP_REG_26__SCAN_IN), .ZN(n14945)
         );
  XNOR2_X1 U16824 ( .A(keyinput_58), .B(P1_REIP_REG_25__SCAN_IN), .ZN(n14944)
         );
  NOR3_X1 U16825 ( .A1(n14946), .A2(n14945), .A3(n14944), .ZN(n14949) );
  XNOR2_X1 U16826 ( .A(keyinput_59), .B(P1_REIP_REG_24__SCAN_IN), .ZN(n14948)
         );
  XNOR2_X1 U16827 ( .A(keyinput_60), .B(P1_REIP_REG_23__SCAN_IN), .ZN(n14947)
         );
  OAI21_X1 U16828 ( .B1(n14949), .B2(n14948), .A(n14947), .ZN(n14952) );
  XOR2_X1 U16829 ( .A(keyinput_61), .B(P1_REIP_REG_22__SCAN_IN), .Z(n14951) );
  XOR2_X1 U16830 ( .A(keyinput_62), .B(P1_REIP_REG_21__SCAN_IN), .Z(n14950) );
  AOI21_X1 U16831 ( .B1(n14952), .B2(n14951), .A(n14950), .ZN(n14955) );
  XOR2_X1 U16832 ( .A(keyinput_63), .B(P1_REIP_REG_20__SCAN_IN), .Z(n14954) );
  XNOR2_X1 U16833 ( .A(keyinput_64), .B(P1_REIP_REG_19__SCAN_IN), .ZN(n14953)
         );
  NOR3_X1 U16834 ( .A1(n14955), .A2(n14954), .A3(n14953), .ZN(n14958) );
  XOR2_X1 U16835 ( .A(keyinput_66), .B(P1_REIP_REG_17__SCAN_IN), .Z(n14957) );
  XOR2_X1 U16836 ( .A(keyinput_65), .B(P1_REIP_REG_18__SCAN_IN), .Z(n14956) );
  NOR3_X1 U16837 ( .A1(n14958), .A2(n14957), .A3(n14956), .ZN(n14961) );
  XOR2_X1 U16838 ( .A(keyinput_67), .B(P1_REIP_REG_16__SCAN_IN), .Z(n14960) );
  XNOR2_X1 U16839 ( .A(keyinput_68), .B(P1_REIP_REG_15__SCAN_IN), .ZN(n14959)
         );
  NOR3_X1 U16840 ( .A1(n14961), .A2(n14960), .A3(n14959), .ZN(n14964) );
  XNOR2_X1 U16841 ( .A(P1_REIP_REG_14__SCAN_IN), .B(keyinput_69), .ZN(n14963)
         );
  XNOR2_X1 U16842 ( .A(keyinput_70), .B(P1_REIP_REG_13__SCAN_IN), .ZN(n14962)
         );
  NOR3_X1 U16843 ( .A1(n14964), .A2(n14963), .A3(n14962), .ZN(n14968) );
  XOR2_X1 U16844 ( .A(keyinput_73), .B(P1_REIP_REG_10__SCAN_IN), .Z(n14967) );
  XOR2_X1 U16845 ( .A(keyinput_71), .B(P1_REIP_REG_12__SCAN_IN), .Z(n14966) );
  XOR2_X1 U16846 ( .A(keyinput_72), .B(P1_REIP_REG_11__SCAN_IN), .Z(n14965) );
  NOR4_X1 U16847 ( .A1(n14968), .A2(n14967), .A3(n14966), .A4(n14965), .ZN(
        n14971) );
  XOR2_X1 U16848 ( .A(keyinput_75), .B(P1_REIP_REG_8__SCAN_IN), .Z(n14970) );
  XOR2_X1 U16849 ( .A(keyinput_74), .B(P1_REIP_REG_9__SCAN_IN), .Z(n14969) );
  NOR3_X1 U16850 ( .A1(n14971), .A2(n14970), .A3(n14969), .ZN(n14974) );
  XOR2_X1 U16851 ( .A(keyinput_76), .B(P1_REIP_REG_7__SCAN_IN), .Z(n14973) );
  XOR2_X1 U16852 ( .A(keyinput_77), .B(P1_REIP_REG_6__SCAN_IN), .Z(n14972) );
  NOR3_X1 U16853 ( .A1(n14974), .A2(n14973), .A3(n14972), .ZN(n14977) );
  XOR2_X1 U16854 ( .A(keyinput_78), .B(P1_REIP_REG_5__SCAN_IN), .Z(n14976) );
  XOR2_X1 U16855 ( .A(keyinput_79), .B(P1_REIP_REG_4__SCAN_IN), .Z(n14975) );
  NOR3_X1 U16856 ( .A1(n14977), .A2(n14976), .A3(n14975), .ZN(n14981) );
  XOR2_X1 U16857 ( .A(keyinput_81), .B(P1_REIP_REG_2__SCAN_IN), .Z(n14980) );
  XOR2_X1 U16858 ( .A(keyinput_82), .B(P1_REIP_REG_1__SCAN_IN), .Z(n14979) );
  XNOR2_X1 U16859 ( .A(keyinput_80), .B(P1_REIP_REG_3__SCAN_IN), .ZN(n14978)
         );
  NOR4_X1 U16860 ( .A1(n14981), .A2(n14980), .A3(n14979), .A4(n14978), .ZN(
        n14985) );
  XOR2_X1 U16861 ( .A(keyinput_84), .B(P1_EBX_REG_31__SCAN_IN), .Z(n14984) );
  XOR2_X1 U16862 ( .A(keyinput_83), .B(P1_REIP_REG_0__SCAN_IN), .Z(n14983) );
  XOR2_X1 U16863 ( .A(keyinput_85), .B(P1_EBX_REG_30__SCAN_IN), .Z(n14982) );
  NOR4_X1 U16864 ( .A1(n14985), .A2(n14984), .A3(n14983), .A4(n14982), .ZN(
        n14988) );
  XOR2_X1 U16865 ( .A(keyinput_86), .B(P1_EBX_REG_29__SCAN_IN), .Z(n14987) );
  XOR2_X1 U16866 ( .A(keyinput_87), .B(P1_EBX_REG_28__SCAN_IN), .Z(n14986) );
  NOR3_X1 U16867 ( .A1(n14988), .A2(n14987), .A3(n14986), .ZN(n14992) );
  XOR2_X1 U16868 ( .A(keyinput_88), .B(P1_EBX_REG_27__SCAN_IN), .Z(n14991) );
  XOR2_X1 U16869 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_90), .Z(n14990) );
  XNOR2_X1 U16870 ( .A(keyinput_89), .B(P1_EBX_REG_26__SCAN_IN), .ZN(n14989)
         );
  OAI211_X1 U16871 ( .C1(n14992), .C2(n14991), .A(n14990), .B(n14989), .ZN(
        n14995) );
  XNOR2_X1 U16872 ( .A(keyinput_91), .B(P1_EBX_REG_24__SCAN_IN), .ZN(n14994)
         );
  XNOR2_X1 U16873 ( .A(keyinput_92), .B(P1_EBX_REG_23__SCAN_IN), .ZN(n14993)
         );
  AOI21_X1 U16874 ( .B1(n14995), .B2(n14994), .A(n14993), .ZN(n14998) );
  XOR2_X1 U16875 ( .A(keyinput_93), .B(P1_EBX_REG_22__SCAN_IN), .Z(n14997) );
  XOR2_X1 U16876 ( .A(keyinput_94), .B(P1_EBX_REG_21__SCAN_IN), .Z(n14996) );
  NOR3_X1 U16877 ( .A1(n14998), .A2(n14997), .A3(n14996), .ZN(n15005) );
  XOR2_X1 U16878 ( .A(P1_EBX_REG_20__SCAN_IN), .B(keyinput_95), .Z(n15002) );
  XOR2_X1 U16879 ( .A(P1_EBX_REG_18__SCAN_IN), .B(keyinput_97), .Z(n15001) );
  XNOR2_X1 U16880 ( .A(keyinput_98), .B(P1_EBX_REG_17__SCAN_IN), .ZN(n15000)
         );
  XNOR2_X1 U16881 ( .A(keyinput_96), .B(P1_EBX_REG_19__SCAN_IN), .ZN(n14999)
         );
  NAND4_X1 U16882 ( .A1(n15002), .A2(n15001), .A3(n15000), .A4(n14999), .ZN(
        n15004) );
  XNOR2_X1 U16883 ( .A(keyinput_99), .B(P1_EBX_REG_16__SCAN_IN), .ZN(n15003)
         );
  OAI21_X1 U16884 ( .B1(n15005), .B2(n15004), .A(n15003), .ZN(n15008) );
  XOR2_X1 U16885 ( .A(keyinput_100), .B(P1_EBX_REG_15__SCAN_IN), .Z(n15007) );
  XOR2_X1 U16886 ( .A(keyinput_101), .B(P1_EBX_REG_14__SCAN_IN), .Z(n15006) );
  AOI21_X1 U16887 ( .B1(n15008), .B2(n15007), .A(n15006), .ZN(n15011) );
  XOR2_X1 U16888 ( .A(keyinput_102), .B(P1_EBX_REG_13__SCAN_IN), .Z(n15010) );
  XNOR2_X1 U16889 ( .A(keyinput_103), .B(P1_EBX_REG_12__SCAN_IN), .ZN(n15009)
         );
  OAI21_X1 U16890 ( .B1(n15011), .B2(n15010), .A(n15009), .ZN(n15015) );
  XOR2_X1 U16891 ( .A(keyinput_104), .B(P1_EBX_REG_11__SCAN_IN), .Z(n15014) );
  XOR2_X1 U16892 ( .A(keyinput_106), .B(P1_EBX_REG_9__SCAN_IN), .Z(n15013) );
  XNOR2_X1 U16893 ( .A(keyinput_105), .B(P1_EBX_REG_10__SCAN_IN), .ZN(n15012)
         );
  AOI211_X1 U16894 ( .C1(n15015), .C2(n15014), .A(n15013), .B(n15012), .ZN(
        n15019) );
  XOR2_X1 U16895 ( .A(keyinput_107), .B(P1_EBX_REG_8__SCAN_IN), .Z(n15018) );
  XOR2_X1 U16896 ( .A(keyinput_108), .B(P1_EBX_REG_7__SCAN_IN), .Z(n15017) );
  XNOR2_X1 U16897 ( .A(P1_EBX_REG_6__SCAN_IN), .B(keyinput_109), .ZN(n15016)
         );
  NOR4_X1 U16898 ( .A1(n15019), .A2(n15018), .A3(n15017), .A4(n15016), .ZN(
        n15025) );
  AOI22_X1 U16899 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(keyinput_114), .B1(n15459), 
        .B2(keyinput_113), .ZN(n15020) );
  OAI221_X1 U16900 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(keyinput_114), .C1(n15459), .C2(keyinput_113), .A(n15020), .ZN(n15024) );
  AOI22_X1 U16901 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(keyinput_112), .B1(
        P1_EBX_REG_5__SCAN_IN), .B2(keyinput_110), .ZN(n15021) );
  OAI221_X1 U16902 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(keyinput_112), .C1(
        P1_EBX_REG_5__SCAN_IN), .C2(keyinput_110), .A(n15021), .ZN(n15023) );
  XNOR2_X1 U16903 ( .A(P1_EBX_REG_4__SCAN_IN), .B(keyinput_111), .ZN(n15022)
         );
  OR4_X1 U16904 ( .A1(n15025), .A2(n15024), .A3(n15023), .A4(n15022), .ZN(
        n15029) );
  XNOR2_X1 U16905 ( .A(keyinput_117), .B(P1_EAX_REG_30__SCAN_IN), .ZN(n15028)
         );
  XNOR2_X1 U16906 ( .A(keyinput_115), .B(P1_EBX_REG_0__SCAN_IN), .ZN(n15027)
         );
  XNOR2_X1 U16907 ( .A(keyinput_116), .B(P1_EAX_REG_31__SCAN_IN), .ZN(n15026)
         );
  NAND4_X1 U16908 ( .A1(n15029), .A2(n15028), .A3(n15027), .A4(n15026), .ZN(
        n15031) );
  XOR2_X1 U16909 ( .A(keyinput_118), .B(P1_EAX_REG_29__SCAN_IN), .Z(n15030) );
  NAND2_X1 U16910 ( .A1(n15031), .A2(n15030), .ZN(n15037) );
  OAI22_X1 U16911 ( .A1(n13533), .A2(keyinput_119), .B1(keyinput_120), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n15032) );
  AOI221_X1 U16912 ( .B1(n13533), .B2(keyinput_119), .C1(
        P1_EAX_REG_27__SCAN_IN), .C2(keyinput_120), .A(n15032), .ZN(n15036) );
  XOR2_X1 U16913 ( .A(keyinput_122), .B(P1_EAX_REG_25__SCAN_IN), .Z(n15035) );
  OAI22_X1 U16914 ( .A1(n13488), .A2(keyinput_121), .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput_123), .ZN(n15033) );
  AOI221_X1 U16915 ( .B1(n13488), .B2(keyinput_121), .C1(keyinput_123), .C2(
        P1_EAX_REG_24__SCAN_IN), .A(n15033), .ZN(n15034) );
  NAND4_X1 U16916 ( .A1(n15037), .A2(n15036), .A3(n15035), .A4(n15034), .ZN(
        n15041) );
  XOR2_X1 U16917 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_125), .Z(n15040) );
  XOR2_X1 U16918 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_124), .Z(n15039) );
  XNOR2_X1 U16919 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_126), .ZN(n15038)
         );
  NAND4_X1 U16920 ( .A1(n15041), .A2(n15040), .A3(n15039), .A4(n15038), .ZN(
        n15044) );
  XOR2_X1 U16921 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_127), .Z(n15043) );
  XOR2_X1 U16922 ( .A(keyinput_255), .B(P1_EAX_REG_20__SCAN_IN), .Z(n15042) );
  AOI21_X1 U16923 ( .B1(n15044), .B2(n15043), .A(n15042), .ZN(n15045) );
  INV_X1 U16924 ( .A(n15045), .ZN(n15046) );
  NOR4_X1 U16925 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n15051) );
  NOR4_X1 U16926 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n15050) );
  NOR4_X1 U16927 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n15049) );
  NOR4_X1 U16928 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n15048) );
  NAND4_X1 U16929 ( .A1(n15051), .A2(n15050), .A3(n15049), .A4(n15048), .ZN(
        n15056) );
  NOR4_X1 U16930 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n15054) );
  NOR4_X1 U16931 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n15053) );
  NOR4_X1 U16932 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n15052) );
  INV_X1 U16933 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20441) );
  NAND4_X1 U16934 ( .A1(n15054), .A2(n15053), .A3(n15052), .A4(n20441), .ZN(
        n15055) );
  AOI22_X1 U16935 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n20264), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n20263), .ZN(n20411) );
  INV_X1 U16936 ( .A(n15061), .ZN(n15063) );
  NAND2_X1 U16937 ( .A1(n15063), .A2(n14367), .ZN(n15064) );
  NAND2_X1 U16938 ( .A1(n11354), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n15067) );
  NAND4_X1 U16939 ( .A1(n14353), .A2(n15067), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n14346), .ZN(n15068) );
  NAND2_X1 U16940 ( .A1(n15070), .A2(n14346), .ZN(n19941) );
  NAND3_X1 U16941 ( .A1(n12216), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19861) );
  NOR2_X1 U16942 ( .A1(n19861), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20271) );
  INV_X1 U16943 ( .A(n20271), .ZN(n15081) );
  NAND2_X1 U16944 ( .A1(n19932), .A2(n19846), .ZN(n19985) );
  OAI211_X1 U16945 ( .C1(n15078), .C2(n19941), .A(n15081), .B(n19985), .ZN(
        n15077) );
  OAI21_X1 U16946 ( .B1(n20172), .B2(n20339), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n15075) );
  INV_X1 U16947 ( .A(n15071), .ZN(n15073) );
  AND2_X1 U16948 ( .A1(n15073), .A2(n15072), .ZN(n19969) );
  NAND2_X1 U16949 ( .A1(n19969), .A2(n19967), .ZN(n15074) );
  AOI21_X1 U16950 ( .B1(n15075), .B2(n15074), .A(n20259), .ZN(n15076) );
  NAND2_X1 U16951 ( .A1(n15077), .A2(n15076), .ZN(n20273) );
  AOI21_X1 U16952 ( .B1(n15078), .B2(n15081), .A(n19916), .ZN(n15079) );
  AOI21_X1 U16953 ( .B1(n19969), .B2(n15080), .A(n15079), .ZN(n19869) );
  MUX2_X1 U16954 ( .A(BUF1_REG_0__SCAN_IN), .B(BUF2_REG_0__SCAN_IN), .S(n15306), .Z(n20314) );
  INV_X1 U16955 ( .A(n20434), .ZN(n15082) );
  INV_X1 U16956 ( .A(n20261), .ZN(n16030) );
  NAND2_X1 U16957 ( .A1(n11156), .A2(n16030), .ZN(n20403) );
  OAI22_X1 U16958 ( .A1(n19869), .A2(n15082), .B1(n20403), .B2(n15081), .ZN(
        n15084) );
  AOI22_X1 U16959 ( .A1(n20264), .A2(BUF2_REG_16__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n20426) );
  NOR2_X1 U16960 ( .A1(n20426), .A2(n20215), .ZN(n15083) );
  AOI211_X1 U16961 ( .C1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .C2(n20273), .A(
        n15084), .B(n15083), .ZN(n15085) );
  OAI21_X1 U16962 ( .B1(n20411), .B2(n20349), .A(n15085), .ZN(n15086) );
  XNOR2_X1 U16963 ( .A(n15087), .B(n15086), .ZN(P2_U3144) );
  NOR4_X1 U16964 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20779), .A4(n22779), .ZN(n15089) );
  NOR4_X1 U16965 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n15088) );
  NAND3_X1 U16966 ( .A1(n16731), .A2(n15089), .A3(n15088), .ZN(U214) );
  NOR2_X1 U16967 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n15091) );
  NOR4_X1 U16968 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n15090) );
  NAND4_X1 U16969 ( .A1(n15091), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n15090), .ZN(n15092) );
  OR2_X1 U16970 ( .A1(n16354), .A2(n15092), .ZN(n20711) );
  INV_X2 U16971 ( .A(U214), .ZN(n20764) );
  NAND2_X1 U16972 ( .A1(n19194), .A2(n11173), .ZN(n19029) );
  AOI211_X1 U16973 ( .C1(n17509), .C2(n15093), .A(n19125), .B(n19029), .ZN(
        n15105) );
  INV_X1 U16974 ( .A(n19092), .ZN(n19160) );
  AOI22_X1 U16975 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n19207), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19163), .ZN(n15094) );
  OAI211_X1 U16976 ( .C1(n15095), .C2(n19160), .A(n15094), .B(n19325), .ZN(
        n15104) );
  INV_X1 U16977 ( .A(n15096), .ZN(n15097) );
  OAI22_X1 U16978 ( .A1(n15097), .A2(n19147), .B1(n17511), .B2(n19182), .ZN(
        n15103) );
  AOI21_X1 U16979 ( .B1(n15098), .B2(n17278), .A(n17264), .ZN(n17668) );
  INV_X1 U16980 ( .A(n17668), .ZN(n15101) );
  XNOR2_X1 U16981 ( .A(n15100), .B(n15099), .ZN(n17666) );
  OAI22_X1 U16982 ( .A1(n15101), .A2(n19165), .B1(n17666), .B2(n19222), .ZN(
        n15102) );
  INV_X1 U16983 ( .A(n16065), .ZN(n19040) );
  INV_X1 U16984 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n18045) );
  NOR2_X1 U16985 ( .A1(n18021), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15108) );
  INV_X1 U16986 ( .A(n15108), .ZN(n15106) );
  OAI211_X1 U16987 ( .C1(n19040), .C2(n18045), .A(n15106), .B(n15111), .ZN(
        P2_U2814) );
  INV_X1 U16988 ( .A(n15107), .ZN(n19013) );
  OAI21_X1 U16989 ( .B1(n15108), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19013), 
        .ZN(n15109) );
  OAI21_X1 U16990 ( .B1(n19009), .B2(n19013), .A(n15109), .ZN(P2_U3612) );
  MUX2_X1 U16991 ( .A(n12028), .B(n19023), .S(n17281), .Z(n15110) );
  OAI21_X1 U16992 ( .B1(n18018), .B2(n17272), .A(n15110), .ZN(P2_U2887) );
  NOR2_X1 U16993 ( .A1(n15111), .A2(n22317), .ZN(n15112) );
  AOI22_X1 U16994 ( .A1(n15262), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n15303), .ZN(n15114) );
  INV_X1 U16995 ( .A(n15112), .ZN(n15113) );
  AOI22_X1 U16996 ( .A1(n16353), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16354), .ZN(n20205) );
  INV_X1 U16997 ( .A(n20205), .ZN(n17380) );
  NAND2_X1 U16998 ( .A1(n11291), .A2(n17380), .ZN(n15277) );
  NAND2_X1 U16999 ( .A1(n15114), .A2(n15277), .ZN(P2_U2969) );
  AOI22_X1 U17000 ( .A1(n15262), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n15303), .ZN(n15115) );
  INV_X1 U17001 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20721) );
  INV_X1 U17002 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n21325) );
  OAI22_X1 U17003 ( .A1(n16354), .A2(n20721), .B1(n21325), .B2(n16353), .ZN(
        n20109) );
  NAND2_X1 U17004 ( .A1(n11291), .A2(n20109), .ZN(n15268) );
  NAND2_X1 U17005 ( .A1(n15115), .A2(n15268), .ZN(P2_U2971) );
  AOI22_X1 U17006 ( .A1(n15262), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n15303), .ZN(n15116) );
  AOI22_X1 U17007 ( .A1(n16353), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16354), .ZN(n20022) );
  INV_X1 U17008 ( .A(n20022), .ZN(n17348) );
  NAND2_X1 U17009 ( .A1(n11291), .A2(n17348), .ZN(n15286) );
  NAND2_X1 U17010 ( .A1(n15116), .A2(n15286), .ZN(P2_U2973) );
  AOI22_X1 U17011 ( .A1(n15262), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n15303), .ZN(n15118) );
  AOI22_X1 U17012 ( .A1(n16353), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15306), .ZN(n19833) );
  INV_X1 U17013 ( .A(n19833), .ZN(n15117) );
  NAND2_X1 U17014 ( .A1(n11291), .A2(n15117), .ZN(n15266) );
  NAND2_X1 U17015 ( .A1(n15118), .A2(n15266), .ZN(P2_U2974) );
  AOI22_X1 U17016 ( .A1(n15262), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n15303), .ZN(n15119) );
  AOI22_X1 U17017 ( .A1(n16353), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15306), .ZN(n20069) );
  INV_X1 U17018 ( .A(n20069), .ZN(n17351) );
  NAND2_X1 U17019 ( .A1(n11291), .A2(n17351), .ZN(n15270) );
  NAND2_X1 U17020 ( .A1(n15119), .A2(n15270), .ZN(P2_U2972) );
  AOI22_X1 U17021 ( .A1(n15262), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n15296), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n15120) );
  AOI22_X1 U17022 ( .A1(n16353), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16354), .ZN(n20163) );
  INV_X1 U17023 ( .A(n20163), .ZN(n17371) );
  NAND2_X1 U17024 ( .A1(n11291), .A2(n17371), .ZN(n15279) );
  NAND2_X1 U17025 ( .A1(n15120), .A2(n15279), .ZN(P2_U2970) );
  INV_X1 U17026 ( .A(n15370), .ZN(n15122) );
  NAND2_X1 U17027 ( .A1(n15121), .A2(n12888), .ZN(n17862) );
  INV_X1 U17028 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20527) );
  OR2_X1 U17029 ( .A1(n21956), .A2(n22248), .ZN(n15123) );
  NOR2_X1 U17030 ( .A1(n16731), .A2(n14682), .ZN(n15124) );
  AOI21_X1 U17031 ( .B1(n16731), .B2(BUF1_REG_15__SCAN_IN), .A(n15124), .ZN(
        n16783) );
  INV_X1 U17032 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n15125) );
  OAI222_X1 U17033 ( .A1(n22379), .A2(n20527), .B1(n22373), .B2(n16783), .C1(
        n15261), .C2(n15125), .ZN(P1_U2967) );
  INV_X1 U17034 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n17378) );
  NOR2_X1 U17035 ( .A1(n15126), .A2(n15634), .ZN(n15657) );
  NAND2_X1 U17036 ( .A1(n15657), .A2(n19341), .ZN(n15128) );
  NAND2_X1 U17037 ( .A1(n15303), .A2(n22312), .ZN(n15127) );
  INV_X1 U17038 ( .A(n15129), .ZN(n15130) );
  INV_X1 U17039 ( .A(n15131), .ZN(n18016) );
  NOR2_X1 U17040 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18016), .ZN(n15414) );
  CLKBUF_X2 U17041 ( .A(n15414), .Z(n19016) );
  NOR2_X4 U17042 ( .A1(n19016), .A2(n18048), .ZN(n18068) );
  AOI22_X1 U17043 ( .A1(n15414), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n15132) );
  OAI21_X1 U17044 ( .B1(n17378), .B2(n15420), .A(n15132), .ZN(P2_U2933) );
  INV_X1 U17045 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n17384) );
  AOI22_X1 U17046 ( .A1(n19016), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n15133) );
  OAI21_X1 U17047 ( .B1(n17384), .B2(n15420), .A(n15133), .ZN(P2_U2934) );
  INV_X1 U17048 ( .A(n20706), .ZN(n15868) );
  NOR2_X1 U17049 ( .A1(n15136), .A2(n15868), .ZN(n22780) );
  INV_X1 U17050 ( .A(n22780), .ZN(n15137) );
  NAND2_X1 U17051 ( .A1(n15134), .A2(n15813), .ZN(n16370) );
  INV_X1 U17052 ( .A(n16369), .ZN(n15135) );
  OAI33_X1 U17053 ( .A1(n15137), .A2(n22782), .A3(P1_READREQUEST_REG_SCAN_IN), 
        .B1(n16376), .B2(n15798), .B3(n16400), .ZN(n15138) );
  INV_X1 U17054 ( .A(n15138), .ZN(P1_U3487) );
  AOI21_X1 U17055 ( .B1(n15206), .B2(n15140), .A(n15139), .ZN(n15210) );
  INV_X1 U17056 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15141) );
  AOI22_X1 U17057 ( .A1(n15210), .A2(n17983), .B1(n18002), .B2(n15141), .ZN(
        n15146) );
  XNOR2_X1 U17058 ( .A(n15142), .B(n15206), .ZN(n15209) );
  NAND2_X1 U17059 ( .A1(n18010), .A2(n15209), .ZN(n15143) );
  NAND2_X1 U17060 ( .A1(n19282), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15205) );
  OAI211_X1 U17061 ( .C1(n17987), .C2(n15141), .A(n15143), .B(n15205), .ZN(
        n15144) );
  INV_X1 U17062 ( .A(n15144), .ZN(n15145) );
  OAI211_X1 U17063 ( .C1(n17188), .C2(n15057), .A(n15146), .B(n15145), .ZN(
        P2_U3013) );
  OR2_X1 U17064 ( .A1(n15148), .A2(n15147), .ZN(n15150) );
  AND2_X1 U17065 ( .A1(n15150), .A2(n15149), .ZN(n19020) );
  XNOR2_X1 U17066 ( .A(n19027), .B(n19020), .ZN(n15166) );
  INV_X1 U17067 ( .A(n15650), .ZN(n15151) );
  NAND2_X1 U17068 ( .A1(n15151), .A2(n15641), .ZN(n15155) );
  INV_X1 U17069 ( .A(n15699), .ZN(n15152) );
  NAND4_X1 U17070 ( .A1(n15153), .A2(n15152), .A3(n15635), .A4(n19342), .ZN(
        n15154) );
  NAND2_X1 U17071 ( .A1(n15155), .A2(n15154), .ZN(n15661) );
  AND2_X1 U17072 ( .A1(n15157), .A2(n15156), .ZN(n15158) );
  NAND2_X1 U17073 ( .A1(n20153), .A2(n15160), .ZN(n20253) );
  AOI22_X1 U17074 ( .A1(n20319), .A2(n19020), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n20313), .ZN(n15165) );
  INV_X1 U17075 ( .A(n15161), .ZN(n15162) );
  NOR2_X2 U17076 ( .A1(n20313), .A2(n15162), .ZN(n20315) );
  NAND2_X1 U17077 ( .A1(n11997), .A2(n12006), .ZN(n15163) );
  OR2_X1 U17078 ( .A1(n20315), .A2(n16355), .ZN(n16084) );
  NAND2_X1 U17079 ( .A1(n16084), .A2(n20314), .ZN(n15164) );
  OAI211_X1 U17080 ( .C1(n15166), .C2(n20253), .A(n15165), .B(n15164), .ZN(
        P2_U2919) );
  INV_X1 U17081 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15172) );
  NOR2_X1 U17082 ( .A1(n16370), .A2(n12888), .ZN(n17058) );
  INV_X1 U17083 ( .A(n17862), .ZN(n15167) );
  OR2_X1 U17084 ( .A1(n17058), .A2(n15167), .ZN(n15170) );
  NAND2_X1 U17085 ( .A1(n15168), .A2(n22302), .ZN(n22297) );
  INV_X1 U17086 ( .A(n22297), .ZN(n16375) );
  AND2_X1 U17087 ( .A1(n15370), .A2(n16375), .ZN(n15169) );
  NAND2_X1 U17088 ( .A1(n20504), .A2(n12895), .ZN(n15485) );
  NAND2_X1 U17089 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n22255) );
  NOR2_X1 U17090 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22255), .ZN(n20521) );
  NOR2_X4 U17091 ( .A1(n20504), .A2(n21955), .ZN(n20514) );
  AOI22_X1 U17092 ( .A1(n21955), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n15171) );
  OAI21_X1 U17093 ( .B1(n15172), .B2(n15485), .A(n15171), .ZN(P1_U2914) );
  AOI22_X1 U17094 ( .A1(n21955), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n15173) );
  OAI21_X1 U17095 ( .B1(n13442), .B2(n15485), .A(n15173), .ZN(P1_U2912) );
  AOI22_X1 U17096 ( .A1(n21955), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n15174) );
  OAI21_X1 U17097 ( .B1(n15175), .B2(n15485), .A(n15174), .ZN(P1_U2915) );
  AOI22_X1 U17098 ( .A1(n21955), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n15176) );
  OAI21_X1 U17099 ( .B1(n15250), .B2(n15485), .A(n15176), .ZN(P1_U2913) );
  AOI22_X1 U17100 ( .A1(n21955), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n15177) );
  OAI21_X1 U17101 ( .B1(n13465), .B2(n15485), .A(n15177), .ZN(P1_U2911) );
  INV_X1 U17102 ( .A(n15178), .ZN(n15181) );
  OAI21_X1 U17103 ( .B1(n15181), .B2(n15180), .A(n15179), .ZN(n20634) );
  NAND2_X1 U17104 ( .A1(n12900), .A2(n12842), .ZN(n15182) );
  NAND2_X2 U17105 ( .A1(n16789), .A2(n15182), .ZN(n16782) );
  INV_X1 U17106 ( .A(n15182), .ZN(n15183) );
  MUX2_X1 U17107 ( .A(DATAI_0_), .B(BUF1_REG_0__SCAN_IN), .S(n16731), .Z(
        n16777) );
  INV_X1 U17108 ( .A(n16777), .ZN(n15184) );
  INV_X1 U17109 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20506) );
  OAI222_X1 U17110 ( .A1(n20634), .A2(n16782), .B1(n16791), .B2(n15184), .C1(
        n16789), .C2(n20506), .ZN(P1_U2904) );
  NAND2_X1 U17111 ( .A1(n15254), .A2(n16777), .ZN(n15187) );
  AOI22_X1 U17112 ( .A1(n22377), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n15257), 
        .B2(P1_EAX_REG_0__SCAN_IN), .ZN(n15185) );
  NAND2_X1 U17113 ( .A1(n15187), .A2(n15185), .ZN(P1_U2952) );
  AOI22_X1 U17114 ( .A1(n22377), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n15257), 
        .B2(P1_EAX_REG_16__SCAN_IN), .ZN(n15186) );
  NAND2_X1 U17115 ( .A1(n15187), .A2(n15186), .ZN(P1_U2937) );
  OR2_X1 U17116 ( .A1(n15189), .A2(n15188), .ZN(n15190) );
  NAND2_X1 U17117 ( .A1(n15191), .A2(n15190), .ZN(n19303) );
  NAND2_X1 U17118 ( .A1(n20253), .A2(n20154), .ZN(n20064) );
  INV_X1 U17119 ( .A(n20064), .ZN(n15793) );
  INV_X1 U17120 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n18062) );
  OAI222_X1 U17121 ( .A1(n19303), .A2(n15793), .B1(n20022), .B2(n20257), .C1(
        n18062), .C2(n20153), .ZN(P2_U2913) );
  INV_X1 U17122 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20715) );
  NOR2_X1 U17123 ( .A1(n16731), .A2(DATAI_1_), .ZN(n15192) );
  AOI21_X1 U17124 ( .B1(n16731), .B2(n20715), .A(n15192), .ZN(n16771) );
  NAND2_X1 U17125 ( .A1(n15254), .A2(n16771), .ZN(n15237) );
  AOI22_X1 U17126 ( .A1(n22377), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n15257), 
        .B2(P1_EAX_REG_1__SCAN_IN), .ZN(n15193) );
  NAND2_X1 U17127 ( .A1(n15237), .A2(n15193), .ZN(P1_U2953) );
  MUX2_X1 U17128 ( .A(DATAI_2_), .B(BUF1_REG_2__SCAN_IN), .S(n16731), .Z(
        n16768) );
  NAND2_X1 U17129 ( .A1(n15254), .A2(n16768), .ZN(n15252) );
  AOI22_X1 U17130 ( .A1(n22377), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n15257), 
        .B2(P1_EAX_REG_2__SCAN_IN), .ZN(n15194) );
  NAND2_X1 U17131 ( .A1(n15252), .A2(n15194), .ZN(P1_U2954) );
  MUX2_X1 U17132 ( .A(DATAI_6_), .B(BUF1_REG_6__SCAN_IN), .S(n16731), .Z(
        n16753) );
  NAND2_X1 U17133 ( .A1(n15254), .A2(n16753), .ZN(n15243) );
  AOI22_X1 U17134 ( .A1(n22377), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n15257), 
        .B2(P1_EAX_REG_6__SCAN_IN), .ZN(n15195) );
  NAND2_X1 U17135 ( .A1(n15243), .A2(n15195), .ZN(P1_U2958) );
  INV_X1 U17136 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20727) );
  NOR2_X1 U17137 ( .A1(n16731), .A2(DATAI_7_), .ZN(n15196) );
  AOI21_X1 U17138 ( .B1(n16731), .B2(n20727), .A(n15196), .ZN(n16750) );
  NAND2_X1 U17139 ( .A1(n15254), .A2(n16750), .ZN(n15249) );
  AOI22_X1 U17140 ( .A1(n22377), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n15257), 
        .B2(P1_EAX_REG_7__SCAN_IN), .ZN(n15197) );
  NAND2_X1 U17141 ( .A1(n15249), .A2(n15197), .ZN(P1_U2959) );
  INV_X1 U17142 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20719) );
  NOR2_X1 U17143 ( .A1(n16731), .A2(DATAI_3_), .ZN(n15198) );
  AOI21_X1 U17144 ( .B1(n16731), .B2(n20719), .A(n15198), .ZN(n16764) );
  NAND2_X1 U17145 ( .A1(n15254), .A2(n16764), .ZN(n15240) );
  AOI22_X1 U17146 ( .A1(n22377), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n15257), 
        .B2(P1_EAX_REG_3__SCAN_IN), .ZN(n15199) );
  NAND2_X1 U17147 ( .A1(n15240), .A2(n15199), .ZN(P1_U2955) );
  MUX2_X1 U17148 ( .A(DATAI_5_), .B(BUF1_REG_5__SCAN_IN), .S(n16731), .Z(
        n16756) );
  NAND2_X1 U17149 ( .A1(n15254), .A2(n16756), .ZN(n15246) );
  AOI22_X1 U17150 ( .A1(n22377), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n15257), 
        .B2(P1_EAX_REG_5__SCAN_IN), .ZN(n15200) );
  NAND2_X1 U17151 ( .A1(n15246), .A2(n15200), .ZN(P1_U2957) );
  NAND2_X1 U17152 ( .A1(n15202), .A2(n15201), .ZN(n15203) );
  NAND2_X1 U17153 ( .A1(n15204), .A2(n15203), .ZN(n20249) );
  OAI21_X1 U17154 ( .B1(n19225), .B2(n15206), .A(n15205), .ZN(n15208) );
  AOI211_X1 U17155 ( .C1(n19224), .C2(n15206), .A(n16157), .B(n19237), .ZN(
        n15207) );
  AOI211_X1 U17156 ( .C1(n19281), .C2(n20249), .A(n15208), .B(n15207), .ZN(
        n15212) );
  AOI22_X1 U17157 ( .A1(n19335), .A2(n15210), .B1(n19271), .B2(n15209), .ZN(
        n15211) );
  OAI211_X1 U17158 ( .C1(n17188), .C2(n19285), .A(n15212), .B(n15211), .ZN(
        P2_U3045) );
  OAI21_X1 U17159 ( .B1(n15215), .B2(n15214), .A(n15213), .ZN(n20199) );
  INV_X1 U17160 ( .A(n20199), .ZN(n16074) );
  NAND2_X1 U17161 ( .A1(n15217), .A2(n15216), .ZN(n15218) );
  NAND2_X1 U17162 ( .A1(n15219), .A2(n15218), .ZN(n17908) );
  XNOR2_X1 U17163 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n16157), .ZN(
        n15220) );
  INV_X1 U17164 ( .A(n15220), .ZN(n15221) );
  OAI22_X1 U17165 ( .A1(n15221), .A2(n17759), .B1(n17756), .B2(n15220), .ZN(
        n15224) );
  NAND2_X1 U17166 ( .A1(n19282), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n17910) );
  OAI21_X1 U17167 ( .B1(n19225), .B2(n15222), .A(n17910), .ZN(n15223) );
  NOR2_X1 U17168 ( .A1(n15224), .A2(n15223), .ZN(n15230) );
  OAI21_X1 U17169 ( .B1(n15227), .B2(n15226), .A(n15225), .ZN(n15228) );
  INV_X1 U17170 ( .A(n15228), .ZN(n17904) );
  NAND2_X1 U17171 ( .A1(n19271), .A2(n17904), .ZN(n15229) );
  OAI211_X1 U17172 ( .C1(n17908), .C2(n19304), .A(n15230), .B(n15229), .ZN(
        n15231) );
  AOI21_X1 U17173 ( .B1(n17905), .B2(n19329), .A(n15231), .ZN(n15232) );
  OAI21_X1 U17174 ( .B1(n16074), .B2(n19327), .A(n15232), .ZN(P2_U3044) );
  OR2_X1 U17175 ( .A1(n15234), .A2(n15233), .ZN(n15235) );
  NAND2_X1 U17176 ( .A1(n15235), .A2(n16101), .ZN(n19065) );
  INV_X1 U17177 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n18066) );
  AOI22_X1 U17178 ( .A1(n16353), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16354), .ZN(n15274) );
  OAI222_X1 U17179 ( .A1(n19065), .A2(n15793), .B1(n20153), .B2(n18066), .C1(
        n20257), .C2(n15274), .ZN(P2_U2911) );
  INV_X1 U17180 ( .A(P1_UWORD_REG_1__SCAN_IN), .ZN(n15238) );
  NAND2_X1 U17181 ( .A1(n15257), .A2(P1_EAX_REG_17__SCAN_IN), .ZN(n15236) );
  OAI211_X1 U17182 ( .C1(n15261), .C2(n15238), .A(n15237), .B(n15236), .ZN(
        P1_U2938) );
  NAND2_X1 U17183 ( .A1(n22377), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n15239) );
  OAI211_X1 U17184 ( .C1(n22379), .C2(n15241), .A(n15240), .B(n15239), .ZN(
        P1_U2940) );
  INV_X1 U17185 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n15244) );
  NAND2_X1 U17186 ( .A1(n15257), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n15242) );
  OAI211_X1 U17187 ( .C1(n15261), .C2(n15244), .A(n15243), .B(n15242), .ZN(
        P1_U2943) );
  INV_X1 U17188 ( .A(P1_UWORD_REG_5__SCAN_IN), .ZN(n15247) );
  NAND2_X1 U17189 ( .A1(n15257), .A2(P1_EAX_REG_21__SCAN_IN), .ZN(n15245) );
  OAI211_X1 U17190 ( .C1(n15261), .C2(n15247), .A(n15246), .B(n15245), .ZN(
        P1_U2942) );
  NAND2_X1 U17191 ( .A1(n22377), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n15248) );
  OAI211_X1 U17192 ( .C1(n22379), .C2(n15250), .A(n15249), .B(n15248), .ZN(
        P1_U2944) );
  INV_X1 U17193 ( .A(P1_UWORD_REG_2__SCAN_IN), .ZN(n15253) );
  NAND2_X1 U17194 ( .A1(n15257), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n15251) );
  OAI211_X1 U17195 ( .C1(n15261), .C2(n15253), .A(n15252), .B(n15251), .ZN(
        P1_U2939) );
  INV_X1 U17196 ( .A(P1_LWORD_REG_4__SCAN_IN), .ZN(n15256) );
  MUX2_X1 U17197 ( .A(DATAI_4_), .B(BUF1_REG_4__SCAN_IN), .S(n16731), .Z(
        n16760) );
  NAND2_X1 U17198 ( .A1(n15254), .A2(n16760), .ZN(n15259) );
  NAND2_X1 U17199 ( .A1(n15257), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n15255) );
  OAI211_X1 U17200 ( .C1(n15261), .C2(n15256), .A(n15259), .B(n15255), .ZN(
        P1_U2956) );
  INV_X1 U17201 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n15260) );
  NAND2_X1 U17202 ( .A1(n15257), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n15258) );
  OAI211_X1 U17203 ( .C1(n15261), .C2(n15260), .A(n15259), .B(n15258), .ZN(
        P1_U2941) );
  AOI22_X1 U17204 ( .A1(n15313), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n15303), .ZN(n15265) );
  INV_X1 U17205 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20737) );
  OR2_X1 U17206 ( .A1(n15306), .A2(n20737), .ZN(n15264) );
  NAND2_X1 U17207 ( .A1(n15306), .A2(BUF2_REG_12__SCAN_IN), .ZN(n15263) );
  NAND2_X1 U17208 ( .A1(n15264), .A2(n15263), .ZN(n17293) );
  NAND2_X1 U17209 ( .A1(n11291), .A2(n17293), .ZN(n15297) );
  NAND2_X1 U17210 ( .A1(n15265), .A2(n15297), .ZN(P2_U2964) );
  AOI22_X1 U17211 ( .A1(n15313), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n15303), .ZN(n15267) );
  NAND2_X1 U17212 ( .A1(n15267), .A2(n15266), .ZN(P2_U2959) );
  AOI22_X1 U17213 ( .A1(n15313), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n15296), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n15269) );
  NAND2_X1 U17214 ( .A1(n15269), .A2(n15268), .ZN(P2_U2956) );
  AOI22_X1 U17215 ( .A1(n15313), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n15303), .ZN(n15271) );
  NAND2_X1 U17216 ( .A1(n15271), .A2(n15270), .ZN(P2_U2957) );
  AOI22_X1 U17217 ( .A1(n15313), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n15303), .ZN(n15272) );
  AOI22_X1 U17218 ( .A1(n16353), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n15306), .ZN(n15792) );
  INV_X1 U17219 ( .A(n15792), .ZN(n16356) );
  NAND2_X1 U17220 ( .A1(n11291), .A2(n16356), .ZN(n15294) );
  NAND2_X1 U17221 ( .A1(n15272), .A2(n15294), .ZN(P2_U2966) );
  AOI22_X1 U17222 ( .A1(n15313), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n15296), 
        .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n15273) );
  AOI22_X1 U17223 ( .A1(n16353), .A2(BUF1_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n15306), .ZN(n15427) );
  INV_X1 U17224 ( .A(n15427), .ZN(n17314) );
  NAND2_X1 U17225 ( .A1(n11291), .A2(n17314), .ZN(n15301) );
  NAND2_X1 U17226 ( .A1(n15273), .A2(n15301), .ZN(P2_U2962) );
  AOI22_X1 U17227 ( .A1(n15313), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n15303), .ZN(n15275) );
  INV_X1 U17228 ( .A(n15274), .ZN(n17327) );
  NAND2_X1 U17229 ( .A1(n11291), .A2(n17327), .ZN(n15288) );
  NAND2_X1 U17230 ( .A1(n15275), .A2(n15288), .ZN(P2_U2960) );
  AOI22_X1 U17231 ( .A1(n15313), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n15296), .ZN(n15276) );
  AOI22_X1 U17232 ( .A1(n16353), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16354), .ZN(n20258) );
  INV_X1 U17233 ( .A(n20258), .ZN(n17390) );
  NAND2_X1 U17234 ( .A1(n11291), .A2(n17390), .ZN(n15290) );
  NAND2_X1 U17235 ( .A1(n15276), .A2(n15290), .ZN(P2_U2953) );
  AOI22_X1 U17236 ( .A1(n15313), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n15296), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n15278) );
  NAND2_X1 U17237 ( .A1(n15278), .A2(n15277), .ZN(P2_U2954) );
  AOI22_X1 U17238 ( .A1(n15313), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n15296), .ZN(n15280) );
  NAND2_X1 U17239 ( .A1(n15280), .A2(n15279), .ZN(P2_U2955) );
  AOI22_X1 U17240 ( .A1(n15313), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n15296), .ZN(n15283) );
  INV_X1 U17241 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20739) );
  OR2_X1 U17242 ( .A1(n16354), .A2(n20739), .ZN(n15282) );
  NAND2_X1 U17243 ( .A1(n15306), .A2(BUF2_REG_13__SCAN_IN), .ZN(n15281) );
  AND2_X1 U17244 ( .A1(n15282), .A2(n15281), .ZN(n19825) );
  INV_X1 U17245 ( .A(n19825), .ZN(n17282) );
  NAND2_X1 U17246 ( .A1(n11291), .A2(n17282), .ZN(n15299) );
  NAND2_X1 U17247 ( .A1(n15283), .A2(n15299), .ZN(P2_U2980) );
  AOI22_X1 U17248 ( .A1(n15313), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n15303), .ZN(n15285) );
  AOI22_X1 U17249 ( .A1(n16353), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n15306), .ZN(n19828) );
  INV_X1 U17250 ( .A(n19828), .ZN(n15284) );
  NAND2_X1 U17251 ( .A1(n11291), .A2(n15284), .ZN(n15292) );
  NAND2_X1 U17252 ( .A1(n15285), .A2(n15292), .ZN(P2_U2976) );
  AOI22_X1 U17253 ( .A1(n15313), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n15303), .ZN(n15287) );
  NAND2_X1 U17254 ( .A1(n15287), .A2(n15286), .ZN(P2_U2958) );
  AOI22_X1 U17255 ( .A1(n15313), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n15303), .ZN(n15289) );
  NAND2_X1 U17256 ( .A1(n15289), .A2(n15288), .ZN(P2_U2975) );
  AOI22_X1 U17257 ( .A1(n15313), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n15303), .ZN(n15291) );
  NAND2_X1 U17258 ( .A1(n15291), .A2(n15290), .ZN(P2_U2968) );
  AOI22_X1 U17259 ( .A1(n15313), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n15303), .ZN(n15293) );
  NAND2_X1 U17260 ( .A1(n15293), .A2(n15292), .ZN(P2_U2961) );
  AOI22_X1 U17261 ( .A1(n15313), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n15296), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n15295) );
  NAND2_X1 U17262 ( .A1(n15295), .A2(n15294), .ZN(P2_U2981) );
  AOI22_X1 U17263 ( .A1(n15313), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n15296), .ZN(n15298) );
  NAND2_X1 U17264 ( .A1(n15298), .A2(n15297), .ZN(P2_U2979) );
  AOI22_X1 U17265 ( .A1(n15313), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n15303), .ZN(n15300) );
  NAND2_X1 U17266 ( .A1(n15300), .A2(n15299), .ZN(P2_U2965) );
  AOI22_X1 U17267 ( .A1(n15313), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_10__SCAN_IN), .B2(n15303), .ZN(n15302) );
  NAND2_X1 U17268 ( .A1(n15302), .A2(n15301), .ZN(P2_U2977) );
  AOI22_X1 U17269 ( .A1(n16353), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16354), .ZN(n19822) );
  INV_X1 U17270 ( .A(n19822), .ZN(n15304) );
  AOI222_X1 U17271 ( .A1(n15313), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n11291), 
        .B2(n15304), .C1(P2_EAX_REG_15__SCAN_IN), .C2(n15303), .ZN(n15305) );
  INV_X1 U17272 ( .A(n15305), .ZN(P2_U2982) );
  INV_X1 U17273 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n18072) );
  NAND2_X1 U17274 ( .A1(n15313), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n15309) );
  INV_X1 U17275 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20735) );
  OR2_X1 U17276 ( .A1(n15306), .A2(n20735), .ZN(n15308) );
  NAND2_X1 U17277 ( .A1(n15306), .A2(BUF2_REG_11__SCAN_IN), .ZN(n15307) );
  NAND2_X1 U17278 ( .A1(n15308), .A2(n15307), .ZN(n17300) );
  NAND2_X1 U17279 ( .A1(n11291), .A2(n17300), .ZN(n15310) );
  OAI211_X1 U17280 ( .C1(n18072), .C2(n15316), .A(n15309), .B(n15310), .ZN(
        P2_U2978) );
  INV_X1 U17281 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15410) );
  NAND2_X1 U17282 ( .A1(n15313), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n15311) );
  OAI211_X1 U17283 ( .C1(n15410), .C2(n15316), .A(n15311), .B(n15310), .ZN(
        P2_U2963) );
  NAND2_X1 U17284 ( .A1(n15313), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n15312) );
  NAND2_X1 U17285 ( .A1(n11291), .A2(n20314), .ZN(n15314) );
  OAI211_X1 U17286 ( .C1(n15401), .C2(n15316), .A(n15312), .B(n15314), .ZN(
        P2_U2952) );
  INV_X1 U17287 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n18050) );
  NAND2_X1 U17288 ( .A1(n15313), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n15315) );
  OAI211_X1 U17289 ( .C1(n18050), .C2(n15316), .A(n15315), .B(n15314), .ZN(
        P2_U2967) );
  INV_X1 U17290 ( .A(n19860), .ZN(n18027) );
  NOR2_X1 U17291 ( .A1(n17188), .A2(n14651), .ZN(n15317) );
  AOI21_X1 U17292 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n14651), .A(n15317), .ZN(
        n15318) );
  OAI21_X1 U17293 ( .B1(n18027), .B2(n17272), .A(n15318), .ZN(P2_U2886) );
  OAI211_X1 U17294 ( .C1(n12847), .C2(n12895), .A(n15320), .B(n15319), .ZN(
        n15321) );
  NAND2_X1 U17295 ( .A1(n15321), .A2(n12891), .ZN(n15327) );
  AOI21_X1 U17296 ( .B1(n12899), .B2(n12891), .A(n15813), .ZN(n15322) );
  NAND2_X1 U17297 ( .A1(n15323), .A2(n15322), .ZN(n15342) );
  NAND2_X1 U17298 ( .A1(n12914), .A2(n16376), .ZN(n15326) );
  NAND2_X1 U17299 ( .A1(n15324), .A2(n12895), .ZN(n15325) );
  AND4_X1 U17300 ( .A1(n15327), .A2(n15342), .A3(n15326), .A4(n15325), .ZN(
        n15391) );
  AND3_X1 U17301 ( .A1(n13660), .A2(n15328), .A3(n12917), .ZN(n15329) );
  AND3_X1 U17302 ( .A1(n15391), .A2(n15329), .A3(n11164), .ZN(n17063) );
  XNOR2_X1 U17303 ( .A(n17059), .B(n11312), .ZN(n15337) );
  AND2_X1 U17304 ( .A1(n17062), .A2(n15337), .ZN(n15333) );
  NAND2_X1 U17305 ( .A1(n15330), .A2(n16419), .ZN(n15331) );
  OR2_X1 U17306 ( .A1(n16366), .A2(n15373), .ZN(n17052) );
  INV_X1 U17307 ( .A(n15337), .ZN(n15332) );
  AOI22_X1 U17308 ( .A1(n17063), .A2(n15333), .B1(n17052), .B2(n15332), .ZN(
        n15336) );
  NAND2_X1 U17309 ( .A1(n17058), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15334) );
  NAND2_X1 U17310 ( .A1(n17058), .A2(n11623), .ZN(n17066) );
  MUX2_X1 U17311 ( .A(n15334), .B(n17066), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n15335) );
  OAI211_X1 U17312 ( .C1(n16674), .C2(n17063), .A(n15336), .B(n15335), .ZN(
        n17866) );
  INV_X1 U17313 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15393) );
  AOI22_X1 U17314 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n16934), .B2(n15393), .ZN(
        n17042) );
  INV_X1 U17315 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n22123) );
  NOR2_X1 U17316 ( .A1(n22250), .A2(n22123), .ZN(n17044) );
  AOI222_X1 U17317 ( .A1(n17866), .A2(n17824), .B1(n17042), .B2(n17044), .C1(
        n22259), .C2(n15337), .ZN(n15352) );
  OAI21_X1 U17318 ( .B1(n17058), .B2(n13659), .A(n16375), .ZN(n15338) );
  NAND2_X1 U17319 ( .A1(n15338), .A2(n15378), .ZN(n15340) );
  NOR2_X1 U17320 ( .A1(n16371), .A2(n22296), .ZN(n15339) );
  NAND2_X1 U17321 ( .A1(n15340), .A2(n15339), .ZN(n15350) );
  INV_X1 U17322 ( .A(n15341), .ZN(n15343) );
  NAND2_X1 U17323 ( .A1(n15343), .A2(n15342), .ZN(n15344) );
  NAND2_X1 U17324 ( .A1(n16370), .A2(n15344), .ZN(n15365) );
  NOR2_X1 U17325 ( .A1(n12883), .A2(n12895), .ZN(n15345) );
  AOI22_X1 U17326 ( .A1(n16366), .A2(n16371), .B1(n15345), .B2(n12891), .ZN(
        n15346) );
  NAND2_X1 U17327 ( .A1(n15365), .A2(n15346), .ZN(n15347) );
  NOR2_X1 U17328 ( .A1(n15348), .A2(n15347), .ZN(n15349) );
  NAND2_X1 U17329 ( .A1(n15350), .A2(n15349), .ZN(n17888) );
  INV_X1 U17330 ( .A(n17888), .ZN(n17870) );
  OR2_X1 U17331 ( .A1(n22256), .A2(n22255), .ZN(n15433) );
  OAI22_X1 U17332 ( .A1(n17870), .A2(n22265), .B1(n15433), .B2(n22246), .ZN(
        n17823) );
  AOI21_X1 U17333 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22256), .A(n17823), 
        .ZN(n17047) );
  NAND2_X1 U17334 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n17047), .ZN(
        n15351) );
  OAI21_X1 U17335 ( .B1(n15352), .B2(n17047), .A(n15351), .ZN(P1_U3472) );
  INV_X1 U17336 ( .A(n17063), .ZN(n17068) );
  NAND2_X1 U17337 ( .A1(n13083), .A2(n17068), .ZN(n15355) );
  NAND2_X1 U17338 ( .A1(n12846), .A2(n15353), .ZN(n15354) );
  NAND2_X1 U17339 ( .A1(n15355), .A2(n15354), .ZN(n17869) );
  INV_X1 U17340 ( .A(n22259), .ZN(n17070) );
  OAI22_X1 U17341 ( .A1(n22250), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n17070), .ZN(n15356) );
  AOI21_X1 U17342 ( .B1(n17869), .B2(n17824), .A(n15356), .ZN(n15358) );
  AND2_X1 U17343 ( .A1(n17058), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17868) );
  AOI22_X1 U17344 ( .A1(n17868), .A2(n17824), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n17047), .ZN(n15357) );
  OAI21_X1 U17345 ( .B1(n15358), .B2(n17047), .A(n15357), .ZN(P1_U3474) );
  XNOR2_X1 U17346 ( .A(n11163), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15528) );
  NAND2_X1 U17347 ( .A1(n12891), .A2(n22297), .ZN(n15362) );
  INV_X1 U17348 ( .A(n15360), .ZN(n15361) );
  NAND3_X1 U17349 ( .A1(n15362), .A2(n12883), .A3(n15361), .ZN(n15364) );
  NAND3_X1 U17350 ( .A1(n16371), .A2(n12846), .A3(n12891), .ZN(n15363) );
  NAND3_X1 U17351 ( .A1(n15365), .A2(n15364), .A3(n15363), .ZN(n15366) );
  NAND2_X1 U17352 ( .A1(n15366), .A2(n20704), .ZN(n15372) );
  OAI21_X1 U17353 ( .B1(n12891), .B2(n16375), .A(n22248), .ZN(n15802) );
  INV_X1 U17354 ( .A(n15802), .ZN(n15367) );
  NAND2_X1 U17355 ( .A1(n13659), .A2(n15367), .ZN(n15368) );
  NAND3_X1 U17356 ( .A1(n15368), .A2(n12895), .A3(n12884), .ZN(n15369) );
  NAND3_X1 U17357 ( .A1(n15370), .A2(n15598), .A3(n15369), .ZN(n15371) );
  INV_X1 U17358 ( .A(n15373), .ZN(n15374) );
  NAND2_X1 U17359 ( .A1(n15375), .A2(n15374), .ZN(n16364) );
  INV_X1 U17360 ( .A(n16364), .ZN(n15379) );
  INV_X1 U17361 ( .A(n15382), .ZN(n15376) );
  NAND2_X1 U17362 ( .A1(n15376), .A2(n15381), .ZN(n15377) );
  NAND4_X1 U17363 ( .A1(n15379), .A2(n11164), .A3(n15378), .A4(n15377), .ZN(
        n15380) );
  OAI21_X1 U17364 ( .B1(n15382), .B2(n15381), .A(n17862), .ZN(n15383) );
  INV_X1 U17365 ( .A(n15384), .ZN(n15564) );
  NAND2_X1 U17366 ( .A1(n16178), .A2(n15393), .ZN(n15385) );
  NAND2_X1 U17367 ( .A1(n16400), .A2(n22129), .ZN(n15386) );
  NAND2_X1 U17368 ( .A1(n15387), .A2(n15386), .ZN(n15462) );
  MUX2_X1 U17369 ( .A(n11165), .B(n16178), .S(P1_EBX_REG_0__SCAN_IN), .Z(
        n15516) );
  XNOR2_X1 U17370 ( .A(n15462), .B(n15516), .ZN(n15388) );
  NAND2_X1 U17371 ( .A1(n15388), .A2(n16419), .ZN(n15463) );
  OAI21_X1 U17372 ( .B1(n15388), .B2(n16419), .A(n15463), .ZN(n22125) );
  INV_X1 U17373 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20592) );
  NOR2_X1 U17374 ( .A1(n22093), .A2(n20592), .ZN(n15524) );
  NAND2_X1 U17375 ( .A1(n15395), .A2(n17058), .ZN(n22122) );
  NAND2_X1 U17376 ( .A1(n15389), .A2(n15813), .ZN(n15390) );
  NAND2_X1 U17377 ( .A1(n15391), .A2(n15390), .ZN(n15392) );
  NAND2_X1 U17378 ( .A1(n15395), .A2(n15392), .ZN(n22111) );
  INV_X1 U17379 ( .A(n17025), .ZN(n22039) );
  NAND2_X1 U17380 ( .A1(n22123), .A2(n22122), .ZN(n15466) );
  AND3_X1 U17381 ( .A1(n22039), .A2(n15393), .A3(n15466), .ZN(n15394) );
  AOI211_X1 U17382 ( .C1(n22106), .C2(n22125), .A(n15524), .B(n15394), .ZN(
        n15399) );
  OR2_X1 U17383 ( .A1(n22111), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15396) );
  OR2_X1 U17384 ( .A1(n15395), .A2(n22102), .ZN(n22121) );
  OAI21_X1 U17385 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n22112), .A(
        n22016), .ZN(n15397) );
  NAND2_X1 U17386 ( .A1(n15397), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15398) );
  OAI211_X1 U17387 ( .C1(n15528), .C2(n22043), .A(n15399), .B(n15398), .ZN(
        P1_U3030) );
  AOI22_X1 U17388 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n18068), .B1(n19016), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n15400) );
  OAI21_X1 U17389 ( .B1(n15401), .B2(n15420), .A(n15400), .ZN(P2_U2935) );
  INV_X1 U17390 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n17344) );
  AOI22_X1 U17391 ( .A1(n15414), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n15402) );
  OAI21_X1 U17392 ( .B1(n17344), .B2(n15420), .A(n15402), .ZN(P2_U2929) );
  INV_X1 U17393 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15404) );
  AOI22_X1 U17394 ( .A1(n15414), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n15403) );
  OAI21_X1 U17395 ( .B1(n15404), .B2(n15420), .A(n15403), .ZN(P2_U2930) );
  INV_X1 U17396 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n15406) );
  AOI22_X1 U17397 ( .A1(n15414), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n15405) );
  OAI21_X1 U17398 ( .B1(n15406), .B2(n15420), .A(n15405), .ZN(P2_U2923) );
  INV_X1 U17399 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n15408) );
  AOI22_X1 U17400 ( .A1(n15414), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n15407) );
  OAI21_X1 U17401 ( .B1(n15408), .B2(n15420), .A(n15407), .ZN(P2_U2927) );
  AOI22_X1 U17402 ( .A1(n15414), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n15409) );
  OAI21_X1 U17403 ( .B1(n15410), .B2(n15420), .A(n15409), .ZN(P2_U2924) );
  INV_X1 U17404 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n17366) );
  AOI22_X1 U17405 ( .A1(n15414), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n15411) );
  OAI21_X1 U17406 ( .B1(n17366), .B2(n15420), .A(n15411), .ZN(P2_U2932) );
  INV_X1 U17407 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n17321) );
  AOI22_X1 U17408 ( .A1(n15414), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n15412) );
  OAI21_X1 U17409 ( .B1(n17321), .B2(n15420), .A(n15412), .ZN(P2_U2926) );
  INV_X1 U17410 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n17310) );
  AOI22_X1 U17411 ( .A1(n15414), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n15413) );
  OAI21_X1 U17412 ( .B1(n17310), .B2(n15420), .A(n15413), .ZN(P2_U2925) );
  INV_X1 U17413 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U17414 ( .A1(n15414), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n15415) );
  OAI21_X1 U17415 ( .B1(n17357), .B2(n15420), .A(n15415), .ZN(P2_U2931) );
  INV_X1 U17416 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n17333) );
  AOI22_X1 U17417 ( .A1(n19016), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n15416) );
  OAI21_X1 U17418 ( .B1(n17333), .B2(n15420), .A(n15416), .ZN(P2_U2928) );
  INV_X1 U17419 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15418) );
  AOI22_X1 U17420 ( .A1(n19016), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n15417) );
  OAI21_X1 U17421 ( .B1(n15418), .B2(n15420), .A(n15417), .ZN(P2_U2922) );
  INV_X1 U17422 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n15421) );
  AOI22_X1 U17423 ( .A1(n19016), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n15419) );
  OAI21_X1 U17424 ( .B1(n15421), .B2(n15420), .A(n15419), .ZN(P2_U2921) );
  MUX2_X1 U17425 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n17905), .S(n17281), .Z(
        n15422) );
  AOI21_X1 U17426 ( .B1(n18023), .B2(n17274), .A(n15422), .ZN(n15423) );
  INV_X1 U17427 ( .A(n15423), .ZN(P2_U2885) );
  OR2_X1 U17428 ( .A1(n15425), .A2(n15424), .ZN(n15426) );
  NAND2_X1 U17429 ( .A1(n15426), .A2(n15492), .ZN(n19077) );
  INV_X1 U17430 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n18070) );
  OAI222_X1 U17431 ( .A1(n19077), .A2(n15793), .B1(n15427), .B2(n20257), .C1(
        n18070), .C2(n20153), .ZN(P2_U2909) );
  NAND2_X1 U17432 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22489), .ZN(n22253) );
  INV_X1 U17433 ( .A(n15429), .ZN(n15431) );
  OAI21_X1 U17434 ( .B1(n15431), .B2(n15430), .A(n17889), .ZN(n15432) );
  NAND2_X1 U17435 ( .A1(n15432), .A2(n22246), .ZN(n17034) );
  AOI21_X1 U17436 ( .B1(n17034), .B2(n22246), .A(n15433), .ZN(n15434) );
  OR2_X1 U17437 ( .A1(n15593), .A2(n15434), .ZN(n17898) );
  NAND2_X1 U17438 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22452), .ZN(n17036) );
  NAND2_X1 U17439 ( .A1(n17898), .A2(n17036), .ZN(n16352) );
  INV_X1 U17440 ( .A(n17898), .ZN(n16350) );
  NAND2_X1 U17441 ( .A1(n16350), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15438) );
  XNOR2_X1 U17442 ( .A(n15961), .B(n22416), .ZN(n15436) );
  NAND3_X1 U17443 ( .A1(n15436), .A2(n22497), .A3(n17898), .ZN(n15437) );
  OAI211_X1 U17444 ( .C1(n16352), .C2(n16674), .A(n15438), .B(n15437), .ZN(
        P1_U3476) );
  INV_X1 U17445 ( .A(n19982), .ZN(n19876) );
  NAND2_X1 U17446 ( .A1(n19330), .A2(n17281), .ZN(n15441) );
  NAND2_X1 U17447 ( .A1(n14651), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n15440) );
  OAI211_X1 U17448 ( .C1(n19876), .C2(n17272), .A(n15441), .B(n15440), .ZN(
        P2_U2884) );
  INV_X1 U17449 ( .A(n16771), .ZN(n15445) );
  INV_X1 U17450 ( .A(n15442), .ZN(n15443) );
  XNOR2_X1 U17451 ( .A(n15444), .B(n15443), .ZN(n22135) );
  INV_X1 U17452 ( .A(n22135), .ZN(n15451) );
  OAI222_X1 U17453 ( .A1(n15445), .A2(n16791), .B1(n16789), .B2(n13076), .C1(
        n16782), .C2(n15451), .ZN(P1_U2903) );
  NAND3_X1 U17454 ( .A1(n16366), .A2(n20704), .A3(n16371), .ZN(n15449) );
  INV_X1 U17455 ( .A(n15446), .ZN(n15447) );
  NAND4_X1 U17456 ( .A1(n15447), .A2(n16726), .A3(n17062), .A4(n16419), .ZN(
        n15448) );
  INV_X1 U17457 ( .A(n20621), .ZN(n16703) );
  AOI22_X1 U17458 ( .A1(n20617), .A2(n22125), .B1(n16703), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n15450) );
  OAI21_X1 U17459 ( .B1(n15451), .B2(n16723), .A(n15450), .ZN(P1_U2871) );
  INV_X1 U17460 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15453) );
  AOI22_X1 U17461 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20514), .B1(n21955), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n15452) );
  OAI21_X1 U17462 ( .B1(n15453), .B2(n15485), .A(n15452), .ZN(P1_U2920) );
  XNOR2_X1 U17463 ( .A(n15455), .B(n15454), .ZN(n15523) );
  NAND2_X1 U17464 ( .A1(n16178), .A2(n15456), .ZN(n15458) );
  NAND2_X1 U17465 ( .A1(n16419), .A2(n15459), .ZN(n15457) );
  NAND3_X1 U17466 ( .A1(n15458), .A2(n15457), .A3(n11165), .ZN(n15461) );
  NAND2_X1 U17467 ( .A1(n16400), .A2(n15459), .ZN(n15460) );
  AND2_X1 U17468 ( .A1(n15461), .A2(n15460), .ZN(n15465) );
  NAND2_X1 U17469 ( .A1(n15463), .A2(n15462), .ZN(n15464) );
  AOI21_X1 U17470 ( .B1(n15465), .B2(n15464), .A(n15825), .ZN(n16675) );
  NAND2_X1 U17471 ( .A1(n21982), .A2(n15466), .ZN(n22022) );
  NOR2_X1 U17472 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n22022), .ZN(
        n15467) );
  AOI21_X1 U17473 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n16174) );
  INV_X1 U17474 ( .A(n16174), .ZN(n16016) );
  NOR2_X1 U17475 ( .A1(n22112), .A2(n16016), .ZN(n21981) );
  INV_X1 U17476 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20529) );
  NOR2_X1 U17477 ( .A1(n22093), .A2(n20529), .ZN(n15518) );
  AOI211_X1 U17478 ( .C1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n15467), .A(
        n21981), .B(n15518), .ZN(n15468) );
  INV_X1 U17479 ( .A(n15468), .ZN(n15469) );
  AOI21_X1 U17480 ( .B1(n16675), .B2(n22106), .A(n15469), .ZN(n15473) );
  NAND2_X1 U17481 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15470) );
  OAI22_X1 U17482 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n22018), .B1(
        n15470), .B2(n22112), .ZN(n15471) );
  OAI21_X1 U17483 ( .B1(n15471), .B2(n21980), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15472) );
  OAI211_X1 U17484 ( .C1(n15523), .C2(n22043), .A(n15473), .B(n15472), .ZN(
        P1_U3029) );
  INV_X1 U17485 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n15475) );
  AOI22_X1 U17486 ( .A1(n21955), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n15474) );
  OAI21_X1 U17487 ( .B1(n15475), .B2(n15485), .A(n15474), .ZN(P1_U2918) );
  AOI22_X1 U17488 ( .A1(n21955), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n15476) );
  OAI21_X1 U17489 ( .B1(n15241), .B2(n15485), .A(n15476), .ZN(P1_U2917) );
  AOI22_X1 U17490 ( .A1(n21955), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n15477) );
  OAI21_X1 U17491 ( .B1(n22369), .B2(n15485), .A(n15477), .ZN(P1_U2907) );
  AOI22_X1 U17492 ( .A1(n21955), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n15478) );
  OAI21_X1 U17493 ( .B1(n13533), .B2(n15485), .A(n15478), .ZN(P1_U2908) );
  AOI22_X1 U17494 ( .A1(n21955), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n15479) );
  OAI21_X1 U17495 ( .B1(n22375), .B2(n15485), .A(n15479), .ZN(P1_U2906) );
  AOI22_X1 U17496 ( .A1(n21955), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n15480) );
  OAI21_X1 U17497 ( .B1(n13511), .B2(n15485), .A(n15480), .ZN(P1_U2909) );
  AOI22_X1 U17498 ( .A1(n21955), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n15481) );
  OAI21_X1 U17499 ( .B1(n13488), .B2(n15485), .A(n15481), .ZN(P1_U2910) );
  AOI22_X1 U17500 ( .A1(n21955), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n15482) );
  OAI21_X1 U17501 ( .B1(n15483), .B2(n15485), .A(n15482), .ZN(P1_U2916) );
  AOI22_X1 U17502 ( .A1(n21955), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n15484) );
  OAI21_X1 U17503 ( .B1(n13304), .B2(n15485), .A(n15484), .ZN(P1_U2919) );
  XNOR2_X1 U17504 ( .A(n15486), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15490) );
  OR2_X1 U17505 ( .A1(n15487), .A2(n15496), .ZN(n15488) );
  NAND2_X1 U17506 ( .A1(n15488), .A2(n15529), .ZN(n19286) );
  MUX2_X1 U17507 ( .A(n12081), .B(n19286), .S(n17281), .Z(n15489) );
  OAI21_X1 U17508 ( .B1(n15490), .B2(n17272), .A(n15489), .ZN(P2_U2880) );
  AOI21_X1 U17509 ( .B1(n15493), .B2(n15492), .A(n15491), .ZN(n19238) );
  INV_X1 U17510 ( .A(n19238), .ZN(n15495) );
  INV_X1 U17511 ( .A(n17300), .ZN(n15494) );
  OAI222_X1 U17512 ( .A1(n15495), .A2(n15793), .B1(n15494), .B2(n20257), .C1(
        n18072), .C2(n20153), .ZN(P2_U2908) );
  AOI21_X1 U17513 ( .B1(n15497), .B2(n16121), .A(n15496), .ZN(n19298) );
  INV_X1 U17514 ( .A(n19298), .ZN(n17533) );
  NOR2_X1 U17515 ( .A1(n15498), .A2(n20108), .ZN(n15500) );
  INV_X1 U17516 ( .A(n15486), .ZN(n15499) );
  OAI211_X1 U17517 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n15500), .A(
        n15499), .B(n17274), .ZN(n15502) );
  NAND2_X1 U17518 ( .A1(n14651), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n15501) );
  OAI211_X1 U17519 ( .C1(n17533), .C2(n14651), .A(n15502), .B(n15501), .ZN(
        P2_U2881) );
  OR2_X1 U17520 ( .A1(n15503), .A2(n15491), .ZN(n15504) );
  NAND2_X1 U17521 ( .A1(n15504), .A2(n17689), .ZN(n19089) );
  INV_X1 U17522 ( .A(n17293), .ZN(n15505) );
  INV_X1 U17523 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n18074) );
  OAI222_X1 U17524 ( .A1(n19089), .A2(n15793), .B1(n15505), .B2(n20257), .C1(
        n18074), .C2(n20153), .ZN(P2_U2907) );
  INV_X1 U17525 ( .A(n22384), .ZN(n15510) );
  AOI21_X1 U17526 ( .B1(n15913), .B2(n22416), .A(n22506), .ZN(n15904) );
  INV_X1 U17527 ( .A(n22416), .ZN(n15734) );
  OAI21_X1 U17528 ( .B1(n15961), .B2(n15734), .A(n15962), .ZN(n15507) );
  NAND3_X1 U17529 ( .A1(n15904), .A2(n17898), .A3(n15507), .ZN(n15509) );
  NAND2_X1 U17530 ( .A1(n16350), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15508) );
  OAI211_X1 U17531 ( .C1(n15510), .C2(n16352), .A(n15509), .B(n15508), .ZN(
        P1_U3475) );
  INV_X1 U17532 ( .A(n15511), .ZN(n15512) );
  AOI21_X1 U17533 ( .B1(n15514), .B2(n15513), .A(n15512), .ZN(n15521) );
  INV_X1 U17534 ( .A(n15521), .ZN(n16685) );
  AOI22_X1 U17535 ( .A1(n16675), .A2(n20617), .B1(n16703), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n15515) );
  OAI21_X1 U17536 ( .B1(n16685), .B2(n16723), .A(n15515), .ZN(P1_U2870) );
  OAI21_X1 U17537 ( .B1(n16440), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n15516), .ZN(n22114) );
  INV_X1 U17538 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n15808) );
  OAI222_X1 U17539 ( .A1(n22114), .A2(n16724), .B1(n15808), .B2(n20621), .C1(
        n20623), .C2(n20634), .ZN(P1_U2872) );
  INV_X1 U17540 ( .A(n16768), .ZN(n15517) );
  OAI222_X1 U17541 ( .A1(n16685), .A2(n16782), .B1(n16791), .B2(n15517), .C1(
        n16789), .C2(n13067), .ZN(P1_U2902) );
  AOI21_X1 U17542 ( .B1(n20694), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n15518), .ZN(n15519) );
  OAI21_X1 U17543 ( .B1(n20703), .B2(n16677), .A(n15519), .ZN(n15520) );
  AOI21_X1 U17544 ( .B1(n15521), .B2(n20689), .A(n15520), .ZN(n15522) );
  OAI21_X1 U17545 ( .B1(n20696), .B2(n15523), .A(n15522), .ZN(P1_U2997) );
  AOI21_X1 U17546 ( .B1(n20694), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15524), .ZN(n15525) );
  OAI21_X1 U17547 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15525), .ZN(n15526) );
  AOI21_X1 U17548 ( .B1(n22135), .B2(n20689), .A(n15526), .ZN(n15527) );
  OAI21_X1 U17549 ( .B1(n15528), .B2(n20696), .A(n15527), .ZN(P1_U2998) );
  NAND2_X1 U17550 ( .A1(n15530), .A2(n15529), .ZN(n15533) );
  INV_X1 U17551 ( .A(n15531), .ZN(n15532) );
  INV_X1 U17552 ( .A(n19061), .ZN(n17764) );
  INV_X1 U17553 ( .A(n15534), .ZN(n15536) );
  OAI211_X1 U17554 ( .C1(n11181), .C2(n15536), .A(n17274), .B(n15535), .ZN(
        n15538) );
  NAND2_X1 U17555 ( .A1(n14651), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n15537) );
  OAI211_X1 U17556 ( .C1(n17764), .C2(n14651), .A(n15538), .B(n15537), .ZN(
        P2_U2879) );
  NAND3_X1 U17557 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n22409), .A3(
        n22476), .ZN(n15968) );
  INV_X1 U17558 ( .A(n15968), .ZN(n15546) );
  INV_X1 U17559 ( .A(n16347), .ZN(n15540) );
  NAND2_X1 U17560 ( .A1(n15540), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22492) );
  NOR2_X1 U17561 ( .A1(n16674), .A2(n15874), .ZN(n22432) );
  INV_X1 U17562 ( .A(n15842), .ZN(n22488) );
  NOR2_X1 U17563 ( .A1(n22487), .A2(n15968), .ZN(n15600) );
  AOI21_X1 U17564 ( .B1(n22432), .B2(n22488), .A(n15600), .ZN(n15544) );
  OAI211_X1 U17565 ( .C1(n15621), .C2(n22492), .A(n22497), .B(n15544), .ZN(
        n15541) );
  OAI211_X1 U17566 ( .C1(n22497), .C2(n15546), .A(n22495), .B(n15541), .ZN(
        n15542) );
  INV_X1 U17567 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15554) );
  OR2_X1 U17568 ( .A1(n16731), .A2(n20697), .ZN(n15596) );
  INV_X1 U17569 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20745) );
  NAND2_X1 U17570 ( .A1(n15593), .A2(n16777), .ZN(n22485) );
  INV_X1 U17571 ( .A(n15544), .ZN(n15545) );
  NAND2_X1 U17572 ( .A1(n15545), .A2(n22497), .ZN(n15548) );
  NAND2_X1 U17573 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15546), .ZN(n15547) );
  NAND2_X1 U17574 ( .A1(n15548), .A2(n15547), .ZN(n15594) );
  AOI22_X1 U17575 ( .A1(n22727), .A2(n22477), .B1(n22507), .B2(n15594), .ZN(
        n15553) );
  INV_X1 U17576 ( .A(n15596), .ZN(n15580) );
  NAND2_X1 U17577 ( .A1(n15580), .A2(DATAI_24_), .ZN(n15550) );
  INV_X1 U17578 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20761) );
  OR2_X1 U17579 ( .A1(n15595), .A2(n20761), .ZN(n15549) );
  AND2_X1 U17580 ( .A1(n15550), .A2(n15549), .ZN(n22386) );
  INV_X1 U17581 ( .A(n22386), .ZN(n22515) );
  NOR2_X2 U17582 ( .A1(n15599), .A2(n15813), .ZN(n22508) );
  AOI22_X1 U17583 ( .A1(n15985), .A2(n22515), .B1(n15600), .B2(n22508), .ZN(
        n15552) );
  OAI211_X1 U17584 ( .C1(n15604), .C2(n15554), .A(n15553), .B(n15552), .ZN(
        P1_U3073) );
  INV_X1 U17585 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15560) );
  INV_X1 U17586 ( .A(DATAI_23_), .ZN(n15555) );
  INV_X1 U17587 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20759) );
  NAND2_X1 U17588 ( .A1(n15593), .A2(n16750), .ZN(n22758) );
  INV_X1 U17589 ( .A(n22758), .ZN(n22768) );
  AOI22_X1 U17590 ( .A1(n22727), .A2(n22753), .B1(n22768), .B2(n15594), .ZN(
        n15559) );
  INV_X1 U17591 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20776) );
  OAI22_X1 U17592 ( .A1(n15556), .A2(n15596), .B1(n20776), .B2(n15595), .ZN(
        n22771) );
  NOR2_X2 U17593 ( .A1(n15599), .A2(n15557), .ZN(n22770) );
  AOI22_X1 U17594 ( .A1(n15985), .A2(n11308), .B1(n22770), .B2(n15600), .ZN(
        n15558) );
  OAI211_X1 U17595 ( .C1(n15604), .C2(n15560), .A(n15559), .B(n15558), .ZN(
        P1_U3080) );
  INV_X1 U17596 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15567) );
  INV_X1 U17597 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20751) );
  NAND2_X1 U17598 ( .A1(n15593), .A2(n16764), .ZN(n22600) );
  INV_X1 U17599 ( .A(n22600), .ZN(n22603) );
  AOI22_X1 U17600 ( .A1(n22727), .A2(n22597), .B1(n22603), .B2(n15594), .ZN(
        n15566) );
  NAND2_X1 U17601 ( .A1(n15580), .A2(DATAI_27_), .ZN(n15563) );
  INV_X1 U17602 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20768) );
  OR2_X1 U17603 ( .A1(n15595), .A2(n20768), .ZN(n15562) );
  INV_X1 U17604 ( .A(n22581), .ZN(n22605) );
  NOR2_X2 U17605 ( .A1(n15599), .A2(n15564), .ZN(n22604) );
  AOI22_X1 U17606 ( .A1(n15985), .A2(n22605), .B1(n15600), .B2(n22604), .ZN(
        n15565) );
  OAI211_X1 U17607 ( .C1(n15604), .C2(n15567), .A(n15566), .B(n15565), .ZN(
        P1_U3076) );
  INV_X1 U17608 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15573) );
  INV_X1 U17609 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20753) );
  OAI22_X1 U17610 ( .A1(n15568), .A2(n15596), .B1(n20753), .B2(n15595), .ZN(
        n22627) );
  NAND2_X1 U17611 ( .A1(n15593), .A2(n16760), .ZN(n22630) );
  INV_X1 U17612 ( .A(n22630), .ZN(n22633) );
  AOI22_X1 U17613 ( .A1(n22727), .A2(n22627), .B1(n22633), .B2(n15594), .ZN(
        n15572) );
  INV_X1 U17614 ( .A(DATAI_28_), .ZN(n15569) );
  INV_X1 U17615 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20770) );
  OAI22_X1 U17616 ( .A1(n15569), .A2(n15596), .B1(n20770), .B2(n15595), .ZN(
        n22635) );
  NOR2_X2 U17617 ( .A1(n15599), .A2(n15570), .ZN(n22634) );
  AOI22_X1 U17618 ( .A1(n15985), .A2(n11310), .B1(n22634), .B2(n15600), .ZN(
        n15571) );
  OAI211_X1 U17619 ( .C1(n15604), .C2(n15573), .A(n15572), .B(n15571), .ZN(
        P1_U3077) );
  INV_X1 U17620 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15578) );
  INV_X1 U17621 ( .A(DATAI_21_), .ZN(n15574) );
  INV_X1 U17622 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20755) );
  NAND2_X1 U17623 ( .A1(n15593), .A2(n16756), .ZN(n22660) );
  INV_X1 U17624 ( .A(n22660), .ZN(n22663) );
  AOI22_X1 U17625 ( .A1(n22727), .A2(n22657), .B1(n22663), .B2(n15594), .ZN(
        n15577) );
  INV_X1 U17626 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20772) );
  OAI22_X1 U17627 ( .A1(n15575), .A2(n15596), .B1(n20772), .B2(n15595), .ZN(
        n22665) );
  NOR2_X2 U17628 ( .A1(n15599), .A2(n16726), .ZN(n22664) );
  AOI22_X1 U17629 ( .A1(n15985), .A2(n11306), .B1(n22664), .B2(n15600), .ZN(
        n15576) );
  OAI211_X1 U17630 ( .C1(n15604), .C2(n15578), .A(n15577), .B(n15576), .ZN(
        P1_U3078) );
  INV_X1 U17631 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15586) );
  INV_X1 U17632 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20757) );
  OAI22_X1 U17633 ( .A1(n15579), .A2(n15596), .B1(n20757), .B2(n15595), .ZN(
        n22686) );
  NAND2_X1 U17634 ( .A1(n15593), .A2(n16753), .ZN(n22689) );
  INV_X1 U17635 ( .A(n22689), .ZN(n22692) );
  AOI22_X1 U17636 ( .A1(n22727), .A2(n22686), .B1(n22692), .B2(n15594), .ZN(
        n15585) );
  NAND2_X1 U17637 ( .A1(n15580), .A2(DATAI_30_), .ZN(n15582) );
  INV_X1 U17638 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20774) );
  OR2_X1 U17639 ( .A1(n15595), .A2(n20774), .ZN(n15581) );
  AND2_X1 U17640 ( .A1(n15582), .A2(n15581), .ZN(n22670) );
  INV_X1 U17641 ( .A(n22670), .ZN(n22694) );
  NOR2_X2 U17642 ( .A1(n15599), .A2(n15583), .ZN(n22693) );
  AOI22_X1 U17643 ( .A1(n15985), .A2(n22694), .B1(n15600), .B2(n22693), .ZN(
        n15584) );
  OAI211_X1 U17644 ( .C1(n15604), .C2(n15586), .A(n15585), .B(n15584), .ZN(
        P1_U3079) );
  INV_X1 U17645 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15591) );
  INV_X1 U17646 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20747) );
  OAI22_X1 U17647 ( .A1(n15587), .A2(n15596), .B1(n20747), .B2(n15595), .ZN(
        n22538) );
  NAND2_X1 U17648 ( .A1(n15593), .A2(n16771), .ZN(n22541) );
  INV_X1 U17649 ( .A(n22541), .ZN(n22544) );
  AOI22_X1 U17650 ( .A1(n22727), .A2(n11302), .B1(n22544), .B2(n15594), .ZN(
        n15590) );
  INV_X1 U17651 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20763) );
  OAI22_X1 U17652 ( .A1(n15588), .A2(n15596), .B1(n20763), .B2(n15595), .ZN(
        n22546) );
  NOR2_X2 U17653 ( .A1(n15599), .A2(n12888), .ZN(n22545) );
  AOI22_X1 U17654 ( .A1(n15985), .A2(n11304), .B1(n22545), .B2(n15600), .ZN(
        n15589) );
  OAI211_X1 U17655 ( .C1(n15604), .C2(n15591), .A(n15590), .B(n15589), .ZN(
        P1_U3074) );
  INV_X1 U17656 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15603) );
  INV_X1 U17657 ( .A(DATAI_18_), .ZN(n15592) );
  INV_X1 U17658 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20749) );
  OAI22_X1 U17659 ( .A1(n15592), .A2(n15596), .B1(n20749), .B2(n15595), .ZN(
        n22568) );
  NAND2_X1 U17660 ( .A1(n15593), .A2(n16768), .ZN(n22571) );
  INV_X1 U17661 ( .A(n22571), .ZN(n22574) );
  AOI22_X1 U17662 ( .A1(n22727), .A2(n22568), .B1(n22574), .B2(n15594), .ZN(
        n15602) );
  INV_X1 U17663 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20766) );
  NOR2_X2 U17664 ( .A1(n15599), .A2(n15598), .ZN(n22575) );
  AOI22_X1 U17665 ( .A1(n15985), .A2(n22576), .B1(n22575), .B2(n15600), .ZN(
        n15601) );
  OAI211_X1 U17666 ( .C1(n15604), .C2(n15603), .A(n15602), .B(n15601), .ZN(
        P1_U3075) );
  INV_X1 U17667 ( .A(n16764), .ZN(n15608) );
  OAI21_X1 U17668 ( .B1(n15607), .B2(n15606), .A(n15605), .ZN(n20604) );
  OAI222_X1 U17669 ( .A1(n16791), .A2(n15608), .B1(n16789), .B2(n13098), .C1(
        n16782), .C2(n20604), .ZN(P1_U2901) );
  NAND3_X1 U17670 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n22409), .ZN(n22435) );
  INV_X1 U17671 ( .A(n22435), .ZN(n15618) );
  INV_X1 U17672 ( .A(n15609), .ZN(n15610) );
  NAND2_X1 U17673 ( .A1(n15610), .A2(n13083), .ZN(n22418) );
  INV_X1 U17674 ( .A(n22418), .ZN(n15906) );
  NOR2_X1 U17675 ( .A1(n15611), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15727) );
  AOI21_X1 U17676 ( .B1(n22432), .B2(n15906), .A(n15727), .ZN(n15616) );
  OAI211_X1 U17677 ( .C1(n15621), .C2(n15734), .A(n22497), .B(n15616), .ZN(
        n15612) );
  OAI211_X1 U17678 ( .C1(n22497), .C2(n15618), .A(n22495), .B(n15612), .ZN(
        n15613) );
  INV_X1 U17679 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15624) );
  INV_X1 U17680 ( .A(n15616), .ZN(n15617) );
  NAND2_X1 U17681 ( .A1(n15617), .A2(n22497), .ZN(n15620) );
  NAND2_X1 U17682 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15618), .ZN(n15619) );
  NAND2_X1 U17683 ( .A1(n15620), .A2(n15619), .ZN(n15726) );
  AOI22_X1 U17684 ( .A1(n22735), .A2(n22753), .B1(n22768), .B2(n15726), .ZN(
        n15623) );
  AOI22_X1 U17685 ( .A1(n22728), .A2(n11308), .B1(n22770), .B2(n15727), .ZN(
        n15622) );
  OAI211_X1 U17686 ( .C1(n15731), .C2(n15624), .A(n15623), .B(n15622), .ZN(
        P1_U3096) );
  INV_X1 U17687 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15627) );
  AOI22_X1 U17688 ( .A1(n22735), .A2(n22657), .B1(n22663), .B2(n15726), .ZN(
        n15626) );
  AOI22_X1 U17689 ( .A1(n22728), .A2(n11306), .B1(n22664), .B2(n15727), .ZN(
        n15625) );
  OAI211_X1 U17690 ( .C1(n15731), .C2(n15627), .A(n15626), .B(n15625), .ZN(
        P1_U3094) );
  INV_X1 U17691 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15630) );
  AOI22_X1 U17692 ( .A1(n22728), .A2(n22605), .B1(n22603), .B2(n15726), .ZN(
        n15629) );
  AOI22_X1 U17693 ( .A1(n22735), .A2(n22597), .B1(n22604), .B2(n15727), .ZN(
        n15628) );
  OAI211_X1 U17694 ( .C1(n15731), .C2(n15630), .A(n15629), .B(n15628), .ZN(
        P1_U3092) );
  INV_X1 U17695 ( .A(n15631), .ZN(n15642) );
  NAND2_X1 U17696 ( .A1(n14120), .A2(n15632), .ZN(n15633) );
  NOR2_X1 U17697 ( .A1(n15634), .A2(n15633), .ZN(n17818) );
  AOI22_X1 U17698 ( .A1(n15641), .A2(n15648), .B1(n15635), .B2(n15699), .ZN(
        n15640) );
  OAI22_X1 U17699 ( .A1(n17843), .A2(n12003), .B1(n15636), .B2(n15708), .ZN(
        n15638) );
  NAND2_X1 U17700 ( .A1(n15638), .A2(n15637), .ZN(n15639) );
  OAI211_X1 U17701 ( .C1(n15650), .C2(n15641), .A(n15640), .B(n15639), .ZN(
        n19352) );
  NOR3_X1 U17702 ( .A1(n15642), .A2(n17818), .A3(n19352), .ZN(n15705) );
  NOR2_X1 U17704 ( .A1(n11792), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15671) );
  OAI21_X1 U17705 ( .B1(n15644), .B2(n14202), .A(n15643), .ZN(n15670) );
  INV_X1 U17706 ( .A(n14071), .ZN(n15645) );
  NAND2_X1 U17707 ( .A1(n14180), .A2(n15645), .ZN(n15646) );
  NAND2_X1 U17708 ( .A1(n15670), .A2(n15646), .ZN(n15647) );
  NOR2_X1 U17709 ( .A1(n15671), .A2(n15647), .ZN(n15653) );
  INV_X1 U17710 ( .A(n15648), .ZN(n15649) );
  NAND2_X1 U17711 ( .A1(n15650), .A2(n15649), .ZN(n15666) );
  INV_X1 U17712 ( .A(n15671), .ZN(n15651) );
  AOI22_X1 U17713 ( .A1(n15666), .A2(n15651), .B1(n14071), .B2(n14180), .ZN(
        n15652) );
  MUX2_X1 U17714 ( .A(n15653), .B(n15652), .S(n11936), .Z(n15655) );
  NAND2_X1 U17715 ( .A1(n15655), .A2(n15654), .ZN(n15656) );
  AOI21_X1 U17716 ( .B1(n19330), .B2(n15681), .A(n15656), .ZN(n17786) );
  NAND2_X1 U17717 ( .A1(n15657), .A2(n19342), .ZN(n15663) );
  NAND2_X1 U17718 ( .A1(n15659), .A2(n15658), .ZN(n15660) );
  NOR2_X1 U17719 ( .A1(n15661), .A2(n15660), .ZN(n15662) );
  INV_X1 U17720 ( .A(n17773), .ZN(n15687) );
  NAND2_X1 U17721 ( .A1(n17786), .A2(n15687), .ZN(n15665) );
  NAND2_X1 U17722 ( .A1(n17773), .A2(n11936), .ZN(n15664) );
  NAND2_X1 U17723 ( .A1(n15665), .A2(n15664), .ZN(n15695) );
  INV_X1 U17724 ( .A(n15695), .ZN(n15697) );
  OAI21_X1 U17725 ( .B1(n11786), .B2(n15671), .A(n15666), .ZN(n15669) );
  NAND2_X1 U17726 ( .A1(n14180), .A2(n15667), .ZN(n15668) );
  OAI211_X1 U17727 ( .C1(n15671), .C2(n15670), .A(n15669), .B(n15668), .ZN(
        n15672) );
  AOI21_X1 U17728 ( .B1(n17905), .B2(n15681), .A(n15672), .ZN(n17781) );
  AND2_X1 U17729 ( .A1(n17773), .A2(n15673), .ZN(n15674) );
  AOI21_X1 U17730 ( .B1(n17781), .B2(n15687), .A(n15674), .ZN(n15693) );
  AOI22_X1 U17731 ( .A1(n15697), .A2(n15693), .B1(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n17773), .ZN(n15704) );
  INV_X1 U17732 ( .A(n14180), .ZN(n15684) );
  NAND2_X1 U17733 ( .A1(n11171), .A2(n15681), .ZN(n15680) );
  INV_X1 U17734 ( .A(n14212), .ZN(n15676) );
  NAND2_X1 U17735 ( .A1(n15676), .A2(n15675), .ZN(n15682) );
  OAI21_X1 U17736 ( .B1(n15678), .B2(n15677), .A(n15682), .ZN(n15679) );
  OAI211_X1 U17737 ( .C1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n15684), .A(
        n15680), .B(n15679), .ZN(n17777) );
  INV_X1 U17738 ( .A(n17777), .ZN(n15691) );
  INV_X1 U17739 ( .A(n15681), .ZN(n15686) );
  INV_X1 U17740 ( .A(n15682), .ZN(n15683) );
  MUX2_X1 U17741 ( .A(n15684), .B(n15683), .S(n11761), .Z(n15685) );
  OAI21_X1 U17742 ( .B1(n19023), .B2(n15686), .A(n15685), .ZN(n17770) );
  AOI211_X1 U17743 ( .C1(n12216), .C2(n17777), .A(n20000), .B(n17770), .ZN(
        n15690) );
  INV_X1 U17744 ( .A(n17781), .ZN(n15688) );
  OAI21_X1 U17745 ( .B1(n15688), .B2(n19884), .A(n15687), .ZN(n15689) );
  AOI211_X1 U17746 ( .C1(n15691), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15690), .B(n15689), .ZN(n15692) );
  AOI21_X1 U17747 ( .B1(n15693), .B2(n19884), .A(n15692), .ZN(n15694) );
  OAI21_X1 U17748 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15695), .A(
        n15694), .ZN(n15696) );
  OAI211_X1 U17749 ( .C1(n15697), .C2(n18034), .A(n17845), .B(n15696), .ZN(
        n15703) );
  INV_X1 U17750 ( .A(n22312), .ZN(n15698) );
  AOI21_X1 U17751 ( .B1(n19009), .B2(n15698), .A(n22317), .ZN(n15700) );
  NOR3_X1 U17752 ( .A1(n15701), .A2(n15700), .A3(n15699), .ZN(n19351) );
  OAI21_X1 U17753 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19351), .ZN(n15702) );
  NAND4_X1 U17754 ( .A1(n15705), .A2(n15704), .A3(n15703), .A4(n15702), .ZN(
        n17809) );
  OR2_X1 U17755 ( .A1(n15706), .A2(n17809), .ZN(n15711) );
  NOR3_X1 U17756 ( .A1(n15709), .A2(n15708), .A3(n15707), .ZN(n15710) );
  OAI21_X1 U17757 ( .B1(n19345), .B2(n17901), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n15713) );
  NOR2_X1 U17758 ( .A1(n17901), .A2(n18016), .ZN(n17808) );
  INV_X1 U17759 ( .A(n17808), .ZN(n17844) );
  NAND2_X1 U17760 ( .A1(n15713), .A2(n17844), .ZN(P2_U3593) );
  INV_X1 U17761 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15716) );
  AOI22_X1 U17762 ( .A1(n22735), .A2(n11302), .B1(n22544), .B2(n15726), .ZN(
        n15715) );
  AOI22_X1 U17763 ( .A1(n22728), .A2(n11304), .B1(n22545), .B2(n15727), .ZN(
        n15714) );
  OAI211_X1 U17764 ( .C1(n15731), .C2(n15716), .A(n15715), .B(n15714), .ZN(
        P1_U3090) );
  INV_X1 U17765 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15719) );
  AOI22_X1 U17766 ( .A1(n22735), .A2(n22627), .B1(n22633), .B2(n15726), .ZN(
        n15718) );
  AOI22_X1 U17767 ( .A1(n22728), .A2(n11310), .B1(n22634), .B2(n15727), .ZN(
        n15717) );
  OAI211_X1 U17768 ( .C1(n15731), .C2(n15719), .A(n15718), .B(n15717), .ZN(
        P1_U3093) );
  INV_X1 U17769 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15722) );
  AOI22_X1 U17770 ( .A1(n22735), .A2(n22568), .B1(n22574), .B2(n15726), .ZN(
        n15721) );
  AOI22_X1 U17771 ( .A1(n22728), .A2(n22576), .B1(n22575), .B2(n15727), .ZN(
        n15720) );
  OAI211_X1 U17772 ( .C1(n15731), .C2(n15722), .A(n15721), .B(n15720), .ZN(
        P1_U3091) );
  INV_X1 U17773 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15725) );
  AOI22_X1 U17774 ( .A1(n22735), .A2(n22477), .B1(n22507), .B2(n15726), .ZN(
        n15724) );
  AOI22_X1 U17775 ( .A1(n22728), .A2(n22515), .B1(n15727), .B2(n22508), .ZN(
        n15723) );
  OAI211_X1 U17776 ( .C1(n15731), .C2(n15725), .A(n15724), .B(n15723), .ZN(
        P1_U3089) );
  INV_X1 U17777 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15730) );
  AOI22_X1 U17778 ( .A1(n22728), .A2(n22694), .B1(n22692), .B2(n15726), .ZN(
        n15729) );
  AOI22_X1 U17779 ( .A1(n22735), .A2(n22686), .B1(n22693), .B2(n15727), .ZN(
        n15728) );
  OAI211_X1 U17780 ( .C1(n15731), .C2(n15730), .A(n15729), .B(n15728), .ZN(
        P1_U3095) );
  INV_X1 U17781 ( .A(n22746), .ZN(n15765) );
  NOR3_X1 U17782 ( .A1(n15846), .A2(n22506), .A3(n15734), .ZN(n15735) );
  NAND3_X1 U17783 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n22408), .ZN(n22461) );
  INV_X1 U17784 ( .A(n22461), .ZN(n15736) );
  NAND2_X1 U17785 ( .A1(n15759), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n15740) );
  NAND2_X1 U17786 ( .A1(n15841), .A2(n15963), .ZN(n22472) );
  INV_X1 U17787 ( .A(n22604), .ZN(n22580) );
  OR2_X1 U17788 ( .A1(n22487), .A2(n22461), .ZN(n15761) );
  NAND2_X1 U17789 ( .A1(n22384), .A2(n16674), .ZN(n22456) );
  OAI21_X1 U17790 ( .B1(n22456), .B2(n22418), .A(n15761), .ZN(n15737) );
  AOI22_X1 U17791 ( .A1(n15737), .A2(n22497), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15736), .ZN(n15760) );
  OAI22_X1 U17792 ( .A1(n22580), .A2(n15761), .B1(n22600), .B2(n15760), .ZN(
        n15738) );
  AOI21_X1 U17793 ( .B1(n22754), .B2(n22597), .A(n15738), .ZN(n15739) );
  OAI211_X1 U17794 ( .C1(n22581), .C2(n15765), .A(n15740), .B(n15739), .ZN(
        P1_U3124) );
  NAND2_X1 U17795 ( .A1(n15759), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n15743) );
  INV_X1 U17796 ( .A(n22693), .ZN(n22669) );
  OAI22_X1 U17797 ( .A1(n22669), .A2(n15761), .B1(n22689), .B2(n15760), .ZN(
        n15741) );
  AOI21_X1 U17798 ( .B1(n22754), .B2(n22686), .A(n15741), .ZN(n15742) );
  OAI211_X1 U17799 ( .C1(n22670), .C2(n15765), .A(n15743), .B(n15742), .ZN(
        P1_U3127) );
  NAND2_X1 U17800 ( .A1(n15759), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n15746) );
  INV_X1 U17801 ( .A(n22634), .ZN(n22609) );
  OAI22_X1 U17802 ( .A1(n22609), .A2(n15761), .B1(n22630), .B2(n15760), .ZN(
        n15744) );
  AOI21_X1 U17803 ( .B1(n22754), .B2(n22627), .A(n15744), .ZN(n15745) );
  OAI211_X1 U17804 ( .C1(n15765), .C2(n11309), .A(n15746), .B(n15745), .ZN(
        P1_U3125) );
  NAND2_X1 U17805 ( .A1(n15759), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n15749) );
  INV_X1 U17806 ( .A(n22770), .ZN(n22699) );
  OAI22_X1 U17807 ( .A1(n22699), .A2(n15761), .B1(n22758), .B2(n15760), .ZN(
        n15747) );
  AOI21_X1 U17808 ( .B1(n22754), .B2(n22753), .A(n15747), .ZN(n15748) );
  OAI211_X1 U17809 ( .C1(n15765), .C2(n11307), .A(n15749), .B(n15748), .ZN(
        P1_U3128) );
  NAND2_X1 U17810 ( .A1(n15759), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n15752) );
  INV_X1 U17811 ( .A(n22508), .ZN(n22385) );
  OAI22_X1 U17812 ( .A1(n22385), .A2(n15761), .B1(n22485), .B2(n15760), .ZN(
        n15750) );
  AOI21_X1 U17813 ( .B1(n22754), .B2(n22477), .A(n15750), .ZN(n15751) );
  OAI211_X1 U17814 ( .C1(n22386), .C2(n15765), .A(n15752), .B(n15751), .ZN(
        P1_U3121) );
  NAND2_X1 U17815 ( .A1(n15759), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n15755) );
  INV_X1 U17816 ( .A(n22545), .ZN(n22519) );
  OAI22_X1 U17817 ( .A1(n22519), .A2(n15761), .B1(n22541), .B2(n15760), .ZN(
        n15753) );
  AOI21_X1 U17818 ( .B1(n22754), .B2(n11302), .A(n15753), .ZN(n15754) );
  OAI211_X1 U17819 ( .C1(n15765), .C2(n11303), .A(n15755), .B(n15754), .ZN(
        P1_U3122) );
  INV_X1 U17820 ( .A(n22576), .ZN(n22565) );
  NAND2_X1 U17821 ( .A1(n15759), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n15758) );
  INV_X1 U17822 ( .A(n22575), .ZN(n22549) );
  OAI22_X1 U17823 ( .A1(n22549), .A2(n15761), .B1(n22571), .B2(n15760), .ZN(
        n15756) );
  AOI21_X1 U17824 ( .B1(n22754), .B2(n22568), .A(n15756), .ZN(n15757) );
  OAI211_X1 U17825 ( .C1(n15765), .C2(n22565), .A(n15758), .B(n15757), .ZN(
        P1_U3123) );
  NAND2_X1 U17826 ( .A1(n15759), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n15764) );
  INV_X1 U17827 ( .A(n22664), .ZN(n22639) );
  OAI22_X1 U17828 ( .A1(n22639), .A2(n15761), .B1(n22660), .B2(n15760), .ZN(
        n15762) );
  AOI21_X1 U17829 ( .B1(n22754), .B2(n22657), .A(n15762), .ZN(n15763) );
  OAI211_X1 U17830 ( .C1(n15765), .C2(n11305), .A(n15764), .B(n15763), .ZN(
        P1_U3126) );
  AOI21_X1 U17831 ( .B1(n15767), .B2(n15605), .A(n15766), .ZN(n15788) );
  INV_X1 U17832 ( .A(n15788), .ZN(n15879) );
  INV_X1 U17833 ( .A(n16178), .ZN(n15768) );
  NAND2_X1 U17834 ( .A1(n16178), .A2(n21986), .ZN(n15770) );
  INV_X1 U17835 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n15871) );
  NAND2_X1 U17836 ( .A1(n16419), .A2(n15871), .ZN(n15769) );
  NAND3_X1 U17837 ( .A1(n15770), .A2(n15769), .A3(n11166), .ZN(n15772) );
  NAND2_X1 U17838 ( .A1(n16400), .A2(n15871), .ZN(n15771) );
  MUX2_X1 U17839 ( .A(n16430), .B(n11165), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n15774) );
  OR2_X1 U17840 ( .A1(n16440), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15773) );
  AND2_X1 U17841 ( .A1(n15774), .A2(n15773), .ZN(n15824) );
  NAND2_X1 U17842 ( .A1(n15825), .A2(n15824), .ZN(n15894) );
  XOR2_X1 U17843 ( .A(n15893), .B(n15894), .Z(n21990) );
  AOI22_X1 U17844 ( .A1(n21990), .A2(n20617), .B1(n16703), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n15775) );
  OAI21_X1 U17845 ( .B1(n15879), .B2(n20623), .A(n15775), .ZN(P1_U2868) );
  INV_X1 U17846 ( .A(n15535), .ZN(n15778) );
  OAI211_X1 U17847 ( .C1(n15778), .C2(n14381), .A(n17274), .B(n15777), .ZN(
        n15782) );
  OR2_X1 U17848 ( .A1(n15779), .A2(n15531), .ZN(n15780) );
  NAND2_X1 U17849 ( .A1(n15780), .A2(n15953), .ZN(n17952) );
  INV_X1 U17850 ( .A(n17952), .ZN(n17738) );
  NAND2_X1 U17851 ( .A1(n17738), .A2(n17281), .ZN(n15781) );
  OAI211_X1 U17852 ( .C1(n17281), .C2(n12091), .A(n15782), .B(n15781), .ZN(
        P2_U2878) );
  INV_X1 U17853 ( .A(n16760), .ZN(n15783) );
  INV_X1 U17854 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20511) );
  OAI222_X1 U17855 ( .A1(n15879), .A2(n16782), .B1(n16791), .B2(n15783), .C1(
        n20511), .C2(n16789), .ZN(P1_U2900) );
  XNOR2_X1 U17856 ( .A(n15785), .B(n15784), .ZN(n21987) );
  INV_X1 U17857 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20532) );
  NOR2_X1 U17858 ( .A1(n22093), .A2(n20532), .ZN(n21984) );
  AOI21_X1 U17859 ( .B1(n20694), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21984), .ZN(n15786) );
  OAI21_X1 U17860 ( .B1(n20703), .B2(n15866), .A(n15786), .ZN(n15787) );
  AOI21_X1 U17861 ( .B1(n15788), .B2(n20689), .A(n15787), .ZN(n15789) );
  OAI21_X1 U17862 ( .B1(n20696), .B2(n21987), .A(n15789), .ZN(P1_U2995) );
  OR2_X1 U17863 ( .A1(n15790), .A2(n17688), .ZN(n15791) );
  NAND2_X1 U17864 ( .A1(n15791), .A2(n16209), .ZN(n19256) );
  INV_X1 U17865 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n18077) );
  OAI222_X1 U17866 ( .A1(n19256), .A2(n15793), .B1(n15792), .B2(n20257), .C1(
        n18077), .C2(n20153), .ZN(P2_U2905) );
  NOR2_X1 U17867 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22260) );
  NAND2_X1 U17868 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n22260), .ZN(n17895) );
  NAND2_X1 U17869 ( .A1(n13053), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15794) );
  MUX2_X1 U17870 ( .A(n17895), .B(n15794), .S(n22256), .Z(n15795) );
  INV_X1 U17871 ( .A(n15795), .ZN(n15796) );
  NOR2_X1 U17872 ( .A1(n15796), .A2(n22102), .ZN(n15797) );
  NOR2_X1 U17873 ( .A1(n15805), .A2(n22250), .ZN(n15799) );
  OR2_X1 U17874 ( .A1(n15815), .A2(n12915), .ZN(n15800) );
  NOR2_X1 U17875 ( .A1(n15815), .A2(n15813), .ZN(n15812) );
  NAND2_X1 U17876 ( .A1(n22248), .A2(n22268), .ZN(n17861) );
  AND3_X1 U17877 ( .A1(n12891), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n17861), .ZN(
        n15801) );
  INV_X1 U17878 ( .A(n22114), .ZN(n15810) );
  NOR2_X1 U17879 ( .A1(n15802), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15811) );
  AND2_X1 U17880 ( .A1(n12891), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n15803) );
  NOR2_X1 U17881 ( .A1(n15811), .A2(n15803), .ZN(n15804) );
  AND2_X2 U17882 ( .A1(n22190), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22242) );
  AND2_X1 U17883 ( .A1(n15805), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15806) );
  OAI21_X1 U17884 ( .B1(n22242), .B2(n22216), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15807) );
  OAI21_X1 U17885 ( .B1(n22235), .B2(n15808), .A(n15807), .ZN(n15809) );
  AOI21_X1 U17886 ( .B1(n22199), .B2(n15810), .A(n15809), .ZN(n15817) );
  NAND2_X1 U17887 ( .A1(n15813), .A2(n12891), .ZN(n15814) );
  NOR2_X1 U17888 ( .A1(n15815), .A2(n15814), .ZN(n22127) );
  AOI22_X1 U17889 ( .A1(n22161), .A2(P1_REIP_REG_0__SCAN_IN), .B1(n13083), 
        .B2(n22127), .ZN(n15816) );
  OAI211_X1 U17890 ( .C1(n20634), .C2(n22124), .A(n15817), .B(n15816), .ZN(
        P1_U2840) );
  XOR2_X1 U17891 ( .A(n15818), .B(n15819), .Z(n21997) );
  NAND2_X1 U17892 ( .A1(n21997), .A2(n13804), .ZN(n15823) );
  INV_X1 U17893 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n15820) );
  NOR2_X1 U17894 ( .A1(n22093), .A2(n15820), .ZN(n21994) );
  NOR2_X1 U17895 ( .A1(n20703), .A2(n15827), .ZN(n15821) );
  AOI211_X1 U17896 ( .C1(n20694), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n21994), .B(n15821), .ZN(n15822) );
  OAI211_X1 U17897 ( .C1(n20697), .C2(n20604), .A(n15823), .B(n15822), .ZN(
        P1_U2996) );
  OR2_X1 U17898 ( .A1(n15825), .A2(n15824), .ZN(n15826) );
  AND2_X1 U17899 ( .A1(n15894), .A2(n15826), .ZN(n21995) );
  INV_X1 U17900 ( .A(n22190), .ZN(n22162) );
  AOI22_X1 U17901 ( .A1(n22242), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n22162), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n15830) );
  INV_X1 U17902 ( .A(n15827), .ZN(n15828) );
  NAND2_X1 U17903 ( .A1(n22216), .A2(n15828), .ZN(n15829) );
  OAI211_X1 U17904 ( .C1(n22235), .C2(n20607), .A(n15830), .B(n15829), .ZN(
        n15832) );
  NAND2_X1 U17905 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n16679) );
  NOR2_X1 U17906 ( .A1(n15820), .A2(n16679), .ZN(n15865) );
  AOI211_X1 U17907 ( .C1(n16679), .C2(n15820), .A(n15865), .B(n22197), .ZN(
        n15831) );
  AOI211_X1 U17908 ( .C1(n21995), .C2(n22199), .A(n15832), .B(n15831), .ZN(
        n15834) );
  NAND2_X1 U17909 ( .A1(n22384), .A2(n22127), .ZN(n15833) );
  OAI211_X1 U17910 ( .C1(n20604), .C2(n22124), .A(n15834), .B(n15833), .ZN(
        P1_U2837) );
  INV_X1 U17911 ( .A(n15835), .ZN(n15839) );
  INV_X1 U17912 ( .A(n15766), .ZN(n15838) );
  AOI21_X1 U17913 ( .B1(n15839), .B2(n15838), .A(n15837), .ZN(n20636) );
  INV_X1 U17914 ( .A(n20636), .ZN(n15941) );
  INV_X1 U17915 ( .A(n16756), .ZN(n15840) );
  INV_X1 U17916 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20513) );
  OAI222_X1 U17917 ( .A1(n15941), .A2(n16782), .B1(n16791), .B2(n15840), .C1(
        n16789), .C2(n20513), .ZN(P1_U2899) );
  NAND3_X1 U17918 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n22408), .A3(
        n22476), .ZN(n22443) );
  INV_X1 U17919 ( .A(n22443), .ZN(n15848) );
  OR2_X1 U17920 ( .A1(n22456), .A2(n15842), .ZN(n15843) );
  NOR2_X1 U17921 ( .A1(n22487), .A2(n22443), .ZN(n22739) );
  INV_X1 U17922 ( .A(n22739), .ZN(n15857) );
  NAND2_X1 U17923 ( .A1(n15843), .A2(n15857), .ZN(n15847) );
  INV_X1 U17924 ( .A(n15847), .ZN(n15844) );
  OAI21_X1 U17925 ( .B1(n15846), .B2(n22492), .A(n15844), .ZN(n15845) );
  OAI221_X1 U17926 ( .B1(n22497), .B2(n15848), .C1(n22506), .C2(n15845), .A(
        n22495), .ZN(n22741) );
  NAND2_X1 U17927 ( .A1(n22741), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n15853) );
  NAND2_X1 U17928 ( .A1(n15847), .A2(n22497), .ZN(n15850) );
  NAND2_X1 U17929 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15848), .ZN(n15849) );
  AND2_X1 U17930 ( .A1(n15850), .A2(n15849), .ZN(n22533) );
  OAI22_X1 U17931 ( .A1(n22385), .A2(n15857), .B1(n22485), .B2(n22533), .ZN(
        n15851) );
  AOI21_X1 U17932 ( .B1(n22747), .B2(n22477), .A(n15851), .ZN(n15852) );
  OAI211_X1 U17933 ( .C1(n22386), .C2(n22744), .A(n15853), .B(n15852), .ZN(
        P1_U3105) );
  NAND2_X1 U17934 ( .A1(n22741), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n15856) );
  OAI22_X1 U17935 ( .A1(n22669), .A2(n15857), .B1(n22533), .B2(n22689), .ZN(
        n15854) );
  AOI21_X1 U17936 ( .B1(n22747), .B2(n22686), .A(n15854), .ZN(n15855) );
  OAI211_X1 U17937 ( .C1(n22670), .C2(n22744), .A(n15856), .B(n15855), .ZN(
        P1_U3111) );
  NAND2_X1 U17938 ( .A1(n22741), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n15860) );
  OAI22_X1 U17939 ( .A1(n22580), .A2(n15857), .B1(n22533), .B2(n22600), .ZN(
        n15858) );
  AOI21_X1 U17940 ( .B1(n22747), .B2(n22597), .A(n15858), .ZN(n15859) );
  OAI211_X1 U17941 ( .C1(n22581), .C2(n22744), .A(n15860), .B(n15859), .ZN(
        P1_U3108) );
  OAI21_X1 U17942 ( .B1(n15837), .B2(n15861), .A(n15863), .ZN(n15943) );
  INV_X1 U17943 ( .A(n16753), .ZN(n15864) );
  OAI222_X1 U17944 ( .A1(n15943), .A2(n16782), .B1(n16791), .B2(n15864), .C1(
        n16789), .C2(n13127), .ZN(P1_U2898) );
  NAND2_X1 U17945 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n15865), .ZN(n16444) );
  AOI21_X1 U17946 ( .B1(n22222), .B2(n16444), .A(n22162), .ZN(n15887) );
  AOI21_X1 U17947 ( .B1(n22222), .B2(n15865), .A(P1_REIP_REG_4__SCAN_IN), .ZN(
        n15870) );
  INV_X1 U17948 ( .A(n15866), .ZN(n15867) );
  AOI22_X1 U17949 ( .A1(n15867), .A2(n22216), .B1(n22242), .B2(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n15869) );
  NAND2_X1 U17950 ( .A1(n22190), .A2(n15868), .ZN(n22232) );
  OAI211_X1 U17951 ( .C1(n15887), .C2(n15870), .A(n15869), .B(n22232), .ZN(
        n15873) );
  NOR2_X1 U17952 ( .A1(n22235), .A2(n15871), .ZN(n15872) );
  AOI211_X1 U17953 ( .C1(n22199), .C2(n21990), .A(n15873), .B(n15872), .ZN(
        n15878) );
  INV_X1 U17954 ( .A(n15874), .ZN(n15905) );
  NOR2_X1 U17955 ( .A1(n15875), .A2(n15905), .ZN(n15876) );
  XNOR2_X1 U17956 ( .A(n15876), .B(n17889), .ZN(n17884) );
  NAND2_X1 U17957 ( .A1(n17884), .A2(n22127), .ZN(n15877) );
  OAI211_X1 U17958 ( .C1(n15879), .C2(n22124), .A(n15878), .B(n15877), .ZN(
        P1_U2836) );
  OAI211_X1 U17959 ( .C1(n15880), .C2(n15882), .A(n15881), .B(n17274), .ZN(
        n15886) );
  OAI21_X1 U17960 ( .B1(n15884), .B2(n15883), .A(n16036), .ZN(n19240) );
  INV_X1 U17961 ( .A(n19240), .ZN(n17973) );
  NAND2_X1 U17962 ( .A1(n17973), .A2(n17281), .ZN(n15885) );
  OAI211_X1 U17963 ( .C1(n17281), .C2(n12101), .A(n15886), .B(n15885), .ZN(
        P2_U2876) );
  NOR2_X1 U17964 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n16444), .ZN(n15902) );
  INV_X1 U17965 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n15942) );
  INV_X1 U17966 ( .A(n15887), .ZN(n15888) );
  NAND2_X1 U17967 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n15888), .ZN(n15889) );
  AND2_X1 U17968 ( .A1(n22232), .A2(n15889), .ZN(n15892) );
  INV_X1 U17969 ( .A(n15890), .ZN(n20635) );
  AOI22_X1 U17970 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n22242), .B1(
        n22216), .B2(n20635), .ZN(n15891) );
  OAI211_X1 U17971 ( .C1(n22235), .C2(n15942), .A(n15892), .B(n15891), .ZN(
        n15901) );
  MUX2_X1 U17972 ( .A(n11166), .B(n16430), .S(n15942), .Z(n15896) );
  OR2_X1 U17973 ( .A1(n16440), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15895) );
  NAND2_X1 U17974 ( .A1(n15896), .A2(n15895), .ZN(n15897) );
  NAND2_X1 U17975 ( .A1(n15898), .A2(n15897), .ZN(n15899) );
  NAND2_X1 U17976 ( .A1(n15949), .A2(n15899), .ZN(n16018) );
  NOR2_X1 U17977 ( .A1(n22237), .A2(n16018), .ZN(n15900) );
  AOI211_X1 U17978 ( .C1(n22222), .C2(n15902), .A(n15901), .B(n15900), .ZN(
        n15903) );
  OAI21_X1 U17979 ( .B1(n15941), .B2(n22124), .A(n15903), .ZN(P1_U2835) );
  NAND3_X1 U17980 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22500) );
  AOI21_X1 U17981 ( .B1(n22506), .B2(n22500), .A(n15904), .ZN(n15908) );
  NOR2_X1 U17982 ( .A1(n16674), .A2(n15905), .ZN(n22502) );
  NAND2_X1 U17983 ( .A1(n22502), .A2(n15906), .ZN(n15907) );
  AOI21_X1 U17984 ( .B1(n15907), .B2(n15936), .A(n22506), .ZN(n15909) );
  OAI21_X1 U17985 ( .B1(n15908), .B2(n15909), .A(n22495), .ZN(n15939) );
  INV_X1 U17986 ( .A(n15909), .ZN(n15912) );
  INV_X1 U17987 ( .A(n22500), .ZN(n15910) );
  NAND2_X1 U17988 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15910), .ZN(n15911) );
  AND2_X1 U17989 ( .A1(n15912), .A2(n15911), .ZN(n15935) );
  OAI22_X1 U17990 ( .A1(n22700), .A2(n11301), .B1(n22541), .B2(n15935), .ZN(
        n15915) );
  OAI22_X1 U17991 ( .A1(n22776), .A2(n11303), .B1(n15936), .B2(n22519), .ZN(
        n15914) );
  AOI211_X1 U17992 ( .C1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .C2(n15939), .A(
        n15915), .B(n15914), .ZN(n15916) );
  INV_X1 U17993 ( .A(n15916), .ZN(P1_U3154) );
  INV_X1 U17994 ( .A(n22686), .ZN(n22697) );
  OAI22_X1 U17995 ( .A1(n22700), .A2(n22697), .B1(n22689), .B2(n15935), .ZN(
        n15918) );
  OAI22_X1 U17996 ( .A1(n22776), .A2(n22670), .B1(n15936), .B2(n22669), .ZN(
        n15917) );
  AOI211_X1 U17997 ( .C1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .C2(n15939), .A(
        n15918), .B(n15917), .ZN(n15919) );
  INV_X1 U17998 ( .A(n15919), .ZN(P1_U3159) );
  INV_X1 U17999 ( .A(n22597), .ZN(n22608) );
  OAI22_X1 U18000 ( .A1(n22700), .A2(n22608), .B1(n22600), .B2(n15935), .ZN(
        n15921) );
  OAI22_X1 U18001 ( .A1(n22776), .A2(n22581), .B1(n15936), .B2(n22580), .ZN(
        n15920) );
  AOI211_X1 U18002 ( .C1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .C2(n15939), .A(
        n15921), .B(n15920), .ZN(n15922) );
  INV_X1 U18003 ( .A(n15922), .ZN(P1_U3156) );
  INV_X1 U18004 ( .A(n22568), .ZN(n22579) );
  OAI22_X1 U18005 ( .A1(n22700), .A2(n22579), .B1(n22571), .B2(n15935), .ZN(
        n15924) );
  OAI22_X1 U18006 ( .A1(n22776), .A2(n22565), .B1(n15936), .B2(n22549), .ZN(
        n15923) );
  AOI211_X1 U18007 ( .C1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .C2(n15939), .A(
        n15924), .B(n15923), .ZN(n15925) );
  INV_X1 U18008 ( .A(n15925), .ZN(P1_U3155) );
  INV_X1 U18009 ( .A(n22753), .ZN(n22777) );
  OAI22_X1 U18010 ( .A1(n22700), .A2(n22777), .B1(n22758), .B2(n15935), .ZN(
        n15927) );
  OAI22_X1 U18011 ( .A1(n22776), .A2(n11307), .B1(n15936), .B2(n22699), .ZN(
        n15926) );
  AOI211_X1 U18012 ( .C1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .C2(n15939), .A(
        n15927), .B(n15926), .ZN(n15928) );
  INV_X1 U18013 ( .A(n15928), .ZN(P1_U3160) );
  INV_X1 U18014 ( .A(n22627), .ZN(n22638) );
  OAI22_X1 U18015 ( .A1(n22700), .A2(n22638), .B1(n22630), .B2(n15935), .ZN(
        n15930) );
  OAI22_X1 U18016 ( .A1(n22776), .A2(n11309), .B1(n15936), .B2(n22609), .ZN(
        n15929) );
  AOI211_X1 U18017 ( .C1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .C2(n15939), .A(
        n15930), .B(n15929), .ZN(n15931) );
  INV_X1 U18018 ( .A(n15931), .ZN(P1_U3157) );
  INV_X1 U18019 ( .A(n22657), .ZN(n22668) );
  OAI22_X1 U18020 ( .A1(n22700), .A2(n22668), .B1(n22660), .B2(n15935), .ZN(
        n15933) );
  OAI22_X1 U18021 ( .A1(n22776), .A2(n11305), .B1(n15936), .B2(n22639), .ZN(
        n15932) );
  AOI211_X1 U18022 ( .C1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .C2(n15939), .A(
        n15933), .B(n15932), .ZN(n15934) );
  INV_X1 U18023 ( .A(n15934), .ZN(P1_U3158) );
  INV_X1 U18024 ( .A(n22477), .ZN(n22518) );
  OAI22_X1 U18025 ( .A1(n22700), .A2(n22518), .B1(n22485), .B2(n15935), .ZN(
        n15938) );
  OAI22_X1 U18026 ( .A1(n22776), .A2(n22386), .B1(n15936), .B2(n22385), .ZN(
        n15937) );
  AOI211_X1 U18027 ( .C1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .C2(n15939), .A(
        n15938), .B(n15937), .ZN(n15940) );
  INV_X1 U18028 ( .A(n15940), .ZN(P1_U3153) );
  OAI222_X1 U18029 ( .A1(n16018), .A2(n16724), .B1(n20621), .B2(n15942), .C1(
        n16723), .C2(n15941), .ZN(P1_U2867) );
  INV_X1 U18030 ( .A(n15943), .ZN(n22143) );
  INV_X1 U18031 ( .A(n16723), .ZN(n20618) );
  NAND2_X1 U18032 ( .A1(n16178), .A2(n22006), .ZN(n15945) );
  NAND2_X1 U18033 ( .A1(n16419), .A2(n22138), .ZN(n15944) );
  NAND3_X1 U18034 ( .A1(n15945), .A2(n15944), .A3(n11165), .ZN(n15947) );
  NAND2_X1 U18035 ( .A1(n16400), .A2(n22138), .ZN(n15946) );
  AND2_X1 U18036 ( .A1(n15949), .A2(n15948), .ZN(n15950) );
  OR2_X1 U18037 ( .A1(n15950), .A2(n16177), .ZN(n22139) );
  OAI22_X1 U18038 ( .A1(n22139), .A2(n16724), .B1(n22138), .B2(n20621), .ZN(
        n15951) );
  AOI21_X1 U18039 ( .B1(n22143), .B2(n20618), .A(n15951), .ZN(n15952) );
  INV_X1 U18040 ( .A(n15952), .ZN(P1_U2866) );
  NAND2_X1 U18041 ( .A1(n15954), .A2(n15953), .ZN(n15956) );
  INV_X1 U18042 ( .A(n15883), .ZN(n15955) );
  AND2_X1 U18043 ( .A1(n15956), .A2(n15955), .ZN(n19073) );
  INV_X1 U18044 ( .A(n19073), .ZN(n17724) );
  NOR2_X1 U18045 ( .A1(n17724), .A2(n14651), .ZN(n15959) );
  AOI211_X1 U18046 ( .C1(n15957), .C2(n15777), .A(n17272), .B(n15880), .ZN(
        n15958) );
  AOI211_X1 U18047 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n14651), .A(n15959), .B(
        n15958), .ZN(n15960) );
  INV_X1 U18048 ( .A(n15960), .ZN(P2_U2877) );
  OAI21_X1 U18049 ( .B1(n22720), .B2(n15985), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15967) );
  NAND2_X1 U18050 ( .A1(n22432), .A2(n15965), .ZN(n15966) );
  AOI21_X1 U18051 ( .B1(n15967), .B2(n15966), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n15970) );
  NOR2_X1 U18052 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15968), .ZN(
        n16009) );
  INV_X1 U18053 ( .A(n15973), .ZN(n15969) );
  NOR2_X1 U18054 ( .A1(n15969), .A2(n22489), .ZN(n22459) );
  INV_X1 U18055 ( .A(n22432), .ZN(n15972) );
  NAND2_X1 U18056 ( .A1(n15965), .A2(n22497), .ZN(n15971) );
  OR2_X1 U18057 ( .A1(n15972), .A2(n15971), .ZN(n15975) );
  INV_X1 U18058 ( .A(n22445), .ZN(n22457) );
  NOR2_X1 U18059 ( .A1(n22446), .A2(n22457), .ZN(n22393) );
  NOR2_X1 U18060 ( .A1(n15973), .A2(n22489), .ZN(n22503) );
  NAND2_X1 U18061 ( .A1(n22393), .A2(n22503), .ZN(n15974) );
  NAND2_X1 U18062 ( .A1(n15975), .A2(n15974), .ZN(n15986) );
  AOI22_X1 U18063 ( .A1(n15985), .A2(n22477), .B1(n22507), .B2(n15986), .ZN(
        n15977) );
  NAND2_X1 U18064 ( .A1(n22508), .A2(n16009), .ZN(n15976) );
  OAI211_X1 U18065 ( .C1(n22386), .C2(n16012), .A(n15977), .B(n15976), .ZN(
        n15978) );
  AOI21_X1 U18066 ( .B1(n16005), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n15978), .ZN(n15979) );
  INV_X1 U18067 ( .A(n15979), .ZN(P1_U3065) );
  XNOR2_X1 U18068 ( .A(n11160), .B(n15980), .ZN(n22001) );
  NOR2_X1 U18069 ( .A1(n22093), .A2(n20536), .ZN(n22003) );
  AOI21_X1 U18070 ( .B1(n20694), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n22003), .ZN(n15982) );
  OAI21_X1 U18071 ( .B1(n20703), .B2(n22141), .A(n15982), .ZN(n15983) );
  AOI21_X1 U18072 ( .B1(n22143), .B2(n20689), .A(n15983), .ZN(n15984) );
  OAI21_X1 U18073 ( .B1(n22001), .B2(n20696), .A(n15984), .ZN(P1_U2993) );
  NAND2_X1 U18074 ( .A1(n16005), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n15989) );
  INV_X1 U18075 ( .A(n15985), .ZN(n16007) );
  INV_X1 U18076 ( .A(n15986), .ZN(n16006) );
  OAI22_X1 U18077 ( .A1(n16007), .A2(n11301), .B1(n16006), .B2(n22541), .ZN(
        n15987) );
  AOI21_X1 U18078 ( .B1(n16009), .B2(n22545), .A(n15987), .ZN(n15988) );
  OAI211_X1 U18079 ( .C1(n16012), .C2(n11303), .A(n15989), .B(n15988), .ZN(
        P1_U3066) );
  NAND2_X1 U18080 ( .A1(n16005), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n15992) );
  OAI22_X1 U18081 ( .A1(n16007), .A2(n22697), .B1(n22689), .B2(n16006), .ZN(
        n15990) );
  AOI21_X1 U18082 ( .B1(n22693), .B2(n16009), .A(n15990), .ZN(n15991) );
  OAI211_X1 U18083 ( .C1(n22670), .C2(n16012), .A(n15992), .B(n15991), .ZN(
        P1_U3071) );
  NAND2_X1 U18084 ( .A1(n16005), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n15995) );
  OAI22_X1 U18085 ( .A1(n16007), .A2(n22777), .B1(n16006), .B2(n22758), .ZN(
        n15993) );
  AOI21_X1 U18086 ( .B1(n16009), .B2(n22770), .A(n15993), .ZN(n15994) );
  OAI211_X1 U18087 ( .C1(n16012), .C2(n11307), .A(n15995), .B(n15994), .ZN(
        P1_U3072) );
  NAND2_X1 U18088 ( .A1(n16005), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n15998) );
  OAI22_X1 U18089 ( .A1(n16007), .A2(n22579), .B1(n16006), .B2(n22571), .ZN(
        n15996) );
  AOI21_X1 U18090 ( .B1(n16009), .B2(n22575), .A(n15996), .ZN(n15997) );
  OAI211_X1 U18091 ( .C1(n16012), .C2(n22565), .A(n15998), .B(n15997), .ZN(
        P1_U3067) );
  NAND2_X1 U18092 ( .A1(n16005), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n16001) );
  OAI22_X1 U18093 ( .A1(n16007), .A2(n22668), .B1(n16006), .B2(n22660), .ZN(
        n15999) );
  AOI21_X1 U18094 ( .B1(n16009), .B2(n22664), .A(n15999), .ZN(n16000) );
  OAI211_X1 U18095 ( .C1(n16012), .C2(n11305), .A(n16001), .B(n16000), .ZN(
        P1_U3070) );
  NAND2_X1 U18096 ( .A1(n16005), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n16004) );
  OAI22_X1 U18097 ( .A1(n16007), .A2(n22638), .B1(n16006), .B2(n22630), .ZN(
        n16002) );
  AOI21_X1 U18098 ( .B1(n16009), .B2(n22634), .A(n16002), .ZN(n16003) );
  OAI211_X1 U18099 ( .C1(n16012), .C2(n11309), .A(n16004), .B(n16003), .ZN(
        P1_U3069) );
  NAND2_X1 U18100 ( .A1(n16005), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n16011) );
  OAI22_X1 U18101 ( .A1(n16007), .A2(n22608), .B1(n22600), .B2(n16006), .ZN(
        n16008) );
  AOI21_X1 U18102 ( .B1(n22604), .B2(n16009), .A(n16008), .ZN(n16010) );
  OAI211_X1 U18103 ( .C1(n22581), .C2(n16012), .A(n16011), .B(n16010), .ZN(
        P1_U3068) );
  XOR2_X1 U18104 ( .A(n16014), .B(n11161), .Z(n20637) );
  INV_X1 U18105 ( .A(n20637), .ZN(n16021) );
  NOR2_X1 U18106 ( .A1(n21986), .A2(n13719), .ZN(n21993) );
  NAND2_X1 U18107 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21993), .ZN(
        n16173) );
  NOR2_X1 U18108 ( .A1(n16174), .A2(n16173), .ZN(n16918) );
  NAND3_X1 U18109 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n21993), .ZN(n16921) );
  AOI21_X1 U18110 ( .B1(n21982), .B2(n16921), .A(n21980), .ZN(n16015) );
  OAI21_X1 U18111 ( .B1(n16918), .B2(n22112), .A(n16015), .ZN(n16171) );
  NAND4_X1 U18112 ( .A1(n22021), .A2(n16016), .A3(n21993), .A4(n16923), .ZN(
        n16017) );
  NAND2_X1 U18113 ( .A1(n22102), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n20638) );
  OAI211_X1 U18114 ( .C1(n16018), .C2(n22115), .A(n16017), .B(n20638), .ZN(
        n16019) );
  NOR3_X1 U18115 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16921), .A3(
        n22022), .ZN(n16172) );
  AOI211_X1 U18116 ( .C1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n16171), .A(
        n16019), .B(n16172), .ZN(n16020) );
  OAI21_X1 U18117 ( .B1(n16021), .B2(n22043), .A(n16020), .ZN(P1_U3026) );
  INV_X1 U18118 ( .A(n19924), .ZN(n16022) );
  NAND2_X1 U18119 ( .A1(n19884), .A2(n18034), .ZN(n20004) );
  NOR2_X1 U18120 ( .A1(n19939), .A2(n20004), .ZN(n16023) );
  AOI221_X1 U18121 ( .B1(n20415), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n20414), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n16023), .ZN(n16026) );
  NAND2_X1 U18122 ( .A1(n13947), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16024) );
  NOR3_X2 U18123 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12216), .A3(
        n20004), .ZN(n20412) );
  AOI21_X1 U18124 ( .B1(n16024), .B2(n14346), .A(n20412), .ZN(n16025) );
  AOI22_X1 U18125 ( .A1(n20264), .A2(BUF2_REG_27__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n20191) );
  INV_X1 U18126 ( .A(n20191), .ZN(n20195) );
  AOI22_X1 U18127 ( .A1(n20264), .A2(BUF2_REG_19__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n20198) );
  AOI22_X1 U18128 ( .A1(n20414), .A2(n20195), .B1(n20415), .B2(n20188), .ZN(
        n16033) );
  OAI21_X1 U18129 ( .B1(n16027), .B2(n20412), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16028) );
  OAI21_X1 U18130 ( .B1(n20004), .B2(n19939), .A(n16028), .ZN(n20413) );
  AOI22_X1 U18131 ( .A1(n20413), .A2(n16029), .B1(n20194), .B2(n20412), .ZN(
        n16032) );
  OAI211_X1 U18132 ( .C1(n20419), .C2(n16034), .A(n16033), .B(n16032), .ZN(
        P2_U3067) );
  NAND2_X1 U18133 ( .A1(n16036), .A2(n16035), .ZN(n16037) );
  AND2_X1 U18134 ( .A1(n16230), .A2(n16037), .ZN(n19085) );
  INV_X1 U18135 ( .A(n19085), .ZN(n17710) );
  INV_X1 U18136 ( .A(n15881), .ZN(n16040) );
  OAI211_X1 U18137 ( .C1(n16040), .C2(n14382), .A(n17274), .B(n16039), .ZN(
        n16042) );
  NAND2_X1 U18138 ( .A1(n14651), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n16041) );
  OAI211_X1 U18139 ( .C1(n17710), .C2(n14651), .A(n16042), .B(n16041), .ZN(
        P2_U2875) );
  MUX2_X1 U18140 ( .A(n16430), .B(n11166), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n16044) );
  OR2_X1 U18141 ( .A1(n16440), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16043) );
  XOR2_X1 U18142 ( .A(n16176), .B(n16177), .Z(n22150) );
  INV_X1 U18143 ( .A(n22150), .ZN(n16049) );
  INV_X1 U18144 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n16048) );
  NAND2_X1 U18145 ( .A1(n15863), .A2(n16046), .ZN(n16047) );
  AND2_X1 U18146 ( .A1(n16045), .A2(n16047), .ZN(n22155) );
  INV_X1 U18147 ( .A(n22155), .ZN(n16050) );
  OAI222_X1 U18148 ( .A1(n16049), .A2(n16724), .B1(n20621), .B2(n16048), .C1(
        n16723), .C2(n16050), .ZN(P1_U2865) );
  INV_X1 U18149 ( .A(n16750), .ZN(n16051) );
  OAI222_X1 U18150 ( .A1(n16791), .A2(n16051), .B1(n16789), .B2(n13140), .C1(
        n16782), .C2(n16050), .ZN(P1_U2897) );
  NAND2_X1 U18151 ( .A1(n11173), .A2(n16052), .ZN(n16053) );
  XNOR2_X1 U18152 ( .A(n17912), .B(n16053), .ZN(n16054) );
  NAND2_X1 U18153 ( .A1(n16054), .A2(n19194), .ZN(n16064) );
  AOI22_X1 U18154 ( .A1(n19163), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_EBX_REG_3__SCAN_IN), .B2(n19207), .ZN(n16055) );
  OAI21_X1 U18155 ( .B1(n16056), .B2(n19147), .A(n16055), .ZN(n16062) );
  NAND2_X1 U18156 ( .A1(n16058), .A2(n16057), .ZN(n16060) );
  INV_X1 U18157 ( .A(n16078), .ZN(n16059) );
  NAND2_X1 U18158 ( .A1(n16060), .A2(n16059), .ZN(n20155) );
  OAI22_X1 U18159 ( .A1(n17923), .A2(n19182), .B1(n19222), .B2(n20155), .ZN(
        n16061) );
  AOI211_X1 U18160 ( .C1(n19217), .C2(n19330), .A(n16062), .B(n16061), .ZN(
        n16063) );
  OAI211_X1 U18161 ( .C1(n19876), .C2(n16065), .A(n16064), .B(n16063), .ZN(
        P2_U2852) );
  INV_X1 U18162 ( .A(n16066), .ZN(n16067) );
  NAND2_X1 U18163 ( .A1(n16068), .A2(n16067), .ZN(n16069) );
  OAI21_X1 U18164 ( .B1(n16070), .B2(n16069), .A(n15498), .ZN(n19038) );
  NOR2_X1 U18165 ( .A1(n19860), .A2(n20249), .ZN(n16073) );
  INV_X1 U18166 ( .A(n20249), .ZN(n16072) );
  INV_X1 U18167 ( .A(n16073), .ZN(n16071) );
  OAI21_X1 U18168 ( .B1(n18027), .B2(n16072), .A(n16071), .ZN(n20251) );
  INV_X1 U18169 ( .A(n19020), .ZN(n19226) );
  NOR2_X1 U18170 ( .A1(n18018), .A2(n19226), .ZN(n20252) );
  NOR2_X1 U18171 ( .A1(n20251), .A2(n20252), .ZN(n20250) );
  NOR2_X1 U18172 ( .A1(n16073), .A2(n20250), .ZN(n16075) );
  XNOR2_X1 U18173 ( .A(n16074), .B(n16075), .ZN(n20201) );
  INV_X1 U18174 ( .A(n20201), .ZN(n16077) );
  NAND2_X1 U18175 ( .A1(n16075), .A2(n20199), .ZN(n16076) );
  OAI21_X1 U18176 ( .B1(n16077), .B2(n20200), .A(n16076), .ZN(n20158) );
  XOR2_X1 U18177 ( .A(n20155), .B(n19982), .Z(n20159) );
  NOR2_X1 U18178 ( .A1(n20158), .A2(n20159), .ZN(n20157) );
  INV_X1 U18179 ( .A(n20155), .ZN(n18030) );
  NOR2_X1 U18180 ( .A1(n19982), .A2(n18030), .ZN(n16082) );
  OR2_X1 U18181 ( .A1(n16079), .A2(n16078), .ZN(n16081) );
  NAND2_X1 U18182 ( .A1(n16081), .A2(n16080), .ZN(n19312) );
  OAI21_X1 U18183 ( .B1(n20157), .B2(n16082), .A(n19312), .ZN(n20066) );
  XOR2_X1 U18184 ( .A(n19038), .B(n20066), .Z(n16087) );
  INV_X1 U18185 ( .A(n19312), .ZN(n16083) );
  AOI22_X1 U18186 ( .A1(n20319), .A2(n16083), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n20313), .ZN(n16086) );
  NAND2_X1 U18187 ( .A1(n16084), .A2(n20109), .ZN(n16085) );
  OAI211_X1 U18188 ( .C1(n16087), .C2(n20253), .A(n16086), .B(n16085), .ZN(
        P2_U2915) );
  OR2_X1 U18189 ( .A1(n16090), .A2(n16089), .ZN(n16091) );
  AND2_X1 U18190 ( .A1(n16092), .A2(n16091), .ZN(n19320) );
  NAND2_X1 U18191 ( .A1(n19320), .A2(n17983), .ZN(n16100) );
  INV_X1 U18192 ( .A(n16094), .ZN(n16095) );
  OAI21_X1 U18193 ( .B1(n16096), .B2(n12078), .A(n16095), .ZN(n19039) );
  NOR2_X1 U18194 ( .A1(n19039), .A2(n15057), .ZN(n16098) );
  OAI22_X1 U18195 ( .A1(n12076), .A2(n19325), .B1(n18001), .B2(n19032), .ZN(
        n16097) );
  AOI211_X1 U18196 ( .C1(n18003), .C2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16098), .B(n16097), .ZN(n16099) );
  OAI211_X1 U18197 ( .C1(n19323), .C2(n17996), .A(n16100), .B(n16099), .ZN(
        P2_U3010) );
  AOI21_X1 U18198 ( .B1(n16102), .B2(n16101), .A(n15424), .ZN(n19826) );
  NAND2_X1 U18199 ( .A1(n11173), .A2(n16103), .ZN(n16104) );
  XNOR2_X1 U18200 ( .A(n17951), .B(n16104), .ZN(n16105) );
  AOI22_X1 U18201 ( .A1(n19826), .A2(n19140), .B1(n19194), .B2(n16105), .ZN(
        n16110) );
  AOI22_X1 U18202 ( .A1(n16106), .A2(n19218), .B1(n19208), .B2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16107) );
  OAI211_X1 U18203 ( .C1(n12091), .C2(n19199), .A(n16107), .B(n19325), .ZN(
        n16108) );
  AOI21_X1 U18204 ( .B1(P2_REIP_REG_9__SCAN_IN), .B2(n19163), .A(n16108), .ZN(
        n16109) );
  OAI211_X1 U18205 ( .C1(n17952), .C2(n19165), .A(n16110), .B(n16109), .ZN(
        P2_U2846) );
  NAND2_X1 U18206 ( .A1(n11173), .A2(n16111), .ZN(n16112) );
  XNOR2_X1 U18207 ( .A(n17964), .B(n16112), .ZN(n16113) );
  AOI22_X1 U18208 ( .A1(n19238), .A2(n19140), .B1(n19194), .B2(n16113), .ZN(
        n16119) );
  OAI21_X1 U18209 ( .B1(n12101), .B2(n19199), .A(n19325), .ZN(n16114) );
  AOI21_X1 U18210 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19208), .A(
        n16114), .ZN(n16115) );
  OAI21_X1 U18211 ( .B1(n19210), .B2(n16116), .A(n16115), .ZN(n16117) );
  AOI21_X1 U18212 ( .B1(n17973), .B2(n19217), .A(n16117), .ZN(n16118) );
  OAI211_X1 U18213 ( .C1(n16120), .C2(n19147), .A(n16119), .B(n16118), .ZN(
        P2_U2844) );
  OAI21_X1 U18214 ( .B1(n16122), .B2(n16094), .A(n16121), .ZN(n17926) );
  INV_X1 U18215 ( .A(n16123), .ZN(n16126) );
  INV_X1 U18216 ( .A(n16124), .ZN(n16125) );
  AOI21_X1 U18217 ( .B1(n16126), .B2(n16080), .A(n16125), .ZN(n20063) );
  NAND2_X1 U18218 ( .A1(n11173), .A2(n16127), .ZN(n16128) );
  XNOR2_X1 U18219 ( .A(n17924), .B(n16128), .ZN(n16129) );
  AOI22_X1 U18220 ( .A1(n19140), .A2(n20063), .B1(n19194), .B2(n16129), .ZN(
        n16137) );
  INV_X1 U18221 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n16134) );
  INV_X1 U18222 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n16130) );
  OAI22_X1 U18223 ( .A1(n16131), .A2(n19147), .B1(n19210), .B2(n16130), .ZN(
        n16132) );
  INV_X1 U18224 ( .A(n16132), .ZN(n16133) );
  OAI211_X1 U18225 ( .C1(n16134), .C2(n19199), .A(n16133), .B(n19325), .ZN(
        n16135) );
  AOI21_X1 U18226 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19124), .A(
        n16135), .ZN(n16136) );
  OAI211_X1 U18227 ( .C1(n17926), .C2(n19165), .A(n16137), .B(n16136), .ZN(
        P2_U2850) );
  AOI21_X1 U18228 ( .B1(n16139), .B2(n16138), .A(n15233), .ZN(n19829) );
  NAND2_X1 U18229 ( .A1(n11173), .A2(n16140), .ZN(n16141) );
  XNOR2_X1 U18230 ( .A(n17933), .B(n16141), .ZN(n16142) );
  AOI22_X1 U18231 ( .A1(n19140), .A2(n19829), .B1(n19194), .B2(n16142), .ZN(
        n16149) );
  OAI22_X1 U18232 ( .A1(n16144), .A2(n19147), .B1(n16143), .B2(n19182), .ZN(
        n16145) );
  INV_X1 U18233 ( .A(n16145), .ZN(n16146) );
  OAI211_X1 U18234 ( .C1(n12081), .C2(n19199), .A(n16146), .B(n19325), .ZN(
        n16147) );
  AOI21_X1 U18235 ( .B1(P2_REIP_REG_7__SCAN_IN), .B2(n19163), .A(n16147), .ZN(
        n16148) );
  OAI211_X1 U18236 ( .C1(n19286), .C2(n19165), .A(n16149), .B(n16148), .ZN(
        P2_U2848) );
  OAI21_X1 U18237 ( .B1(n16152), .B2(n16151), .A(n16150), .ZN(n17925) );
  NAND2_X1 U18238 ( .A1(n16154), .A2(n16153), .ZN(n16156) );
  XNOR2_X1 U18239 ( .A(n16156), .B(n16155), .ZN(n17928) );
  AOI21_X1 U18240 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n16157), .A(
        n17756), .ZN(n16158) );
  OR2_X1 U18241 ( .A1(n16160), .A2(n16158), .ZN(n17758) );
  NOR2_X1 U18242 ( .A1(n19339), .A2(n17758), .ZN(n19340) );
  INV_X1 U18243 ( .A(n19340), .ZN(n16159) );
  OAI21_X1 U18244 ( .B1(n16161), .B2(n16160), .A(n16159), .ZN(n19318) );
  NAND2_X1 U18245 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17760), .ZN(
        n19313) );
  AOI221_X1 U18246 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n16166), .C2(n19317), .A(
        n19313), .ZN(n16162) );
  AOI21_X1 U18247 ( .B1(n19282), .B2(P2_REIP_REG_5__SCAN_IN), .A(n16162), .ZN(
        n16163) );
  OAI21_X1 U18248 ( .B1(n19285), .B2(n17926), .A(n16163), .ZN(n16164) );
  AOI21_X1 U18249 ( .B1(n19281), .B2(n20063), .A(n16164), .ZN(n16165) );
  OAI21_X1 U18250 ( .B1(n19318), .B2(n16166), .A(n16165), .ZN(n16167) );
  AOI21_X1 U18251 ( .B1(n17928), .B2(n19271), .A(n16167), .ZN(n16168) );
  OAI21_X1 U18252 ( .B1(n17925), .B2(n19304), .A(n16168), .ZN(P2_U3041) );
  XNOR2_X1 U18253 ( .A(n16170), .B(n16169), .ZN(n16195) );
  NOR2_X1 U18254 ( .A1(n16172), .A2(n16171), .ZN(n22005) );
  AOI22_X1 U18255 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n22005), .B1(
        n17025), .B2(n22016), .ZN(n16205) );
  INV_X1 U18256 ( .A(n16173), .ZN(n16175) );
  NAND2_X1 U18257 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21983) );
  OAI22_X1 U18258 ( .A1(n22112), .A2(n16174), .B1(n21983), .B2(n22022), .ZN(
        n21996) );
  NAND2_X1 U18259 ( .A1(n16175), .A2(n21996), .ZN(n22007) );
  OR2_X1 U18260 ( .A1(n22006), .A2(n22007), .ZN(n16252) );
  NAND2_X1 U18261 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16253) );
  OAI21_X1 U18262 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16253), .ZN(n16187) );
  NAND2_X1 U18263 ( .A1(n16177), .A2(n16176), .ZN(n16184) );
  NAND2_X1 U18264 ( .A1(n16178), .A2(n16179), .ZN(n16180) );
  OAI211_X1 U18265 ( .C1(P1_EBX_REG_8__SCAN_IN), .C2(n16439), .A(n16180), .B(
        n11166), .ZN(n16182) );
  OR2_X1 U18266 ( .A1(n11166), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n16181) );
  NAND2_X1 U18267 ( .A1(n16184), .A2(n16183), .ZN(n16185) );
  AND2_X1 U18268 ( .A1(n16258), .A2(n16185), .ZN(n16196) );
  NOR2_X1 U18269 ( .A1(n22093), .A2(n22164), .ZN(n16191) );
  AOI21_X1 U18270 ( .B1(n16196), .B2(n22106), .A(n16191), .ZN(n16186) );
  OAI21_X1 U18271 ( .B1(n16252), .B2(n16187), .A(n16186), .ZN(n16188) );
  AOI21_X1 U18272 ( .B1(n16205), .B2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n16188), .ZN(n16189) );
  OAI21_X1 U18273 ( .B1(n16195), .B2(n22043), .A(n16189), .ZN(P1_U3023) );
  XOR2_X1 U18274 ( .A(n16190), .B(n16045), .Z(n22168) );
  AOI21_X1 U18275 ( .B1(n20694), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16191), .ZN(n16192) );
  OAI21_X1 U18276 ( .B1(n20703), .B2(n22166), .A(n16192), .ZN(n16193) );
  AOI21_X1 U18277 ( .B1(n22168), .B2(n20689), .A(n16193), .ZN(n16194) );
  OAI21_X1 U18278 ( .B1(n16195), .B2(n20696), .A(n16194), .ZN(P1_U2991) );
  INV_X1 U18279 ( .A(n16196), .ZN(n22163) );
  INV_X1 U18280 ( .A(n22168), .ZN(n16200) );
  OAI222_X1 U18281 ( .A1(n22163), .A2(n16724), .B1(n16723), .B2(n16200), .C1(
        n20621), .C2(n16197), .ZN(P1_U2864) );
  INV_X1 U18282 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20729) );
  NOR2_X1 U18283 ( .A1(n16731), .A2(DATAI_8_), .ZN(n16198) );
  AOI21_X1 U18284 ( .B1(n16731), .B2(n20729), .A(n16198), .ZN(n16746) );
  INV_X1 U18285 ( .A(n16746), .ZN(n22343) );
  OAI222_X1 U18286 ( .A1(n16791), .A2(n22343), .B1(n16782), .B2(n16200), .C1(
        n16199), .C2(n16789), .ZN(P1_U2896) );
  XOR2_X1 U18287 ( .A(n16202), .B(n16201), .Z(n20642) );
  INV_X1 U18288 ( .A(n20642), .ZN(n16207) );
  NAND2_X1 U18289 ( .A1(n22150), .A2(n22106), .ZN(n16203) );
  OR2_X1 U18290 ( .A1(n22093), .A2(n22158), .ZN(n20643) );
  OAI211_X1 U18291 ( .C1(n16252), .C2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n16203), .B(n20643), .ZN(n16204) );
  AOI21_X1 U18292 ( .B1(n16205), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n16204), .ZN(n16206) );
  OAI21_X1 U18293 ( .B1(n16207), .B2(n22043), .A(n16206), .ZN(P1_U3024) );
  AOI21_X1 U18294 ( .B1(n16210), .B2(n16209), .A(n16208), .ZN(n19820) );
  NAND2_X1 U18295 ( .A1(n11173), .A2(n16211), .ZN(n16212) );
  XNOR2_X1 U18296 ( .A(n17526), .B(n16212), .ZN(n16213) );
  AOI22_X1 U18297 ( .A1(n19820), .A2(n19140), .B1(n19194), .B2(n16213), .ZN(
        n16221) );
  NAND2_X1 U18298 ( .A1(n16214), .A2(n16215), .ZN(n16216) );
  NAND2_X1 U18299 ( .A1(n17276), .A2(n16216), .ZN(n17678) );
  INV_X1 U18300 ( .A(n17678), .ZN(n16246) );
  INV_X1 U18301 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n17522) );
  OAI21_X1 U18302 ( .B1(n12119), .B2(n19199), .A(n19325), .ZN(n16217) );
  AOI21_X1 U18303 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19124), .A(
        n16217), .ZN(n16218) );
  OAI21_X1 U18304 ( .B1(n19210), .B2(n17522), .A(n16218), .ZN(n16219) );
  AOI21_X1 U18305 ( .B1(n16246), .B2(n19217), .A(n16219), .ZN(n16220) );
  OAI211_X1 U18306 ( .C1(n16222), .C2(n19147), .A(n16221), .B(n16220), .ZN(
        P2_U2840) );
  AND2_X1 U18307 ( .A1(n16224), .A2(n16223), .ZN(n16226) );
  OR2_X1 U18308 ( .A1(n16226), .A2(n16225), .ZN(n22179) );
  INV_X1 U18309 ( .A(n16791), .ZN(n16295) );
  INV_X1 U18310 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20731) );
  NOR2_X1 U18311 ( .A1(n16731), .A2(DATAI_9_), .ZN(n16227) );
  AOI21_X1 U18312 ( .B1(n16731), .B2(n20731), .A(n16227), .ZN(n22347) );
  AOI22_X1 U18313 ( .A1(n16295), .A2(n22347), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n16775), .ZN(n16228) );
  OAI21_X1 U18314 ( .B1(n22179), .B2(n16782), .A(n16228), .ZN(P1_U2895) );
  AND2_X1 U18315 ( .A1(n16230), .A2(n16229), .ZN(n16231) );
  NOR2_X1 U18316 ( .A1(n17281), .A2(n12110), .ZN(n16235) );
  AOI211_X1 U18317 ( .C1(n16233), .C2(n16039), .A(n17272), .B(n16232), .ZN(
        n16234) );
  AOI211_X1 U18318 ( .C1(n11273), .C2(n17281), .A(n16235), .B(n16234), .ZN(
        n16236) );
  INV_X1 U18319 ( .A(n16236), .ZN(P2_U2874) );
  OAI21_X1 U18320 ( .B1(n16238), .B2(n16237), .A(n16214), .ZN(n17989) );
  INV_X1 U18321 ( .A(n16239), .ZN(n16240) );
  OAI211_X1 U18322 ( .C1(n16232), .C2(n16241), .A(n16240), .B(n17274), .ZN(
        n16243) );
  NAND2_X1 U18323 ( .A1(n14651), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n16242) );
  OAI211_X1 U18324 ( .C1(n17989), .C2(n14651), .A(n16243), .B(n16242), .ZN(
        P2_U2873) );
  OAI211_X1 U18325 ( .C1(n16239), .C2(n16245), .A(n16244), .B(n17274), .ZN(
        n16248) );
  NAND2_X1 U18326 ( .A1(n16246), .A2(n17281), .ZN(n16247) );
  OAI211_X1 U18327 ( .C1(n17281), .C2(n12119), .A(n16248), .B(n16247), .ZN(
        P2_U2872) );
  OAI21_X1 U18328 ( .B1(n16250), .B2(n16249), .A(n20647), .ZN(n16268) );
  NOR2_X1 U18329 ( .A1(n22006), .A2(n16253), .ZN(n16251) );
  OAI21_X1 U18330 ( .B1(n17025), .B2(n16251), .A(n22005), .ZN(n22009) );
  NOR3_X1 U18331 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16253), .A3(
        n16252), .ZN(n22010) );
  AOI21_X1 U18332 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n22009), .A(
        n22010), .ZN(n16261) );
  OR2_X1 U18333 ( .A1(n16430), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n16256) );
  NAND2_X1 U18334 ( .A1(n11166), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16254) );
  OAI211_X1 U18335 ( .C1(P1_EBX_REG_9__SCAN_IN), .C2(n16439), .A(n16178), .B(
        n16254), .ZN(n16255) );
  NAND2_X1 U18336 ( .A1(n16256), .A2(n16255), .ZN(n16257) );
  AND2_X1 U18337 ( .A1(n16258), .A2(n16257), .ZN(n16259) );
  NOR2_X1 U18338 ( .A1(n20609), .A2(n16259), .ZN(n22173) );
  INV_X1 U18339 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n22183) );
  NOR2_X1 U18340 ( .A1(n22093), .A2(n22183), .ZN(n16262) );
  AOI21_X1 U18341 ( .B1(n22173), .B2(n22106), .A(n16262), .ZN(n16260) );
  OAI211_X1 U18342 ( .C1(n16268), .C2(n22043), .A(n16261), .B(n16260), .ZN(
        P1_U3022) );
  AOI21_X1 U18343 ( .B1(n20694), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16262), .ZN(n16265) );
  NAND2_X1 U18344 ( .A1(n20676), .A2(n16263), .ZN(n16264) );
  OAI211_X1 U18345 ( .C1(n22179), .C2(n20697), .A(n16265), .B(n16264), .ZN(
        n16266) );
  INV_X1 U18346 ( .A(n16266), .ZN(n16267) );
  OAI21_X1 U18347 ( .B1(n16268), .B2(n20696), .A(n16267), .ZN(P1_U2990) );
  MUX2_X1 U18348 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n16731), .Z(
        n16740) );
  INV_X1 U18349 ( .A(n16740), .ZN(n22353) );
  XOR2_X1 U18350 ( .A(n16269), .B(n16225), .Z(n22192) );
  INV_X1 U18351 ( .A(n22192), .ZN(n16270) );
  OAI222_X1 U18352 ( .A1(n16789), .A2(n16271), .B1(n16791), .B2(n22353), .C1(
        n16782), .C2(n16270), .ZN(P1_U2894) );
  NAND2_X1 U18353 ( .A1(n16273), .A2(n16274), .ZN(n16275) );
  NAND2_X1 U18354 ( .A1(n16272), .A2(n16275), .ZN(n16292) );
  XNOR2_X1 U18355 ( .A(n16292), .B(n13203), .ZN(n22206) );
  INV_X1 U18356 ( .A(n22206), .ZN(n20661) );
  NOR2_X1 U18357 ( .A1(n16277), .A2(BUF1_REG_11__SCAN_IN), .ZN(n16276) );
  AOI21_X1 U18358 ( .B1(n16278), .B2(n16277), .A(n16276), .ZN(n16737) );
  INV_X1 U18359 ( .A(n16737), .ZN(n22357) );
  OAI222_X1 U18360 ( .A1(n20661), .A2(n16782), .B1(n16789), .B2(n16279), .C1(
        n16791), .C2(n22357), .ZN(P1_U2893) );
  MUX2_X1 U18361 ( .A(n16430), .B(n11166), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n16281) );
  OR2_X1 U18362 ( .A1(n16440), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16280) );
  NAND2_X1 U18363 ( .A1(n16281), .A2(n16280), .ZN(n16286) );
  NAND2_X1 U18364 ( .A1(n11166), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16282) );
  NAND2_X1 U18365 ( .A1(n16178), .A2(n16282), .ZN(n16283) );
  OAI21_X1 U18366 ( .B1(P1_EBX_REG_10__SCAN_IN), .B2(n16439), .A(n16283), .ZN(
        n16285) );
  OR2_X1 U18367 ( .A1(n11165), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n16284) );
  INV_X1 U18368 ( .A(n20608), .ZN(n16288) );
  INV_X1 U18369 ( .A(n16286), .ZN(n16287) );
  AOI21_X1 U18370 ( .B1(n20609), .B2(n16288), .A(n16287), .ZN(n16289) );
  OR2_X1 U18371 ( .A1(n16722), .A2(n16289), .ZN(n22030) );
  OAI222_X1 U18372 ( .A1(n20661), .A2(n16723), .B1(n16724), .B2(n22030), .C1(
        n20621), .C2(n16290), .ZN(P1_U2861) );
  OAI21_X1 U18373 ( .B1(n16292), .B2(n16291), .A(n16272), .ZN(n16294) );
  NAND2_X1 U18374 ( .A1(n16294), .A2(n16293), .ZN(n16662) );
  OAI21_X1 U18375 ( .B1(n16294), .B2(n16293), .A(n16662), .ZN(n20665) );
  MUX2_X1 U18376 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n16731), .Z(
        n22361) );
  AOI22_X1 U18377 ( .A1(n16295), .A2(n22361), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n16775), .ZN(n16296) );
  OAI21_X1 U18378 ( .B1(n20665), .B2(n16782), .A(n16296), .ZN(P1_U2892) );
  INV_X1 U18379 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16297) );
  OAI21_X1 U18380 ( .B1(n16298), .B2(n21492), .A(n16297), .ZN(n17813) );
  NAND2_X1 U18381 ( .A1(n16299), .A2(n17813), .ZN(n21923) );
  NAND2_X1 U18382 ( .A1(n21481), .A2(n21937), .ZN(n21507) );
  NOR2_X1 U18383 ( .A1(n21923), .A2(n21507), .ZN(n16305) );
  NAND2_X1 U18384 ( .A1(n21901), .A2(n16300), .ZN(n18109) );
  INV_X1 U18385 ( .A(n18109), .ZN(n16304) );
  NAND2_X1 U18386 ( .A1(n20851), .A2(n16301), .ZN(n17833) );
  INV_X1 U18387 ( .A(n22332), .ZN(n22285) );
  AOI211_X1 U18388 ( .C1(n21282), .C2(n17833), .A(n22285), .B(n21897), .ZN(
        n16303) );
  NOR2_X1 U18389 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21937), .ZN(n19385) );
  INV_X1 U18390 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21951) );
  NAND2_X1 U18391 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18497) );
  NOR2_X1 U18392 ( .A1(n20846), .A2(n18497), .ZN(n17830) );
  INV_X1 U18393 ( .A(n17830), .ZN(n21935) );
  NOR2_X1 U18394 ( .A1(n21951), .A2(n21935), .ZN(n17815) );
  AOI211_X2 U18395 ( .C1(n21926), .C2(n21912), .A(n19385), .B(n17815), .ZN(
        n21508) );
  MUX2_X1 U18396 ( .A(n16305), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n21508), .Z(P3_U3284) );
  OAI21_X1 U18397 ( .B1(n18003), .B2(n16306), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16315) );
  AND2_X1 U18398 ( .A1(n16307), .A2(n19224), .ZN(n16308) );
  NOR2_X1 U18399 ( .A1(n16309), .A2(n16308), .ZN(n19228) );
  OR2_X1 U18400 ( .A1(n19019), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16310) );
  NAND2_X1 U18401 ( .A1(n16311), .A2(n16310), .ZN(n19233) );
  INV_X1 U18402 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18037) );
  NOR2_X1 U18403 ( .A1(n19325), .A2(n18037), .ZN(n19229) );
  NOR2_X1 U18404 ( .A1(n19229), .A2(n11753), .ZN(n16312) );
  OAI21_X1 U18405 ( .B1(n18008), .B2(n19233), .A(n16312), .ZN(n16313) );
  AOI21_X1 U18406 ( .B1(n18010), .B2(n19228), .A(n16313), .ZN(n16314) );
  NAND2_X1 U18407 ( .A1(n16315), .A2(n16314), .ZN(P2_U3014) );
  NAND2_X1 U18408 ( .A1(n18002), .A2(n16316), .ZN(n16318) );
  OAI211_X1 U18409 ( .C1(n16319), .C2(n17987), .A(n16318), .B(n16317), .ZN(
        n16322) );
  NOR2_X1 U18410 ( .A1(n16320), .A2(n17996), .ZN(n16321) );
  OAI21_X1 U18411 ( .B1(n16325), .B2(n18008), .A(n16324), .ZN(P2_U2984) );
  INV_X1 U18412 ( .A(n16326), .ZN(n16328) );
  XNOR2_X1 U18413 ( .A(n11667), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16794) );
  OAI211_X1 U18414 ( .C1(n16328), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16794), .B(n16327), .ZN(n16329) );
  XNOR2_X1 U18415 ( .A(n16329), .B(n16933), .ZN(n16954) );
  AOI21_X1 U18416 ( .B1(n16331), .B2(n16463), .A(n16330), .ZN(n16452) );
  NAND2_X1 U18417 ( .A1(n20676), .A2(n16457), .ZN(n16332) );
  NAND2_X1 U18418 ( .A1(n22102), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16948) );
  OAI211_X1 U18419 ( .C1(n16333), .C2(n20646), .A(n16332), .B(n16948), .ZN(
        n16334) );
  AOI21_X1 U18420 ( .B1(n16452), .B2(n20689), .A(n16334), .ZN(n16335) );
  OAI21_X1 U18421 ( .B1(n16954), .B2(n20696), .A(n16335), .ZN(P1_U2969) );
  XOR2_X1 U18422 ( .A(n15498), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n16338)
         );
  NOR2_X1 U18423 ( .A1(n17926), .A2(n14651), .ZN(n16336) );
  AOI21_X1 U18424 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n14651), .A(n16336), .ZN(
        n16337) );
  OAI21_X1 U18425 ( .B1(n16338), .B2(n17272), .A(n16337), .ZN(P2_U2882) );
  MUX2_X1 U18426 ( .A(n11860), .B(n19039), .S(n17281), .Z(n16339) );
  OAI21_X1 U18427 ( .B1(n19038), .B2(n17272), .A(n16339), .ZN(P2_U2883) );
  NOR2_X1 U18428 ( .A1(n18001), .A2(n17095), .ZN(n16340) );
  AOI211_X1 U18429 ( .C1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n18003), .A(
        n16341), .B(n16340), .ZN(n16342) );
  OAI21_X1 U18430 ( .B1(n17206), .B2(n15057), .A(n16342), .ZN(n16343) );
  AOI21_X1 U18431 ( .B1(n16344), .B2(n18010), .A(n16343), .ZN(n16345) );
  OAI21_X1 U18432 ( .B1(n16346), .B2(n18008), .A(n16345), .ZN(P2_U2986) );
  NAND2_X1 U18433 ( .A1(n16347), .A2(n22268), .ZN(n16348) );
  AOI211_X1 U18434 ( .C1(n22492), .C2(n16348), .A(n22506), .B(n16350), .ZN(
        n16349) );
  AOI21_X1 U18435 ( .B1(n16350), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16349), .ZN(n16351) );
  OAI21_X1 U18436 ( .B1(n15965), .B2(n16352), .A(n16351), .ZN(P1_U3477) );
  INV_X1 U18437 ( .A(n20316), .ZN(n17386) );
  INV_X1 U18438 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n16358) );
  AOI22_X1 U18439 ( .A1(n20315), .A2(n16356), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n20313), .ZN(n16357) );
  OAI21_X1 U18440 ( .B1(n17386), .B2(n16358), .A(n16357), .ZN(n16361) );
  NOR2_X1 U18441 ( .A1(n16359), .A2(n20154), .ZN(n16360) );
  AOI211_X1 U18442 ( .C1(BUF1_REG_30__SCAN_IN), .C2(n20317), .A(n16361), .B(
        n16360), .ZN(n16362) );
  OAI21_X1 U18443 ( .B1(n16363), .B2(n20253), .A(n16362), .ZN(P2_U2889) );
  OAI21_X1 U18444 ( .B1(n16364), .B2(n15121), .A(n16371), .ZN(n16368) );
  NAND2_X1 U18445 ( .A1(n16366), .A2(n16365), .ZN(n16367) );
  OAI211_X1 U18446 ( .C1(n16370), .C2(n16369), .A(n16368), .B(n16367), .ZN(
        n17880) );
  INV_X1 U18447 ( .A(n15121), .ZN(n16373) );
  AND2_X1 U18448 ( .A1(n16371), .A2(n12915), .ZN(n16372) );
  AOI21_X1 U18449 ( .B1(n16374), .B2(n16373), .A(n16372), .ZN(n20705) );
  OR3_X1 U18450 ( .A1(n16419), .A2(n16376), .A3(n16375), .ZN(n16377) );
  NAND2_X1 U18451 ( .A1(n16377), .A2(n22248), .ZN(n21958) );
  AND2_X1 U18452 ( .A1(n20705), .A2(n21958), .ZN(n17883) );
  NOR2_X1 U18453 ( .A1(n17883), .A2(n22265), .ZN(n22247) );
  MUX2_X1 U18454 ( .A(P1_MORE_REG_SCAN_IN), .B(n17880), .S(n22247), .Z(
        P1_U3484) );
  INV_X1 U18455 ( .A(n16378), .ZN(n16451) );
  NAND2_X1 U18456 ( .A1(n16178), .A2(n22025), .ZN(n16379) );
  OAI211_X1 U18457 ( .C1(P1_EBX_REG_12__SCAN_IN), .C2(n16439), .A(n16379), .B(
        n11165), .ZN(n16381) );
  OR2_X1 U18458 ( .A1(n11165), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n16380) );
  NAND2_X1 U18459 ( .A1(n16381), .A2(n16380), .ZN(n16721) );
  MUX2_X1 U18460 ( .A(n16430), .B(n11166), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n16383) );
  OR2_X1 U18461 ( .A1(n16440), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16382) );
  NAND2_X1 U18462 ( .A1(n16383), .A2(n16382), .ZN(n16668) );
  MUX2_X1 U18463 ( .A(n16430), .B(n11165), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n16385) );
  OR2_X1 U18464 ( .A1(n16440), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16384) );
  AND2_X1 U18465 ( .A1(n16385), .A2(n16384), .ZN(n16638) );
  NAND2_X1 U18466 ( .A1(n16178), .A2(n16386), .ZN(n16388) );
  OR2_X1 U18467 ( .A1(n16439), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n16387) );
  NAND3_X1 U18468 ( .A1(n16388), .A2(n11165), .A3(n16387), .ZN(n16390) );
  OR2_X1 U18469 ( .A1(n11165), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n16389) );
  NAND2_X1 U18470 ( .A1(n16390), .A2(n16389), .ZN(n16650) );
  NAND2_X1 U18471 ( .A1(n16638), .A2(n16650), .ZN(n16391) );
  INV_X1 U18472 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n20682) );
  NAND2_X1 U18473 ( .A1(n16178), .A2(n20682), .ZN(n16392) );
  OAI211_X1 U18474 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n16439), .A(n16392), .B(
        n11166), .ZN(n16394) );
  OR2_X1 U18475 ( .A1(n11166), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n16393) );
  OR2_X1 U18476 ( .A1(n16430), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n16397) );
  NAND2_X1 U18477 ( .A1(n11165), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16395) );
  OAI211_X1 U18478 ( .C1(P1_EBX_REG_17__SCAN_IN), .C2(n16439), .A(n16178), .B(
        n16395), .ZN(n16396) );
  AND2_X1 U18479 ( .A1(n16397), .A2(n16396), .ZN(n16623) );
  NAND2_X1 U18480 ( .A1(n16178), .A2(n22048), .ZN(n16399) );
  INV_X1 U18481 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n16707) );
  NAND2_X1 U18482 ( .A1(n16419), .A2(n16707), .ZN(n16398) );
  NAND3_X1 U18483 ( .A1(n16399), .A2(n16398), .A3(n11165), .ZN(n16402) );
  NAND2_X1 U18484 ( .A1(n16400), .A2(n16707), .ZN(n16401) );
  MUX2_X1 U18485 ( .A(n16430), .B(n11165), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n16404) );
  OR2_X1 U18486 ( .A1(n16440), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16403) );
  NAND2_X1 U18487 ( .A1(n16404), .A2(n16403), .ZN(n16596) );
  NAND2_X1 U18488 ( .A1(n16178), .A2(n16857), .ZN(n16406) );
  INV_X1 U18489 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n16586) );
  NAND2_X1 U18490 ( .A1(n16419), .A2(n16586), .ZN(n16405) );
  NAND3_X1 U18491 ( .A1(n16406), .A2(n16405), .A3(n11166), .ZN(n16408) );
  NAND2_X1 U18492 ( .A1(n16400), .A2(n16586), .ZN(n16407) );
  NAND2_X1 U18493 ( .A1(n16408), .A2(n16407), .ZN(n16582) );
  OR2_X1 U18494 ( .A1(n16430), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n16411) );
  NAND2_X1 U18495 ( .A1(n11166), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16409) );
  OAI211_X1 U18496 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n16439), .A(n16178), .B(
        n16409), .ZN(n16410) );
  NAND2_X1 U18497 ( .A1(n16411), .A2(n16410), .ZN(n16563) );
  INV_X1 U18498 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16992) );
  NAND2_X1 U18499 ( .A1(n16178), .A2(n16992), .ZN(n16412) );
  OAI211_X1 U18500 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n16439), .A(n16412), .B(
        n11166), .ZN(n16415) );
  INV_X1 U18501 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n16413) );
  NAND2_X1 U18502 ( .A1(n16400), .A2(n16413), .ZN(n16414) );
  MUX2_X1 U18503 ( .A(n16430), .B(n11166), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n16417) );
  OR2_X1 U18504 ( .A1(n16440), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16416) );
  AND2_X1 U18505 ( .A1(n16417), .A2(n16416), .ZN(n16538) );
  NAND2_X1 U18506 ( .A1(n11165), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16418) );
  NAND2_X1 U18507 ( .A1(n16178), .A2(n16418), .ZN(n16421) );
  INV_X1 U18508 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n16698) );
  NAND2_X1 U18509 ( .A1(n16419), .A2(n16698), .ZN(n16420) );
  NAND2_X1 U18510 ( .A1(n16421), .A2(n16420), .ZN(n16423) );
  NAND2_X1 U18511 ( .A1(n16400), .A2(n16698), .ZN(n16422) );
  NAND2_X1 U18512 ( .A1(n16423), .A2(n16422), .ZN(n16527) );
  OR2_X1 U18513 ( .A1(n16430), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n16426) );
  NAND2_X1 U18514 ( .A1(n11165), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16424) );
  OAI211_X1 U18515 ( .C1(n16439), .C2(P1_EBX_REG_25__SCAN_IN), .A(n16178), .B(
        n16424), .ZN(n16425) );
  NAND2_X1 U18516 ( .A1(n16426), .A2(n16425), .ZN(n16516) );
  INV_X1 U18517 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16971) );
  NAND2_X1 U18518 ( .A1(n16178), .A2(n16971), .ZN(n16427) );
  OAI211_X1 U18519 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n16439), .A(n16427), .B(
        n11165), .ZN(n16429) );
  INV_X1 U18520 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n16695) );
  NAND2_X1 U18521 ( .A1(n16400), .A2(n16695), .ZN(n16428) );
  AND2_X1 U18522 ( .A1(n16429), .A2(n16428), .ZN(n16501) );
  MUX2_X1 U18523 ( .A(n16430), .B(n11165), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n16432) );
  OR2_X1 U18524 ( .A1(n16440), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16431) );
  NAND2_X1 U18525 ( .A1(n16432), .A2(n16431), .ZN(n16489) );
  NOR2_X1 U18526 ( .A1(n15768), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16434) );
  OAI21_X1 U18527 ( .B1(n16439), .B2(P1_EBX_REG_28__SCAN_IN), .A(n11166), .ZN(
        n16433) );
  OAI22_X1 U18528 ( .A1(n16434), .A2(n16433), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n11165), .ZN(n16478) );
  OAI22_X1 U18529 ( .A1(n16440), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n16439), .ZN(n16453) );
  MUX2_X1 U18530 ( .A(P1_EBX_REG_29__SCAN_IN), .B(n16453), .S(n11166), .Z(
        n16467) );
  AND2_X1 U18531 ( .A1(n16439), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16436) );
  AOI21_X1 U18532 ( .B1(n16440), .B2(P1_EBX_REG_30__SCAN_IN), .A(n16436), .ZN(
        n16454) );
  AOI22_X1 U18533 ( .A1(n16440), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16439), .ZN(n16441) );
  INV_X1 U18534 ( .A(n16441), .ZN(n16442) );
  INV_X1 U18535 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20653) );
  NOR2_X1 U18536 ( .A1(n20535), .A2(n16444), .ZN(n22137) );
  NAND2_X1 U18537 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n22137), .ZN(n22147) );
  NOR2_X1 U18538 ( .A1(n22158), .A2(n22147), .ZN(n22159) );
  NAND2_X1 U18539 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n22159), .ZN(n22172) );
  NOR2_X1 U18540 ( .A1(n22183), .A2(n22172), .ZN(n22186) );
  NAND2_X1 U18541 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n22186), .ZN(n22185) );
  NOR2_X1 U18542 ( .A1(n20653), .A2(n22185), .ZN(n22221) );
  NAND2_X1 U18543 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n22221), .ZN(n16664) );
  NOR2_X1 U18544 ( .A1(n21966), .A2(n16664), .ZN(n16663) );
  INV_X1 U18545 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20554) );
  NOR4_X1 U18546 ( .A1(n20551), .A2(n20554), .A3(n22227), .A4(n20549), .ZN(
        n16445) );
  NAND2_X1 U18547 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n16445), .ZN(n16603) );
  NOR2_X1 U18548 ( .A1(n22067), .A2(n16603), .ZN(n16577) );
  NAND3_X1 U18549 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n16663), .A3(n16577), 
        .ZN(n16569) );
  NAND2_X1 U18550 ( .A1(n16535), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n16496) );
  INV_X1 U18551 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20573) );
  INV_X1 U18552 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20570) );
  NOR2_X1 U18553 ( .A1(n16446), .A2(n22228), .ZN(n16456) );
  MUX2_X1 U18554 ( .A(n16446), .B(n16456), .S(P1_REIP_REG_31__SCAN_IN), .Z(
        n16449) );
  INV_X1 U18555 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16447) );
  OAI22_X1 U18556 ( .A1(n22235), .A2(n16686), .B1(n16447), .B2(n22204), .ZN(
        n16448) );
  AOI211_X1 U18557 ( .C1(n16940), .C2(n22199), .A(n16449), .B(n16448), .ZN(
        n16450) );
  OAI21_X1 U18558 ( .B1(n16451), .B2(n22238), .A(n16450), .ZN(P1_U2809) );
  INV_X1 U18559 ( .A(n16452), .ZN(n16730) );
  OAI22_X1 U18560 ( .A1(n16466), .A2(n11165), .B1(n16453), .B2(n16477), .ZN(
        n16455) );
  XNOR2_X1 U18561 ( .A(n16455), .B(n16454), .ZN(n16952) );
  INV_X1 U18562 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n16689) );
  OAI21_X1 U18563 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n11321), .A(n16456), 
        .ZN(n16459) );
  AOI22_X1 U18564 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n22242), .B1(
        n22216), .B2(n16457), .ZN(n16458) );
  OAI211_X1 U18565 ( .C1(n22235), .C2(n16689), .A(n16459), .B(n16458), .ZN(
        n16460) );
  AOI21_X1 U18566 ( .B1(n16952), .B2(n22199), .A(n16460), .ZN(n16461) );
  OAI21_X1 U18567 ( .B1(n16730), .B2(n22238), .A(n16461), .ZN(P1_U2810) );
  INV_X1 U18568 ( .A(n16463), .ZN(n16464) );
  INV_X1 U18569 ( .A(n16795), .ZN(n16734) );
  OAI22_X1 U18570 ( .A1(n16492), .A2(n20570), .B1(n22228), .B2(n20573), .ZN(
        n16471) );
  AOI21_X1 U18571 ( .B1(n16467), .B2(n16477), .A(n16466), .ZN(n16958) );
  NAND2_X1 U18572 ( .A1(n16958), .A2(n22199), .ZN(n16469) );
  AOI22_X1 U18573 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n22242), .B1(
        n22216), .B2(n16798), .ZN(n16468) );
  OAI211_X1 U18574 ( .C1(n22235), .C2(n16691), .A(n16469), .B(n16468), .ZN(
        n16470) );
  AOI21_X1 U18575 ( .B1(n16472), .B2(n16471), .A(n16470), .ZN(n16473) );
  OAI21_X1 U18576 ( .B1(n16734), .B2(n22238), .A(n16473), .ZN(P1_U2811) );
  OAI22_X1 U18577 ( .A1(n16476), .A2(n22204), .B1(n22244), .B2(n16801), .ZN(
        n16480) );
  OAI21_X1 U18578 ( .B1(n16488), .B2(n16478), .A(n16477), .ZN(n16970) );
  NOR2_X1 U18579 ( .A1(n16970), .A2(n22237), .ZN(n16479) );
  AOI211_X1 U18580 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n22201), .A(n16480), .B(
        n16479), .ZN(n16483) );
  NAND2_X1 U18581 ( .A1(n16492), .A2(n22161), .ZN(n16481) );
  MUX2_X1 U18582 ( .A(n16492), .B(n16481), .S(P1_REIP_REG_28__SCAN_IN), .Z(
        n16482) );
  OAI211_X1 U18583 ( .C1(n16810), .C2(n22238), .A(n16483), .B(n16482), .ZN(
        P1_U2812) );
  INV_X1 U18584 ( .A(n16474), .ZN(n16487) );
  NAND2_X2 U18585 ( .A1(n16487), .A2(n16486), .ZN(n16814) );
  AOI21_X1 U18586 ( .B1(n16489), .B2(n16503), .A(n16488), .ZN(n22082) );
  INV_X1 U18587 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n16694) );
  AOI22_X1 U18588 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n22242), .B1(
        n22216), .B2(n16817), .ZN(n16490) );
  OAI21_X1 U18589 ( .B1(n22235), .B2(n16694), .A(n16490), .ZN(n16491) );
  AOI21_X1 U18590 ( .B1(n22082), .B2(n22199), .A(n16491), .ZN(n16495) );
  NOR2_X1 U18591 ( .A1(n22228), .A2(n22085), .ZN(n16493) );
  OAI21_X1 U18592 ( .B1(n16509), .B2(n16493), .A(n16492), .ZN(n16494) );
  OAI211_X1 U18593 ( .C1(n16814), .C2(n22238), .A(n16495), .B(n16494), .ZN(
        P1_U2813) );
  INV_X1 U18594 ( .A(n16496), .ZN(n16523) );
  AOI21_X1 U18595 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n22161), .A(n16523), 
        .ZN(n16508) );
  BUF_X1 U18596 ( .A(n16497), .Z(n16498) );
  AOI21_X1 U18597 ( .B1(n16499), .B2(n16498), .A(n16484), .ZN(n16825) );
  NAND2_X1 U18598 ( .A1(n16825), .A2(n22215), .ZN(n16507) );
  OAI22_X1 U18599 ( .A1(n16500), .A2(n22204), .B1(n22244), .B2(n16823), .ZN(
        n16505) );
  NAND2_X1 U18600 ( .A1(n16514), .A2(n16501), .ZN(n16502) );
  NAND2_X1 U18601 ( .A1(n16503), .A2(n16502), .ZN(n16976) );
  NOR2_X1 U18602 ( .A1(n16976), .A2(n22237), .ZN(n16504) );
  AOI211_X1 U18603 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n22201), .A(n16505), .B(
        n16504), .ZN(n16506) );
  OAI211_X1 U18604 ( .C1(n16509), .C2(n16508), .A(n16507), .B(n16506), .ZN(
        P1_U2814) );
  AOI21_X1 U18605 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n22161), .A(n16535), 
        .ZN(n16522) );
  INV_X1 U18606 ( .A(n16498), .ZN(n16512) );
  AOI21_X1 U18607 ( .B1(n16513), .B2(n16511), .A(n16512), .ZN(n16696) );
  NAND2_X1 U18608 ( .A1(n16696), .A2(n22215), .ZN(n16521) );
  INV_X1 U18609 ( .A(n16514), .ZN(n16515) );
  AOI21_X1 U18610 ( .B1(n16516), .B2(n16529), .A(n16515), .ZN(n22099) );
  AOI22_X1 U18611 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n22242), .B1(
        n22216), .B2(n16835), .ZN(n16517) );
  OAI21_X1 U18612 ( .B1(n22235), .B2(n16518), .A(n16517), .ZN(n16519) );
  AOI21_X1 U18613 ( .B1(n22099), .B2(n22199), .A(n16519), .ZN(n16520) );
  OAI211_X1 U18614 ( .C1(n16523), .C2(n16522), .A(n16521), .B(n16520), .ZN(
        P1_U2815) );
  AOI21_X1 U18615 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n22161), .A(n16542), 
        .ZN(n16534) );
  OAI21_X1 U18616 ( .B1(n16524), .B2(n16525), .A(n16511), .ZN(n16749) );
  INV_X1 U18617 ( .A(n16749), .ZN(n16847) );
  NAND2_X1 U18618 ( .A1(n16847), .A2(n22215), .ZN(n16533) );
  OAI22_X1 U18619 ( .A1(n16526), .A2(n22204), .B1(n22244), .B2(n16845), .ZN(
        n16531) );
  OR2_X1 U18620 ( .A1(n16540), .A2(n16527), .ZN(n16528) );
  NAND2_X1 U18621 ( .A1(n16529), .A2(n16528), .ZN(n16980) );
  NOR2_X1 U18622 ( .A1(n16980), .A2(n22237), .ZN(n16530) );
  AOI211_X1 U18623 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n22201), .A(n16531), .B(
        n16530), .ZN(n16532) );
  OAI211_X1 U18624 ( .C1(n16535), .C2(n16534), .A(n16533), .B(n16532), .ZN(
        P1_U2816) );
  INV_X1 U18625 ( .A(n16524), .ZN(n16536) );
  OAI21_X1 U18626 ( .B1(n16537), .B2(n11219), .A(n16536), .ZN(n16852) );
  NOR2_X1 U18627 ( .A1(n16552), .A2(n16538), .ZN(n16539) );
  OR2_X1 U18628 ( .A1(n16540), .A2(n16539), .ZN(n16699) );
  INV_X1 U18629 ( .A(n16699), .ZN(n22105) );
  AOI22_X1 U18630 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n22242), .B1(
        n22216), .B2(n16855), .ZN(n16541) );
  OAI21_X1 U18631 ( .B1(n22235), .B2(n16700), .A(n16541), .ZN(n16545) );
  AOI211_X1 U18632 ( .C1(n20563), .C2(n16543), .A(n22228), .B(n16542), .ZN(
        n16544) );
  AOI211_X1 U18633 ( .C1(n22199), .C2(n22105), .A(n16545), .B(n16544), .ZN(
        n16546) );
  OAI21_X1 U18634 ( .B1(n16852), .B2(n22238), .A(n16546), .ZN(P1_U2817) );
  NOR2_X1 U18635 ( .A1(n16547), .A2(n16548), .ZN(n16549) );
  OR2_X1 U18636 ( .A1(n11219), .A2(n16549), .ZN(n20698) );
  AND2_X1 U18637 ( .A1(n16565), .A2(n16550), .ZN(n16551) );
  NOR2_X1 U18638 ( .A1(n16552), .A2(n16551), .ZN(n16995) );
  INV_X1 U18639 ( .A(n16569), .ZN(n16553) );
  AND2_X1 U18640 ( .A1(n22190), .A2(n16553), .ZN(n16554) );
  OR2_X1 U18641 ( .A1(n22228), .A2(n16554), .ZN(n16590) );
  OAI21_X1 U18642 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n22197), .A(n16590), 
        .ZN(n16555) );
  MUX2_X1 U18643 ( .A(n16556), .B(n16555), .S(P1_REIP_REG_22__SCAN_IN), .Z(
        n16559) );
  INV_X1 U18644 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16557) );
  NOR2_X1 U18645 ( .A1(n22204), .A2(n16557), .ZN(n16558) );
  AOI211_X1 U18646 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n22201), .A(n16559), .B(
        n16558), .ZN(n16560) );
  OAI21_X1 U18647 ( .B1(n20702), .B2(n22244), .A(n16560), .ZN(n16561) );
  AOI21_X1 U18648 ( .B1(n16995), .B2(n22199), .A(n16561), .ZN(n16562) );
  OAI21_X1 U18649 ( .B1(n20698), .B2(n22238), .A(n16562), .ZN(P1_U2818) );
  NAND2_X1 U18650 ( .A1(n16581), .A2(n16563), .ZN(n16564) );
  NAND2_X1 U18651 ( .A1(n16565), .A2(n16564), .ZN(n22075) );
  AOI21_X1 U18652 ( .B1(n16568), .B2(n16567), .A(n16547), .ZN(n16865) );
  NAND2_X1 U18653 ( .A1(n16865), .A2(n22215), .ZN(n16576) );
  INV_X1 U18654 ( .A(n16590), .ZN(n16574) );
  NOR3_X1 U18655 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n22197), .A3(n16569), 
        .ZN(n16570) );
  AOI21_X1 U18656 ( .B1(n22242), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16570), .ZN(n16572) );
  NAND2_X1 U18657 ( .A1(n22216), .A2(n16861), .ZN(n16571) );
  OAI211_X1 U18658 ( .C1(n22235), .C2(n16702), .A(n16572), .B(n16571), .ZN(
        n16573) );
  AOI21_X1 U18659 ( .B1(n16574), .B2(P1_REIP_REG_21__SCAN_IN), .A(n16573), 
        .ZN(n16575) );
  OAI211_X1 U18660 ( .C1(n22237), .C2(n22075), .A(n16576), .B(n16575), .ZN(
        P1_U2819) );
  NAND2_X1 U18661 ( .A1(n22222), .A2(n16663), .ZN(n16602) );
  INV_X1 U18662 ( .A(n16602), .ZN(n16651) );
  AOI21_X1 U18663 ( .B1(n16577), .B2(n16651), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n16591) );
  INV_X1 U18664 ( .A(n16567), .ZN(n16579) );
  AOI21_X1 U18665 ( .B1(n16580), .B2(n16593), .A(n16579), .ZN(n20690) );
  NAND2_X1 U18666 ( .A1(n20690), .A2(n22215), .ZN(n16589) );
  OAI21_X1 U18667 ( .B1(n16595), .B2(n16582), .A(n16581), .ZN(n16583) );
  INV_X1 U18668 ( .A(n16583), .ZN(n17013) );
  INV_X1 U18669 ( .A(n20693), .ZN(n16584) );
  AOI22_X1 U18670 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n22242), .B1(
        n22216), .B2(n16584), .ZN(n16585) );
  OAI21_X1 U18671 ( .B1(n22235), .B2(n16586), .A(n16585), .ZN(n16587) );
  AOI21_X1 U18672 ( .B1(n17013), .B2(n22199), .A(n16587), .ZN(n16588) );
  OAI211_X1 U18673 ( .C1(n16591), .C2(n16590), .A(n16589), .B(n16588), .ZN(
        P1_U2820) );
  AOI21_X1 U18674 ( .B1(n16594), .B2(n16592), .A(n16578), .ZN(n16873) );
  INV_X1 U18675 ( .A(n16873), .ZN(n16767) );
  NAND2_X1 U18676 ( .A1(n16615), .A2(n16596), .ZN(n16597) );
  NAND2_X1 U18677 ( .A1(n11629), .A2(n16597), .ZN(n16705) );
  INV_X1 U18678 ( .A(n16705), .ZN(n22065) );
  NAND2_X1 U18679 ( .A1(n22201), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n16601) );
  NAND2_X1 U18680 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n16651), .ZN(n16643) );
  NOR2_X1 U18681 ( .A1(n20549), .A2(n16643), .ZN(n22231) );
  NAND2_X1 U18682 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n22231), .ZN(n22229) );
  NOR2_X1 U18683 ( .A1(n20551), .A2(n22229), .ZN(n16598) );
  NOR2_X1 U18684 ( .A1(n22228), .A2(n16598), .ZN(n16627) );
  AND2_X1 U18685 ( .A1(n20554), .A2(n16598), .ZN(n16609) );
  OAI21_X1 U18686 ( .B1(n16627), .B2(n16609), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n16600) );
  AOI22_X1 U18687 ( .A1(n22242), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n22216), .B2(n16869), .ZN(n16599) );
  NAND4_X1 U18688 ( .A1(n16601), .A2(n16600), .A3(n16599), .A4(n22232), .ZN(
        n16605) );
  NOR3_X1 U18689 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n16603), .A3(n16602), 
        .ZN(n16604) );
  AOI211_X1 U18690 ( .C1(n22065), .C2(n22199), .A(n16605), .B(n16604), .ZN(
        n16606) );
  OAI21_X1 U18691 ( .B1(n16767), .B2(n22238), .A(n16606), .ZN(P1_U2821) );
  OAI21_X1 U18692 ( .B1(n16607), .B2(n16608), .A(n16592), .ZN(n16877) );
  INV_X1 U18693 ( .A(n22232), .ZN(n22213) );
  NOR2_X1 U18694 ( .A1(n22213), .A2(n16609), .ZN(n16612) );
  INV_X1 U18695 ( .A(n16879), .ZN(n16610) );
  AOI22_X1 U18696 ( .A1(n16610), .A2(n22216), .B1(n22242), .B2(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16611) );
  OAI211_X1 U18697 ( .C1(n22235), .C2(n16707), .A(n16612), .B(n16611), .ZN(
        n16617) );
  NAND2_X1 U18698 ( .A1(n16624), .A2(n16613), .ZN(n16614) );
  NAND2_X1 U18699 ( .A1(n16615), .A2(n16614), .ZN(n22042) );
  NOR2_X1 U18700 ( .A1(n22042), .A2(n22237), .ZN(n16616) );
  AOI211_X1 U18701 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n16627), .A(n16617), 
        .B(n16616), .ZN(n16618) );
  OAI21_X1 U18702 ( .B1(n16877), .B2(n22238), .A(n16618), .ZN(P1_U2822) );
  INV_X1 U18703 ( .A(n16619), .ZN(n16622) );
  INV_X1 U18704 ( .A(n16620), .ZN(n16621) );
  AOI21_X1 U18705 ( .B1(n16622), .B2(n16621), .A(n16607), .ZN(n16892) );
  INV_X1 U18706 ( .A(n16892), .ZN(n16774) );
  OR2_X1 U18707 ( .A1(n16714), .A2(n16623), .ZN(n16625) );
  AND2_X1 U18708 ( .A1(n16625), .A2(n16624), .ZN(n22051) );
  NAND2_X1 U18709 ( .A1(n20551), .A2(n22229), .ZN(n16626) );
  NAND2_X1 U18710 ( .A1(n16627), .A2(n16626), .ZN(n16633) );
  NAND2_X1 U18711 ( .A1(n22242), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16630) );
  INV_X1 U18712 ( .A(n16890), .ZN(n16628) );
  NAND2_X1 U18713 ( .A1(n22216), .A2(n16628), .ZN(n16629) );
  NAND3_X1 U18714 ( .A1(n16630), .A2(n16629), .A3(n22232), .ZN(n16631) );
  AOI21_X1 U18715 ( .B1(n22201), .B2(P1_EBX_REG_17__SCAN_IN), .A(n16631), .ZN(
        n16632) );
  NAND2_X1 U18716 ( .A1(n16633), .A2(n16632), .ZN(n16634) );
  AOI21_X1 U18717 ( .B1(n22051), .B2(n22199), .A(n16634), .ZN(n16635) );
  OAI21_X1 U18718 ( .B1(n16774), .B2(n22238), .A(n16635), .ZN(P1_U2823) );
  XNOR2_X1 U18719 ( .A(n16636), .B(n13272), .ZN(n20614) );
  INV_X1 U18720 ( .A(n20614), .ZN(n16784) );
  INV_X1 U18721 ( .A(n16650), .ZN(n16640) );
  INV_X1 U18722 ( .A(n16638), .ZN(n16639) );
  OAI21_X1 U18723 ( .B1(n11180), .B2(n16640), .A(n16639), .ZN(n16641) );
  NAND2_X1 U18724 ( .A1(n16641), .A2(n16716), .ZN(n20612) );
  INV_X1 U18725 ( .A(n20612), .ZN(n17027) );
  OAI22_X1 U18726 ( .A1(n22235), .A2(n20616), .B1(n16900), .B2(n22244), .ZN(
        n16645) );
  NAND2_X1 U18727 ( .A1(n22161), .A2(n16643), .ZN(n16657) );
  AOI21_X1 U18728 ( .B1(n22242), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n22213), .ZN(n16642) );
  OAI221_X1 U18729 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n16643), .C1(n20549), 
        .C2(n16657), .A(n16642), .ZN(n16644) );
  AOI211_X1 U18730 ( .C1(n17027), .C2(n22199), .A(n16645), .B(n16644), .ZN(
        n16646) );
  OAI21_X1 U18731 ( .B1(n16784), .B2(n22238), .A(n16646), .ZN(P1_U2825) );
  OR2_X1 U18732 ( .A1(n16647), .A2(n16648), .ZN(n16649) );
  AND2_X1 U18733 ( .A1(n16636), .A2(n16649), .ZN(n20677) );
  INV_X1 U18734 ( .A(n20677), .ZN(n16787) );
  XNOR2_X1 U18735 ( .A(n11180), .B(n16650), .ZN(n21976) );
  NOR2_X1 U18736 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n16651), .ZN(n16656) );
  NAND2_X1 U18737 ( .A1(n22216), .A2(n20675), .ZN(n16652) );
  OAI211_X1 U18738 ( .C1(n22204), .C2(n16653), .A(n22232), .B(n16652), .ZN(
        n16654) );
  AOI21_X1 U18739 ( .B1(n22201), .B2(P1_EBX_REG_14__SCAN_IN), .A(n16654), .ZN(
        n16655) );
  OAI21_X1 U18740 ( .B1(n16657), .B2(n16656), .A(n16655), .ZN(n16658) );
  AOI21_X1 U18741 ( .B1(n21976), .B2(n22199), .A(n16658), .ZN(n16659) );
  OAI21_X1 U18742 ( .B1(n16787), .B2(n22238), .A(n16659), .ZN(P1_U2826) );
  INV_X1 U18743 ( .A(n16660), .ZN(n16661) );
  AOI21_X1 U18744 ( .B1(n16662), .B2(n16661), .A(n16647), .ZN(n16914) );
  INV_X1 U18745 ( .A(n16914), .ZN(n16792) );
  AOI211_X1 U18746 ( .C1(n21966), .C2(n16664), .A(n16663), .B(n22197), .ZN(
        n16672) );
  OAI22_X1 U18747 ( .A1(n22235), .A2(n16720), .B1(n16665), .B2(n22204), .ZN(
        n16666) );
  INV_X1 U18748 ( .A(n16666), .ZN(n16667) );
  OAI211_X1 U18749 ( .C1(n22190), .C2(n21966), .A(n16667), .B(n22232), .ZN(
        n16671) );
  NAND2_X1 U18750 ( .A1(n11274), .A2(n16668), .ZN(n16669) );
  AND2_X1 U18751 ( .A1(n11180), .A2(n16669), .ZN(n21964) );
  INV_X1 U18752 ( .A(n21964), .ZN(n16719) );
  OAI22_X1 U18753 ( .A1(n16719), .A2(n22237), .B1(n16912), .B2(n22244), .ZN(
        n16670) );
  NOR3_X1 U18754 ( .A1(n16672), .A2(n16671), .A3(n16670), .ZN(n16673) );
  OAI21_X1 U18755 ( .B1(n16792), .B2(n22238), .A(n16673), .ZN(P1_U2827) );
  INV_X1 U18756 ( .A(n16674), .ZN(n22383) );
  INV_X1 U18757 ( .A(n16675), .ZN(n16682) );
  AOI22_X1 U18758 ( .A1(n22242), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n22162), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n16676) );
  OAI21_X1 U18759 ( .B1(n22244), .B2(n16677), .A(n16676), .ZN(n16678) );
  AOI21_X1 U18760 ( .B1(n22201), .B2(P1_EBX_REG_2__SCAN_IN), .A(n16678), .ZN(
        n16681) );
  OAI211_X1 U18761 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), 
        .A(n22222), .B(n16679), .ZN(n16680) );
  OAI211_X1 U18762 ( .C1(n16682), .C2(n22237), .A(n16681), .B(n16680), .ZN(
        n16683) );
  AOI21_X1 U18763 ( .B1(n22383), .B2(n22127), .A(n16683), .ZN(n16684) );
  OAI21_X1 U18764 ( .B1(n16685), .B2(n22124), .A(n16684), .ZN(P1_U2838) );
  INV_X1 U18765 ( .A(n16940), .ZN(n16687) );
  OAI22_X1 U18766 ( .A1(n16687), .A2(n16724), .B1(n16686), .B2(n20621), .ZN(
        P1_U2841) );
  INV_X1 U18767 ( .A(n16952), .ZN(n16688) );
  OAI222_X1 U18768 ( .A1(n16723), .A2(n16730), .B1(n20621), .B2(n16689), .C1(
        n16688), .C2(n16724), .ZN(P1_U2842) );
  INV_X1 U18769 ( .A(n16958), .ZN(n16690) );
  OAI222_X1 U18770 ( .A1(n16691), .A2(n20621), .B1(n16724), .B2(n16690), .C1(
        n16734), .C2(n16723), .ZN(P1_U2843) );
  OAI222_X1 U18771 ( .A1(n16692), .A2(n20621), .B1(n16724), .B2(n16970), .C1(
        n16810), .C2(n16723), .ZN(P1_U2844) );
  INV_X1 U18772 ( .A(n22082), .ZN(n16693) );
  OAI222_X1 U18773 ( .A1(n16694), .A2(n20621), .B1(n16724), .B2(n16693), .C1(
        n16814), .C2(n20623), .ZN(P1_U2845) );
  INV_X1 U18774 ( .A(n16825), .ZN(n16743) );
  OAI222_X1 U18775 ( .A1(n16695), .A2(n20621), .B1(n16724), .B2(n16976), .C1(
        n16743), .C2(n20623), .ZN(P1_U2846) );
  INV_X1 U18776 ( .A(n16696), .ZN(n16837) );
  AOI22_X1 U18777 ( .A1(n22099), .A2(n20617), .B1(n16703), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n16697) );
  OAI21_X1 U18778 ( .B1(n16837), .B2(n16723), .A(n16697), .ZN(P1_U2847) );
  OAI222_X1 U18779 ( .A1(n16698), .A2(n20621), .B1(n16724), .B2(n16980), .C1(
        n16749), .C2(n16723), .ZN(P1_U2848) );
  OAI222_X1 U18780 ( .A1(n16700), .A2(n20621), .B1(n16724), .B2(n16699), .C1(
        n16852), .C2(n16723), .ZN(P1_U2849) );
  AOI22_X1 U18781 ( .A1(n16995), .A2(n20617), .B1(n16703), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n16701) );
  OAI21_X1 U18782 ( .B1(n20698), .B2(n20623), .A(n16701), .ZN(P1_U2850) );
  INV_X1 U18783 ( .A(n16865), .ZN(n16759) );
  OAI222_X1 U18784 ( .A1(n16702), .A2(n20621), .B1(n16724), .B2(n22075), .C1(
        n16759), .C2(n16723), .ZN(P1_U2851) );
  INV_X1 U18785 ( .A(n20690), .ZN(n16763) );
  AOI22_X1 U18786 ( .A1(n17013), .A2(n20617), .B1(n16703), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n16704) );
  OAI21_X1 U18787 ( .B1(n16763), .B2(n20623), .A(n16704), .ZN(P1_U2852) );
  INV_X1 U18788 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n16706) );
  OAI222_X1 U18789 ( .A1(n16706), .A2(n20621), .B1(n16724), .B2(n16705), .C1(
        n16767), .C2(n16723), .ZN(P1_U2853) );
  OAI22_X1 U18790 ( .A1(n22042), .A2(n16724), .B1(n16707), .B2(n20621), .ZN(
        n16708) );
  INV_X1 U18791 ( .A(n16708), .ZN(n16709) );
  OAI21_X1 U18792 ( .B1(n16877), .B2(n20623), .A(n16709), .ZN(P1_U2854) );
  INV_X1 U18793 ( .A(n22051), .ZN(n16710) );
  OAI222_X1 U18794 ( .A1(n16711), .A2(n20621), .B1(n16724), .B2(n16710), .C1(
        n16774), .C2(n16723), .ZN(P1_U2855) );
  AOI21_X1 U18795 ( .B1(n16713), .B2(n16712), .A(n16620), .ZN(n20685) );
  INV_X1 U18796 ( .A(n20685), .ZN(n22239) );
  INV_X1 U18797 ( .A(n16714), .ZN(n16718) );
  NAND2_X1 U18798 ( .A1(n16716), .A2(n16715), .ZN(n16717) );
  NAND2_X1 U18799 ( .A1(n16718), .A2(n16717), .ZN(n22236) );
  OAI222_X1 U18800 ( .A1(n22234), .A2(n20621), .B1(n16723), .B2(n22239), .C1(
        n22236), .C2(n16724), .ZN(P1_U2856) );
  OAI222_X1 U18801 ( .A1(n16720), .A2(n20621), .B1(n16724), .B2(n16719), .C1(
        n16792), .C2(n16723), .ZN(P1_U2859) );
  OAI21_X1 U18802 ( .B1(n16722), .B2(n16721), .A(n11274), .ZN(n22211) );
  OAI222_X1 U18803 ( .A1(n22211), .A2(n16724), .B1(n22210), .B2(n20621), .C1(
        n16723), .C2(n20665), .ZN(P1_U2860) );
  AOI22_X1 U18804 ( .A1(n16776), .A2(DATAI_30_), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n16775), .ZN(n16729) );
  AND2_X1 U18805 ( .A1(n16726), .A2(n12842), .ZN(n16727) );
  MUX2_X1 U18806 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n16731), .Z(
        n16785) );
  AOI22_X1 U18807 ( .A1(n16779), .A2(BUF1_REG_30__SCAN_IN), .B1(n16778), .B2(
        n16785), .ZN(n16728) );
  OAI211_X1 U18808 ( .C1(n16730), .C2(n16782), .A(n16729), .B(n16728), .ZN(
        P1_U2874) );
  AOI22_X1 U18809 ( .A1(n16776), .A2(DATAI_29_), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n16775), .ZN(n16733) );
  MUX2_X1 U18810 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n16731), .Z(
        n16788) );
  AOI22_X1 U18811 ( .A1(n16779), .A2(BUF1_REG_29__SCAN_IN), .B1(n16778), .B2(
        n16788), .ZN(n16732) );
  OAI211_X1 U18812 ( .C1(n16734), .C2(n16782), .A(n16733), .B(n16732), .ZN(
        P1_U2875) );
  AOI22_X1 U18813 ( .A1(n16776), .A2(DATAI_28_), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n16775), .ZN(n16736) );
  AOI22_X1 U18814 ( .A1(n16779), .A2(BUF1_REG_28__SCAN_IN), .B1(n16778), .B2(
        n22361), .ZN(n16735) );
  OAI211_X1 U18815 ( .C1(n16810), .C2(n16782), .A(n16736), .B(n16735), .ZN(
        P1_U2876) );
  AOI22_X1 U18816 ( .A1(n16776), .A2(DATAI_27_), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n16775), .ZN(n16739) );
  AOI22_X1 U18817 ( .A1(n16779), .A2(BUF1_REG_27__SCAN_IN), .B1(n16778), .B2(
        n16737), .ZN(n16738) );
  OAI211_X1 U18818 ( .C1(n16814), .C2(n16782), .A(n16739), .B(n16738), .ZN(
        P1_U2877) );
  AOI22_X1 U18819 ( .A1(n16776), .A2(DATAI_26_), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n16775), .ZN(n16742) );
  AOI22_X1 U18820 ( .A1(n16779), .A2(BUF1_REG_26__SCAN_IN), .B1(n16778), .B2(
        n16740), .ZN(n16741) );
  OAI211_X1 U18821 ( .C1(n16743), .C2(n16782), .A(n16742), .B(n16741), .ZN(
        P1_U2878) );
  AOI22_X1 U18822 ( .A1(n16776), .A2(DATAI_25_), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n16775), .ZN(n16745) );
  AOI22_X1 U18823 ( .A1(n16779), .A2(BUF1_REG_25__SCAN_IN), .B1(n16778), .B2(
        n22347), .ZN(n16744) );
  OAI211_X1 U18824 ( .C1(n16837), .C2(n16782), .A(n16745), .B(n16744), .ZN(
        P1_U2879) );
  AOI22_X1 U18825 ( .A1(n16776), .A2(DATAI_24_), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n16775), .ZN(n16748) );
  AOI22_X1 U18826 ( .A1(n16779), .A2(BUF1_REG_24__SCAN_IN), .B1(n16778), .B2(
        n16746), .ZN(n16747) );
  OAI211_X1 U18827 ( .C1(n16749), .C2(n16782), .A(n16748), .B(n16747), .ZN(
        P1_U2880) );
  AOI22_X1 U18828 ( .A1(n16776), .A2(DATAI_23_), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n16775), .ZN(n16752) );
  AOI22_X1 U18829 ( .A1(n16779), .A2(BUF1_REG_23__SCAN_IN), .B1(n16778), .B2(
        n16750), .ZN(n16751) );
  OAI211_X1 U18830 ( .C1(n16852), .C2(n16782), .A(n16752), .B(n16751), .ZN(
        P1_U2881) );
  AOI22_X1 U18831 ( .A1(n16776), .A2(DATAI_22_), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n16775), .ZN(n16755) );
  AOI22_X1 U18832 ( .A1(n16779), .A2(BUF1_REG_22__SCAN_IN), .B1(n16778), .B2(
        n16753), .ZN(n16754) );
  OAI211_X1 U18833 ( .C1(n20698), .C2(n16782), .A(n16755), .B(n16754), .ZN(
        P1_U2882) );
  AOI22_X1 U18834 ( .A1(n16776), .A2(DATAI_21_), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n16775), .ZN(n16758) );
  AOI22_X1 U18835 ( .A1(n16779), .A2(BUF1_REG_21__SCAN_IN), .B1(n16778), .B2(
        n16756), .ZN(n16757) );
  OAI211_X1 U18836 ( .C1(n16759), .C2(n16782), .A(n16758), .B(n16757), .ZN(
        P1_U2883) );
  AOI22_X1 U18837 ( .A1(n16776), .A2(DATAI_20_), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n16775), .ZN(n16762) );
  AOI22_X1 U18838 ( .A1(n16779), .A2(BUF1_REG_20__SCAN_IN), .B1(n16778), .B2(
        n16760), .ZN(n16761) );
  OAI211_X1 U18839 ( .C1(n16763), .C2(n16782), .A(n16762), .B(n16761), .ZN(
        P1_U2884) );
  AOI22_X1 U18840 ( .A1(n16776), .A2(DATAI_19_), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n16775), .ZN(n16766) );
  AOI22_X1 U18841 ( .A1(n16779), .A2(BUF1_REG_19__SCAN_IN), .B1(n16778), .B2(
        n16764), .ZN(n16765) );
  OAI211_X1 U18842 ( .C1(n16767), .C2(n16782), .A(n16766), .B(n16765), .ZN(
        P1_U2885) );
  AOI22_X1 U18843 ( .A1(n16776), .A2(DATAI_18_), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n16775), .ZN(n16770) );
  AOI22_X1 U18844 ( .A1(n16779), .A2(BUF1_REG_18__SCAN_IN), .B1(n16778), .B2(
        n16768), .ZN(n16769) );
  OAI211_X1 U18845 ( .C1(n16877), .C2(n16782), .A(n16770), .B(n16769), .ZN(
        P1_U2886) );
  AOI22_X1 U18846 ( .A1(n16776), .A2(DATAI_17_), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n16775), .ZN(n16773) );
  AOI22_X1 U18847 ( .A1(n16779), .A2(BUF1_REG_17__SCAN_IN), .B1(n16778), .B2(
        n16771), .ZN(n16772) );
  OAI211_X1 U18848 ( .C1(n16774), .C2(n16782), .A(n16773), .B(n16772), .ZN(
        P1_U2887) );
  AOI22_X1 U18849 ( .A1(n16776), .A2(DATAI_16_), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n16775), .ZN(n16781) );
  AOI22_X1 U18850 ( .A1(n16779), .A2(BUF1_REG_16__SCAN_IN), .B1(n16778), .B2(
        n16777), .ZN(n16780) );
  OAI211_X1 U18851 ( .C1(n22239), .C2(n16782), .A(n16781), .B(n16780), .ZN(
        P1_U2888) );
  OAI222_X1 U18852 ( .A1(n16782), .A2(n16784), .B1(n16791), .B2(n16783), .C1(
        n16789), .C2(n20527), .ZN(P1_U2889) );
  INV_X1 U18853 ( .A(n16785), .ZN(n22372) );
  OAI222_X1 U18854 ( .A1(n16787), .A2(n16782), .B1(n16791), .B2(n22372), .C1(
        n16786), .C2(n16789), .ZN(P1_U2890) );
  INV_X1 U18855 ( .A(n16788), .ZN(n22367) );
  OAI222_X1 U18856 ( .A1(n16782), .A2(n16792), .B1(n16791), .B2(n22367), .C1(
        n16790), .C2(n16789), .ZN(P1_U2891) );
  XOR2_X1 U18857 ( .A(n16794), .B(n16793), .Z(n16961) );
  NAND2_X1 U18858 ( .A1(n16795), .A2(n20689), .ZN(n16800) );
  NOR2_X1 U18859 ( .A1(n22093), .A2(n20573), .ZN(n16956) );
  NOR2_X1 U18860 ( .A1(n20646), .A2(n16796), .ZN(n16797) );
  AOI211_X1 U18861 ( .C1(n20676), .C2(n16798), .A(n16956), .B(n16797), .ZN(
        n16799) );
  OAI211_X1 U18862 ( .C1(n16961), .C2(n20696), .A(n16800), .B(n16799), .ZN(
        P1_U2970) );
  NOR2_X1 U18863 ( .A1(n22093), .A2(n20570), .ZN(n16967) );
  NOR2_X1 U18864 ( .A1(n20703), .A2(n16801), .ZN(n16802) );
  AOI211_X1 U18865 ( .C1(n20694), .C2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16967), .B(n16802), .ZN(n16809) );
  INV_X1 U18866 ( .A(n16926), .ZN(n16931) );
  OAI21_X1 U18867 ( .B1(n16931), .B2(n11670), .A(n16850), .ZN(n16806) );
  OAI21_X1 U18868 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n16803), .A(
        n16806), .ZN(n16805) );
  INV_X1 U18869 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n22087) );
  MUX2_X1 U18870 ( .A(n22087), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n11667), .Z(n16804) );
  OAI211_X1 U18871 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n16806), .A(
        n16805), .B(n16804), .ZN(n16807) );
  XNOR2_X1 U18872 ( .A(n16807), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16962) );
  NAND2_X1 U18873 ( .A1(n16962), .A2(n13804), .ZN(n16808) );
  OAI211_X1 U18874 ( .C1(n16810), .C2(n20697), .A(n16809), .B(n16808), .ZN(
        P1_U2971) );
  XNOR2_X1 U18875 ( .A(n11667), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16811) );
  XNOR2_X1 U18876 ( .A(n16812), .B(n16811), .ZN(n22081) );
  INV_X1 U18877 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16813) );
  OAI22_X1 U18878 ( .A1(n20646), .A2(n16813), .B1(n22093), .B2(n22085), .ZN(
        n16816) );
  NOR2_X1 U18879 ( .A1(n16814), .A2(n20697), .ZN(n16815) );
  AOI211_X2 U18880 ( .C1(n20676), .C2(n16817), .A(n16816), .B(n16815), .ZN(
        n16818) );
  OAI21_X1 U18881 ( .B1(n22081), .B2(n20696), .A(n16818), .ZN(P1_U2972) );
  OR2_X1 U18882 ( .A1(n16819), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16820) );
  NAND2_X1 U18883 ( .A1(n16821), .A2(n16820), .ZN(n16979) );
  NOR2_X1 U18884 ( .A1(n22093), .A2(n20568), .ZN(n16973) );
  AOI21_X1 U18885 ( .B1(n20694), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16973), .ZN(n16822) );
  OAI21_X1 U18886 ( .B1(n20703), .B2(n16823), .A(n16822), .ZN(n16824) );
  AOI21_X1 U18887 ( .B1(n16825), .B2(n20689), .A(n16824), .ZN(n16826) );
  OAI21_X1 U18888 ( .B1(n20696), .B2(n16979), .A(n16826), .ZN(P1_U2973) );
  MUX2_X1 U18889 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n16827), .S(
        n13786), .Z(n16830) );
  INV_X1 U18890 ( .A(n16850), .ZN(n16839) );
  NAND2_X1 U18891 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n22094) );
  INV_X1 U18892 ( .A(n22094), .ZN(n16828) );
  AOI21_X1 U18893 ( .B1(n16839), .B2(n16842), .A(n16828), .ZN(n16829) );
  XNOR2_X1 U18894 ( .A(n16831), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n22097) );
  AOI22_X1 U18895 ( .A1(n13804), .A2(n22097), .B1(n22102), .B2(
        P1_REIP_REG_25__SCAN_IN), .ZN(n16832) );
  OAI21_X1 U18896 ( .B1(n16833), .B2(n20646), .A(n16832), .ZN(n16834) );
  OAI21_X1 U18897 ( .B1(n16837), .B2(n20697), .A(n16836), .ZN(P1_U2974) );
  NAND2_X1 U18898 ( .A1(n16850), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16841) );
  NAND2_X1 U18899 ( .A1(n16839), .A2(n16838), .ZN(n16840) );
  MUX2_X1 U18900 ( .A(n16841), .B(n16840), .S(n11670), .Z(n16843) );
  XNOR2_X1 U18901 ( .A(n16843), .B(n16842), .ZN(n16989) );
  AOI22_X1 U18902 ( .A1(n20694), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n22102), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n16844) );
  OAI21_X1 U18903 ( .B1(n20703), .B2(n16845), .A(n16844), .ZN(n16846) );
  AOI21_X1 U18904 ( .B1(n16847), .B2(n20689), .A(n16846), .ZN(n16848) );
  OAI21_X1 U18905 ( .B1(n20696), .B2(n16989), .A(n16848), .ZN(P1_U2975) );
  XNOR2_X1 U18906 ( .A(n13786), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16849) );
  XNOR2_X1 U18907 ( .A(n16850), .B(n16849), .ZN(n22104) );
  INV_X1 U18908 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16851) );
  OAI22_X1 U18909 ( .A1(n20646), .A2(n16851), .B1(n22093), .B2(n20563), .ZN(
        n16854) );
  NOR2_X1 U18910 ( .A1(n16852), .A2(n20697), .ZN(n16853) );
  AOI211_X1 U18911 ( .C1(n20676), .C2(n16855), .A(n16854), .B(n16853), .ZN(
        n16856) );
  OAI21_X1 U18912 ( .B1(n22104), .B2(n20696), .A(n16856), .ZN(P1_U2976) );
  XNOR2_X1 U18913 ( .A(n11667), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16875) );
  AOI22_X1 U18914 ( .A1(n16876), .A2(n16875), .B1(n11670), .B2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16868) );
  INV_X1 U18915 ( .A(n16868), .ZN(n17010) );
  MUX2_X1 U18916 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n16868), .S(
        n11670), .Z(n17009) );
  NAND2_X1 U18917 ( .A1(n16857), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16858) );
  OAI211_X1 U18918 ( .C1(n16857), .C2(n17010), .A(n17009), .B(n16858), .ZN(
        n16860) );
  XNOR2_X1 U18919 ( .A(n16860), .B(n16859), .ZN(n22074) );
  INV_X1 U18920 ( .A(n16861), .ZN(n16863) );
  AOI22_X1 U18921 ( .A1(n20694), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n22102), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n16862) );
  OAI21_X1 U18922 ( .B1(n20703), .B2(n16863), .A(n16862), .ZN(n16864) );
  AOI21_X1 U18923 ( .B1(n16865), .B2(n20689), .A(n16864), .ZN(n16866) );
  OAI21_X1 U18924 ( .B1(n20696), .B2(n22074), .A(n16866), .ZN(P1_U2978) );
  XNOR2_X1 U18925 ( .A(n11670), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16867) );
  XNOR2_X1 U18926 ( .A(n16868), .B(n16867), .ZN(n22064) );
  INV_X1 U18927 ( .A(n16869), .ZN(n16871) );
  AOI22_X1 U18928 ( .A1(n20694), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n22102), .ZN(n16870) );
  OAI21_X1 U18929 ( .B1(n20703), .B2(n16871), .A(n16870), .ZN(n16872) );
  AOI21_X1 U18930 ( .B1(n16873), .B2(n20689), .A(n16872), .ZN(n16874) );
  OAI21_X1 U18931 ( .B1(n22064), .B2(n20696), .A(n16874), .ZN(P1_U2980) );
  XNOR2_X1 U18932 ( .A(n16876), .B(n16875), .ZN(n22044) );
  INV_X1 U18933 ( .A(n16877), .ZN(n16881) );
  AOI22_X1 U18934 ( .A1(n20694), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n22102), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n16878) );
  OAI21_X1 U18935 ( .B1(n20703), .B2(n16879), .A(n16878), .ZN(n16880) );
  AOI21_X1 U18936 ( .B1(n16881), .B2(n20689), .A(n16880), .ZN(n16882) );
  OAI21_X1 U18937 ( .B1(n22044), .B2(n20696), .A(n16882), .ZN(P1_U2981) );
  NAND2_X1 U18938 ( .A1(n13786), .A2(n22049), .ZN(n16886) );
  INV_X1 U18939 ( .A(n16896), .ZN(n16884) );
  NOR2_X1 U18940 ( .A1(n16884), .A2(n16883), .ZN(n16885) );
  MUX2_X1 U18941 ( .A(n16886), .B(n20681), .S(n16885), .Z(n16888) );
  INV_X1 U18942 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16887) );
  XNOR2_X1 U18943 ( .A(n16888), .B(n16887), .ZN(n22050) );
  AOI22_X1 U18944 ( .A1(n20694), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n22102), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16889) );
  OAI21_X1 U18945 ( .B1(n20703), .B2(n16890), .A(n16889), .ZN(n16891) );
  AOI21_X1 U18946 ( .B1(n16892), .B2(n20689), .A(n16891), .ZN(n16893) );
  OAI21_X1 U18947 ( .B1(n20696), .B2(n22050), .A(n16893), .ZN(P1_U2982) );
  MUX2_X1 U18948 ( .A(n17030), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .S(
        n11667), .Z(n16894) );
  NAND3_X1 U18949 ( .A1(n16896), .A2(n16895), .A3(n16894), .ZN(n20680) );
  INV_X1 U18950 ( .A(n20680), .ZN(n16898) );
  AOI21_X1 U18951 ( .B1(n16896), .B2(n16895), .A(n16894), .ZN(n16897) );
  NOR2_X1 U18952 ( .A1(n16898), .A2(n16897), .ZN(n17033) );
  NAND2_X1 U18953 ( .A1(n20694), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16899) );
  NAND2_X1 U18954 ( .A1(n22102), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n17029) );
  OAI211_X1 U18955 ( .C1(n20703), .C2(n16900), .A(n16899), .B(n17029), .ZN(
        n16901) );
  AOI21_X1 U18956 ( .B1(n20614), .B2(n20689), .A(n16901), .ZN(n16902) );
  OAI21_X1 U18957 ( .B1(n17033), .B2(n20696), .A(n16902), .ZN(P1_U2984) );
  INV_X1 U18958 ( .A(n20669), .ZN(n20654) );
  OAI21_X1 U18959 ( .B1(n20654), .B2(n16905), .A(n16904), .ZN(n20664) );
  INV_X1 U18960 ( .A(n16908), .ZN(n16907) );
  NAND2_X1 U18961 ( .A1(n16907), .A2(n16906), .ZN(n20663) );
  NOR2_X1 U18962 ( .A1(n20664), .A2(n20663), .ZN(n20662) );
  NOR2_X1 U18963 ( .A1(n20662), .A2(n16908), .ZN(n16910) );
  XNOR2_X1 U18964 ( .A(n16910), .B(n16909), .ZN(n21965) );
  INV_X1 U18965 ( .A(n21965), .ZN(n16916) );
  AOI22_X1 U18966 ( .A1(n20694), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n22102), .ZN(n16911) );
  OAI21_X1 U18967 ( .B1(n20703), .B2(n16912), .A(n16911), .ZN(n16913) );
  AOI21_X1 U18968 ( .B1(n16914), .B2(n20689), .A(n16913), .ZN(n16915) );
  OAI21_X1 U18969 ( .B1(n16916), .B2(n20696), .A(n16915), .ZN(P1_U2986) );
  NAND4_X1 U18970 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n22049), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n22041) );
  NOR2_X1 U18971 ( .A1(n22048), .A2(n22041), .ZN(n17001) );
  INV_X1 U18972 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16917) );
  NAND4_X1 U18973 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21974) );
  NOR2_X1 U18974 ( .A1(n16917), .A2(n21974), .ZN(n16920) );
  NAND3_X1 U18975 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16920), .A3(
        n16918), .ZN(n22020) );
  NOR2_X1 U18976 ( .A1(n22025), .A2(n22020), .ZN(n17022) );
  NAND2_X1 U18977 ( .A1(n17001), .A2(n17022), .ZN(n16996) );
  NOR3_X1 U18978 ( .A1(n16992), .A2(n16919), .A3(n16996), .ZN(n16928) );
  NOR2_X1 U18979 ( .A1(n16992), .A2(n16919), .ZN(n16925) );
  INV_X1 U18980 ( .A(n17001), .ZN(n16924) );
  INV_X1 U18981 ( .A(n16920), .ZN(n16922) );
  NOR3_X1 U18982 ( .A1(n16923), .A2(n16922), .A3(n16921), .ZN(n22017) );
  NAND3_X1 U18983 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n22017), .ZN(n17020) );
  NOR2_X1 U18984 ( .A1(n16924), .A2(n17020), .ZN(n16998) );
  NAND2_X1 U18985 ( .A1(n16925), .A2(n16998), .ZN(n16930) );
  NOR2_X1 U18986 ( .A1(n16930), .A2(n22022), .ZN(n16982) );
  AOI21_X1 U18987 ( .B1(n16928), .B2(n22021), .A(n16982), .ZN(n22110) );
  NOR2_X1 U18988 ( .A1(n22110), .A2(n16926), .ZN(n16972) );
  NAND2_X1 U18989 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n16972), .ZN(
        n22084) );
  NOR3_X1 U18990 ( .A1(n22084), .A2(n16965), .A3(n16927), .ZN(n16944) );
  NOR2_X1 U18991 ( .A1(n16933), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16939) );
  NOR2_X1 U18992 ( .A1(n22039), .A2(n21980), .ZN(n16935) );
  OAI221_X1 U18993 ( .B1(n22112), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), 
        .C1(n22112), .C2(n16928), .A(n22016), .ZN(n16929) );
  AOI21_X1 U18994 ( .B1(n21982), .B2(n16930), .A(n16929), .ZN(n16981) );
  OAI21_X1 U18995 ( .B1(n16931), .B2(n17025), .A(n16981), .ZN(n22098) );
  NOR2_X1 U18996 ( .A1(n16971), .A2(n22098), .ZN(n16932) );
  NOR2_X1 U18997 ( .A1(n16935), .A2(n16932), .ZN(n22089) );
  NOR2_X1 U18998 ( .A1(n17025), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16947) );
  NOR4_X1 U18999 ( .A1(n22089), .A2(n16947), .A3(n16933), .A4(n16965), .ZN(
        n16936) );
  NOR3_X1 U19000 ( .A1(n16936), .A2(n16935), .A3(n16934), .ZN(n16937) );
  AOI211_X1 U19001 ( .C1(n16944), .C2(n16939), .A(n16938), .B(n16937), .ZN(
        n16942) );
  NAND2_X1 U19002 ( .A1(n16940), .A2(n22106), .ZN(n16941) );
  OAI211_X1 U19003 ( .C1(n16943), .C2(n22043), .A(n16942), .B(n16941), .ZN(
        P1_U3000) );
  INV_X1 U19004 ( .A(n16944), .ZN(n16950) );
  INV_X1 U19005 ( .A(n16965), .ZN(n16946) );
  INV_X1 U19006 ( .A(n22089), .ZN(n16945) );
  OAI21_X1 U19007 ( .B1(n16946), .B2(n17025), .A(n16945), .ZN(n16957) );
  OAI21_X1 U19008 ( .B1(n16957), .B2(n16947), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16949) );
  OAI211_X1 U19009 ( .C1(n16950), .C2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16949), .B(n16948), .ZN(n16951) );
  AOI21_X1 U19010 ( .B1(n16952), .B2(n22106), .A(n16951), .ZN(n16953) );
  OAI21_X1 U19011 ( .B1(n16954), .B2(n22043), .A(n16953), .ZN(P1_U3001) );
  NOR3_X1 U19012 ( .A1(n22084), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n16965), .ZN(n16955) );
  AOI211_X1 U19013 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16957), .A(
        n16956), .B(n16955), .ZN(n16960) );
  NAND2_X1 U19014 ( .A1(n16958), .A2(n22106), .ZN(n16959) );
  OAI211_X1 U19015 ( .C1(n16961), .C2(n22043), .A(n16960), .B(n16959), .ZN(
        P1_U3002) );
  NAND2_X1 U19016 ( .A1(n16962), .A2(n22118), .ZN(n16969) );
  NOR2_X1 U19017 ( .A1(n16963), .A2(n22084), .ZN(n16964) );
  AND2_X1 U19018 ( .A1(n16965), .A2(n16964), .ZN(n16966) );
  AOI211_X1 U19019 ( .C1(n22089), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16967), .B(n16966), .ZN(n16968) );
  OAI211_X1 U19020 ( .C1(n22115), .C2(n16970), .A(n16969), .B(n16968), .ZN(
        P1_U3003) );
  AOI22_X1 U19021 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n22098), .B1(
        n16972), .B2(n16971), .ZN(n16975) );
  INV_X1 U19022 ( .A(n16973), .ZN(n16974) );
  OAI211_X1 U19023 ( .C1(n16976), .C2(n22115), .A(n16975), .B(n16974), .ZN(
        n16977) );
  INV_X1 U19024 ( .A(n16977), .ZN(n16978) );
  OAI21_X1 U19025 ( .B1(n16979), .B2(n22043), .A(n16978), .ZN(P1_U3005) );
  NOR2_X1 U19026 ( .A1(n16980), .A2(n22115), .ZN(n16987) );
  NOR3_X1 U19027 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n22110), .A3(
        n16838), .ZN(n16986) );
  NOR2_X1 U19028 ( .A1(n22093), .A2(n20565), .ZN(n16985) );
  INV_X1 U19029 ( .A(n16981), .ZN(n22103) );
  OAI221_X1 U19030 ( .B1(n22103), .B2(n16982), .C1(n22103), .C2(n16838), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16983) );
  INV_X1 U19031 ( .A(n16983), .ZN(n16984) );
  NOR4_X1 U19032 ( .A1(n16987), .A2(n16986), .A3(n16985), .A4(n16984), .ZN(
        n16988) );
  OAI21_X1 U19033 ( .B1(n16989), .B2(n22043), .A(n16988), .ZN(P1_U3007) );
  NAND2_X1 U19034 ( .A1(n16991), .A2(n16990), .ZN(n16993) );
  XNOR2_X1 U19035 ( .A(n16993), .B(n16992), .ZN(n20695) );
  NOR2_X1 U19036 ( .A1(n22093), .A2(n20561), .ZN(n16994) );
  AOI21_X1 U19037 ( .B1(n16995), .B2(n22106), .A(n16994), .ZN(n17004) );
  NAND2_X1 U19038 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17005) );
  AOI21_X1 U19039 ( .B1(n22021), .B2(n16996), .A(n21980), .ZN(n16997) );
  OAI21_X1 U19040 ( .B1(n22018), .B2(n16998), .A(n16997), .ZN(n22070) );
  OAI22_X1 U19041 ( .A1(n17005), .A2(n22070), .B1(n22039), .B2(n21980), .ZN(
        n22080) );
  INV_X1 U19042 ( .A(n22080), .ZN(n17002) );
  INV_X1 U19043 ( .A(n22122), .ZN(n17000) );
  NOR2_X1 U19044 ( .A1(n22111), .A2(n22123), .ZN(n16999) );
  AOI211_X1 U19045 ( .C1(n22021), .C2(n17022), .A(n17000), .B(n16999), .ZN(
        n21972) );
  AOI21_X1 U19046 ( .B1(n17020), .B2(n22112), .A(n21972), .ZN(n21968) );
  NAND2_X1 U19047 ( .A1(n17001), .A2(n21968), .ZN(n17014) );
  NOR3_X1 U19048 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17005), .A3(
        n17014), .ZN(n22073) );
  OAI21_X1 U19049 ( .B1(n17002), .B2(n22073), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17003) );
  NAND2_X1 U19050 ( .A1(n17004), .A2(n17003), .ZN(n17007) );
  NOR4_X1 U19051 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16859), .A3(
        n17005), .A4(n17014), .ZN(n17006) );
  NOR2_X1 U19052 ( .A1(n17007), .A2(n17006), .ZN(n17008) );
  OAI21_X1 U19053 ( .B1(n20695), .B2(n22043), .A(n17008), .ZN(P1_U3009) );
  OAI21_X1 U19054 ( .B1(n11403), .B2(n17010), .A(n17009), .ZN(n17011) );
  XNOR2_X1 U19055 ( .A(n17011), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n20688) );
  NOR3_X1 U19056 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11403), .A3(
        n17014), .ZN(n17018) );
  INV_X1 U19057 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20557) );
  NOR2_X1 U19058 ( .A1(n22093), .A2(n20557), .ZN(n17012) );
  AOI21_X1 U19059 ( .B1(n17013), .B2(n22106), .A(n17012), .ZN(n17016) );
  NOR2_X1 U19060 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17014), .ZN(
        n22069) );
  OAI21_X1 U19061 ( .B1(n22069), .B2(n22070), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17015) );
  NAND2_X1 U19062 ( .A1(n17016), .A2(n17015), .ZN(n17017) );
  AOI211_X1 U19063 ( .C1(n20688), .C2(n22118), .A(n17018), .B(n17017), .ZN(
        n17019) );
  INV_X1 U19064 ( .A(n17019), .ZN(P1_U3011) );
  NAND2_X1 U19065 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17023) );
  INV_X1 U19066 ( .A(n21968), .ZN(n22040) );
  NOR2_X1 U19067 ( .A1(n17023), .A2(n22040), .ZN(n22061) );
  AOI21_X1 U19068 ( .B1(n21982), .B2(n17020), .A(n21980), .ZN(n17021) );
  OAI21_X1 U19069 ( .B1(n17022), .B2(n22112), .A(n17021), .ZN(n22038) );
  INV_X1 U19070 ( .A(n17023), .ZN(n17024) );
  NOR2_X1 U19071 ( .A1(n17025), .A2(n17024), .ZN(n17026) );
  NOR2_X1 U19072 ( .A1(n22038), .A2(n17026), .ZN(n22057) );
  NAND2_X1 U19073 ( .A1(n17027), .A2(n22106), .ZN(n17028) );
  OAI211_X1 U19074 ( .C1(n22057), .C2(n17030), .A(n17029), .B(n17028), .ZN(
        n17031) );
  AOI21_X1 U19075 ( .B1(n17030), .B2(n22061), .A(n17031), .ZN(n17032) );
  OAI21_X1 U19076 ( .B1(n17033), .B2(n22043), .A(n17032), .ZN(P1_U3016) );
  INV_X1 U19077 ( .A(n17034), .ZN(n17035) );
  NOR2_X1 U19078 ( .A1(n17035), .A2(n22255), .ZN(n22263) );
  AOI21_X1 U19079 ( .B1(n13083), .B2(n17036), .A(n22263), .ZN(n17037) );
  OAI21_X1 U19080 ( .B1(n13696), .B2(n22506), .A(n17037), .ZN(n17038) );
  MUX2_X1 U19081 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n17038), .S(
        n17898), .Z(P1_U3478) );
  INV_X1 U19082 ( .A(n15965), .ZN(n22501) );
  INV_X1 U19083 ( .A(n17066), .ZN(n17041) );
  NOR3_X1 U19084 ( .A1(n17039), .A2(n15430), .A3(n17059), .ZN(n17040) );
  AOI211_X1 U19085 ( .C1(n22501), .C2(n17068), .A(n17041), .B(n17040), .ZN(
        n17871) );
  INV_X1 U19086 ( .A(n17824), .ZN(n17072) );
  INV_X1 U19087 ( .A(n17042), .ZN(n17045) );
  NOR3_X1 U19088 ( .A1(n15430), .A2(n17059), .A3(n17070), .ZN(n17043) );
  AOI21_X1 U19089 ( .B1(n17045), .B2(n17044), .A(n17043), .ZN(n17046) );
  OAI21_X1 U19090 ( .B1(n17871), .B2(n17072), .A(n17046), .ZN(n17048) );
  INV_X1 U19091 ( .A(n17047), .ZN(n17826) );
  MUX2_X1 U19092 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n17048), .S(
        n17826), .Z(P1_U3473) );
  INV_X1 U19093 ( .A(n17051), .ZN(n17050) );
  NAND2_X1 U19094 ( .A1(n17054), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17049) );
  NAND2_X1 U19095 ( .A1(n17050), .A2(n17049), .ZN(n17057) );
  MUX2_X1 U19096 ( .A(n17051), .B(n12757), .S(n17059), .Z(n17053) );
  OAI21_X1 U19097 ( .B1(n17054), .B2(n17053), .A(n17052), .ZN(n17055) );
  INV_X1 U19098 ( .A(n17055), .ZN(n17056) );
  AOI21_X1 U19099 ( .B1(n17058), .B2(n17057), .A(n17056), .ZN(n17065) );
  AOI21_X1 U19100 ( .B1(n17059), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n17060) );
  NOR2_X1 U19101 ( .A1(n17061), .A2(n17060), .ZN(n17069) );
  NAND3_X1 U19102 ( .A1(n17063), .A2(n17062), .A3(n17069), .ZN(n17064) );
  OAI211_X1 U19103 ( .C1(n17066), .C2(n12757), .A(n17065), .B(n17064), .ZN(
        n17067) );
  AOI21_X1 U19104 ( .B1(n22384), .B2(n17068), .A(n17067), .ZN(n17867) );
  INV_X1 U19105 ( .A(n17069), .ZN(n17071) );
  OAI22_X1 U19106 ( .A1(n17867), .A2(n17072), .B1(n17071), .B2(n17070), .ZN(
        n17073) );
  MUX2_X1 U19107 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17073), .S(
        n17826), .Z(P1_U3469) );
  NOR2_X1 U19108 ( .A1(n17074), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n17075) );
  MUX2_X1 U19109 ( .A(n11250), .B(n17075), .S(n11843), .Z(n17397) );
  INV_X1 U19110 ( .A(n17397), .ZN(n17092) );
  INV_X1 U19111 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n17077) );
  AOI22_X1 U19112 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n19124), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n19163), .ZN(n17076) );
  OAI21_X1 U19113 ( .B1(n17077), .B2(n19199), .A(n17076), .ZN(n17078) );
  AOI21_X1 U19114 ( .B1(n17080), .B2(n17079), .A(n17078), .ZN(n17091) );
  AOI22_X1 U19115 ( .A1(n12066), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n17082) );
  NAND2_X1 U19116 ( .A1(n12183), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n17081) );
  OAI211_X1 U19117 ( .C1(n17084), .C2(n17083), .A(n17082), .B(n17081), .ZN(
        n17086) );
  AOI222_X1 U19118 ( .A1(n12321), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12368), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n12192), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n17088) );
  XNOR2_X1 U19119 ( .A(n17089), .B(n17088), .ZN(n17542) );
  AOI22_X1 U19120 ( .A1(n17193), .A2(n19217), .B1(n19140), .B2(n17542), .ZN(
        n17090) );
  OAI211_X1 U19121 ( .C1(n17092), .C2(n19147), .A(n17091), .B(n17090), .ZN(
        P2_U2824) );
  NOR2_X1 U19122 ( .A1(n19193), .A2(n17093), .ZN(n17094) );
  XOR2_X1 U19123 ( .A(n17095), .B(n17094), .Z(n17097) );
  AOI22_X1 U19124 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19207), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19163), .ZN(n17096) );
  OAI21_X1 U19125 ( .B1(n19347), .B2(n17097), .A(n17096), .ZN(n17098) );
  INV_X1 U19126 ( .A(n17098), .ZN(n17103) );
  INV_X1 U19127 ( .A(n17206), .ZN(n17101) );
  OAI22_X1 U19128 ( .A1(n17296), .A2(n19222), .B1(n17099), .B2(n19182), .ZN(
        n17100) );
  AOI21_X1 U19129 ( .B1(n17101), .B2(n19217), .A(n17100), .ZN(n17102) );
  OAI211_X1 U19130 ( .C1(n17104), .C2(n19147), .A(n17103), .B(n17102), .ZN(
        P2_U2827) );
  INV_X1 U19131 ( .A(n17105), .ZN(n17109) );
  NAND2_X1 U19132 ( .A1(n11173), .A2(n17106), .ZN(n17108) );
  OAI21_X1 U19133 ( .B1(n17109), .B2(n17108), .A(n19194), .ZN(n17107) );
  AOI21_X1 U19134 ( .B1(n17109), .B2(n17108), .A(n17107), .ZN(n17110) );
  INV_X1 U19135 ( .A(n17110), .ZN(n17117) );
  INV_X1 U19136 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n18094) );
  OAI22_X1 U19137 ( .A1(n17111), .A2(n19182), .B1(n18094), .B2(n19210), .ZN(
        n17114) );
  OAI22_X1 U19138 ( .A1(n17303), .A2(n19222), .B1(n17112), .B2(n19199), .ZN(
        n17113) );
  AOI211_X1 U19139 ( .C1(n17115), .C2(n19217), .A(n17114), .B(n17113), .ZN(
        n17116) );
  OAI211_X1 U19140 ( .C1(n19147), .C2(n17118), .A(n17117), .B(n17116), .ZN(
        P2_U2828) );
  NOR2_X1 U19141 ( .A1(n19193), .A2(n17119), .ZN(n17121) );
  OAI21_X1 U19142 ( .B1(n17445), .B2(n17121), .A(n19194), .ZN(n17120) );
  AOI21_X1 U19143 ( .B1(n17445), .B2(n17121), .A(n17120), .ZN(n17134) );
  NOR2_X1 U19144 ( .A1(n17122), .A2(n19147), .ZN(n17133) );
  NOR2_X1 U19145 ( .A1(n17124), .A2(n17125), .ZN(n17126) );
  OR2_X1 U19146 ( .A1(n17123), .A2(n17126), .ZN(n17591) );
  INV_X1 U19147 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n18093) );
  OAI22_X1 U19148 ( .A1(n17443), .A2(n19182), .B1(n18093), .B2(n19210), .ZN(
        n17130) );
  XNOR2_X1 U19149 ( .A(n17139), .B(n17127), .ZN(n17586) );
  OAI22_X1 U19150 ( .A1(n17586), .A2(n19222), .B1(n17128), .B2(n19199), .ZN(
        n17129) );
  NOR2_X1 U19151 ( .A1(n17130), .A2(n17129), .ZN(n17131) );
  OAI21_X1 U19152 ( .B1(n17591), .B2(n19165), .A(n17131), .ZN(n17132) );
  OR3_X1 U19153 ( .A1(n17134), .A2(n17133), .A3(n17132), .ZN(P2_U2831) );
  INV_X1 U19154 ( .A(n17124), .ZN(n17135) );
  OAI21_X1 U19155 ( .B1(n17245), .B2(n17136), .A(n17135), .ZN(n17599) );
  NAND2_X1 U19156 ( .A1(n17343), .A2(n17137), .ZN(n17138) );
  NAND2_X1 U19157 ( .A1(n17139), .A2(n17138), .ZN(n17598) );
  INV_X1 U19158 ( .A(n17598), .ZN(n17336) );
  INV_X1 U19159 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n18092) );
  OAI22_X1 U19160 ( .A1(n17454), .A2(n19182), .B1(n18092), .B2(n19210), .ZN(
        n17142) );
  NOR2_X1 U19161 ( .A1(n19199), .A2(n17140), .ZN(n17141) );
  AOI211_X1 U19162 ( .C1(n17336), .C2(n19140), .A(n17142), .B(n17141), .ZN(
        n17143) );
  OAI21_X1 U19163 ( .B1(n17599), .B2(n19165), .A(n17143), .ZN(n17148) );
  AND2_X1 U19164 ( .A1(n11173), .A2(n17144), .ZN(n17146) );
  OAI21_X1 U19165 ( .B1(n17456), .B2(n17146), .A(n19194), .ZN(n17145) );
  AOI21_X1 U19166 ( .B1(n17456), .B2(n17146), .A(n17145), .ZN(n17147) );
  AOI211_X1 U19167 ( .C1(n19218), .C2(n17149), .A(n17148), .B(n17147), .ZN(
        n17150) );
  INV_X1 U19168 ( .A(n17150), .ZN(P2_U2832) );
  AND2_X1 U19169 ( .A1(n11173), .A2(n17151), .ZN(n19155) );
  NAND2_X1 U19170 ( .A1(n19155), .A2(n17479), .ZN(n17152) );
  OAI211_X1 U19171 ( .C1(n17479), .C2(n19155), .A(n17152), .B(n19194), .ZN(
        n17165) );
  NAND2_X1 U19172 ( .A1(n17154), .A2(n17153), .ZN(n17155) );
  NAND2_X1 U19173 ( .A1(n17243), .A2(n17155), .ZN(n17628) );
  INV_X1 U19174 ( .A(n17628), .ZN(n17163) );
  INV_X1 U19175 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n18090) );
  OAI22_X1 U19176 ( .A1(n12144), .A2(n19199), .B1(n18090), .B2(n19210), .ZN(
        n17162) );
  INV_X1 U19177 ( .A(n17156), .ZN(n17159) );
  INV_X1 U19178 ( .A(n17157), .ZN(n17158) );
  NAND2_X1 U19179 ( .A1(n17159), .A2(n17158), .ZN(n17160) );
  NAND2_X1 U19180 ( .A1(n17341), .A2(n17160), .ZN(n17624) );
  OAI22_X1 U19181 ( .A1(n17624), .A2(n19222), .B1(n17477), .B2(n19182), .ZN(
        n17161) );
  AOI211_X1 U19182 ( .C1(n17163), .C2(n19217), .A(n17162), .B(n17161), .ZN(
        n17164) );
  OAI211_X1 U19183 ( .C1(n19147), .C2(n17166), .A(n17165), .B(n17164), .ZN(
        P2_U2834) );
  AOI22_X1 U19184 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19208), .B1(
        n19140), .B2(n20199), .ZN(n17168) );
  NAND2_X1 U19185 ( .A1(n19207), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n17167) );
  OAI211_X1 U19186 ( .C1(n19147), .C2(n17169), .A(n17168), .B(n17167), .ZN(
        n17170) );
  AOI21_X1 U19187 ( .B1(P2_REIP_REG_2__SCAN_IN), .B2(n19163), .A(n17170), .ZN(
        n17171) );
  OAI21_X1 U19188 ( .B1(n17172), .B2(n19165), .A(n17171), .ZN(n17177) );
  INV_X1 U19189 ( .A(n17174), .ZN(n17903) );
  NOR2_X1 U19190 ( .A1(n19193), .A2(n17179), .ZN(n17175) );
  INV_X1 U19191 ( .A(n17175), .ZN(n17173) );
  AOI221_X1 U19192 ( .B1(n17903), .B2(n17175), .C1(n17174), .C2(n17173), .A(
        n19347), .ZN(n17176) );
  AOI211_X1 U19193 ( .C1(n19040), .C2(n18023), .A(n17177), .B(n17176), .ZN(
        n17178) );
  INV_X1 U19194 ( .A(n17178), .ZN(P2_U2853) );
  AOI211_X1 U19195 ( .C1(n17181), .C2(n17180), .A(n19193), .B(n17179), .ZN(
        n17776) );
  INV_X1 U19196 ( .A(n17776), .ZN(n17192) );
  INV_X1 U19197 ( .A(n17182), .ZN(n17183) );
  AOI22_X1 U19198 ( .A1(n19218), .A2(n17183), .B1(P2_EBX_REG_1__SCAN_IN), .B2(
        n19207), .ZN(n17184) );
  OAI21_X1 U19199 ( .B1(n19210), .B2(n17185), .A(n17184), .ZN(n17186) );
  AOI21_X1 U19200 ( .B1(n19140), .B2(n20249), .A(n17186), .ZN(n17187) );
  OAI21_X1 U19201 ( .B1(n17188), .B2(n19165), .A(n17187), .ZN(n17190) );
  MUX2_X1 U19202 ( .A(n19092), .B(n19124), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n17189) );
  AOI211_X1 U19203 ( .C1(n19040), .C2(n19860), .A(n17190), .B(n17189), .ZN(
        n17191) );
  OAI21_X1 U19204 ( .B1(n17192), .B2(n19347), .A(n17191), .ZN(P2_U2854) );
  MUX2_X1 U19205 ( .A(n17193), .B(P2_EBX_REG_31__SCAN_IN), .S(n14651), .Z(
        P2_U2856) );
  XNOR2_X1 U19206 ( .A(n17195), .B(n17194), .ZN(n17196) );
  XNOR2_X1 U19207 ( .A(n17197), .B(n17196), .ZN(n17292) );
  OR2_X1 U19208 ( .A1(n17199), .A2(n17198), .ZN(n17200) );
  NAND2_X1 U19209 ( .A1(n12188), .A2(n17200), .ZN(n17550) );
  NOR2_X1 U19210 ( .A1(n17550), .A2(n14651), .ZN(n17201) );
  AOI21_X1 U19211 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n14651), .A(n17201), .ZN(
        n17202) );
  OAI21_X1 U19212 ( .B1(n17292), .B2(n17272), .A(n17202), .ZN(P2_U2858) );
  NAND2_X1 U19213 ( .A1(n17209), .A2(n17203), .ZN(n17205) );
  XNOR2_X1 U19214 ( .A(n17205), .B(n17204), .ZN(n17299) );
  NOR2_X1 U19215 ( .A1(n17206), .A2(n14651), .ZN(n17207) );
  AOI21_X1 U19216 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n14651), .A(n17207), .ZN(
        n17208) );
  OAI21_X1 U19217 ( .B1(n17299), .B2(n17272), .A(n17208), .ZN(P2_U2859) );
  NOR2_X1 U19218 ( .A1(n17211), .A2(n14651), .ZN(n17212) );
  AOI21_X1 U19219 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n14651), .A(n17212), .ZN(
        n17213) );
  OAI21_X1 U19220 ( .B1(n17306), .B2(n17272), .A(n17213), .ZN(P2_U2860) );
  AOI21_X1 U19221 ( .B1(n17216), .B2(n17215), .A(n17214), .ZN(n17217) );
  INV_X1 U19222 ( .A(n17217), .ZN(n17316) );
  INV_X1 U19223 ( .A(n17219), .ZN(n17220) );
  AOI21_X1 U19224 ( .B1(n17221), .B2(n17218), .A(n17220), .ZN(n19202) );
  NOR2_X1 U19225 ( .A1(n17281), .A2(n12164), .ZN(n17222) );
  AOI21_X1 U19226 ( .B1(n19202), .B2(n17281), .A(n17222), .ZN(n17223) );
  OAI21_X1 U19227 ( .B1(n17316), .B2(n17272), .A(n17223), .ZN(P2_U2861) );
  OAI21_X1 U19228 ( .B1(n17224), .B2(n17226), .A(n17225), .ZN(n17317) );
  OR2_X1 U19229 ( .A1(n17123), .A2(n17227), .ZN(n17228) );
  NAND2_X1 U19230 ( .A1(n17218), .A2(n17228), .ZN(n17573) );
  NOR2_X1 U19231 ( .A1(n17573), .A2(n14651), .ZN(n17229) );
  AOI21_X1 U19232 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n14651), .A(n17229), .ZN(
        n17230) );
  OAI21_X1 U19233 ( .B1(n17317), .B2(n17272), .A(n17230), .ZN(P2_U2862) );
  OAI21_X1 U19234 ( .B1(n17231), .B2(n17233), .A(n17232), .ZN(n17332) );
  NOR2_X1 U19235 ( .A1(n17591), .A2(n14651), .ZN(n17234) );
  AOI21_X1 U19236 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n14651), .A(n17234), .ZN(
        n17235) );
  OAI21_X1 U19237 ( .B1(n17332), .B2(n17272), .A(n17235), .ZN(P2_U2863) );
  XNOR2_X1 U19238 ( .A(n17236), .B(n17237), .ZN(n17339) );
  NOR2_X1 U19239 ( .A1(n17599), .A2(n14651), .ZN(n17238) );
  AOI21_X1 U19240 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n14651), .A(n17238), .ZN(
        n17239) );
  OAI21_X1 U19241 ( .B1(n17339), .B2(n17272), .A(n17239), .ZN(P2_U2864) );
  OAI21_X1 U19242 ( .B1(n17240), .B2(n17241), .A(n17236), .ZN(n17350) );
  AND2_X1 U19243 ( .A1(n17243), .A2(n17242), .ZN(n17244) );
  NOR2_X1 U19244 ( .A1(n17245), .A2(n17244), .ZN(n17468) );
  INV_X1 U19245 ( .A(n17468), .ZN(n19166) );
  MUX2_X1 U19246 ( .A(n12148), .B(n19166), .S(n17281), .Z(n17246) );
  OAI21_X1 U19247 ( .B1(n17350), .B2(n17272), .A(n17246), .ZN(P2_U2865) );
  AOI21_X1 U19248 ( .B1(n17248), .B2(n17247), .A(n17240), .ZN(n17355) );
  NAND2_X1 U19249 ( .A1(n17355), .A2(n17274), .ZN(n17250) );
  NAND2_X1 U19250 ( .A1(n14651), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n17249) );
  OAI211_X1 U19251 ( .C1(n17628), .C2(n14651), .A(n17250), .B(n17249), .ZN(
        P2_U2866) );
  OAI21_X1 U19252 ( .B1(n11582), .B2(n11755), .A(n17247), .ZN(n17362) );
  MUX2_X1 U19253 ( .A(n19149), .B(n19152), .S(n17281), .Z(n17252) );
  OAI21_X1 U19254 ( .B1(n17362), .B2(n17272), .A(n17252), .ZN(P2_U2867) );
  OAI21_X1 U19255 ( .B1(n17253), .B2(n17254), .A(n17251), .ZN(n17373) );
  NOR2_X1 U19256 ( .A1(n17255), .A2(n17256), .ZN(n17257) );
  OR2_X1 U19257 ( .A1(n17258), .A2(n17257), .ZN(n19139) );
  NOR2_X1 U19258 ( .A1(n19139), .A2(n14651), .ZN(n17259) );
  AOI21_X1 U19259 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n14651), .A(n17259), .ZN(
        n17260) );
  OAI21_X1 U19260 ( .B1(n17373), .B2(n17272), .A(n17260), .ZN(P2_U2868) );
  AOI21_X1 U19261 ( .B1(n17261), .B2(n11179), .A(n17253), .ZN(n17262) );
  INV_X1 U19262 ( .A(n17262), .ZN(n17383) );
  INV_X1 U19263 ( .A(n17263), .ZN(n17266) );
  INV_X1 U19264 ( .A(n17264), .ZN(n17265) );
  AOI21_X1 U19265 ( .B1(n17266), .B2(n17265), .A(n17255), .ZN(n19128) );
  NOR2_X1 U19266 ( .A1(n17281), .A2(n12132), .ZN(n17267) );
  AOI21_X1 U19267 ( .B1(n19128), .B2(n17281), .A(n17267), .ZN(n17268) );
  OAI21_X1 U19268 ( .B1(n17383), .B2(n17272), .A(n17268), .ZN(P2_U2869) );
  OAI21_X1 U19269 ( .B1(n11191), .B2(n11299), .A(n11179), .ZN(n17392) );
  NAND2_X1 U19270 ( .A1(n14651), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n17271) );
  NAND2_X1 U19271 ( .A1(n17668), .A2(n17281), .ZN(n17270) );
  OAI211_X1 U19272 ( .C1(n17392), .C2(n17272), .A(n17271), .B(n17270), .ZN(
        P2_U2870) );
  AOI21_X1 U19273 ( .B1(n17273), .B2(n16244), .A(n11191), .ZN(n20321) );
  NAND2_X1 U19274 ( .A1(n20321), .A2(n17274), .ZN(n17280) );
  NAND2_X1 U19275 ( .A1(n17276), .A2(n17275), .ZN(n17277) );
  NAND2_X1 U19276 ( .A1(n17278), .A2(n17277), .ZN(n18007) );
  NAND2_X1 U19277 ( .A1(n19265), .A2(n17281), .ZN(n17279) );
  OAI211_X1 U19278 ( .C1(n17281), .C2(n12124), .A(n17280), .B(n17279), .ZN(
        P2_U2871) );
  INV_X1 U19279 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n17284) );
  AOI22_X1 U19280 ( .A1(n20315), .A2(n17282), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n20313), .ZN(n17283) );
  OAI21_X1 U19281 ( .B1(n17386), .B2(n17284), .A(n17283), .ZN(n17290) );
  OR2_X1 U19282 ( .A1(n17286), .A2(n17285), .ZN(n17287) );
  NOR2_X1 U19283 ( .A1(n19223), .A2(n20154), .ZN(n17289) );
  AOI211_X1 U19284 ( .C1(n20317), .C2(BUF1_REG_29__SCAN_IN), .A(n17290), .B(
        n17289), .ZN(n17291) );
  OAI21_X1 U19285 ( .B1(n17292), .B2(n20253), .A(n17291), .ZN(P2_U2890) );
  AOI22_X1 U19286 ( .A1(n20315), .A2(n17293), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n20313), .ZN(n17295) );
  AOI22_X1 U19287 ( .A1(n20317), .A2(BUF1_REG_28__SCAN_IN), .B1(n20316), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n17294) );
  OAI211_X1 U19288 ( .C1(n17296), .C2(n20154), .A(n17295), .B(n17294), .ZN(
        n17297) );
  INV_X1 U19289 ( .A(n17297), .ZN(n17298) );
  OAI21_X1 U19290 ( .B1(n17299), .B2(n20253), .A(n17298), .ZN(P2_U2891) );
  AOI22_X1 U19291 ( .A1(n20315), .A2(n17300), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n20313), .ZN(n17302) );
  AOI22_X1 U19292 ( .A1(n20317), .A2(BUF1_REG_27__SCAN_IN), .B1(n20316), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n17301) );
  OAI211_X1 U19293 ( .C1(n17303), .C2(n20154), .A(n17302), .B(n17301), .ZN(
        n17304) );
  INV_X1 U19294 ( .A(n17304), .ZN(n17305) );
  OAI21_X1 U19295 ( .B1(n17306), .B2(n20253), .A(n17305), .ZN(P2_U2892) );
  NAND2_X1 U19296 ( .A1(n17307), .A2(n17308), .ZN(n17309) );
  NAND2_X1 U19297 ( .A1(n11209), .A2(n17309), .ZN(n19206) );
  OAI22_X1 U19298 ( .A1(n19206), .A2(n20154), .B1(n17310), .B2(n20153), .ZN(
        n17313) );
  INV_X1 U19299 ( .A(n20317), .ZN(n17387) );
  INV_X1 U19300 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n17311) );
  OAI22_X1 U19301 ( .A1(n17387), .A2(n20766), .B1(n17386), .B2(n17311), .ZN(
        n17312) );
  AOI211_X1 U19302 ( .C1(n20315), .C2(n17314), .A(n17313), .B(n17312), .ZN(
        n17315) );
  OAI21_X1 U19303 ( .B1(n17316), .B2(n20253), .A(n17315), .ZN(P2_U2893) );
  NOR2_X1 U19304 ( .A1(n17317), .A2(n20253), .ZN(n17326) );
  INV_X1 U19305 ( .A(n20315), .ZN(n17334) );
  AOI22_X1 U19306 ( .A1(n20317), .A2(BUF1_REG_25__SCAN_IN), .B1(n20316), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n17324) );
  OR2_X1 U19307 ( .A1(n17319), .A2(n17318), .ZN(n17320) );
  NAND2_X1 U19308 ( .A1(n17307), .A2(n17320), .ZN(n19190) );
  OAI22_X1 U19309 ( .A1(n19190), .A2(n20154), .B1(n20153), .B2(n17321), .ZN(
        n17322) );
  INV_X1 U19310 ( .A(n17322), .ZN(n17323) );
  OAI211_X1 U19311 ( .C1(n19828), .C2(n17334), .A(n17324), .B(n17323), .ZN(
        n17325) );
  OR2_X1 U19312 ( .A1(n17326), .A2(n17325), .ZN(P2_U2894) );
  AOI22_X1 U19313 ( .A1(n20317), .A2(BUF1_REG_24__SCAN_IN), .B1(n20316), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U19314 ( .A1(n20315), .A2(n17327), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n20313), .ZN(n17328) );
  OAI211_X1 U19315 ( .C1(n17586), .C2(n20154), .A(n17329), .B(n17328), .ZN(
        n17330) );
  INV_X1 U19316 ( .A(n17330), .ZN(n17331) );
  OAI21_X1 U19317 ( .B1(n17332), .B2(n20253), .A(n17331), .ZN(P2_U2895) );
  OAI22_X1 U19318 ( .A1(n17334), .A2(n19833), .B1(n20153), .B2(n17333), .ZN(
        n17335) );
  AOI21_X1 U19319 ( .B1(n20319), .B2(n17336), .A(n17335), .ZN(n17338) );
  AOI22_X1 U19320 ( .A1(n20317), .A2(BUF1_REG_23__SCAN_IN), .B1(n20316), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n17337) );
  OAI211_X1 U19321 ( .C1(n17339), .C2(n20253), .A(n17338), .B(n17337), .ZN(
        P2_U2896) );
  NAND2_X1 U19322 ( .A1(n17341), .A2(n17340), .ZN(n17342) );
  NAND2_X1 U19323 ( .A1(n17343), .A2(n17342), .ZN(n19176) );
  OAI22_X1 U19324 ( .A1(n20154), .A2(n19176), .B1(n20153), .B2(n17344), .ZN(
        n17347) );
  INV_X1 U19325 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n17345) );
  OAI22_X1 U19326 ( .A1(n17387), .A2(n20757), .B1(n17386), .B2(n17345), .ZN(
        n17346) );
  AOI211_X1 U19327 ( .C1(n20315), .C2(n17348), .A(n17347), .B(n17346), .ZN(
        n17349) );
  OAI21_X1 U19328 ( .B1(n17350), .B2(n20253), .A(n17349), .ZN(P2_U2897) );
  INV_X1 U19329 ( .A(n20253), .ZN(n20320) );
  AOI22_X1 U19330 ( .A1(n20317), .A2(BUF1_REG_21__SCAN_IN), .B1(n20316), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U19331 ( .A1(n20315), .A2(n17351), .B1(n20313), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n17352) );
  OAI211_X1 U19332 ( .C1(n20154), .C2(n17624), .A(n17353), .B(n17352), .ZN(
        n17354) );
  AOI21_X1 U19333 ( .B1(n17355), .B2(n20320), .A(n17354), .ZN(n17356) );
  INV_X1 U19334 ( .A(n17356), .ZN(P2_U2898) );
  OAI22_X1 U19335 ( .A1(n20154), .A2(n19151), .B1(n20153), .B2(n17357), .ZN(
        n17360) );
  INV_X1 U19336 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n17358) );
  OAI22_X1 U19337 ( .A1(n17387), .A2(n20753), .B1(n17386), .B2(n17358), .ZN(
        n17359) );
  AOI211_X1 U19338 ( .C1(n20315), .C2(n20109), .A(n17360), .B(n17359), .ZN(
        n17361) );
  OAI21_X1 U19339 ( .B1(n17362), .B2(n20253), .A(n17361), .ZN(P2_U2899) );
  AND2_X1 U19340 ( .A1(n17377), .A2(n17363), .ZN(n17364) );
  NOR2_X1 U19341 ( .A1(n17365), .A2(n17364), .ZN(n19141) );
  INV_X1 U19342 ( .A(n19141), .ZN(n17367) );
  OAI22_X1 U19343 ( .A1(n20154), .A2(n17367), .B1(n20153), .B2(n17366), .ZN(
        n17370) );
  INV_X1 U19344 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n17368) );
  OAI22_X1 U19345 ( .A1(n17387), .A2(n20751), .B1(n17386), .B2(n17368), .ZN(
        n17369) );
  AOI211_X1 U19346 ( .C1(n20315), .C2(n17371), .A(n17370), .B(n17369), .ZN(
        n17372) );
  OAI21_X1 U19347 ( .B1(n17373), .B2(n20253), .A(n17372), .ZN(P2_U2900) );
  OR2_X1 U19348 ( .A1(n17375), .A2(n17374), .ZN(n17376) );
  NAND2_X1 U19349 ( .A1(n17377), .A2(n17376), .ZN(n19132) );
  OAI22_X1 U19350 ( .A1(n20154), .A2(n19132), .B1(n20153), .B2(n17378), .ZN(
        n17379) );
  AOI21_X1 U19351 ( .B1(n20315), .B2(n17380), .A(n17379), .ZN(n17382) );
  AOI22_X1 U19352 ( .A1(n20317), .A2(BUF1_REG_18__SCAN_IN), .B1(n20316), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n17381) );
  OAI211_X1 U19353 ( .C1(n17383), .C2(n20253), .A(n17382), .B(n17381), .ZN(
        P2_U2901) );
  OAI22_X1 U19354 ( .A1(n20154), .A2(n17666), .B1(n20153), .B2(n17384), .ZN(
        n17389) );
  INV_X1 U19355 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n17385) );
  OAI22_X1 U19356 ( .A1(n17387), .A2(n20747), .B1(n17386), .B2(n17385), .ZN(
        n17388) );
  AOI211_X1 U19357 ( .C1(n20315), .C2(n17390), .A(n17389), .B(n17388), .ZN(
        n17391) );
  OAI21_X1 U19358 ( .B1(n17392), .B2(n20253), .A(n17391), .ZN(P2_U2902) );
  INV_X1 U19359 ( .A(n17393), .ZN(n17395) );
  NAND2_X1 U19360 ( .A1(n17397), .A2(n14067), .ZN(n17398) );
  XNOR2_X1 U19361 ( .A(n17398), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17399) );
  XNOR2_X1 U19362 ( .A(n17400), .B(n17399), .ZN(n17547) );
  XNOR2_X1 U19363 ( .A(n17401), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17538) );
  NOR2_X1 U19364 ( .A1(n17544), .A2(n15057), .ZN(n17405) );
  NAND2_X1 U19365 ( .A1(n19282), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n17543) );
  NAND2_X1 U19366 ( .A1(n18003), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17402) );
  OAI211_X1 U19367 ( .C1(n18001), .C2(n17403), .A(n17543), .B(n17402), .ZN(
        n17404) );
  AOI211_X1 U19368 ( .C1(n17538), .C2(n18010), .A(n17405), .B(n17404), .ZN(
        n17406) );
  OAI21_X1 U19369 ( .B1(n17547), .B2(n18008), .A(n17406), .ZN(P2_U2983) );
  NAND2_X1 U19370 ( .A1(n17408), .A2(n17407), .ZN(n17410) );
  XOR2_X1 U19371 ( .A(n17410), .B(n17409), .Z(n17560) );
  INV_X1 U19372 ( .A(n17411), .ZN(n17412) );
  AOI21_X1 U19373 ( .B1(n17412), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17414) );
  NOR2_X1 U19374 ( .A1(n17414), .A2(n17413), .ZN(n17558) );
  NAND2_X1 U19375 ( .A1(n19282), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n17551) );
  OAI21_X1 U19376 ( .B1(n17987), .B2(n17415), .A(n17551), .ZN(n17416) );
  AOI21_X1 U19377 ( .B1(n18002), .B2(n17417), .A(n17416), .ZN(n17418) );
  OAI21_X1 U19378 ( .B1(n17550), .B2(n15057), .A(n17418), .ZN(n17419) );
  AOI21_X1 U19379 ( .B1(n17558), .B2(n18010), .A(n17419), .ZN(n17420) );
  OAI21_X1 U19380 ( .B1(n17560), .B2(n18008), .A(n17420), .ZN(P2_U2985) );
  INV_X1 U19381 ( .A(n17435), .ZN(n17422) );
  AOI21_X1 U19382 ( .B1(n17421), .B2(n17434), .A(n17422), .ZN(n17424) );
  MUX2_X1 U19383 ( .A(n17424), .B(n17434), .S(n17423), .Z(n17426) );
  NAND2_X1 U19384 ( .A1(n17426), .A2(n17425), .ZN(n17572) );
  NAND2_X1 U19385 ( .A1(n11183), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17431) );
  AOI21_X1 U19386 ( .B1(n17566), .B2(n17431), .A(n11220), .ZN(n17561) );
  NAND2_X1 U19387 ( .A1(n19202), .A2(n17998), .ZN(n17428) );
  INV_X1 U19388 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19198) );
  NOR2_X1 U19389 ( .A1(n19325), .A2(n19198), .ZN(n17562) );
  AOI21_X1 U19390 ( .B1(n18003), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17562), .ZN(n17427) );
  OAI211_X1 U19391 ( .C1(n19191), .C2(n18001), .A(n17428), .B(n17427), .ZN(
        n17429) );
  AOI21_X1 U19392 ( .B1(n17561), .B2(n18010), .A(n17429), .ZN(n17430) );
  OAI21_X1 U19393 ( .B1(n18008), .B2(n17572), .A(n17430), .ZN(P2_U2988) );
  OAI21_X1 U19394 ( .B1(n11183), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17431), .ZN(n17583) );
  NAND2_X1 U19395 ( .A1(n19282), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n17574) );
  OAI21_X1 U19396 ( .B1(n17987), .B2(n19183), .A(n17574), .ZN(n17433) );
  NOR2_X1 U19397 ( .A1(n17573), .A2(n15057), .ZN(n17432) );
  AOI211_X1 U19398 ( .C1(n18002), .C2(n11751), .A(n17433), .B(n17432), .ZN(
        n17438) );
  NAND2_X1 U19399 ( .A1(n17435), .A2(n17434), .ZN(n17436) );
  XOR2_X1 U19400 ( .A(n17436), .B(n17421), .Z(n17580) );
  NAND2_X1 U19401 ( .A1(n17580), .A2(n17983), .ZN(n17437) );
  OAI211_X1 U19402 ( .C1(n17583), .C2(n17996), .A(n17438), .B(n17437), .ZN(
        P2_U2989) );
  NOR2_X1 U19403 ( .A1(n17440), .A2(n11255), .ZN(n17441) );
  XNOR2_X1 U19404 ( .A(n17439), .B(n17441), .ZN(n17595) );
  AOI21_X1 U19405 ( .B1(n17442), .B2(n11434), .A(n11183), .ZN(n17593) );
  NAND2_X1 U19406 ( .A1(n19282), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n17585) );
  OAI21_X1 U19407 ( .B1(n17987), .B2(n17443), .A(n17585), .ZN(n17444) );
  AOI21_X1 U19408 ( .B1(n18002), .B2(n17445), .A(n17444), .ZN(n17446) );
  OAI21_X1 U19409 ( .B1(n17591), .B2(n15057), .A(n17446), .ZN(n17447) );
  AOI21_X1 U19410 ( .B1(n17593), .B2(n18010), .A(n17447), .ZN(n17448) );
  OAI21_X1 U19411 ( .B1(n17595), .B2(n18008), .A(n17448), .ZN(P2_U2990) );
  NAND2_X1 U19412 ( .A1(n11259), .A2(n17449), .ZN(n17450) );
  XNOR2_X1 U19413 ( .A(n17451), .B(n17450), .ZN(n17608) );
  NAND2_X1 U19414 ( .A1(n17475), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17460) );
  AOI21_X1 U19415 ( .B1(n17453), .B2(n17460), .A(n17452), .ZN(n17606) );
  NAND2_X1 U19416 ( .A1(n19282), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n17597) );
  OAI21_X1 U19417 ( .B1(n17987), .B2(n17454), .A(n17597), .ZN(n17455) );
  AOI21_X1 U19418 ( .B1(n18002), .B2(n17456), .A(n17455), .ZN(n17457) );
  OAI21_X1 U19419 ( .B1(n17599), .B2(n15057), .A(n17457), .ZN(n17458) );
  AOI21_X1 U19420 ( .B1(n17606), .B2(n18010), .A(n17458), .ZN(n17459) );
  OAI21_X1 U19421 ( .B1(n18008), .B2(n17608), .A(n17459), .ZN(P2_U2991) );
  OAI21_X1 U19422 ( .B1(n17475), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n17460), .ZN(n17618) );
  INV_X1 U19423 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n18091) );
  NOR2_X1 U19424 ( .A1(n19325), .A2(n18091), .ZN(n17610) );
  AOI21_X1 U19425 ( .B1(n18003), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17610), .ZN(n17461) );
  OAI21_X1 U19426 ( .B1(n18001), .B2(n19169), .A(n17461), .ZN(n17467) );
  INV_X1 U19427 ( .A(n17462), .ZN(n17463) );
  AOI21_X1 U19428 ( .B1(n17465), .B2(n17464), .A(n17463), .ZN(n17612) );
  NOR2_X1 U19429 ( .A1(n17612), .A2(n18008), .ZN(n17466) );
  AOI211_X1 U19430 ( .C1(n17998), .C2(n17468), .A(n17467), .B(n17466), .ZN(
        n17469) );
  OAI21_X1 U19431 ( .B1(n17618), .B2(n17996), .A(n17469), .ZN(P2_U2992) );
  NAND2_X1 U19432 ( .A1(n17472), .A2(n17471), .ZN(n17473) );
  XNOR2_X1 U19433 ( .A(n17474), .B(n17473), .ZN(n17632) );
  AOI21_X1 U19434 ( .B1(n17488), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17476) );
  NOR2_X1 U19435 ( .A1(n17476), .A2(n17475), .ZN(n17630) );
  NAND2_X1 U19436 ( .A1(n19282), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n17623) );
  OAI21_X1 U19437 ( .B1(n17987), .B2(n17477), .A(n17623), .ZN(n17478) );
  AOI21_X1 U19438 ( .B1(n18002), .B2(n17479), .A(n17478), .ZN(n17480) );
  OAI21_X1 U19439 ( .B1(n17628), .B2(n15057), .A(n17480), .ZN(n17481) );
  AOI21_X1 U19440 ( .B1(n17630), .B2(n18010), .A(n17481), .ZN(n17482) );
  OAI21_X1 U19441 ( .B1(n17632), .B2(n18008), .A(n17482), .ZN(P2_U2993) );
  NAND2_X1 U19442 ( .A1(n14063), .A2(n17484), .ZN(n17487) );
  XOR2_X1 U19443 ( .A(n17487), .B(n17486), .Z(n17643) );
  AOI21_X1 U19444 ( .B1(n17633), .B2(n17494), .A(n17488), .ZN(n17641) );
  NAND2_X1 U19445 ( .A1(n19282), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n17635) );
  OAI21_X1 U19446 ( .B1(n17987), .B2(n17489), .A(n17635), .ZN(n17490) );
  AOI21_X1 U19447 ( .B1(n19135), .B2(n18002), .A(n17490), .ZN(n17491) );
  OAI21_X1 U19448 ( .B1(n19139), .B2(n15057), .A(n17491), .ZN(n17492) );
  AOI21_X1 U19449 ( .B1(n17641), .B2(n18010), .A(n17492), .ZN(n17493) );
  OAI21_X1 U19450 ( .B1(n17643), .B2(n18008), .A(n17493), .ZN(P2_U2995) );
  OAI21_X1 U19451 ( .B1(n11212), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17494), .ZN(n17653) );
  NOR2_X1 U19452 ( .A1(n19126), .A2(n18001), .ZN(n17497) );
  NAND2_X1 U19453 ( .A1(n19282), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n17645) );
  OAI21_X1 U19454 ( .B1(n17987), .B2(n17495), .A(n17645), .ZN(n17496) );
  AOI211_X1 U19455 ( .C1(n19128), .C2(n17998), .A(n17497), .B(n17496), .ZN(
        n17502) );
  NAND2_X1 U19456 ( .A1(n14062), .A2(n17498), .ZN(n17500) );
  XOR2_X1 U19457 ( .A(n17500), .B(n17499), .Z(n17650) );
  NAND2_X1 U19458 ( .A1(n17650), .A2(n17983), .ZN(n17501) );
  OAI211_X1 U19459 ( .C1(n17653), .C2(n17996), .A(n17502), .B(n17501), .ZN(
        P2_U2996) );
  INV_X1 U19460 ( .A(n17504), .ZN(n17507) );
  AND2_X1 U19461 ( .A1(n17504), .A2(n17503), .ZN(n17506) );
  OAI22_X1 U19462 ( .A1(n17508), .A2(n17507), .B1(n17506), .B2(n17505), .ZN(
        n17671) );
  NAND2_X1 U19463 ( .A1(n17509), .A2(n18002), .ZN(n17510) );
  NAND2_X1 U19464 ( .A1(n19282), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n17664) );
  OAI211_X1 U19465 ( .C1(n17511), .C2(n17987), .A(n17510), .B(n17664), .ZN(
        n17513) );
  AOI211_X1 U19466 ( .C1(n17663), .C2(n18011), .A(n17996), .B(n11212), .ZN(
        n17512) );
  AOI211_X1 U19467 ( .C1(n17668), .C2(n17998), .A(n17513), .B(n17512), .ZN(
        n17514) );
  OAI21_X1 U19468 ( .B1(n18008), .B2(n17671), .A(n17514), .ZN(P2_U2997) );
  NAND2_X1 U19469 ( .A1(n17516), .A2(n17515), .ZN(n17520) );
  NAND2_X1 U19470 ( .A1(n17517), .A2(n17686), .ZN(n17995) );
  INV_X1 U19471 ( .A(n17993), .ZN(n17518) );
  AOI21_X1 U19472 ( .B1(n17995), .B2(n17992), .A(n17518), .ZN(n17519) );
  XOR2_X1 U19473 ( .A(n17520), .B(n17519), .Z(n17683) );
  INV_X1 U19474 ( .A(n19274), .ZN(n17673) );
  INV_X1 U19475 ( .A(n17521), .ZN(n17990) );
  NAND2_X1 U19476 ( .A1(n17990), .A2(n17662), .ZN(n17672) );
  NAND3_X1 U19477 ( .A1(n17673), .A2(n18010), .A3(n17672), .ZN(n17528) );
  OAI22_X1 U19478 ( .A1(n17987), .A2(n17523), .B1(n17522), .B2(n19325), .ZN(
        n17525) );
  NOR2_X1 U19479 ( .A1(n17678), .A2(n15057), .ZN(n17524) );
  AOI211_X1 U19480 ( .C1(n18002), .C2(n17526), .A(n17525), .B(n17524), .ZN(
        n17527) );
  OAI211_X1 U19481 ( .C1(n17683), .C2(n18008), .A(n17528), .B(n17527), .ZN(
        P2_U2999) );
  XNOR2_X1 U19482 ( .A(n17529), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19311) );
  OAI21_X1 U19483 ( .B1(n17532), .B2(n17530), .A(n17531), .ZN(n19305) );
  INV_X1 U19484 ( .A(n19305), .ZN(n17536) );
  INV_X1 U19485 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19302) );
  OAI22_X1 U19486 ( .A1(n19302), .A2(n19325), .B1(n18001), .B2(n19050), .ZN(
        n17535) );
  INV_X1 U19487 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19044) );
  OAI22_X1 U19488 ( .A1(n17533), .A2(n15057), .B1(n17987), .B2(n19044), .ZN(
        n17534) );
  AOI211_X1 U19489 ( .C1(n17536), .C2(n17983), .A(n17535), .B(n17534), .ZN(
        n17537) );
  OAI21_X1 U19490 ( .B1(n19311), .B2(n17996), .A(n17537), .ZN(P2_U3008) );
  NAND2_X1 U19491 ( .A1(n17538), .A2(n19271), .ZN(n17546) );
  INV_X1 U19492 ( .A(n17540), .ZN(n17541) );
  OAI211_X1 U19493 ( .C1(n17547), .C2(n19304), .A(n17546), .B(n17545), .ZN(
        P2_U3015) );
  OAI211_X1 U19494 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17548), .ZN(n17555) );
  NAND2_X1 U19495 ( .A1(n17549), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17554) );
  INV_X1 U19496 ( .A(n17550), .ZN(n19216) );
  OAI21_X1 U19497 ( .B1(n19223), .B2(n19327), .A(n17551), .ZN(n17552) );
  AOI21_X1 U19498 ( .B1(n19216), .B2(n19329), .A(n17552), .ZN(n17553) );
  OAI211_X1 U19499 ( .C1(n17556), .C2(n17555), .A(n17554), .B(n17553), .ZN(
        n17557) );
  AOI21_X1 U19500 ( .B1(n17558), .B2(n19271), .A(n17557), .ZN(n17559) );
  OAI21_X1 U19501 ( .B1(n17560), .B2(n19304), .A(n17559), .ZN(P2_U3017) );
  NAND2_X1 U19502 ( .A1(n17561), .A2(n19271), .ZN(n17571) );
  NAND2_X1 U19503 ( .A1(n19202), .A2(n19329), .ZN(n17564) );
  INV_X1 U19504 ( .A(n17562), .ZN(n17563) );
  OAI211_X1 U19505 ( .C1(n19327), .C2(n19206), .A(n17564), .B(n17563), .ZN(
        n17569) );
  AOI211_X1 U19506 ( .C1(n17567), .C2(n17566), .A(n17565), .B(n17577), .ZN(
        n17568) );
  AOI211_X1 U19507 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17579), .A(
        n17569), .B(n17568), .ZN(n17570) );
  OAI211_X1 U19508 ( .C1(n17572), .C2(n19304), .A(n17571), .B(n17570), .ZN(
        P2_U3020) );
  INV_X1 U19509 ( .A(n17573), .ZN(n19186) );
  OAI21_X1 U19510 ( .B1(n19190), .B2(n19327), .A(n17574), .ZN(n17575) );
  AOI21_X1 U19511 ( .B1(n19186), .B2(n19329), .A(n17575), .ZN(n17576) );
  OAI21_X1 U19512 ( .B1(n17577), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17576), .ZN(n17578) );
  AOI21_X1 U19513 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17579), .A(
        n17578), .ZN(n17582) );
  NAND2_X1 U19514 ( .A1(n17580), .A2(n19335), .ZN(n17581) );
  OAI211_X1 U19515 ( .C1(n17583), .C2(n19332), .A(n17582), .B(n17581), .ZN(
        P2_U3021) );
  INV_X1 U19516 ( .A(n17584), .ZN(n17588) );
  OAI21_X1 U19517 ( .B1(n19327), .B2(n17586), .A(n17585), .ZN(n17587) );
  AOI21_X1 U19518 ( .B1(n17588), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n17587), .ZN(n17589) );
  OAI211_X1 U19519 ( .C1(n19285), .C2(n17591), .A(n17590), .B(n17589), .ZN(
        n17592) );
  AOI21_X1 U19520 ( .B1(n17593), .B2(n19271), .A(n17592), .ZN(n17594) );
  OAI21_X1 U19521 ( .B1(n17595), .B2(n19304), .A(n17594), .ZN(P2_U3022) );
  INV_X1 U19522 ( .A(n17616), .ZN(n17604) );
  OAI21_X1 U19523 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17596), .ZN(n17603) );
  OAI21_X1 U19524 ( .B1(n19327), .B2(n17598), .A(n17597), .ZN(n17601) );
  NOR2_X1 U19525 ( .A1(n17599), .A2(n19285), .ZN(n17600) );
  AOI211_X1 U19526 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n17626), .A(
        n17601), .B(n17600), .ZN(n17602) );
  OAI21_X1 U19527 ( .B1(n17604), .B2(n17603), .A(n17602), .ZN(n17605) );
  AOI21_X1 U19528 ( .B1(n17606), .B2(n19271), .A(n17605), .ZN(n17607) );
  OAI21_X1 U19529 ( .B1(n19304), .B2(n17608), .A(n17607), .ZN(P2_U3023) );
  NOR2_X1 U19530 ( .A1(n19327), .A2(n19176), .ZN(n17609) );
  AOI211_X1 U19531 ( .C1(n17626), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n17610), .B(n17609), .ZN(n17611) );
  OAI21_X1 U19532 ( .B1(n19166), .B2(n19285), .A(n17611), .ZN(n17614) );
  NOR2_X1 U19533 ( .A1(n17612), .A2(n19304), .ZN(n17613) );
  AOI211_X1 U19534 ( .C1(n17616), .C2(n17615), .A(n17614), .B(n17613), .ZN(
        n17617) );
  OAI21_X1 U19535 ( .B1(n17618), .B2(n19332), .A(n17617), .ZN(P2_U3024) );
  NOR2_X1 U19536 ( .A1(n17619), .A2(n17675), .ZN(n17620) );
  NAND2_X1 U19537 ( .A1(n17621), .A2(n17620), .ZN(n17622) );
  OAI211_X1 U19538 ( .C1(n19327), .C2(n17624), .A(n17623), .B(n17622), .ZN(
        n17625) );
  AOI21_X1 U19539 ( .B1(n17626), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n17625), .ZN(n17627) );
  OAI21_X1 U19540 ( .B1(n17628), .B2(n19285), .A(n17627), .ZN(n17629) );
  AOI21_X1 U19541 ( .B1(n17630), .B2(n19271), .A(n17629), .ZN(n17631) );
  OAI21_X1 U19542 ( .B1(n17632), .B2(n19304), .A(n17631), .ZN(P2_U3025) );
  NOR2_X1 U19543 ( .A1(n17634), .A2(n17633), .ZN(n17640) );
  OAI21_X1 U19544 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17636), .A(
        n17635), .ZN(n17637) );
  AOI21_X1 U19545 ( .B1(n19281), .B2(n19141), .A(n17637), .ZN(n17638) );
  OAI21_X1 U19546 ( .B1(n19139), .B2(n19285), .A(n17638), .ZN(n17639) );
  AOI211_X1 U19547 ( .C1(n17641), .C2(n19271), .A(n17640), .B(n17639), .ZN(
        n17642) );
  OAI21_X1 U19548 ( .B1(n17643), .B2(n19304), .A(n17642), .ZN(P2_U3027) );
  OAI211_X1 U19549 ( .C1(n19327), .C2(n19132), .A(n17645), .B(n17644), .ZN(
        n17649) );
  NOR2_X1 U19550 ( .A1(n17647), .A2(n17646), .ZN(n17648) );
  AOI211_X1 U19551 ( .C1(n19128), .C2(n19329), .A(n17649), .B(n17648), .ZN(
        n17652) );
  NAND2_X1 U19552 ( .A1(n17650), .A2(n19335), .ZN(n17651) );
  OAI211_X1 U19553 ( .C1(n17653), .C2(n19332), .A(n17652), .B(n17651), .ZN(
        P2_U3028) );
  OR2_X1 U19554 ( .A1(n17655), .A2(n17654), .ZN(n17657) );
  OAI21_X1 U19555 ( .B1(n17657), .B2(n17662), .A(n17656), .ZN(n17658) );
  AND2_X1 U19556 ( .A1(n17659), .A2(n17658), .ZN(n19272) );
  INV_X1 U19557 ( .A(n17759), .ZN(n19270) );
  OAI21_X1 U19558 ( .B1(n19271), .B2(n19270), .A(n18011), .ZN(n17660) );
  OAI211_X1 U19559 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n19237), .A(
        n19272), .B(n17660), .ZN(n17661) );
  NAND2_X1 U19560 ( .A1(n17661), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17670) );
  OAI22_X1 U19561 ( .A1(n17673), .A2(n19332), .B1(n17675), .B2(n17662), .ZN(
        n19269) );
  NAND3_X1 U19562 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19269), .A3(
        n17663), .ZN(n17665) );
  OAI211_X1 U19563 ( .C1(n19327), .C2(n17666), .A(n17665), .B(n17664), .ZN(
        n17667) );
  AOI21_X1 U19564 ( .B1(n17668), .B2(n19329), .A(n17667), .ZN(n17669) );
  OAI211_X1 U19565 ( .C1(n17671), .C2(n19304), .A(n17670), .B(n17669), .ZN(
        P2_U3029) );
  NAND3_X1 U19566 ( .A1(n17673), .A2(n19271), .A3(n17672), .ZN(n17682) );
  INV_X1 U19567 ( .A(n19272), .ZN(n17680) );
  NAND2_X1 U19568 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19282), .ZN(n17674) );
  OAI21_X1 U19569 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n17675), .A(
        n17674), .ZN(n17676) );
  AOI21_X1 U19570 ( .B1(n19281), .B2(n19820), .A(n17676), .ZN(n17677) );
  OAI21_X1 U19571 ( .B1(n17678), .B2(n19285), .A(n17677), .ZN(n17679) );
  AOI21_X1 U19572 ( .B1(n17680), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n17679), .ZN(n17681) );
  OAI211_X1 U19573 ( .C1(n17683), .C2(n19304), .A(n17682), .B(n17681), .ZN(
        P2_U3031) );
  NAND2_X1 U19574 ( .A1(n17686), .A2(n17685), .ZN(n17687) );
  XNOR2_X1 U19575 ( .A(n17684), .B(n17687), .ZN(n17981) );
  INV_X1 U19576 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n19246) );
  NAND3_X1 U19577 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n17716), .ZN(n17972) );
  NAND2_X1 U19578 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17971), .ZN(
        n17701) );
  AND2_X1 U19579 ( .A1(n19254), .A2(n17716), .ZN(n17991) );
  AOI21_X1 U19580 ( .B1(n17696), .B2(n17701), .A(n17991), .ZN(n17984) );
  NAND2_X1 U19581 ( .A1(n17984), .A2(n19271), .ZN(n17700) );
  AOI21_X1 U19582 ( .B1(n17690), .B2(n17689), .A(n17688), .ZN(n19823) );
  INV_X1 U19583 ( .A(n19823), .ZN(n17691) );
  INV_X1 U19584 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19090) );
  OAI22_X1 U19585 ( .A1(n19327), .A2(n17691), .B1(n19090), .B2(n19325), .ZN(
        n17698) );
  INV_X1 U19586 ( .A(n19253), .ZN(n17741) );
  NOR3_X1 U19587 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17693), .A3(
        n17741), .ZN(n17708) );
  INV_X1 U19588 ( .A(n17693), .ZN(n17692) );
  OAI21_X1 U19589 ( .B1(n17692), .B2(n19237), .A(n17743), .ZN(n17709) );
  NOR2_X1 U19590 ( .A1(n17708), .A2(n17709), .ZN(n19252) );
  NOR2_X1 U19591 ( .A1(n17693), .A2(n17741), .ZN(n17694) );
  NAND2_X1 U19592 ( .A1(n17694), .A2(n17696), .ZN(n19251) );
  OAI22_X1 U19593 ( .A1(n19252), .A2(n17696), .B1(n17695), .B2(n19251), .ZN(
        n17697) );
  AOI211_X1 U19594 ( .C1(n11273), .C2(n19329), .A(n17698), .B(n17697), .ZN(
        n17699) );
  OAI211_X1 U19595 ( .C1(n17981), .C2(n19304), .A(n17700), .B(n17699), .ZN(
        P2_U3033) );
  OAI21_X1 U19596 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17971), .A(
        n17701), .ZN(n17977) );
  INV_X1 U19597 ( .A(n17703), .ZN(n17705) );
  AND2_X1 U19598 ( .A1(n17705), .A2(n17704), .ZN(n17706) );
  XNOR2_X1 U19599 ( .A(n17702), .B(n17706), .ZN(n17976) );
  INV_X1 U19600 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19080) );
  NOR2_X1 U19601 ( .A1(n19080), .A2(n19325), .ZN(n17707) );
  AOI211_X1 U19602 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17709), .A(
        n17708), .B(n17707), .ZN(n17713) );
  OAI22_X1 U19603 ( .A1(n19285), .A2(n17710), .B1(n19327), .B2(n19089), .ZN(
        n17711) );
  INV_X1 U19604 ( .A(n17711), .ZN(n17712) );
  OAI211_X1 U19605 ( .C1(n17976), .C2(n19304), .A(n17713), .B(n17712), .ZN(
        n17714) );
  INV_X1 U19606 ( .A(n17714), .ZN(n17715) );
  OAI21_X1 U19607 ( .B1(n17977), .B2(n19332), .A(n17715), .ZN(P2_U3034) );
  INV_X1 U19608 ( .A(n17716), .ZN(n17737) );
  NOR2_X1 U19609 ( .A1(n17737), .A2(n17742), .ZN(n17736) );
  OAI21_X1 U19610 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17736), .A(
        n17972), .ZN(n17960) );
  NAND2_X1 U19611 ( .A1(n17717), .A2(n17730), .ZN(n17722) );
  INV_X1 U19612 ( .A(n17718), .ZN(n17720) );
  NOR2_X1 U19613 ( .A1(n17720), .A2(n17719), .ZN(n17721) );
  XNOR2_X1 U19614 ( .A(n17722), .B(n17721), .ZN(n17959) );
  OAI21_X1 U19615 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19237), .A(
        n17743), .ZN(n19244) );
  NOR3_X1 U19616 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17742), .A3(
        n17741), .ZN(n19245) );
  INV_X1 U19617 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19068) );
  NOR2_X1 U19618 ( .A1(n19068), .A2(n19325), .ZN(n17723) );
  AOI211_X1 U19619 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n19244), .A(
        n19245), .B(n17723), .ZN(n17727) );
  OAI22_X1 U19620 ( .A1(n19285), .A2(n17724), .B1(n19327), .B2(n19077), .ZN(
        n17725) );
  INV_X1 U19621 ( .A(n17725), .ZN(n17726) );
  OAI211_X1 U19622 ( .C1(n17959), .C2(n19304), .A(n17727), .B(n17726), .ZN(
        n17728) );
  INV_X1 U19623 ( .A(n17728), .ZN(n17729) );
  OAI21_X1 U19624 ( .B1(n17960), .B2(n19332), .A(n17729), .ZN(P2_U3036) );
  INV_X1 U19625 ( .A(n17730), .ZN(n17732) );
  OR2_X1 U19626 ( .A1(n17717), .A2(n17732), .ZN(n17735) );
  OAI21_X1 U19627 ( .B1(n17733), .B2(n17732), .A(n17731), .ZN(n17734) );
  NAND2_X1 U19628 ( .A1(n17735), .A2(n17734), .ZN(n17953) );
  AOI21_X1 U19629 ( .B1(n17737), .B2(n17742), .A(n17736), .ZN(n17955) );
  NAND2_X1 U19630 ( .A1(n17955), .A2(n19271), .ZN(n17747) );
  NAND2_X1 U19631 ( .A1(n19329), .A2(n17738), .ZN(n17740) );
  NAND2_X1 U19632 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19282), .ZN(n17739) );
  OAI211_X1 U19633 ( .C1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17741), .A(
        n17740), .B(n17739), .ZN(n17745) );
  NOR2_X1 U19634 ( .A1(n17743), .A2(n17742), .ZN(n17744) );
  AOI211_X1 U19635 ( .C1(n19281), .C2(n19826), .A(n17745), .B(n17744), .ZN(
        n17746) );
  OAI211_X1 U19636 ( .C1(n17953), .C2(n19304), .A(n17747), .B(n17746), .ZN(
        P2_U3037) );
  OAI21_X1 U19637 ( .B1(n17750), .B2(n17749), .A(n17748), .ZN(n17947) );
  INV_X1 U19638 ( .A(n17752), .ZN(n17753) );
  NOR2_X1 U19639 ( .A1(n17754), .A2(n17753), .ZN(n17755) );
  XNOR2_X1 U19640 ( .A(n17751), .B(n17755), .ZN(n17946) );
  OAI22_X1 U19641 ( .A1(n19237), .A2(n19296), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17756), .ZN(n17757) );
  NOR2_X1 U19642 ( .A1(n17758), .A2(n17757), .ZN(n19301) );
  OAI21_X1 U19643 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17759), .A(
        n19301), .ZN(n19280) );
  INV_X1 U19644 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n18084) );
  NOR2_X1 U19645 ( .A1(n18084), .A2(n19325), .ZN(n17763) );
  NAND3_X1 U19646 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n19296), .A3(
        n17760), .ZN(n19295) );
  AOI221_X1 U19647 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n17761), .C2(n19294), .A(
        n19295), .ZN(n17762) );
  AOI211_X1 U19648 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n19280), .A(
        n17763), .B(n17762), .ZN(n17767) );
  OAI22_X1 U19649 ( .A1(n19285), .A2(n17764), .B1(n19327), .B2(n19065), .ZN(
        n17765) );
  INV_X1 U19650 ( .A(n17765), .ZN(n17766) );
  OAI211_X1 U19651 ( .C1(n17946), .C2(n19304), .A(n17767), .B(n17766), .ZN(
        n17768) );
  INV_X1 U19652 ( .A(n17768), .ZN(n17769) );
  OAI21_X1 U19653 ( .B1(n17947), .B2(n19332), .A(n17769), .ZN(P2_U3038) );
  AOI221_X1 U19654 ( .B1(n11173), .B2(n19030), .C1(n19193), .C2(n19224), .A(
        n12085), .ZN(n17780) );
  AOI21_X1 U19655 ( .B1(n17770), .B2(n14346), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n17772) );
  INV_X1 U19656 ( .A(n17803), .ZN(n17787) );
  OAI22_X1 U19657 ( .A1(n17780), .A2(n17772), .B1(n17771), .B2(n17787), .ZN(
        n17775) );
  OAI22_X1 U19658 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14346), .B1(n17773), 
        .B2(n19350), .ZN(n17774) );
  AOI21_X1 U19659 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17808), .A(n17774), .ZN(
        n17788) );
  INV_X1 U19660 ( .A(n17788), .ZN(n17822) );
  MUX2_X1 U19661 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n17775), .S(
        n17822), .Z(P2_U3601) );
  INV_X1 U19662 ( .A(n18021), .ZN(n17819) );
  AOI21_X1 U19663 ( .B1(n19193), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n17776), .ZN(n17782) );
  AOI222_X1 U19664 ( .A1(n17777), .A2(n17819), .B1(n17780), .B2(n17782), .C1(
        n19860), .C2(n17803), .ZN(n17779) );
  NAND2_X1 U19665 ( .A1(n17788), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17778) );
  OAI21_X1 U19666 ( .B1(n17779), .B2(n17788), .A(n17778), .ZN(P2_U3600) );
  INV_X1 U19667 ( .A(n17780), .ZN(n17783) );
  OAI222_X1 U19668 ( .A1(n17787), .A2(n20200), .B1(n17783), .B2(n17782), .C1(
        n18021), .C2(n17781), .ZN(n17784) );
  MUX2_X1 U19669 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17784), .S(
        n17822), .Z(P2_U3599) );
  OAI22_X1 U19670 ( .A1(n19876), .A2(n17787), .B1(n17786), .B2(n18021), .ZN(
        n17789) );
  MUX2_X1 U19671 ( .A(n17789), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n17788), .Z(P2_U3596) );
  NOR3_X1 U19672 ( .A1(n20430), .A2(n20432), .A3(n20002), .ZN(n17790) );
  AND2_X1 U19673 ( .A1(n19846), .A2(n22273), .ZN(n19847) );
  NOR2_X1 U19674 ( .A1(n17790), .A2(n19847), .ZN(n17792) );
  NOR2_X1 U19675 ( .A1(n19965), .A2(n20004), .ZN(n20427) );
  NOR2_X1 U19676 ( .A1(n20325), .A2(n20427), .ZN(n17796) );
  OAI21_X1 U19677 ( .B1(n17793), .B2(n20427), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17791) );
  INV_X1 U19678 ( .A(n17792), .ZN(n17797) );
  OAI21_X1 U19679 ( .B1(n19846), .B2(n20427), .A(n19932), .ZN(n17795) );
  INV_X1 U19680 ( .A(n19941), .ZN(n20008) );
  NAND2_X1 U19681 ( .A1(n17793), .A2(n20008), .ZN(n17794) );
  AOI22_X1 U19682 ( .A1(n20188), .A2(n20432), .B1(n20194), .B2(n20427), .ZN(
        n17799) );
  NAND2_X1 U19683 ( .A1(n20195), .A2(n20430), .ZN(n17798) );
  OAI211_X1 U19684 ( .C1(n20438), .C2(n17800), .A(n17799), .B(n17798), .ZN(
        n17801) );
  AOI21_X1 U19685 ( .B1(n16029), .B2(n20433), .A(n17801), .ZN(n17802) );
  INV_X1 U19686 ( .A(n17802), .ZN(P2_U3051) );
  OAI21_X1 U19687 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n17803), .A(n19010), 
        .ZN(n17806) );
  INV_X1 U19688 ( .A(n19345), .ZN(n17804) );
  NOR2_X1 U19689 ( .A1(n17804), .A2(n12026), .ZN(n19349) );
  NAND2_X1 U19690 ( .A1(n22317), .A2(n19349), .ZN(n17805) );
  NAND2_X1 U19691 ( .A1(n17806), .A2(n17805), .ZN(n17812) );
  NOR2_X1 U19692 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n17901), .ZN(n19344) );
  AND2_X1 U19693 ( .A1(n22317), .A2(n19344), .ZN(n17841) );
  AOI211_X1 U19694 ( .C1(n17843), .C2(n17808), .A(n17807), .B(n17841), .ZN(
        n17811) );
  AOI22_X1 U19695 ( .A1(n19345), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19341), 
        .B2(n17809), .ZN(n17810) );
  NAND3_X1 U19696 ( .A1(n17812), .A2(n17811), .A3(n17810), .ZN(P2_U3176) );
  NOR2_X1 U19697 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21937), .ZN(
        n19380) );
  OR2_X1 U19698 ( .A1(n17813), .A2(n18466), .ZN(n18498) );
  INV_X1 U19699 ( .A(n18497), .ZN(n17814) );
  NOR2_X1 U19700 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21937), .ZN(
        n21938) );
  INV_X1 U19701 ( .A(n19591), .ZN(n19716) );
  AOI211_X1 U19702 ( .C1(n17830), .C2(n18498), .A(n19716), .B(n17815), .ZN(
        n18896) );
  NAND2_X1 U19703 ( .A1(n21937), .A2(n18497), .ZN(n18500) );
  INV_X1 U19704 ( .A(n18500), .ZN(n20786) );
  NAND2_X1 U19705 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18758) );
  NAND2_X1 U19706 ( .A1(n20786), .A2(n18758), .ZN(n17817) );
  NOR2_X1 U19707 ( .A1(n19403), .A2(n19383), .ZN(n19411) );
  AOI21_X1 U19708 ( .B1(n21937), .B2(n17817), .A(n19411), .ZN(n17816) );
  NOR3_X1 U19709 ( .A1(n19380), .A2(n18896), .A3(n17816), .ZN(n18895) );
  INV_X1 U19710 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19392) );
  OAI21_X1 U19711 ( .B1(n19392), .B2(n21937), .A(n17817), .ZN(n18898) );
  INV_X1 U19712 ( .A(n18896), .ZN(n18899) );
  OAI221_X1 U19713 ( .B1(n18897), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18897), .C2(n18898), .A(n18899), .ZN(n18893) );
  AOI22_X1 U19714 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18895), .B1(
        n18893), .B2(n19383), .ZN(P3_U2865) );
  NAND3_X1 U19715 ( .A1(n17822), .A2(n17819), .A3(n17818), .ZN(n17820) );
  OAI21_X1 U19716 ( .B1(n17822), .B2(n17821), .A(n17820), .ZN(P2_U3595) );
  INV_X1 U19717 ( .A(n13601), .ZN(n17885) );
  NAND4_X1 U19718 ( .A1(n17884), .A2(n17824), .A3(n17885), .A4(n17823), .ZN(
        n17825) );
  OAI21_X1 U19719 ( .B1(n17826), .B2(n17889), .A(n17825), .ZN(P1_U3468) );
  INV_X1 U19720 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17827) );
  INV_X1 U19721 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n22324) );
  OAI21_X1 U19722 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n22324), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18960) );
  NAND2_X1 U19723 ( .A1(n22333), .A2(n18960), .ZN(n17829) );
  INV_X1 U19724 ( .A(n17829), .ZN(n22281) );
  INV_X1 U19725 ( .A(BS16), .ZN(n17857) );
  NAND2_X1 U19726 ( .A1(n22335), .A2(n22324), .ZN(n22283) );
  AOI21_X1 U19727 ( .B1(n17857), .B2(n22283), .A(n17828), .ZN(n22277) );
  AOI21_X1 U19728 ( .B1(n17827), .B2(n17828), .A(n22277), .ZN(P3_U3280) );
  AND2_X1 U19729 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n17828), .ZN(P3_U3028) );
  AND2_X1 U19730 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n17828), .ZN(P3_U3027) );
  AND2_X1 U19731 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n17828), .ZN(P3_U3026) );
  AND2_X1 U19732 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n17828), .ZN(P3_U3025) );
  AND2_X1 U19733 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n17828), .ZN(P3_U3024) );
  AND2_X1 U19734 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n17828), .ZN(P3_U3023) );
  AND2_X1 U19735 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n17828), .ZN(P3_U3022) );
  AND2_X1 U19736 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n17828), .ZN(P3_U3021) );
  AND2_X1 U19737 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n17828), .ZN(
        P3_U3020) );
  AND2_X1 U19738 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n17828), .ZN(
        P3_U3019) );
  AND2_X1 U19739 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n17828), .ZN(
        P3_U3018) );
  AND2_X1 U19740 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n17828), .ZN(
        P3_U3017) );
  AND2_X1 U19741 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17828), .ZN(
        P3_U3016) );
  AND2_X1 U19742 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17829), .ZN(
        P3_U3015) );
  AND2_X1 U19743 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17829), .ZN(
        P3_U3014) );
  AND2_X1 U19744 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17829), .ZN(
        P3_U3013) );
  AND2_X1 U19745 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17829), .ZN(
        P3_U3012) );
  AND2_X1 U19746 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n17829), .ZN(
        P3_U3011) );
  AND2_X1 U19747 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n17829), .ZN(
        P3_U3010) );
  AND2_X1 U19748 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n17829), .ZN(
        P3_U3009) );
  AND2_X1 U19749 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n17829), .ZN(
        P3_U3008) );
  AND2_X1 U19750 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n17829), .ZN(
        P3_U3007) );
  AND2_X1 U19751 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n17829), .ZN(
        P3_U3006) );
  AND2_X1 U19752 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n17829), .ZN(
        P3_U3005) );
  AND2_X1 U19753 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n17829), .ZN(
        P3_U3004) );
  AND2_X1 U19754 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n17828), .ZN(
        P3_U3003) );
  AND2_X1 U19755 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n17828), .ZN(
        P3_U3002) );
  AND2_X1 U19756 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n17828), .ZN(
        P3_U3001) );
  AND2_X1 U19757 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n17828), .ZN(
        P3_U3000) );
  AND2_X1 U19758 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n17829), .ZN(
        P3_U2999) );
  AOI21_X1 U19759 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17831)
         );
  NOR4_X1 U19760 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21481), .A3(n20846), 
        .A4(n22332), .ZN(n21932) );
  AOI211_X1 U19761 ( .C1(n18758), .C2(n17831), .A(n17830), .B(n21932), .ZN(
        P3_U2998) );
  NOR2_X1 U19762 ( .A1(n17832), .A2(n18899), .ZN(P3_U2867) );
  NOR2_X1 U19763 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21808), .ZN(n18652) );
  INV_X1 U19764 ( .A(n18652), .ZN(n18888) );
  AND2_X1 U19765 ( .A1(n18949), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U19766 ( .A(n17834), .ZN(n20782) );
  AOI21_X1 U19767 ( .B1(n21939), .B2(n21937), .A(n17836), .ZN(n17837) );
  INV_X1 U19768 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n17835) );
  AOI22_X1 U19769 ( .A1(n20782), .A2(n17836), .B1(n17837), .B2(n17835), .ZN(
        P3_U3298) );
  INV_X1 U19770 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18920) );
  NOR2_X1 U19771 ( .A1(n11381), .A2(n20848), .ZN(n20891) );
  AOI21_X1 U19772 ( .B1(n17837), .B2(n18920), .A(n20891), .ZN(P3_U3299) );
  NAND2_X1 U19773 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n22320), .ZN(n22315) );
  OAI21_X1 U19774 ( .B1(n22323), .B2(n22315), .A(n22305), .ZN(n22276) );
  INV_X1 U19775 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17856) );
  NAND2_X1 U19776 ( .A1(n22320), .A2(n22307), .ZN(n17838) );
  AOI21_X1 U19777 ( .B1(n17857), .B2(n17838), .A(n11150), .ZN(n22272) );
  AOI21_X1 U19778 ( .B1(n11151), .B2(n17856), .A(n22272), .ZN(P2_U3591) );
  AND2_X1 U19779 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n11151), .ZN(P2_U3208) );
  AND2_X1 U19780 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n11150), .ZN(P2_U3207) );
  AND2_X1 U19781 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n11151), .ZN(P2_U3206) );
  AND2_X1 U19782 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n11150), .ZN(P2_U3205) );
  AND2_X1 U19783 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n11151), .ZN(P2_U3204) );
  AND2_X1 U19784 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n11150), .ZN(P2_U3203) );
  AND2_X1 U19785 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n11151), .ZN(P2_U3202) );
  AND2_X1 U19786 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n11150), .ZN(P2_U3201) );
  AND2_X1 U19787 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n11150), .ZN(
        P2_U3200) );
  AND2_X1 U19788 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n11151), .ZN(
        P2_U3199) );
  AND2_X1 U19789 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n11150), .ZN(
        P2_U3198) );
  AND2_X1 U19790 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n11151), .ZN(
        P2_U3197) );
  AND2_X1 U19791 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n11150), .ZN(
        P2_U3196) );
  AND2_X1 U19792 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n11151), .ZN(
        P2_U3195) );
  AND2_X1 U19793 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n11150), .ZN(
        P2_U3194) );
  AND2_X1 U19794 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n11151), .ZN(
        P2_U3193) );
  AND2_X1 U19795 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n11150), .ZN(
        P2_U3192) );
  AND2_X1 U19796 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n11151), .ZN(
        P2_U3191) );
  AND2_X1 U19797 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n11151), .ZN(
        P2_U3190) );
  AND2_X1 U19798 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n11150), .ZN(
        P2_U3189) );
  AND2_X1 U19799 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n11151), .ZN(
        P2_U3188) );
  AND2_X1 U19800 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n11150), .ZN(
        P2_U3187) );
  AND2_X1 U19801 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n11150), .ZN(
        P2_U3186) );
  AND2_X1 U19802 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n11151), .ZN(
        P2_U3185) );
  AND2_X1 U19803 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n11150), .ZN(
        P2_U3184) );
  AND2_X1 U19804 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n11151), .ZN(
        P2_U3183) );
  AND2_X1 U19805 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n11150), .ZN(
        P2_U3182) );
  AND2_X1 U19806 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n11151), .ZN(
        P2_U3181) );
  AND2_X1 U19807 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n11150), .ZN(
        P2_U3180) );
  AND2_X1 U19808 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n11151), .ZN(
        P2_U3179) );
  OAI21_X1 U19809 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n17844), .ZN(n17840) );
  AOI211_X1 U19810 ( .C1(n17842), .C2(n22273), .A(n17841), .B(n17840), .ZN(
        P2_U3178) );
  OAI221_X1 U19811 ( .B1(n14073), .B2(n17844), .C1(n17843), .C2(n17844), .A(
        n20259), .ZN(n18032) );
  NOR2_X1 U19812 ( .A1(n17845), .A2(n18032), .ZN(P2_U3047) );
  AND2_X1 U19813 ( .A1(n18068), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U19814 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17849) );
  NOR4_X1 U19815 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17848) );
  NOR4_X1 U19816 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17847) );
  NOR4_X1 U19817 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17846) );
  NAND4_X1 U19818 ( .A1(n17849), .A2(n17848), .A3(n17847), .A4(n17846), .ZN(
        n17855) );
  NOR4_X1 U19819 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17853) );
  AOI211_X1 U19820 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17852) );
  NOR4_X1 U19821 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17851) );
  NOR4_X1 U19822 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17850) );
  NAND4_X1 U19823 ( .A1(n17853), .A2(n17852), .A3(n17851), .A4(n17850), .ZN(
        n17854) );
  NOR2_X1 U19824 ( .A1(n17855), .A2(n17854), .ZN(n18043) );
  INV_X1 U19825 ( .A(n18043), .ZN(n18042) );
  NOR2_X1 U19826 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18042), .ZN(n18036) );
  INV_X1 U19827 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22275) );
  NAND3_X1 U19828 ( .A1(n18037), .A2(n22275), .A3(n17856), .ZN(n18041) );
  INV_X1 U19829 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18103) );
  AOI22_X1 U19830 ( .A1(n18036), .A2(n18041), .B1(n18042), .B2(n18103), .ZN(
        P2_U2821) );
  INV_X1 U19831 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18101) );
  AOI22_X1 U19832 ( .A1(n18036), .A2(n18037), .B1(n18042), .B2(n18101), .ZN(
        P2_U2820) );
  INV_X1 U19833 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17858) );
  NOR2_X1 U19834 ( .A1(n22299), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n22289) );
  NAND2_X1 U19835 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n22302), .ZN(n22778) );
  OAI21_X1 U19836 ( .B1(n22289), .B2(n22302), .A(n22778), .ZN(n17859) );
  INV_X1 U19837 ( .A(n17859), .ZN(n22271) );
  AOI221_X1 U19838 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n17857), .C1(
        P1_STATE_REG_2__SCAN_IN), .C2(n17857), .A(n17860), .ZN(n22267) );
  AOI21_X1 U19839 ( .B1(n17858), .B2(n17860), .A(n22267), .ZN(P1_U3464) );
  AND2_X1 U19840 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n17860), .ZN(P1_U3193) );
  AND2_X1 U19841 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n17860), .ZN(P1_U3192) );
  AND2_X1 U19842 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n17860), .ZN(P1_U3191) );
  AND2_X1 U19843 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n17860), .ZN(P1_U3190) );
  AND2_X1 U19844 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n17860), .ZN(P1_U3189) );
  AND2_X1 U19845 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n17860), .ZN(P1_U3188) );
  AND2_X1 U19846 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n17860), .ZN(P1_U3187) );
  AND2_X1 U19847 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n17860), .ZN(P1_U3186) );
  AND2_X1 U19848 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n17860), .ZN(
        P1_U3185) );
  AND2_X1 U19849 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n17860), .ZN(
        P1_U3184) );
  AND2_X1 U19850 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n17860), .ZN(
        P1_U3183) );
  AND2_X1 U19851 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n17860), .ZN(
        P1_U3182) );
  AND2_X1 U19852 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n17860), .ZN(
        P1_U3181) );
  AND2_X1 U19853 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n17859), .ZN(
        P1_U3180) );
  AND2_X1 U19854 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n17859), .ZN(
        P1_U3179) );
  AND2_X1 U19855 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n17859), .ZN(
        P1_U3178) );
  AND2_X1 U19856 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n17859), .ZN(
        P1_U3177) );
  AND2_X1 U19857 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n17859), .ZN(
        P1_U3176) );
  AND2_X1 U19858 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n17859), .ZN(
        P1_U3175) );
  AND2_X1 U19859 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n17859), .ZN(
        P1_U3174) );
  AND2_X1 U19860 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n17859), .ZN(
        P1_U3173) );
  AND2_X1 U19861 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n17859), .ZN(
        P1_U3172) );
  AND2_X1 U19862 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n17859), .ZN(
        P1_U3171) );
  AND2_X1 U19863 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n17859), .ZN(
        P1_U3170) );
  AND2_X1 U19864 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n17859), .ZN(
        P1_U3169) );
  AND2_X1 U19865 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n17859), .ZN(
        P1_U3168) );
  AND2_X1 U19866 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n17859), .ZN(
        P1_U3167) );
  AND2_X1 U19867 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n17860), .ZN(
        P1_U3166) );
  AND2_X1 U19868 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n17860), .ZN(
        P1_U3165) );
  AND2_X1 U19869 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n17860), .ZN(
        P1_U3164) );
  NOR3_X1 U19870 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22489), .A3(n22248), 
        .ZN(n17864) );
  OR3_X1 U19871 ( .A1(n17862), .A2(n22297), .A3(n17861), .ZN(n17863) );
  OAI21_X1 U19872 ( .B1(n17865), .B2(n17864), .A(n17863), .ZN(n17897) );
  OAI221_X1 U19873 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n22268), .C1(n22256), 
        .C2(n22296), .A(n22489), .ZN(n17896) );
  MUX2_X1 U19874 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17866), .S(
        n17888), .Z(n17893) );
  MUX2_X1 U19875 ( .A(n12757), .B(n17867), .S(n17888), .Z(n17877) );
  INV_X1 U19876 ( .A(n17877), .ZN(n17892) );
  NOR3_X1 U19877 ( .A1(n17869), .A2(n17868), .A3(n22487), .ZN(n17873) );
  OR2_X1 U19878 ( .A1(n17871), .A2(n17870), .ZN(n17872) );
  AOI222_X1 U19879 ( .A1(n17873), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .B1(n17873), .B2(n17872), .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C2(n17872), .ZN(n17874) );
  AOI222_X1 U19880 ( .A1(n17893), .A2(n22408), .B1(n17893), .B2(n17874), .C1(
        n22408), .C2(n17874), .ZN(n17875) );
  OR2_X1 U19881 ( .A1(n17875), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n17876) );
  AOI221_X1 U19882 ( .B1(n17877), .B2(n17876), .C1(n17875), .C2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17891) );
  NAND2_X1 U19883 ( .A1(n17878), .A2(n22246), .ZN(n17882) );
  OR2_X1 U19884 ( .A1(n17880), .A2(n17879), .ZN(n17881) );
  AOI21_X1 U19885 ( .B1(n17883), .B2(n17882), .A(n17881), .ZN(n17887) );
  NAND2_X1 U19886 ( .A1(n17885), .A2(n17884), .ZN(n17886) );
  OAI211_X1 U19887 ( .C1(n17889), .C2(n17888), .A(n17887), .B(n17886), .ZN(
        n17890) );
  AOI211_X1 U19888 ( .C1(n17893), .C2(n17892), .A(n17891), .B(n17890), .ZN(
        n22266) );
  INV_X1 U19889 ( .A(n22266), .ZN(n17894) );
  AOI221_X1 U19890 ( .B1(n22256), .B2(n22250), .C1(n17894), .C2(n22250), .A(
        n17897), .ZN(n22258) );
  NOR2_X1 U19891 ( .A1(n22258), .A2(n22256), .ZN(n22257) );
  OAI211_X1 U19892 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n22248), .A(n22257), 
        .B(n17895), .ZN(n22262) );
  OAI222_X1 U19893 ( .A1(n22250), .A2(n17897), .B1(n22250), .B2(n17896), .C1(
        P1_STATE2_REG_1__SCAN_IN), .C2(n22262), .ZN(P1_U3162) );
  NOR2_X1 U19894 ( .A1(n17899), .A2(n17898), .ZN(P1_U3032) );
  AND2_X1 U19895 ( .A1(n20514), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U19896 ( .A1(n22289), .A2(n22302), .ZN(n17900) );
  INV_X2 U19897 ( .A(n22778), .ZN(n20780) );
  AOI21_X1 U19898 ( .B1(n17900), .B2(n14726), .A(n20780), .ZN(P1_U2802) );
  NOR2_X1 U19899 ( .A1(n17901), .A2(n18021), .ZN(n19343) );
  AOI22_X1 U19900 ( .A1(P2_CODEFETCH_REG_SCAN_IN), .A2(n19013), .B1(n19343), 
        .B2(n19916), .ZN(n17902) );
  INV_X1 U19901 ( .A(n17902), .ZN(P2_U2816) );
  AOI22_X1 U19902 ( .A1(n17904), .A2(n18010), .B1(n18002), .B2(n17903), .ZN(
        n17907) );
  NAND2_X1 U19903 ( .A1(n17905), .A2(n17998), .ZN(n17906) );
  OAI211_X1 U19904 ( .C1(n17908), .C2(n18008), .A(n17907), .B(n17906), .ZN(
        n17909) );
  INV_X1 U19905 ( .A(n17909), .ZN(n17911) );
  OAI211_X1 U19906 ( .C1(n17987), .C2(n12049), .A(n17911), .B(n17910), .ZN(
        P2_U3012) );
  AOI22_X1 U19907 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19282), .B1(n18002), 
        .B2(n17912), .ZN(n17922) );
  OAI21_X1 U19908 ( .B1(n17914), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n17913), .ZN(n17916) );
  XOR2_X1 U19909 ( .A(n17916), .B(n17915), .Z(n19324) );
  OAI21_X1 U19910 ( .B1(n17919), .B2(n17918), .A(n17917), .ZN(n17920) );
  INV_X1 U19911 ( .A(n17920), .ZN(n19336) );
  AOI222_X1 U19912 ( .A1(n19324), .A2(n18010), .B1(n17983), .B2(n19336), .C1(
        n19330), .C2(n17998), .ZN(n17921) );
  OAI211_X1 U19913 ( .C1(n17923), .C2(n17987), .A(n17922), .B(n17921), .ZN(
        P2_U3011) );
  AOI22_X1 U19914 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19282), .B1(n18002), 
        .B2(n17924), .ZN(n17931) );
  INV_X1 U19915 ( .A(n17925), .ZN(n17929) );
  INV_X1 U19916 ( .A(n17926), .ZN(n17927) );
  AOI222_X1 U19917 ( .A1(n17929), .A2(n17983), .B1(n18010), .B2(n17928), .C1(
        n17998), .C2(n17927), .ZN(n17930) );
  OAI211_X1 U19918 ( .C1(n17932), .C2(n17987), .A(n17931), .B(n17930), .ZN(
        P2_U3009) );
  AOI22_X1 U19919 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19282), .B1(n18002), 
        .B2(n17933), .ZN(n17945) );
  OAI21_X1 U19920 ( .B1(n17936), .B2(n17935), .A(n17934), .ZN(n19290) );
  OR2_X1 U19921 ( .A1(n17938), .A2(n17937), .ZN(n17939) );
  AND2_X1 U19922 ( .A1(n17940), .A2(n17939), .ZN(n19288) );
  INV_X1 U19923 ( .A(n19286), .ZN(n17941) );
  AOI22_X1 U19924 ( .A1(n19288), .A2(n17983), .B1(n17998), .B2(n17941), .ZN(
        n17942) );
  OAI21_X1 U19925 ( .B1(n19290), .B2(n17996), .A(n17942), .ZN(n17943) );
  INV_X1 U19926 ( .A(n17943), .ZN(n17944) );
  OAI211_X1 U19927 ( .C1(n16143), .C2(n17987), .A(n17945), .B(n17944), .ZN(
        P2_U3007) );
  AOI22_X1 U19928 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18003), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19282), .ZN(n17950) );
  OAI22_X1 U19929 ( .A1(n17947), .A2(n17996), .B1(n17946), .B2(n18008), .ZN(
        n17948) );
  AOI21_X1 U19930 ( .B1(n17998), .B2(n19061), .A(n17948), .ZN(n17949) );
  OAI211_X1 U19931 ( .C1(n18001), .C2(n19059), .A(n17950), .B(n17949), .ZN(
        P2_U3006) );
  AOI22_X1 U19932 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19282), .B1(n18002), 
        .B2(n17951), .ZN(n17957) );
  OAI22_X1 U19933 ( .A1(n17953), .A2(n18008), .B1(n15057), .B2(n17952), .ZN(
        n17954) );
  AOI21_X1 U19934 ( .B1(n17955), .B2(n18010), .A(n17954), .ZN(n17956) );
  OAI211_X1 U19935 ( .C1(n17958), .C2(n17987), .A(n17957), .B(n17956), .ZN(
        P2_U3005) );
  AOI22_X1 U19936 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18003), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19282), .ZN(n17963) );
  OAI22_X1 U19937 ( .A1(n17960), .A2(n17996), .B1(n17959), .B2(n18008), .ZN(
        n17961) );
  AOI21_X1 U19938 ( .B1(n17998), .B2(n19073), .A(n17961), .ZN(n17962) );
  OAI211_X1 U19939 ( .C1(n18001), .C2(n19071), .A(n17963), .B(n17962), .ZN(
        P2_U3004) );
  AOI22_X1 U19940 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19282), .B1(n18002), 
        .B2(n17964), .ZN(n17975) );
  NAND2_X1 U19941 ( .A1(n17966), .A2(n17965), .ZN(n17970) );
  NAND2_X1 U19942 ( .A1(n11735), .A2(n17968), .ZN(n17969) );
  XNOR2_X1 U19943 ( .A(n17970), .B(n17969), .ZN(n19239) );
  AOI21_X1 U19944 ( .B1(n19246), .B2(n17972), .A(n17971), .ZN(n19243) );
  AOI222_X1 U19945 ( .A1(n19239), .A2(n17983), .B1(n17998), .B2(n17973), .C1(
        n18010), .C2(n19243), .ZN(n17974) );
  OAI211_X1 U19946 ( .C1(n12100), .C2(n17987), .A(n17975), .B(n17974), .ZN(
        P2_U3003) );
  AOI22_X1 U19947 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18003), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19282), .ZN(n17980) );
  OAI22_X1 U19948 ( .A1(n17977), .A2(n17996), .B1(n17976), .B2(n18008), .ZN(
        n17978) );
  AOI21_X1 U19949 ( .B1(n17998), .B2(n19085), .A(n17978), .ZN(n17979) );
  OAI211_X1 U19950 ( .C1(n18001), .C2(n19083), .A(n17980), .B(n17979), .ZN(
        P2_U3002) );
  AOI22_X1 U19951 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19282), .B1(n18002), 
        .B2(n19095), .ZN(n17986) );
  INV_X1 U19952 ( .A(n17981), .ZN(n17982) );
  AOI222_X1 U19953 ( .A1(n17984), .A2(n18010), .B1(n17983), .B2(n17982), .C1(
        n17998), .C2(n11273), .ZN(n17985) );
  OAI211_X1 U19954 ( .C1(n17988), .C2(n17987), .A(n17986), .B(n17985), .ZN(
        P2_U3001) );
  AOI22_X1 U19955 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18003), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19282), .ZN(n18000) );
  INV_X1 U19956 ( .A(n17989), .ZN(n19260) );
  OAI21_X1 U19957 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17991), .A(
        n17990), .ZN(n19264) );
  NAND2_X1 U19958 ( .A1(n17993), .A2(n17992), .ZN(n17994) );
  XNOR2_X1 U19959 ( .A(n17995), .B(n17994), .ZN(n19259) );
  OAI22_X1 U19960 ( .A1(n19264), .A2(n17996), .B1(n18008), .B2(n19259), .ZN(
        n17997) );
  AOI21_X1 U19961 ( .B1(n17998), .B2(n19260), .A(n17997), .ZN(n17999) );
  OAI211_X1 U19962 ( .C1(n18001), .C2(n19105), .A(n18000), .B(n17999), .ZN(
        P2_U3000) );
  AOI22_X1 U19963 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18003), .B1(
        n18002), .B2(n19112), .ZN(n18014) );
  OAI21_X1 U19964 ( .B1(n18006), .B2(n18005), .A(n18004), .ZN(n19266) );
  OAI22_X1 U19965 ( .A1(n19266), .A2(n18008), .B1(n15057), .B2(n18007), .ZN(
        n18009) );
  INV_X1 U19966 ( .A(n18009), .ZN(n18013) );
  OAI211_X1 U19967 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n19274), .A(
        n18011), .B(n18010), .ZN(n18012) );
  NAND2_X1 U19968 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n19282), .ZN(n19277) );
  NAND4_X1 U19969 ( .A1(n18014), .A2(n18013), .A3(n18012), .A4(n19277), .ZN(
        P2_U2998) );
  INV_X1 U19970 ( .A(n18032), .ZN(n18035) );
  INV_X1 U19971 ( .A(n18015), .ZN(n18017) );
  OAI22_X1 U19972 ( .A1(n18018), .A2(n19014), .B1(n18017), .B2(n18016), .ZN(
        n18019) );
  AOI21_X1 U19973 ( .B1(n20000), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n18019), 
        .ZN(n18020) );
  OAI22_X1 U19974 ( .A1(n20000), .A2(n18032), .B1(n18035), .B2(n18020), .ZN(
        P2_U3605) );
  AND2_X1 U19975 ( .A1(n19860), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19836) );
  OAI21_X1 U19976 ( .B1(n19836), .B2(n20002), .A(n18021), .ZN(n18031) );
  NAND2_X1 U19977 ( .A1(n20200), .A2(n19836), .ZN(n19981) );
  INV_X1 U19978 ( .A(n19981), .ZN(n18022) );
  AOI222_X1 U19979 ( .A1(n18031), .A2(n18023), .B1(n14357), .B2(n18022), .C1(
        n20199), .C2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18024) );
  AOI22_X1 U19980 ( .A1(n18035), .A2(n19884), .B1(n18024), .B2(n18032), .ZN(
        P2_U3603) );
  NOR2_X1 U19981 ( .A1(n20002), .A2(n22273), .ZN(n18028) );
  OR2_X1 U19982 ( .A1(n19860), .A2(n18028), .ZN(n18025) );
  AOI22_X1 U19983 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20249), .B1(n18031), 
        .B2(n18025), .ZN(n18026) );
  AOI22_X1 U19984 ( .A1(n18035), .A2(n12216), .B1(n18026), .B2(n18032), .ZN(
        P2_U3604) );
  OAI21_X1 U19985 ( .B1(n18027), .B2(n19952), .A(n19900), .ZN(n18029) );
  AOI222_X1 U19986 ( .A1(n18031), .A2(n19982), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n18030), .C1(n18029), .C2(n18028), .ZN(n18033) );
  AOI22_X1 U19987 ( .A1(n18035), .A2(n18034), .B1(n18033), .B2(n18032), .ZN(
        P2_U3602) );
  NAND2_X1 U19988 ( .A1(n18036), .A2(n22275), .ZN(n18040) );
  OAI21_X1 U19989 ( .B1(n18037), .B2(n17185), .A(n18043), .ZN(n18038) );
  OAI21_X1 U19990 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18043), .A(n18038), 
        .ZN(n18039) );
  OAI221_X1 U19991 ( .B1(n18040), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18040), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18039), .ZN(P2_U2822) );
  INV_X1 U19992 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18106) );
  OAI221_X1 U19993 ( .B1(n18043), .B2(n18106), .C1(n18042), .C2(n18041), .A(
        n18040), .ZN(P2_U2823) );
  INV_X1 U19994 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n18044) );
  AOI22_X1 U19995 ( .A1(n22306), .A2(n18045), .B1(n18044), .B2(n18104), .ZN(
        P2_U3611) );
  INV_X1 U19996 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n18046) );
  AOI22_X1 U19997 ( .A1(n22306), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n18046), 
        .B2(n18104), .ZN(P2_U3608) );
  INV_X1 U19998 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18047) );
  OAI21_X1 U19999 ( .B1(n22323), .B2(n18047), .A(n11150), .ZN(P2_U2815) );
  AOI22_X1 U20000 ( .A1(n19016), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n18049) );
  OAI21_X1 U20001 ( .B1(n18080), .B2(n18050), .A(n18049), .ZN(P2_U2951) );
  INV_X1 U20002 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n18052) );
  AOI22_X1 U20003 ( .A1(n19016), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n18051) );
  OAI21_X1 U20004 ( .B1(n18080), .B2(n18052), .A(n18051), .ZN(P2_U2950) );
  INV_X1 U20005 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n18054) );
  AOI22_X1 U20006 ( .A1(n19016), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n18053) );
  OAI21_X1 U20007 ( .B1(n18080), .B2(n18054), .A(n18053), .ZN(P2_U2949) );
  INV_X1 U20008 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n18056) );
  AOI22_X1 U20009 ( .A1(n19016), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n18055) );
  OAI21_X1 U20010 ( .B1(n18080), .B2(n18056), .A(n18055), .ZN(P2_U2948) );
  INV_X1 U20011 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n18058) );
  AOI22_X1 U20012 ( .A1(n19016), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n18057) );
  OAI21_X1 U20013 ( .B1(n18080), .B2(n18058), .A(n18057), .ZN(P2_U2947) );
  INV_X1 U20014 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n18060) );
  AOI22_X1 U20015 ( .A1(n19016), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n18059) );
  OAI21_X1 U20016 ( .B1(n18080), .B2(n18060), .A(n18059), .ZN(P2_U2946) );
  AOI22_X1 U20017 ( .A1(n19016), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n18061) );
  OAI21_X1 U20018 ( .B1(n18080), .B2(n18062), .A(n18061), .ZN(P2_U2945) );
  INV_X1 U20019 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n18064) );
  AOI22_X1 U20020 ( .A1(n19016), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n18063) );
  OAI21_X1 U20021 ( .B1(n18080), .B2(n18064), .A(n18063), .ZN(P2_U2944) );
  AOI22_X1 U20022 ( .A1(n19016), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n18065) );
  OAI21_X1 U20023 ( .B1(n18080), .B2(n18066), .A(n18065), .ZN(P2_U2943) );
  AOI22_X1 U20024 ( .A1(n19016), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n18067) );
  OAI21_X1 U20025 ( .B1(n18080), .B2(n12269), .A(n18067), .ZN(P2_U2942) );
  AOI22_X1 U20026 ( .A1(n19016), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18069) );
  OAI21_X1 U20027 ( .B1(n18080), .B2(n18070), .A(n18069), .ZN(P2_U2941) );
  AOI22_X1 U20028 ( .A1(n19016), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n18071) );
  OAI21_X1 U20029 ( .B1(n18080), .B2(n18072), .A(n18071), .ZN(P2_U2940) );
  AOI22_X1 U20030 ( .A1(n19016), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18073) );
  OAI21_X1 U20031 ( .B1(n18080), .B2(n18074), .A(n18073), .ZN(P2_U2939) );
  AOI22_X1 U20032 ( .A1(n19016), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18075) );
  OAI21_X1 U20033 ( .B1(n18080), .B2(n12318), .A(n18075), .ZN(P2_U2938) );
  AOI22_X1 U20034 ( .A1(n19016), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18076) );
  OAI21_X1 U20035 ( .B1(n18080), .B2(n18077), .A(n18076), .ZN(P2_U2937) );
  INV_X1 U20036 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U20037 ( .A1(n19016), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18068), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18078) );
  OAI21_X1 U20038 ( .B1(n18080), .B2(n18079), .A(n18078), .ZN(P2_U2936) );
  INV_X1 U20039 ( .A(n22305), .ZN(n18081) );
  AOI22_X1 U20040 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n18104), .B1(n18081), .B2(
        n22320), .ZN(n18082) );
  OAI21_X1 U20041 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n18104), .A(n18082), 
        .ZN(P2_U2817) );
  OAI222_X1 U20042 ( .A1(n18099), .A2(n12054), .B1(n20441), .B2(n22306), .C1(
        n17185), .C2(n18096), .ZN(P2_U3212) );
  INV_X1 U20043 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20443) );
  OAI222_X1 U20044 ( .A1(n18099), .A2(n19326), .B1(n20443), .B2(n22306), .C1(
        n12054), .C2(n18096), .ZN(P2_U3213) );
  INV_X1 U20045 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20445) );
  OAI222_X1 U20046 ( .A1(n18099), .A2(n12076), .B1(n20445), .B2(n22306), .C1(
        n19326), .C2(n18096), .ZN(P2_U3214) );
  INV_X1 U20047 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20447) );
  OAI222_X1 U20048 ( .A1(n18099), .A2(n16130), .B1(n20447), .B2(n22306), .C1(
        n12076), .C2(n18096), .ZN(P2_U3215) );
  INV_X1 U20049 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20449) );
  OAI222_X1 U20050 ( .A1(n18099), .A2(n19302), .B1(n20449), .B2(n22306), .C1(
        n16130), .C2(n18096), .ZN(P2_U3216) );
  INV_X1 U20051 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n18083) );
  INV_X1 U20052 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20451) );
  OAI222_X1 U20053 ( .A1(n18099), .A2(n18083), .B1(n20451), .B2(n22306), .C1(
        n19302), .C2(n18096), .ZN(P2_U3217) );
  INV_X1 U20054 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20453) );
  OAI222_X1 U20055 ( .A1(n18099), .A2(n18084), .B1(n20453), .B2(n22306), .C1(
        n18083), .C2(n18096), .ZN(P2_U3218) );
  INV_X1 U20056 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n18085) );
  INV_X1 U20057 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20455) );
  OAI222_X1 U20058 ( .A1(n18099), .A2(n18085), .B1(n20455), .B2(n22306), .C1(
        n18084), .C2(n18096), .ZN(P2_U3219) );
  INV_X1 U20059 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20457) );
  OAI222_X1 U20060 ( .A1(n18096), .A2(n18085), .B1(n20457), .B2(n22306), .C1(
        n19068), .C2(n18099), .ZN(P2_U3220) );
  INV_X1 U20061 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20459) );
  OAI222_X1 U20062 ( .A1(n18096), .A2(n19068), .B1(n20459), .B2(n22306), .C1(
        n16116), .C2(n18099), .ZN(P2_U3221) );
  INV_X1 U20063 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20461) );
  OAI222_X1 U20064 ( .A1(n18096), .A2(n16116), .B1(n20461), .B2(n22306), .C1(
        n19080), .C2(n18099), .ZN(P2_U3222) );
  INV_X1 U20065 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20463) );
  OAI222_X1 U20066 ( .A1(n18096), .A2(n19080), .B1(n20463), .B2(n22306), .C1(
        n19090), .C2(n18099), .ZN(P2_U3223) );
  INV_X1 U20067 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20465) );
  INV_X1 U20068 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n18086) );
  OAI222_X1 U20069 ( .A1(n18096), .A2(n19090), .B1(n20465), .B2(n22306), .C1(
        n18086), .C2(n18099), .ZN(P2_U3224) );
  INV_X1 U20070 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20467) );
  OAI222_X1 U20071 ( .A1(n18096), .A2(n18086), .B1(n20467), .B2(n22306), .C1(
        n17522), .C2(n18099), .ZN(P2_U3225) );
  INV_X1 U20072 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20469) );
  OAI222_X1 U20073 ( .A1(n18096), .A2(n17522), .B1(n20469), .B2(n22306), .C1(
        n18087), .C2(n18099), .ZN(P2_U3226) );
  INV_X1 U20074 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20471) );
  INV_X1 U20075 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n18088) );
  OAI222_X1 U20076 ( .A1(n18096), .A2(n18087), .B1(n20471), .B2(n22306), .C1(
        n18088), .C2(n18099), .ZN(P2_U3227) );
  INV_X1 U20077 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20473) );
  INV_X1 U20078 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19120) );
  OAI222_X1 U20079 ( .A1(n18096), .A2(n18088), .B1(n20473), .B2(n22306), .C1(
        n19120), .C2(n18099), .ZN(P2_U3228) );
  INV_X1 U20080 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n18089) );
  INV_X1 U20081 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20475) );
  OAI222_X1 U20082 ( .A1(n18099), .A2(n18089), .B1(n20475), .B2(n22306), .C1(
        n19120), .C2(n18096), .ZN(P2_U3229) );
  INV_X1 U20083 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20477) );
  OAI222_X1 U20084 ( .A1(n18096), .A2(n18089), .B1(n20477), .B2(n22306), .C1(
        n19150), .C2(n18099), .ZN(P2_U3230) );
  INV_X1 U20085 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20479) );
  OAI222_X1 U20086 ( .A1(n18099), .A2(n18090), .B1(n20479), .B2(n22306), .C1(
        n19150), .C2(n18096), .ZN(P2_U3231) );
  INV_X1 U20087 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20481) );
  OAI222_X1 U20088 ( .A1(n18099), .A2(n18091), .B1(n20481), .B2(n22306), .C1(
        n18090), .C2(n18096), .ZN(P2_U3232) );
  INV_X1 U20089 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20483) );
  OAI222_X1 U20090 ( .A1(n18099), .A2(n18092), .B1(n20483), .B2(n22306), .C1(
        n18091), .C2(n18096), .ZN(P2_U3233) );
  INV_X1 U20091 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20485) );
  OAI222_X1 U20092 ( .A1(n18099), .A2(n18093), .B1(n20485), .B2(n22306), .C1(
        n18092), .C2(n18096), .ZN(P2_U3234) );
  INV_X1 U20093 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19181) );
  INV_X1 U20094 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20487) );
  OAI222_X1 U20095 ( .A1(n18099), .A2(n19181), .B1(n20487), .B2(n22306), .C1(
        n18093), .C2(n18096), .ZN(P2_U3235) );
  INV_X1 U20096 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20490) );
  OAI222_X1 U20097 ( .A1(n18096), .A2(n19181), .B1(n20490), .B2(n22306), .C1(
        n19198), .C2(n18099), .ZN(P2_U3236) );
  INV_X1 U20098 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20492) );
  OAI222_X1 U20099 ( .A1(n18099), .A2(n18094), .B1(n20492), .B2(n22306), .C1(
        n19198), .C2(n18096), .ZN(P2_U3237) );
  INV_X1 U20100 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20494) );
  OAI222_X1 U20101 ( .A1(n18096), .A2(n18094), .B1(n20494), .B2(n22306), .C1(
        n18095), .C2(n18099), .ZN(P2_U3238) );
  INV_X1 U20102 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19211) );
  INV_X1 U20103 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20496) );
  OAI222_X1 U20104 ( .A1(n18099), .A2(n19211), .B1(n20496), .B2(n22306), .C1(
        n18095), .C2(n18096), .ZN(P2_U3239) );
  INV_X1 U20105 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20498) );
  INV_X1 U20106 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n18097) );
  OAI222_X1 U20107 ( .A1(n18096), .A2(n19211), .B1(n20498), .B2(n22306), .C1(
        n18097), .C2(n18099), .ZN(P2_U3240) );
  INV_X1 U20108 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n18098) );
  INV_X1 U20109 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20501) );
  OAI222_X1 U20110 ( .A1(n18099), .A2(n18098), .B1(n20501), .B2(n22306), .C1(
        n18097), .C2(n18096), .ZN(P2_U3241) );
  INV_X1 U20111 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n18100) );
  AOI22_X1 U20112 ( .A1(n22306), .A2(n18101), .B1(n18100), .B2(n18104), .ZN(
        P2_U3588) );
  INV_X1 U20113 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n18102) );
  AOI22_X1 U20114 ( .A1(n22306), .A2(n18103), .B1(n18102), .B2(n18104), .ZN(
        P2_U3587) );
  MUX2_X1 U20115 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n22306), .Z(P2_U3586) );
  INV_X1 U20116 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n18105) );
  AOI22_X1 U20117 ( .A1(n22306), .A2(n18106), .B1(n18105), .B2(n18104), .ZN(
        P2_U3585) );
  NAND3_X1 U20118 ( .A1(n21438), .A2(n19550), .A3(n18107), .ZN(n18108) );
  NAND3_X1 U20119 ( .A1(n21277), .A2(n20850), .A3(n11381), .ZN(n18490) );
  INV_X1 U20120 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20882) );
  NAND3_X1 U20121 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n18112) );
  NOR2_X1 U20122 ( .A1(n20882), .A2(n18112), .ZN(n18111) );
  NOR2_X1 U20123 ( .A1(n21371), .A2(n18150), .ZN(n18167) );
  NOR2_X1 U20124 ( .A1(n21371), .A2(n18490), .ZN(n18380) );
  AOI22_X1 U20125 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18487), .B1(n18111), .B2(
        n18380), .ZN(n18110) );
  OAI22_X1 U20126 ( .A1(n18167), .A2(n18110), .B1(n18321), .B2(n18487), .ZN(
        P3_U2699) );
  AND2_X1 U20127 ( .A1(n18111), .A2(n18380), .ZN(n18114) );
  INV_X2 U20128 ( .A(n18491), .ZN(n18487) );
  INV_X1 U20129 ( .A(n18380), .ZN(n18493) );
  NOR2_X1 U20130 ( .A1(n18112), .A2(n18493), .ZN(n18116) );
  AOI21_X1 U20131 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18487), .A(n18116), .ZN(
        n18113) );
  INV_X1 U20132 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18214) );
  OAI22_X1 U20133 ( .A1(n18114), .A2(n18113), .B1(n18214), .B2(n18487), .ZN(
        P3_U2700) );
  NAND2_X1 U20134 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18486) );
  INV_X1 U20135 ( .A(n18486), .ZN(n18115) );
  AOI221_X1 U20136 ( .B1(n18115), .B2(n18489), .C1(n21371), .C2(n18489), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n18117) );
  AOI211_X1 U20137 ( .C1(n18491), .C2(n18309), .A(n18117), .B(n18116), .ZN(
        P3_U2701) );
  AOI22_X1 U20138 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18474), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18121) );
  AOI22_X1 U20139 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18120) );
  AOI22_X1 U20140 ( .A1(n18363), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18119) );
  AOI22_X1 U20141 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18118) );
  NAND4_X1 U20142 ( .A1(n18121), .A2(n18120), .A3(n18119), .A4(n18118), .ZN(
        n18127) );
  AOI22_X1 U20143 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12576), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18125) );
  AOI22_X1 U20144 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18124) );
  AOI22_X1 U20145 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18123) );
  AOI22_X1 U20146 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18122) );
  NAND4_X1 U20147 ( .A1(n18125), .A2(n18124), .A3(n18123), .A4(n18122), .ZN(
        n18126) );
  NOR2_X1 U20148 ( .A1(n18127), .A2(n18126), .ZN(n21439) );
  NAND4_X1 U20149 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .A4(P3_EBX_REG_5__SCAN_IN), .ZN(n18148) );
  NOR2_X1 U20150 ( .A1(n18148), .A2(n18150), .ZN(n18250) );
  AND3_X1 U20151 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n18128) );
  AOI22_X1 U20152 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18487), .B1(n18128), .B2(
        n18167), .ZN(n18129) );
  OAI22_X1 U20153 ( .A1(n21439), .A2(n18487), .B1(n18250), .B2(n18129), .ZN(
        P3_U2695) );
  INV_X1 U20154 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20910) );
  NOR2_X1 U20155 ( .A1(n20910), .A2(n18150), .ZN(n18134) );
  NAND2_X1 U20156 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18134), .ZN(n18132) );
  INV_X1 U20157 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20939) );
  OAI21_X1 U20158 ( .B1(n18491), .B2(n20939), .A(n18132), .ZN(n18130) );
  OAI221_X1 U20159 ( .B1(n21438), .B2(n18132), .C1(n18132), .C2(n20939), .A(
        n18130), .ZN(n18131) );
  OAI21_X1 U20160 ( .B1(n18298), .B2(n18487), .A(n18131), .ZN(P3_U2696) );
  OAI211_X1 U20161 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n18134), .A(n18132), .B(
        n18487), .ZN(n18133) );
  OAI21_X1 U20162 ( .B1(n18487), .B2(n18409), .A(n18133), .ZN(P3_U2697) );
  INV_X1 U20163 ( .A(n18134), .ZN(n18136) );
  AOI21_X1 U20164 ( .B1(n20910), .B2(n18150), .A(n18491), .ZN(n18135) );
  AOI22_X1 U20165 ( .A1(n18136), .A2(n18135), .B1(
        P3_INSTQUEUE_REG_0__5__SCAN_IN), .B2(n18491), .ZN(n18137) );
  INV_X1 U20166 ( .A(n18137), .ZN(P3_U2698) );
  AOI22_X1 U20167 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18141) );
  AOI22_X1 U20168 ( .A1(n18363), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18140) );
  AOI22_X1 U20169 ( .A1(n12576), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18139) );
  AOI22_X1 U20170 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18138) );
  NAND4_X1 U20171 ( .A1(n18141), .A2(n18140), .A3(n18139), .A4(n18138), .ZN(
        n18147) );
  AOI22_X1 U20172 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18145) );
  AOI22_X1 U20173 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18144) );
  AOI22_X1 U20174 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18143) );
  AOI22_X1 U20175 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18142) );
  NAND4_X1 U20176 ( .A1(n18145), .A2(n18144), .A3(n18143), .A4(n18142), .ZN(
        n18146) );
  NOR2_X1 U20177 ( .A1(n18147), .A2(n18146), .ZN(n21423) );
  INV_X1 U20178 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n21043) );
  INV_X1 U20179 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20969) );
  NOR2_X1 U20180 ( .A1(n20969), .A2(n18148), .ZN(n18149) );
  NAND4_X1 U20181 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .A4(n18149), .ZN(n18166) );
  NAND3_X1 U20182 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(n18169), .ZN(n18152) );
  OAI21_X1 U20183 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n18165), .A(n18463), .ZN(
        n18151) );
  AOI22_X1 U20184 ( .A1(n18491), .A2(n21423), .B1(n18151), .B2(n18487), .ZN(
        P3_U2687) );
  INV_X1 U20185 ( .A(n18152), .ZN(n18153) );
  OAI21_X1 U20186 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n18153), .A(n18487), .ZN(
        n18164) );
  AOI22_X1 U20187 ( .A1(n18363), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18157) );
  AOI22_X1 U20188 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12576), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18156) );
  AOI22_X1 U20189 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18155) );
  AOI22_X1 U20190 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18154) );
  NAND4_X1 U20191 ( .A1(n18157), .A2(n18156), .A3(n18155), .A4(n18154), .ZN(
        n18163) );
  AOI22_X1 U20192 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18329), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18161) );
  AOI22_X1 U20193 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18160) );
  AOI22_X1 U20194 ( .A1(n12475), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18159) );
  AOI22_X1 U20195 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18158) );
  NAND4_X1 U20196 ( .A1(n18161), .A2(n18160), .A3(n18159), .A4(n18158), .ZN(
        n18162) );
  NOR2_X1 U20197 ( .A1(n18163), .A2(n18162), .ZN(n21434) );
  OAI22_X1 U20198 ( .A1(n18165), .A2(n18164), .B1(n21434), .B2(n18487), .ZN(
        P3_U2688) );
  INV_X1 U20199 ( .A(n18166), .ZN(n18168) );
  NAND2_X1 U20200 ( .A1(n18168), .A2(n18167), .ZN(n18193) );
  NOR2_X1 U20201 ( .A1(n18491), .A2(n18169), .ZN(n18209) );
  AOI22_X1 U20202 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18329), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18181) );
  AOI22_X1 U20203 ( .A1(n18476), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18180) );
  INV_X1 U20204 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18171) );
  AOI22_X1 U20205 ( .A1(n12576), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18170) );
  OAI21_X1 U20206 ( .B1(n18172), .B2(n18171), .A(n18170), .ZN(n18178) );
  AOI22_X1 U20207 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18176) );
  AOI22_X1 U20208 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18474), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18175) );
  AOI22_X1 U20209 ( .A1(n12476), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18174) );
  AOI22_X1 U20210 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18173) );
  NAND4_X1 U20211 ( .A1(n18176), .A2(n18175), .A3(n18174), .A4(n18173), .ZN(
        n18177) );
  AOI211_X1 U20212 ( .C1(n18198), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n18178), .B(n18177), .ZN(n18179) );
  NAND3_X1 U20213 ( .A1(n18181), .A2(n18180), .A3(n18179), .ZN(n21285) );
  AOI22_X1 U20214 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18209), .B1(n18491), 
        .B2(n21285), .ZN(n18182) );
  OAI21_X1 U20215 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n18193), .A(n18182), .ZN(
        P3_U2690) );
  INV_X1 U20216 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n21013) );
  AOI21_X1 U20217 ( .B1(n18380), .B2(n21013), .A(n18209), .ZN(n18197) );
  INV_X1 U20218 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18196) );
  AOI22_X1 U20219 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18192) );
  AOI22_X1 U20220 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18191) );
  AOI22_X1 U20221 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18183) );
  OAI21_X1 U20222 ( .B1(n11205), .B2(n18409), .A(n18183), .ZN(n18189) );
  AOI22_X1 U20223 ( .A1(n18476), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18187) );
  AOI22_X1 U20224 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18186) );
  AOI22_X1 U20225 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18185) );
  AOI22_X1 U20226 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18184) );
  NAND4_X1 U20227 ( .A1(n18187), .A2(n18186), .A3(n18185), .A4(n18184), .ZN(
        n18188) );
  AOI211_X1 U20228 ( .C1(n18466), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n18189), .B(n18188), .ZN(n18190) );
  NAND3_X1 U20229 ( .A1(n18192), .A2(n18191), .A3(n18190), .ZN(n21425) );
  NOR3_X1 U20230 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n21013), .A3(n18193), .ZN(
        n18194) );
  AOI21_X1 U20231 ( .B1(n18491), .B2(n21425), .A(n18194), .ZN(n18195) );
  OAI21_X1 U20232 ( .B1(n18197), .B2(n18196), .A(n18195), .ZN(P3_U2689) );
  AOI22_X1 U20233 ( .A1(n18477), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18202) );
  AOI22_X1 U20234 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18201) );
  AOI22_X1 U20235 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18200) );
  AOI22_X1 U20236 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18199) );
  NAND4_X1 U20237 ( .A1(n18202), .A2(n18201), .A3(n18200), .A4(n18199), .ZN(
        n18208) );
  AOI22_X1 U20238 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18329), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18206) );
  AOI22_X1 U20239 ( .A1(n12576), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18205) );
  AOI22_X1 U20240 ( .A1(n12476), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18204) );
  AOI22_X1 U20241 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18203) );
  NAND4_X1 U20242 ( .A1(n18206), .A2(n18205), .A3(n18204), .A4(n18203), .ZN(
        n18207) );
  NOR2_X1 U20243 ( .A1(n18208), .A2(n18207), .ZN(n21290) );
  NAND2_X1 U20244 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18209), .ZN(n18212) );
  INV_X1 U20245 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n20973) );
  NAND2_X1 U20246 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n18250), .ZN(n18249) );
  NOR2_X1 U20247 ( .A1(n20973), .A2(n18249), .ZN(n18238) );
  INV_X1 U20248 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n18210) );
  NAND4_X1 U20249 ( .A1(n21438), .A2(P3_EBX_REG_11__SCAN_IN), .A3(n18238), 
        .A4(n18210), .ZN(n18211) );
  OAI211_X1 U20250 ( .C1(n21290), .C2(n18487), .A(n18212), .B(n18211), .ZN(
        P3_U2691) );
  AOI22_X1 U20251 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18223) );
  AOI22_X1 U20252 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18319), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18222) );
  AOI22_X1 U20253 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18213) );
  OAI21_X1 U20254 ( .B1(n11205), .B2(n18214), .A(n18213), .ZN(n18220) );
  AOI22_X1 U20255 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18218) );
  AOI22_X1 U20256 ( .A1(n18476), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18217) );
  AOI22_X1 U20257 ( .A1(n18363), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18216) );
  AOI22_X1 U20258 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18215) );
  NAND4_X1 U20259 ( .A1(n18218), .A2(n18217), .A3(n18216), .A4(n18215), .ZN(
        n18219) );
  AOI211_X1 U20260 ( .C1(n18474), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n18220), .B(n18219), .ZN(n18221) );
  NAND3_X1 U20261 ( .A1(n18223), .A2(n18222), .A3(n18221), .ZN(n21293) );
  INV_X1 U20262 ( .A(n21293), .ZN(n18225) );
  XNOR2_X1 U20263 ( .A(P3_EBX_REG_11__SCAN_IN), .B(n18238), .ZN(n18224) );
  AOI22_X1 U20264 ( .A1(n18491), .A2(n18225), .B1(n18224), .B2(n18487), .ZN(
        P3_U2692) );
  AOI22_X1 U20265 ( .A1(n12576), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18229) );
  AOI22_X1 U20266 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18228) );
  AOI22_X1 U20267 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18227) );
  AOI22_X1 U20268 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18226) );
  NAND4_X1 U20269 ( .A1(n18229), .A2(n18228), .A3(n18227), .A4(n18226), .ZN(
        n18235) );
  AOI22_X1 U20270 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18233) );
  AOI22_X1 U20271 ( .A1(n12476), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18232) );
  AOI22_X1 U20272 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18231) );
  AOI22_X1 U20273 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18230) );
  NAND4_X1 U20274 ( .A1(n18233), .A2(n18232), .A3(n18231), .A4(n18230), .ZN(
        n18234) );
  NOR2_X1 U20275 ( .A1(n18235), .A2(n18234), .ZN(n21297) );
  INV_X1 U20276 ( .A(n18249), .ZN(n18236) );
  OAI21_X1 U20277 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18236), .A(n18487), .ZN(
        n18237) );
  OAI22_X1 U20278 ( .A1(n21297), .A2(n18487), .B1(n18238), .B2(n18237), .ZN(
        P3_U2693) );
  AOI22_X1 U20279 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18242) );
  AOI22_X1 U20280 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n18476), .ZN(n18241) );
  AOI22_X1 U20281 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12577), .ZN(n18240) );
  AOI22_X1 U20282 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18469), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n18468), .ZN(n18239) );
  NAND4_X1 U20283 ( .A1(n18242), .A2(n18241), .A3(n18240), .A4(n18239), .ZN(
        n18248) );
  AOI22_X1 U20284 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18474), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n18465), .ZN(n18246) );
  AOI22_X1 U20285 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n12476), .ZN(n18245) );
  AOI22_X1 U20286 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12576), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18244) );
  AOI22_X1 U20287 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18363), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18243) );
  NAND4_X1 U20288 ( .A1(n18246), .A2(n18245), .A3(n18244), .A4(n18243), .ZN(
        n18247) );
  NOR2_X1 U20289 ( .A1(n18248), .A2(n18247), .ZN(n21303) );
  OAI21_X1 U20290 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18250), .A(n18249), .ZN(
        n18251) );
  AOI22_X1 U20291 ( .A1(n18491), .A2(n21303), .B1(n18251), .B2(n18487), .ZN(
        P3_U2694) );
  INV_X1 U20292 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n21233) );
  INV_X1 U20293 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n21102) );
  INV_X1 U20294 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n21072) );
  NAND4_X1 U20295 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n18253)
         );
  NAND4_X1 U20296 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(P3_EBX_REG_26__SCAN_IN), .A4(P3_EBX_REG_25__SCAN_IN), .ZN(n18252)
         );
  NOR2_X1 U20297 ( .A1(n18253), .A2(n18252), .ZN(n18376) );
  INV_X1 U20298 ( .A(n18376), .ZN(n18254) );
  NOR3_X1 U20299 ( .A1(n21233), .A2(n18370), .A3(n18254), .ZN(n18357) );
  NAND2_X1 U20300 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n18357), .ZN(n18356) );
  INV_X1 U20301 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n20854) );
  INV_X1 U20302 ( .A(n18356), .ZN(n18255) );
  OAI33_X1 U20303 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18356), .A3(n21371), 
        .B1(n20854), .B2(n18491), .B3(n18255), .ZN(P3_U2672) );
  AOI22_X1 U20304 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18259) );
  AOI22_X1 U20305 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18258) );
  AOI22_X1 U20306 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18257) );
  AOI22_X1 U20307 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18256) );
  NAND4_X1 U20308 ( .A1(n18259), .A2(n18258), .A3(n18257), .A4(n18256), .ZN(
        n18265) );
  AOI22_X1 U20309 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18263) );
  AOI22_X1 U20310 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18262) );
  AOI22_X1 U20311 ( .A1(n12475), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18261) );
  AOI22_X1 U20312 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18260) );
  NAND4_X1 U20313 ( .A1(n18263), .A2(n18262), .A3(n18261), .A4(n18260), .ZN(
        n18264) );
  NOR2_X1 U20314 ( .A1(n18265), .A2(n18264), .ZN(n18385) );
  AOI22_X1 U20315 ( .A1(n18477), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18269) );
  AOI22_X1 U20316 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18474), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18268) );
  AOI22_X1 U20317 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18267) );
  AOI22_X1 U20318 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18266) );
  NAND4_X1 U20319 ( .A1(n18269), .A2(n18268), .A3(n18267), .A4(n18266), .ZN(
        n18275) );
  AOI22_X1 U20320 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18273) );
  AOI22_X1 U20321 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18272) );
  AOI22_X1 U20322 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18271) );
  AOI22_X1 U20323 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18270) );
  NAND4_X1 U20324 ( .A1(n18273), .A2(n18272), .A3(n18271), .A4(n18270), .ZN(
        n18274) );
  NOR2_X1 U20325 ( .A1(n18275), .A2(n18274), .ZN(n18389) );
  AOI22_X1 U20326 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18279) );
  AOI22_X1 U20327 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18329), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n18416), .ZN(n18278) );
  AOI22_X1 U20328 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18277) );
  AOI22_X1 U20329 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18469), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n12577), .ZN(n18276) );
  NAND4_X1 U20330 ( .A1(n18279), .A2(n18278), .A3(n18277), .A4(n18276), .ZN(
        n18285) );
  AOI22_X1 U20331 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n11158), .ZN(n18283) );
  AOI22_X1 U20332 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18477), .ZN(n18282) );
  AOI22_X1 U20333 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18467), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n18465), .ZN(n18281) );
  AOI22_X1 U20334 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18363), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n18454), .ZN(n18280) );
  NAND4_X1 U20335 ( .A1(n18283), .A2(n18282), .A3(n18281), .A4(n18280), .ZN(
        n18284) );
  NOR2_X1 U20336 ( .A1(n18285), .A2(n18284), .ZN(n18398) );
  AOI22_X1 U20337 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18416), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18296) );
  AOI22_X1 U20338 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18295) );
  AOI22_X1 U20339 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18286) );
  OAI21_X1 U20340 ( .B1(n18322), .B2(n18287), .A(n18286), .ZN(n18293) );
  AOI22_X1 U20341 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18291) );
  AOI22_X1 U20342 ( .A1(n18363), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18290) );
  AOI22_X1 U20343 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18289) );
  AOI22_X1 U20344 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18288) );
  NAND4_X1 U20345 ( .A1(n18291), .A2(n18290), .A3(n18289), .A4(n18288), .ZN(
        n18292) );
  AOI211_X1 U20346 ( .C1(n18439), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n18293), .B(n18292), .ZN(n18294) );
  NAND3_X1 U20347 ( .A1(n18296), .A2(n18295), .A3(n18294), .ZN(n18403) );
  AOI22_X1 U20348 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18307) );
  AOI22_X1 U20349 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18474), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18306) );
  AOI22_X1 U20350 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18297) );
  OAI21_X1 U20351 ( .B1(n11238), .B2(n18298), .A(n18297), .ZN(n18304) );
  AOI22_X1 U20352 ( .A1(n18477), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18302) );
  AOI22_X1 U20353 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18301) );
  AOI22_X1 U20354 ( .A1(n18363), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18300) );
  AOI22_X1 U20355 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18299) );
  NAND4_X1 U20356 ( .A1(n18302), .A2(n18301), .A3(n18300), .A4(n18299), .ZN(
        n18303) );
  AOI211_X1 U20357 ( .C1(n18416), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n18304), .B(n18303), .ZN(n18305) );
  NAND3_X1 U20358 ( .A1(n18307), .A2(n18306), .A3(n18305), .ZN(n18404) );
  NAND2_X1 U20359 ( .A1(n18403), .A2(n18404), .ZN(n18402) );
  NOR2_X1 U20360 ( .A1(n18398), .A2(n18402), .ZN(n18395) );
  AOI22_X1 U20361 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18318) );
  AOI22_X1 U20362 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18317) );
  AOI22_X1 U20363 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18308) );
  OAI21_X1 U20364 ( .B1(n18322), .B2(n18309), .A(n18308), .ZN(n18315) );
  AOI22_X1 U20365 ( .A1(n18363), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18313) );
  AOI22_X1 U20366 ( .A1(n18477), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18312) );
  AOI22_X1 U20367 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18311) );
  AOI22_X1 U20368 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18310) );
  NAND4_X1 U20369 ( .A1(n18313), .A2(n18312), .A3(n18311), .A4(n18310), .ZN(
        n18314) );
  AOI211_X1 U20370 ( .C1(n18466), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n18315), .B(n18314), .ZN(n18316) );
  NAND3_X1 U20371 ( .A1(n18318), .A2(n18317), .A3(n18316), .ZN(n18394) );
  NAND2_X1 U20372 ( .A1(n18395), .A2(n18394), .ZN(n18393) );
  NOR2_X1 U20373 ( .A1(n18389), .A2(n18393), .ZN(n18373) );
  AOI22_X1 U20374 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18332) );
  AOI22_X1 U20375 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18331) );
  AOI22_X1 U20376 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18320) );
  OAI21_X1 U20377 ( .B1(n18322), .B2(n18321), .A(n18320), .ZN(n18328) );
  AOI22_X1 U20378 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18326) );
  AOI22_X1 U20379 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18325) );
  AOI22_X1 U20380 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18324) );
  AOI22_X1 U20381 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18323) );
  NAND4_X1 U20382 ( .A1(n18326), .A2(n18325), .A3(n18324), .A4(n18323), .ZN(
        n18327) );
  AOI211_X1 U20383 ( .C1(n18329), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n18328), .B(n18327), .ZN(n18330) );
  NAND3_X1 U20384 ( .A1(n18332), .A2(n18331), .A3(n18330), .ZN(n18372) );
  NAND2_X1 U20385 ( .A1(n18373), .A2(n18372), .ZN(n18384) );
  NOR2_X1 U20386 ( .A1(n18385), .A2(n18384), .ZN(n18383) );
  INV_X1 U20387 ( .A(n18383), .ZN(n18343) );
  AOI22_X1 U20388 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18336) );
  AOI22_X1 U20389 ( .A1(n12476), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18335) );
  AOI22_X1 U20390 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18334) );
  AOI22_X1 U20391 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18333) );
  NAND4_X1 U20392 ( .A1(n18336), .A2(n18335), .A3(n18334), .A4(n18333), .ZN(
        n18342) );
  AOI22_X1 U20393 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18340) );
  AOI22_X1 U20394 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18339) );
  AOI22_X1 U20395 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18338) );
  AOI22_X1 U20396 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18329), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18337) );
  NAND4_X1 U20397 ( .A1(n18340), .A2(n18339), .A3(n18338), .A4(n18337), .ZN(
        n18341) );
  NOR2_X1 U20398 ( .A1(n18342), .A2(n18341), .ZN(n18375) );
  NOR2_X1 U20399 ( .A1(n18343), .A2(n18375), .ZN(n18355) );
  AOI22_X1 U20400 ( .A1(n12475), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18347) );
  AOI22_X1 U20401 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18477), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18346) );
  AOI22_X1 U20402 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18345) );
  AOI22_X1 U20403 ( .A1(n12476), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18344) );
  NAND4_X1 U20404 ( .A1(n18347), .A2(n18346), .A3(n18345), .A4(n18344), .ZN(
        n18353) );
  AOI22_X1 U20405 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18319), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18351) );
  AOI22_X1 U20406 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18350) );
  AOI22_X1 U20407 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18349) );
  AOI22_X1 U20408 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18348) );
  NAND4_X1 U20409 ( .A1(n18351), .A2(n18350), .A3(n18349), .A4(n18348), .ZN(
        n18352) );
  NOR2_X1 U20410 ( .A1(n18353), .A2(n18352), .ZN(n18354) );
  XOR2_X1 U20411 ( .A(n18355), .B(n18354), .Z(n21383) );
  OAI211_X1 U20412 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n18357), .A(n18356), .B(
        n18487), .ZN(n18358) );
  OAI21_X1 U20413 ( .B1(n21383), .B2(n18487), .A(n18358), .ZN(P3_U2673) );
  AOI22_X1 U20414 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18362) );
  AOI22_X1 U20415 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18361) );
  AOI22_X1 U20416 ( .A1(n18477), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18360) );
  AOI22_X1 U20417 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18359) );
  NAND4_X1 U20418 ( .A1(n18362), .A2(n18361), .A3(n18360), .A4(n18359), .ZN(
        n18369) );
  AOI22_X1 U20419 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18367) );
  AOI22_X1 U20420 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18366) );
  AOI22_X1 U20421 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18329), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18365) );
  AOI22_X1 U20422 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18364) );
  NAND4_X1 U20423 ( .A1(n18367), .A2(n18366), .A3(n18365), .A4(n18364), .ZN(
        n18368) );
  NOR2_X1 U20424 ( .A1(n18369), .A2(n18368), .ZN(n21338) );
  AND2_X1 U20425 ( .A1(n18487), .A2(n18370), .ZN(n18433) );
  INV_X1 U20426 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n21129) );
  AOI22_X1 U20427 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18433), .B1(n18377), 
        .B2(n21129), .ZN(n18371) );
  OAI21_X1 U20428 ( .B1(n21338), .B2(n18487), .A(n18371), .ZN(P3_U2682) );
  INV_X1 U20429 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n21186) );
  INV_X1 U20430 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n21161) );
  NAND2_X1 U20431 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n18406), .ZN(n18392) );
  NAND2_X1 U20432 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n18391), .ZN(n18388) );
  AOI21_X1 U20433 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n18487), .A(n18391), .ZN(
        n18374) );
  OAI21_X1 U20434 ( .B1(n18373), .B2(n18372), .A(n18384), .ZN(n21407) );
  OAI22_X1 U20435 ( .A1(n18378), .A2(n18374), .B1(n18487), .B2(n21407), .ZN(
        P3_U2676) );
  XOR2_X1 U20436 ( .A(n18383), .B(n18375), .Z(n21395) );
  NAND3_X1 U20437 ( .A1(n18377), .A2(n18376), .A3(n21233), .ZN(n18382) );
  NOR2_X1 U20438 ( .A1(n18491), .A2(n18378), .ZN(n18386) );
  INV_X1 U20439 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n18379) );
  OAI221_X1 U20440 ( .B1(n18386), .B2(n18380), .C1(n11159), .C2(n18379), .A(
        P3_EBX_REG_29__SCAN_IN), .ZN(n18381) );
  OAI211_X1 U20441 ( .C1(n18487), .C2(n21395), .A(n18382), .B(n18381), .ZN(
        P3_U2674) );
  AOI21_X1 U20442 ( .B1(n18385), .B2(n18384), .A(n18383), .ZN(n21396) );
  AOI22_X1 U20443 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n11159), .B1(n18491), 
        .B2(n21396), .ZN(n18387) );
  OAI21_X1 U20444 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n18388), .A(n18387), .ZN(
        P3_U2675) );
  AOI21_X1 U20445 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18487), .A(n18397), .ZN(
        n18390) );
  XNOR2_X1 U20446 ( .A(n18389), .B(n18393), .ZN(n21381) );
  OAI22_X1 U20447 ( .A1(n18391), .A2(n18390), .B1(n18487), .B2(n21381), .ZN(
        P3_U2677) );
  INV_X1 U20448 ( .A(n18392), .ZN(n18400) );
  AOI21_X1 U20449 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18487), .A(n18400), .ZN(
        n18396) );
  OAI21_X1 U20450 ( .B1(n18395), .B2(n18394), .A(n18393), .ZN(n21375) );
  OAI22_X1 U20451 ( .A1(n18397), .A2(n18396), .B1(n18487), .B2(n21375), .ZN(
        P3_U2678) );
  AOI21_X1 U20452 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18487), .A(n18406), .ZN(
        n18399) );
  XNOR2_X1 U20453 ( .A(n18398), .B(n18402), .ZN(n21412) );
  OAI22_X1 U20454 ( .A1(n18400), .A2(n18399), .B1(n18487), .B2(n21412), .ZN(
        P3_U2679) );
  INV_X1 U20455 ( .A(n18401), .ZN(n18422) );
  AOI21_X1 U20456 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18487), .A(n18422), .ZN(
        n18405) );
  OAI21_X1 U20457 ( .B1(n18404), .B2(n18403), .A(n18402), .ZN(n21417) );
  OAI22_X1 U20458 ( .A1(n18406), .A2(n18405), .B1(n18487), .B2(n21417), .ZN(
        P3_U2680) );
  AOI21_X1 U20459 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18487), .A(n18407), .ZN(
        n18421) );
  AOI22_X1 U20460 ( .A1(n18198), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18419) );
  AOI22_X1 U20461 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18329), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18418) );
  AOI22_X1 U20462 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18408) );
  OAI21_X1 U20463 ( .B1(n11238), .B2(n18409), .A(n18408), .ZN(n18415) );
  AOI22_X1 U20464 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18413) );
  AOI22_X1 U20465 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18449), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18412) );
  AOI22_X1 U20466 ( .A1(n12476), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12577), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18411) );
  AOI22_X1 U20467 ( .A1(n18468), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18410) );
  NAND4_X1 U20468 ( .A1(n18413), .A2(n18412), .A3(n18411), .A4(n18410), .ZN(
        n18414) );
  AOI211_X1 U20469 ( .C1(n18416), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n18415), .B(n18414), .ZN(n18417) );
  NAND3_X1 U20470 ( .A1(n18419), .A2(n18418), .A3(n18417), .ZN(n21347) );
  INV_X1 U20471 ( .A(n21347), .ZN(n18420) );
  OAI22_X1 U20472 ( .A1(n18422), .A2(n18421), .B1(n18420), .B2(n18487), .ZN(
        P3_U2681) );
  AOI22_X1 U20473 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18426) );
  AOI22_X1 U20474 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18449), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18425) );
  AOI22_X1 U20475 ( .A1(n12609), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18424) );
  AOI22_X1 U20476 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18423) );
  NAND4_X1 U20477 ( .A1(n18426), .A2(n18425), .A3(n18424), .A4(n18423), .ZN(
        n18432) );
  AOI22_X1 U20478 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18430) );
  AOI22_X1 U20479 ( .A1(n18467), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18429) );
  AOI22_X1 U20480 ( .A1(n18475), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18319), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18428) );
  AOI22_X1 U20481 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18427) );
  NAND4_X1 U20482 ( .A1(n18430), .A2(n18429), .A3(n18428), .A4(n18427), .ZN(
        n18431) );
  NOR2_X1 U20483 ( .A1(n18432), .A2(n18431), .ZN(n21344) );
  OAI21_X1 U20484 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18462), .A(n18433), .ZN(
        n18434) );
  OAI21_X1 U20485 ( .B1(n21344), .B2(n18487), .A(n18434), .ZN(P3_U2683) );
  AOI22_X1 U20486 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18474), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18438) );
  AOI22_X1 U20487 ( .A1(n18477), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18437) );
  AOI22_X1 U20488 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18436) );
  AOI22_X1 U20489 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11167), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18435) );
  NAND4_X1 U20490 ( .A1(n18438), .A2(n18437), .A3(n18436), .A4(n18435), .ZN(
        n18445) );
  AOI22_X1 U20491 ( .A1(n12475), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18363), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18443) );
  AOI22_X1 U20492 ( .A1(n11158), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18442) );
  AOI22_X1 U20493 ( .A1(n18475), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18441) );
  AOI22_X1 U20494 ( .A1(n12609), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18440) );
  NAND4_X1 U20495 ( .A1(n18443), .A2(n18442), .A3(n18441), .A4(n18440), .ZN(
        n18444) );
  NOR2_X1 U20496 ( .A1(n18445), .A2(n18444), .ZN(n21363) );
  OAI21_X1 U20497 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n18485), .A(n18447), .ZN(
        n18446) );
  AOI22_X1 U20498 ( .A1(n18491), .A2(n21363), .B1(n18446), .B2(n18487), .ZN(
        P3_U2685) );
  INV_X1 U20499 ( .A(n18447), .ZN(n18448) );
  OAI21_X1 U20500 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18448), .A(n18487), .ZN(
        n18461) );
  AOI22_X1 U20501 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18453) );
  AOI22_X1 U20502 ( .A1(n18319), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18449), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18452) );
  AOI22_X1 U20503 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18468), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18451) );
  AOI22_X1 U20504 ( .A1(n12577), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18469), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18450) );
  NAND4_X1 U20505 ( .A1(n18453), .A2(n18452), .A3(n18451), .A4(n18450), .ZN(
        n18460) );
  AOI22_X1 U20506 ( .A1(n18475), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18467), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18458) );
  AOI22_X1 U20507 ( .A1(n18474), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11158), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18457) );
  AOI22_X1 U20508 ( .A1(n18329), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18454), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18456) );
  AOI22_X1 U20509 ( .A1(n18363), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18465), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18455) );
  NAND4_X1 U20510 ( .A1(n18458), .A2(n18457), .A3(n18456), .A4(n18455), .ZN(
        n18459) );
  NOR2_X1 U20511 ( .A1(n18460), .A2(n18459), .ZN(n21356) );
  OAI22_X1 U20512 ( .A1(n18462), .A2(n18461), .B1(n21356), .B2(n18487), .ZN(
        P3_U2684) );
  INV_X1 U20513 ( .A(n18463), .ZN(n18464) );
  OAI21_X1 U20514 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n18464), .A(n18487), .ZN(
        n18484) );
  AOI22_X1 U20515 ( .A1(n18466), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n18465), .ZN(n18473) );
  AOI22_X1 U20516 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18467), .B1(
        n18319), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18472) );
  AOI22_X1 U20517 ( .A1(n12609), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n18468), .ZN(n18471) );
  AOI22_X1 U20518 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12577), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n18469), .ZN(n18470) );
  NAND4_X1 U20519 ( .A1(n18473), .A2(n18472), .A3(n18471), .A4(n18470), .ZN(
        n18483) );
  AOI22_X1 U20520 ( .A1(n18416), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n12476), .ZN(n18481) );
  AOI22_X1 U20521 ( .A1(n18475), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n18474), .ZN(n18480) );
  AOI22_X1 U20522 ( .A1(n18477), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18476), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18479) );
  AOI22_X1 U20523 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11158), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n18363), .ZN(n18478) );
  NAND4_X1 U20524 ( .A1(n18481), .A2(n18480), .A3(n18479), .A4(n18478), .ZN(
        n18482) );
  NOR2_X1 U20525 ( .A1(n18483), .A2(n18482), .ZN(n21368) );
  OAI22_X1 U20526 ( .A1(n18485), .A2(n18484), .B1(n21368), .B2(n18487), .ZN(
        P3_U2686) );
  OAI21_X1 U20527 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n18486), .ZN(n20861) );
  INV_X1 U20528 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20855) );
  OAI222_X1 U20529 ( .A1(n20861), .A2(n18493), .B1(n20855), .B2(n18489), .C1(
        n18488), .C2(n18487), .ZN(P3_U2702) );
  AOI22_X1 U20530 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18491), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n18490), .ZN(n18492) );
  OAI21_X1 U20531 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18493), .A(n18492), .ZN(
        P3_U2703) );
  NAND2_X1 U20532 ( .A1(n21808), .A2(n21937), .ZN(n18496) );
  OAI21_X1 U20533 ( .B1(n18494), .B2(n20789), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18495) );
  OAI21_X1 U20534 ( .B1(n18496), .B2(n21929), .A(n18495), .ZN(P3_U2634) );
  AOI21_X1 U20535 ( .B1(n21951), .B2(n18498), .A(n18497), .ZN(n21942) );
  OAI21_X1 U20536 ( .B1(n21942), .B2(n19380), .A(n18899), .ZN(n18499) );
  OAI221_X1 U20537 ( .B1(n19392), .B2(n18500), .C1(n19392), .C2(n18899), .A(
        n18499), .ZN(P3_U2863) );
  INV_X1 U20538 ( .A(n18757), .ZN(n21616) );
  INV_X1 U20539 ( .A(n21817), .ZN(n21667) );
  INV_X1 U20540 ( .A(n18518), .ZN(n21655) );
  OAI22_X1 U20541 ( .A1(n21667), .A2(n18892), .B1(n21655), .B2(n18756), .ZN(
        n18547) );
  AOI21_X1 U20542 ( .B1(n18731), .B2(n18511), .A(n18547), .ZN(n18735) );
  INV_X1 U20543 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18516) );
  INV_X1 U20544 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n21086) );
  NAND3_X1 U20545 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20959) );
  NAND2_X1 U20546 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n21020) );
  NAND2_X1 U20547 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18541) );
  NOR2_X1 U20548 ( .A1(n18504), .A2(n20857), .ZN(n18505) );
  INV_X1 U20549 ( .A(n18505), .ZN(n21089) );
  NOR2_X1 U20550 ( .A1(n18521), .A2(n20857), .ZN(n21088) );
  AOI21_X1 U20551 ( .B1(n21086), .B2(n21089), .A(n21088), .ZN(n21093) );
  INV_X1 U20552 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21833) );
  NOR2_X1 U20553 ( .A1(n21868), .A2(n21833), .ZN(n18509) );
  NAND3_X1 U20554 ( .A1(n18503), .A2(n21086), .A3(n18655), .ZN(n18507) );
  INV_X1 U20555 ( .A(n18758), .ZN(n18841) );
  AOI21_X1 U20556 ( .B1(n18841), .B2(n18504), .A(n18840), .ZN(n18739) );
  OAI211_X1 U20557 ( .C1(n18505), .C2(n18888), .A(n18507), .B(n18739), .ZN(
        n18520) );
  INV_X1 U20558 ( .A(n18520), .ZN(n18506) );
  AOI21_X1 U20559 ( .B1(n21086), .B2(n18507), .A(n18506), .ZN(n18508) );
  AOI211_X1 U20560 ( .C1(n11148), .C2(n21093), .A(n18509), .B(n18508), .ZN(
        n18513) );
  AOI21_X1 U20561 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18793), .A(
        n18598), .ZN(n18510) );
  XNOR2_X1 U20562 ( .A(n18510), .B(n18514), .ZN(n21831) );
  NOR2_X1 U20563 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18511), .ZN(
        n21830) );
  AOI22_X1 U20564 ( .A1(n18802), .A2(n21831), .B1(n18731), .B2(n21830), .ZN(
        n18512) );
  OAI211_X1 U20565 ( .C1(n18735), .C2(n18516), .A(n18513), .B(n18512), .ZN(
        P3_U2812) );
  INV_X1 U20566 ( .A(n18514), .ZN(n18584) );
  NOR3_X1 U20567 ( .A1(n21762), .A2(n18516), .A3(n18515), .ZN(n18597) );
  AOI21_X1 U20568 ( .B1(n18598), .B2(n18584), .A(n18597), .ZN(n18517) );
  XNOR2_X1 U20569 ( .A(n18517), .B(n21800), .ZN(n21804) );
  NOR2_X1 U20570 ( .A1(n21510), .A2(n18639), .ZN(n18606) );
  NOR3_X1 U20571 ( .A1(n21510), .A2(n21800), .A3(n18518), .ZN(n21795) );
  NOR3_X1 U20572 ( .A1(n21510), .A2(n21800), .A3(n21817), .ZN(n21793) );
  OAI22_X1 U20573 ( .A1(n21795), .A2(n18756), .B1(n21793), .B2(n18892), .ZN(
        n18607) );
  NOR2_X1 U20574 ( .A1(n18600), .A2(n20857), .ZN(n21116) );
  INV_X1 U20575 ( .A(n21116), .ZN(n18601) );
  OAI21_X1 U20576 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n21088), .A(
        n18601), .ZN(n21099) );
  INV_X1 U20577 ( .A(n18732), .ZN(n18709) );
  AOI22_X1 U20578 ( .A1(n21886), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18520), .ZN(n18523) );
  INV_X1 U20579 ( .A(n18655), .ZN(n18692) );
  OR3_X1 U20580 ( .A1(n18521), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(
        n18692), .ZN(n18522) );
  OAI211_X1 U20581 ( .C1(n21099), .C2(n18709), .A(n18523), .B(n18522), .ZN(
        n18524) );
  AOI221_X1 U20582 ( .B1(n18606), .B2(n21800), .C1(n18607), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n18524), .ZN(n18525) );
  OAI21_X1 U20583 ( .B1(n21804), .B2(n18765), .A(n18525), .ZN(P3_U2811) );
  INV_X1 U20584 ( .A(n18526), .ZN(n18532) );
  NAND2_X1 U20585 ( .A1(n18532), .A2(n18655), .ZN(n18540) );
  NAND2_X1 U20586 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18527) );
  NOR3_X1 U20587 ( .A1(n18528), .A2(n21762), .A3(n18527), .ZN(n18780) );
  NAND2_X1 U20588 ( .A1(n21664), .A2(n18780), .ZN(n18530) );
  NAND3_X1 U20589 ( .A1(n18742), .A2(n18741), .A3(n21661), .ZN(n18529) );
  NAND2_X1 U20590 ( .A1(n18530), .A2(n18529), .ZN(n18531) );
  XOR2_X1 U20591 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18531), .Z(
        n21673) );
  INV_X1 U20592 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n21054) );
  NOR2_X1 U20593 ( .A1(n21868), .A2(n21054), .ZN(n21671) );
  NAND2_X1 U20594 ( .A1(n18532), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18745) );
  OAI21_X1 U20595 ( .B1(n18532), .B2(n18758), .A(n18887), .ZN(n18747) );
  AOI21_X1 U20596 ( .B1(n18652), .B2(n18745), .A(n18747), .ZN(n18545) );
  INV_X1 U20597 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n21051) );
  INV_X1 U20598 ( .A(n18745), .ZN(n18533) );
  NAND2_X1 U20599 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18533), .ZN(
        n21058) );
  OAI21_X1 U20600 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18533), .A(
        n21058), .ZN(n21041) );
  OAI22_X1 U20601 ( .A1(n18545), .A2(n21051), .B1(n18709), .B2(n21041), .ZN(
        n18534) );
  AOI211_X1 U20602 ( .C1(n18802), .C2(n21673), .A(n21671), .B(n18534), .ZN(
        n18537) );
  OAI221_X1 U20603 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n21664), 
        .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18535), .A(n18547), .ZN(
        n18536) );
  OAI211_X1 U20604 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18540), .A(
        n18537), .B(n18536), .ZN(P3_U2815) );
  AOI22_X1 U20605 ( .A1(n18793), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n21844), .B2(n21762), .ZN(n18538) );
  XNOR2_X1 U20606 ( .A(n18539), .B(n18538), .ZN(n21850) );
  INV_X1 U20607 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18544) );
  INV_X1 U20608 ( .A(n18728), .ZN(n21067) );
  NOR2_X1 U20609 ( .A1(n21067), .A2(n20857), .ZN(n18733) );
  AOI21_X1 U20610 ( .B1(n18544), .B2(n21058), .A(n18733), .ZN(n21060) );
  AOI21_X1 U20611 ( .B1(n21051), .B2(n18544), .A(n18540), .ZN(n18542) );
  AOI22_X1 U20612 ( .A1(n21060), .A2(n18732), .B1(n18542), .B2(n18541), .ZN(
        n18543) );
  INV_X1 U20613 ( .A(n21868), .ZN(n21801) );
  NAND2_X1 U20614 ( .A1(n21801), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n21847) );
  OAI211_X1 U20615 ( .C1(n18545), .C2(n18544), .A(n18543), .B(n21847), .ZN(
        n18546) );
  AOI221_X1 U20616 ( .B1(n18731), .B2(n21844), .C1(n18547), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n18546), .ZN(n18548) );
  OAI21_X1 U20617 ( .B1(n18765), .B2(n21850), .A(n18548), .ZN(P3_U2814) );
  NOR2_X1 U20618 ( .A1(n18549), .A2(n20857), .ZN(n18759) );
  NAND2_X1 U20619 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18759), .ZN(
        n21012) );
  OAI21_X1 U20620 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18759), .A(
        n21012), .ZN(n21003) );
  NOR2_X1 U20621 ( .A1(n18692), .A2(n18549), .ZN(n18569) );
  INV_X1 U20622 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n21008) );
  AOI21_X1 U20623 ( .B1(n18841), .B2(n18549), .A(n18840), .ZN(n18550) );
  OAI21_X1 U20624 ( .B1(n18759), .B2(n18888), .A(n18550), .ZN(n18562) );
  INV_X1 U20625 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n21005) );
  NOR2_X1 U20626 ( .A1(n21868), .A2(n21005), .ZN(n18551) );
  AOI221_X1 U20627 ( .B1(n18569), .B2(n21008), .C1(n18562), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18551), .ZN(n18560) );
  INV_X1 U20628 ( .A(n21635), .ZN(n21630) );
  NAND2_X1 U20629 ( .A1(n21762), .A2(n18552), .ZN(n18564) );
  OAI221_X1 U20630 ( .B1(n21762), .B2(n21630), .C1(n21762), .C2(n18553), .A(
        n18564), .ZN(n18554) );
  XNOR2_X1 U20631 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18554), .ZN(
        n21628) );
  NOR2_X1 U20632 ( .A1(n18790), .A2(n21635), .ZN(n18557) );
  INV_X1 U20633 ( .A(n21629), .ZN(n18563) );
  NOR2_X1 U20634 ( .A1(n21511), .A2(n18563), .ZN(n21632) );
  INV_X1 U20635 ( .A(n21632), .ZN(n18555) );
  NAND2_X1 U20636 ( .A1(n18757), .A2(n21629), .ZN(n21634) );
  AOI22_X1 U20637 ( .A1(n18878), .A2(n18555), .B1(n18803), .B2(n21634), .ZN(
        n18567) );
  INV_X1 U20638 ( .A(n18567), .ZN(n18556) );
  MUX2_X1 U20639 ( .A(n18557), .B(n18556), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n18558) );
  AOI21_X1 U20640 ( .B1(n18802), .B2(n21628), .A(n18558), .ZN(n18559) );
  OAI211_X1 U20641 ( .C1(n18709), .C2(n21003), .A(n18560), .B(n18559), .ZN(
        P3_U2818) );
  INV_X1 U20642 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18561) );
  AOI22_X1 U20643 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n11297), .B1(
        n18561), .B2(n21012), .ZN(n21021) );
  AOI22_X1 U20644 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18562), .B1(
        n11148), .B2(n21021), .ZN(n18573) );
  OAI22_X1 U20645 ( .A1(n18793), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n18771), .B2(n18563), .ZN(n18565) );
  NAND2_X1 U20646 ( .A1(n18565), .A2(n18564), .ZN(n18566) );
  XNOR2_X1 U20647 ( .A(n18566), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n21851) );
  NAND2_X1 U20648 ( .A1(n21629), .A2(n12552), .ZN(n21861) );
  OAI22_X1 U20649 ( .A1(n18790), .A2(n21861), .B1(n18567), .B2(n12552), .ZN(
        n18568) );
  AOI21_X1 U20650 ( .B1(n18802), .B2(n21851), .A(n18568), .ZN(n18572) );
  NAND2_X1 U20651 ( .A1(n21886), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18571) );
  OAI211_X1 U20652 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18569), .B(n21020), .ZN(n18570) );
  NAND4_X1 U20653 ( .A1(n18573), .A2(n18572), .A3(n18571), .A4(n18570), .ZN(
        P3_U2817) );
  INV_X1 U20654 ( .A(n18596), .ZN(n18574) );
  AOI21_X1 U20655 ( .B1(n18576), .B2(n18575), .A(n18574), .ZN(n18617) );
  XNOR2_X1 U20656 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18617), .ZN(
        n21686) );
  NOR2_X1 U20657 ( .A1(n18640), .A2(n18639), .ZN(n18582) );
  OAI22_X1 U20658 ( .A1(n21519), .A2(n18892), .B1(n21515), .B2(n18756), .ZN(
        n18593) );
  AOI21_X1 U20659 ( .B1(n18652), .B2(n18601), .A(n18840), .ZN(n18577) );
  OAI21_X1 U20660 ( .B1(n11249), .B2(n18758), .A(n18577), .ZN(n18605) );
  AOI21_X1 U20661 ( .B1(n18684), .B2(n21123), .A(n18605), .ZN(n18589) );
  INV_X1 U20662 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21149) );
  NAND3_X1 U20663 ( .A1(n11249), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18578) );
  NOR2_X1 U20664 ( .A1(n18615), .A2(n20857), .ZN(n18612) );
  AOI21_X1 U20665 ( .B1(n21149), .B2(n18578), .A(n18612), .ZN(n21143) );
  AOI22_X1 U20666 ( .A1(n21886), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n18732), 
        .B2(n21143), .ZN(n18580) );
  INV_X1 U20667 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21132) );
  AND2_X1 U20668 ( .A1(n18655), .A2(n11249), .ZN(n18591) );
  OAI221_X1 U20669 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n21149), .C2(n21132), .A(
        n18591), .ZN(n18579) );
  OAI211_X1 U20670 ( .C1(n18589), .C2(n21149), .A(n18580), .B(n18579), .ZN(
        n18581) );
  AOI221_X1 U20671 ( .B1(n18582), .B2(n21770), .C1(n18593), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18581), .ZN(n18583) );
  OAI21_X1 U20672 ( .B1(n18765), .B2(n21686), .A(n18583), .ZN(P3_U2808) );
  INV_X1 U20673 ( .A(n18592), .ZN(n21523) );
  AOI22_X1 U20674 ( .A1(n21523), .A2(n18597), .B1(n18585), .B2(n18584), .ZN(
        n18587) );
  XNOR2_X1 U20675 ( .A(n18587), .B(n18586), .ZN(n21527) );
  INV_X1 U20676 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n21140) );
  NOR2_X1 U20677 ( .A1(n21868), .A2(n21140), .ZN(n21513) );
  NAND2_X1 U20678 ( .A1(n11249), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18588) );
  XOR2_X1 U20679 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n18588), .Z(
        n21125) );
  OAI22_X1 U20680 ( .A1(n18589), .A2(n21132), .B1(n18709), .B2(n21125), .ZN(
        n18590) );
  AOI211_X1 U20681 ( .C1(n18591), .C2(n21132), .A(n21513), .B(n18590), .ZN(
        n18595) );
  NOR2_X1 U20682 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18592), .ZN(
        n21514) );
  AOI22_X1 U20683 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18593), .B1(
        n18606), .B2(n21514), .ZN(n18594) );
  OAI211_X1 U20684 ( .C1(n21527), .C2(n18765), .A(n18595), .B(n18594), .ZN(
        P3_U2809) );
  OAI221_X1 U20685 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18598), 
        .C1(n21800), .C2(n18597), .A(n18596), .ZN(n18599) );
  XOR2_X1 U20686 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18599), .Z(
        n21814) );
  OAI21_X1 U20687 ( .B1(n18600), .B2(n19549), .A(n21123), .ZN(n18604) );
  AOI22_X1 U20688 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n11249), .B1(
        n21123), .B2(n18601), .ZN(n21118) );
  INV_X1 U20689 ( .A(n21118), .ZN(n18602) );
  AOI21_X1 U20690 ( .B1(n18709), .B2(n18693), .A(n18602), .ZN(n18603) );
  INV_X1 U20691 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n21120) );
  NOR2_X1 U20692 ( .A1(n21868), .A2(n21120), .ZN(n21805) );
  AOI211_X1 U20693 ( .C1(n18605), .C2(n18604), .A(n18603), .B(n21805), .ZN(
        n18609) );
  NOR2_X1 U20694 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21800), .ZN(
        n21807) );
  AOI22_X1 U20695 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18607), .B1(
        n18606), .B2(n21807), .ZN(n18608) );
  OAI211_X1 U20696 ( .C1(n18765), .C2(n21814), .A(n18609), .B(n18608), .ZN(
        P3_U2810) );
  AND2_X1 U20697 ( .A1(n21772), .A2(n18803), .ZN(n18611) );
  AND2_X1 U20698 ( .A1(n21771), .A2(n18878), .ZN(n18610) );
  AOI22_X1 U20699 ( .A1(n21515), .A2(n18611), .B1(n21519), .B2(n18610), .ZN(
        n18623) );
  INV_X1 U20700 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18628) );
  OR2_X1 U20701 ( .A1(n19549), .A2(n18642), .ZN(n18616) );
  OAI211_X1 U20702 ( .C1(n18612), .C2(n18888), .A(n18887), .B(n18616), .ZN(
        n18627) );
  NAND2_X1 U20703 ( .A1(n21886), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n21781) );
  INV_X1 U20704 ( .A(n18612), .ZN(n18613) );
  AOI22_X1 U20705 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18642), .B1(
        n18628), .B2(n18613), .ZN(n21157) );
  OAI21_X1 U20706 ( .B1(n11148), .B2(n18684), .A(n21157), .ZN(n18614) );
  OAI211_X1 U20707 ( .C1(n18616), .C2(n18615), .A(n21781), .B(n18614), .ZN(
        n18621) );
  AOI22_X1 U20708 ( .A1(n18878), .A2(n21771), .B1(n18803), .B2(n21772), .ZN(
        n18641) );
  INV_X1 U20709 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21776) );
  OAI221_X1 U20710 ( .B1(n18618), .B2(n18793), .C1(n18618), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18617), .ZN(n18619) );
  XNOR2_X1 U20711 ( .A(n21776), .B(n18619), .ZN(n21782) );
  OAI22_X1 U20712 ( .A1(n18641), .A2(n21776), .B1(n18765), .B2(n21782), .ZN(
        n18620) );
  AOI211_X1 U20713 ( .C1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n18627), .A(
        n18621), .B(n18620), .ZN(n18622) );
  OAI21_X1 U20714 ( .B1(n18623), .B2(n21770), .A(n18622), .ZN(P3_U2807) );
  XNOR2_X1 U20715 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18624), .ZN(
        n21694) );
  INV_X1 U20716 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n21183) );
  NAND3_X1 U20717 ( .A1(n18642), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18626) );
  INV_X1 U20718 ( .A(n18653), .ZN(n18681) );
  NAND2_X1 U20719 ( .A1(n18681), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18683) );
  INV_X1 U20720 ( .A(n18683), .ZN(n18625) );
  AOI21_X1 U20721 ( .B1(n21183), .B2(n18626), .A(n18625), .ZN(n21180) );
  INV_X1 U20722 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18646) );
  NAND2_X1 U20723 ( .A1(n18642), .A2(n18655), .ZN(n18647) );
  AOI221_X1 U20724 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n21183), .C2(n18646), .A(
        n18647), .ZN(n18630) );
  AOI21_X1 U20725 ( .B1(n18684), .B2(n18628), .A(n18627), .ZN(n18645) );
  INV_X1 U20726 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n21192) );
  OAI22_X1 U20727 ( .A1(n18645), .A2(n21183), .B1(n21868), .B2(n21192), .ZN(
        n18629) );
  AOI211_X1 U20728 ( .C1(n21180), .C2(n11148), .A(n18630), .B(n18629), .ZN(
        n18636) );
  XNOR2_X1 U20729 ( .A(n18631), .B(n21695), .ZN(n21698) );
  OAI21_X1 U20730 ( .B1(n21762), .B2(n18633), .A(n11231), .ZN(n18634) );
  XNOR2_X1 U20731 ( .A(n18634), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n21699) );
  AOI22_X1 U20732 ( .A1(n18803), .A2(n21698), .B1(n18802), .B2(n21699), .ZN(
        n18635) );
  OAI211_X1 U20733 ( .C1(n18892), .C2(n21694), .A(n18636), .B(n18635), .ZN(
        P3_U2805) );
  AOI21_X1 U20734 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18638), .A(
        n18637), .ZN(n21791) );
  INV_X1 U20735 ( .A(n18641), .ZN(n18649) );
  NAND2_X1 U20736 ( .A1(n18642), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18643) );
  XNOR2_X1 U20737 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n18643), .ZN(
        n21168) );
  AOI22_X1 U20738 ( .A1(n21886), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18732), 
        .B2(n21168), .ZN(n18644) );
  OAI221_X1 U20739 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18647), .C1(
        n18646), .C2(n18645), .A(n18644), .ZN(n18648) );
  AOI221_X1 U20740 ( .B1(n18659), .B2(n21690), .C1(n18649), .C2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n18648), .ZN(n18650) );
  OAI21_X1 U20741 ( .B1(n21791), .B2(n18765), .A(n18650), .ZN(P3_U2806) );
  INV_X1 U20742 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n21229) );
  INV_X1 U20743 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n21203) );
  INV_X1 U20744 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n21209) );
  NAND2_X1 U20745 ( .A1(n18651), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18672) );
  NAND2_X1 U20746 ( .A1(n18726), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18718) );
  INV_X1 U20747 ( .A(n18718), .ZN(n18696) );
  AOI21_X1 U20748 ( .B1(n21229), .B2(n18672), .A(n18696), .ZN(n21222) );
  AND3_X1 U20749 ( .A1(n21229), .A2(n18655), .A3(n18651), .ZN(n18658) );
  OAI21_X1 U20750 ( .B1(n18653), .B2(n20857), .A(n18652), .ZN(n18654) );
  OAI211_X1 U20751 ( .C1(n18656), .C2(n18758), .A(n18654), .B(n18887), .ZN(
        n18680) );
  AOI21_X1 U20752 ( .B1(n18684), .B2(n21203), .A(n18680), .ZN(n18678) );
  NAND3_X1 U20753 ( .A1(n18656), .A2(n21209), .A3(n18655), .ZN(n18673) );
  NAND2_X1 U20754 ( .A1(n21886), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n21767) );
  OAI221_X1 U20755 ( .B1(n21229), .B2(n18678), .C1(n21229), .C2(n18673), .A(
        n21767), .ZN(n18657) );
  AOI211_X1 U20756 ( .C1(n11148), .C2(n21222), .A(n18658), .B(n18657), .ZN(
        n18668) );
  AOI22_X1 U20757 ( .A1(n18878), .A2(n21707), .B1(n18803), .B2(n21719), .ZN(
        n18689) );
  NAND2_X1 U20758 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18689), .ZN(
        n18675) );
  OAI211_X1 U20759 ( .C1(n18878), .C2(n18803), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18675), .ZN(n18667) );
  NAND3_X1 U20760 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n18659), .ZN(n18690) );
  NOR2_X1 U20761 ( .A1(n21711), .A2(n18690), .ZN(n18705) );
  INV_X1 U20762 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18660) );
  NAND3_X1 U20763 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18705), .A3(
        n18660), .ZN(n18666) );
  AOI21_X1 U20764 ( .B1(n18793), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18661), .ZN(n21764) );
  NAND2_X1 U20765 ( .A1(n18793), .A2(n18670), .ZN(n18669) );
  NAND2_X1 U20766 ( .A1(n21765), .A2(n18669), .ZN(n18664) );
  NAND2_X1 U20767 ( .A1(n18664), .A2(n21764), .ZN(n21750) );
  OAI211_X1 U20768 ( .C1(n21764), .C2(n18664), .A(n18802), .B(n21750), .ZN(
        n18665) );
  NAND4_X1 U20769 ( .A1(n18668), .A2(n18667), .A3(n18666), .A4(n18665), .ZN(
        P3_U2802) );
  OAI21_X1 U20770 ( .B1(n18793), .B2(n18670), .A(n18669), .ZN(n21727) );
  NOR2_X1 U20771 ( .A1(n18671), .A2(n20857), .ZN(n18682) );
  OAI21_X1 U20772 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18682), .A(
        n18672), .ZN(n21204) );
  NAND2_X1 U20773 ( .A1(n21886), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n21728) );
  OAI211_X1 U20774 ( .C1(n18709), .C2(n21204), .A(n21728), .B(n18673), .ZN(
        n18674) );
  AOI21_X1 U20775 ( .B1(n18802), .B2(n21727), .A(n18674), .ZN(n18677) );
  OAI21_X1 U20776 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18705), .A(
        n18675), .ZN(n18676) );
  OAI211_X1 U20777 ( .C1(n18678), .C2(n21209), .A(n18677), .B(n18676), .ZN(
        P3_U2803) );
  OAI221_X1 U20778 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21762), 
        .C1(n21695), .C2(n18633), .A(n11231), .ZN(n18679) );
  XNOR2_X1 U20779 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n18679), .ZN(
        n21714) );
  INV_X1 U20780 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n21716) );
  OAI221_X1 U20781 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18681), .C1(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .C2(n19715), .A(n18680), .ZN(
        n18686) );
  INV_X1 U20782 ( .A(n18693), .ZN(n18684) );
  AOI21_X1 U20783 ( .B1(n21203), .B2(n18683), .A(n18682), .ZN(n21198) );
  OAI21_X1 U20784 ( .B1(n11148), .B2(n18684), .A(n21198), .ZN(n18685) );
  OAI211_X1 U20785 ( .C1(n21716), .C2(n21868), .A(n18686), .B(n18685), .ZN(
        n18687) );
  AOI21_X1 U20786 ( .B1(n18802), .B2(n21714), .A(n18687), .ZN(n18688) );
  OAI221_X1 U20787 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18690), 
        .C1(n21711), .C2(n18689), .A(n18688), .ZN(P3_U2804) );
  OR2_X1 U20788 ( .A1(n18694), .A2(n18692), .ZN(n18712) );
  XOR2_X1 U20789 ( .A(n18691), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n18697) );
  NOR2_X1 U20790 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18693), .ZN(
        n18724) );
  AOI21_X1 U20791 ( .B1(n19715), .B2(n18694), .A(n18840), .ZN(n18695) );
  OAI21_X1 U20792 ( .B1(n18696), .B2(n18888), .A(n18695), .ZN(n18725) );
  NOR2_X1 U20793 ( .A1(n18724), .A2(n18725), .ZN(n18711) );
  OAI22_X1 U20794 ( .A1(n18712), .A2(n18697), .B1(n18711), .B2(n18691), .ZN(
        n18698) );
  AOI211_X1 U20795 ( .C1(n11463), .C2(n11148), .A(n18699), .B(n18698), .ZN(
        n18703) );
  AOI22_X1 U20796 ( .A1(n18701), .A2(n18803), .B1(n18700), .B2(n18802), .ZN(
        n18702) );
  OAI211_X1 U20797 ( .C1(n18704), .C2(n18892), .A(n18703), .B(n18702), .ZN(
        P3_U2799) );
  NAND2_X1 U20798 ( .A1(n18706), .A2(n18705), .ZN(n18716) );
  NAND2_X1 U20799 ( .A1(n21754), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21730) );
  AOI22_X1 U20800 ( .A1(n18803), .A2(n21730), .B1(n18878), .B2(n21731), .ZN(
        n18723) );
  AOI22_X1 U20801 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21758), .B1(
        n18720), .B2(n12570), .ZN(n18707) );
  XNOR2_X1 U20802 ( .A(n12569), .B(n18707), .ZN(n21743) );
  INV_X1 U20803 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18710) );
  OAI21_X1 U20804 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18717), .A(
        n18708), .ZN(n21258) );
  OAI22_X1 U20805 ( .A1(n18711), .A2(n18710), .B1(n18709), .B2(n21258), .ZN(
        n18714) );
  INV_X1 U20806 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n21261) );
  OAI22_X1 U20807 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18712), .B1(
        n21868), .B2(n21261), .ZN(n18713) );
  AOI211_X1 U20808 ( .C1(n18802), .C2(n21743), .A(n18714), .B(n18713), .ZN(
        n18715) );
  OAI221_X1 U20809 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18716), 
        .C1(n12569), .C2(n18723), .A(n18715), .ZN(P3_U2800) );
  INV_X1 U20810 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n21230) );
  INV_X1 U20811 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n18719) );
  AOI21_X1 U20812 ( .B1(n18719), .B2(n18718), .A(n18717), .ZN(n21239) );
  AOI211_X1 U20813 ( .C1(n21753), .C2(n18878), .A(n21754), .B(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n18722) );
  NAND2_X1 U20814 ( .A1(n18720), .A2(n21758), .ZN(n18721) );
  OAI221_X1 U20815 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18726), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n19715), .A(n18725), .ZN(
        n18727) );
  AOI21_X1 U20816 ( .B1(n18728), .B2(n19715), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18740) );
  OAI21_X1 U20817 ( .B1(n18730), .B2(n21837), .A(n18729), .ZN(n21835) );
  AOI21_X1 U20818 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18731), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18734) );
  NOR2_X2 U20819 ( .A1(n18684), .A2(n18732), .ZN(n18885) );
  OAI21_X1 U20820 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18733), .A(
        n21089), .ZN(n21069) );
  OAI22_X1 U20821 ( .A1(n18735), .A2(n18734), .B1(n18885), .B2(n21069), .ZN(
        n18736) );
  AOI21_X1 U20822 ( .B1(n18802), .B2(n21835), .A(n18736), .ZN(n18738) );
  NAND2_X1 U20823 ( .A1(n21886), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18737) );
  OAI211_X1 U20824 ( .C1(n18740), .C2(n18739), .A(n18738), .B(n18737), .ZN(
        P3_U2813) );
  INV_X1 U20825 ( .A(n18780), .ZN(n18769) );
  NAND2_X1 U20826 ( .A1(n18742), .A2(n18741), .ZN(n18743) );
  OAI21_X1 U20827 ( .B1(n18769), .B2(n21645), .A(n18743), .ZN(n18744) );
  XNOR2_X1 U20828 ( .A(n18744), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n21654) );
  AND2_X1 U20829 ( .A1(n11297), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18746) );
  OAI21_X1 U20830 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18746), .A(
        n18745), .ZN(n21026) );
  OAI221_X1 U20831 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n11297), .C1(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n19715), .A(n18747), .ZN(
        n18748) );
  OAI21_X1 U20832 ( .B1(n18885), .B2(n21026), .A(n18748), .ZN(n18749) );
  AOI21_X1 U20833 ( .B1(n21886), .B2(P3_REIP_REG_14__SCAN_IN), .A(n18749), 
        .ZN(n18753) );
  AOI21_X1 U20834 ( .B1(n21661), .B2(n18750), .A(n21657), .ZN(n21650) );
  AOI21_X1 U20835 ( .B1(n21661), .B2(n18751), .A(n21658), .ZN(n21647) );
  AOI22_X1 U20836 ( .A1(n18878), .A2(n21650), .B1(n18803), .B2(n21647), .ZN(
        n18752) );
  OAI211_X1 U20837 ( .C1(n21654), .C2(n18765), .A(n18753), .B(n18752), .ZN(
        P3_U2816) );
  NOR2_X1 U20838 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18754), .ZN(
        n18781) );
  AOI22_X1 U20839 ( .A1(n21621), .A2(n18780), .B1(n18773), .B2(n18781), .ZN(
        n18755) );
  XNOR2_X1 U20840 ( .A(n18755), .B(n21852), .ZN(n21627) );
  OAI22_X1 U20841 ( .A1(n18757), .A2(n18756), .B1(n18892), .B2(n21617), .ZN(
        n18779) );
  INV_X1 U20842 ( .A(n21621), .ZN(n21622) );
  AOI211_X1 U20843 ( .C1(n21622), .C2(n21852), .A(n18790), .B(n21630), .ZN(
        n18763) );
  NOR2_X1 U20844 ( .A1(n18766), .A2(n19549), .ZN(n18785) );
  NAND2_X1 U20845 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18785), .ZN(
        n18774) );
  NAND2_X1 U20846 ( .A1(n18887), .A2(n18758), .ZN(n18881) );
  NAND3_X1 U20847 ( .A1(n18881), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n18774), .ZN(n18761) );
  NAND2_X1 U20848 ( .A1(n20985), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18767) );
  AOI21_X1 U20849 ( .B1(n11470), .B2(n18767), .A(n18759), .ZN(n20989) );
  AOI22_X1 U20850 ( .A1(n21886), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n20989), 
        .B2(n18873), .ZN(n18760) );
  OAI211_X1 U20851 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n18774), .A(
        n18761), .B(n18760), .ZN(n18762) );
  AOI211_X1 U20852 ( .C1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n18779), .A(
        n18763), .B(n18762), .ZN(n18764) );
  OAI21_X1 U20853 ( .B1(n21627), .B2(n18765), .A(n18764), .ZN(P3_U2819) );
  OR2_X1 U20854 ( .A1(n18766), .A2(n20857), .ZN(n18783) );
  INV_X1 U20855 ( .A(n18767), .ZN(n18768) );
  AOI21_X1 U20856 ( .B1(n20974), .B2(n18783), .A(n18768), .ZN(n20968) );
  AOI22_X1 U20857 ( .A1(n21886), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n20968), 
        .B2(n18873), .ZN(n18778) );
  AOI221_X1 U20858 ( .B1(n18793), .B2(n18769), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18769), .A(n21862), .ZN(
        n18772) );
  AOI221_X1 U20859 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18780), .C1(
        n21889), .C2(n18781), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18770) );
  AOI221_X1 U20860 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18772), .C1(
        n18771), .C2(n18772), .A(n18770), .ZN(n21863) );
  AOI22_X1 U20861 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18779), .B1(
        n18802), .B2(n21863), .ZN(n18777) );
  OR3_X1 U20862 ( .A1(n21621), .A2(n18773), .A3(n18790), .ZN(n18776) );
  OAI211_X1 U20863 ( .C1(n18785), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18881), .B(n18774), .ZN(n18775) );
  NAND4_X1 U20864 ( .A1(n18778), .A2(n18777), .A3(n18776), .A4(n18775), .ZN(
        P3_U2820) );
  INV_X1 U20865 ( .A(n18779), .ZN(n18789) );
  NOR2_X1 U20866 ( .A1(n18781), .A2(n18780), .ZN(n18782) );
  XNOR2_X1 U20867 ( .A(n18782), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n21884) );
  INV_X1 U20868 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20954) );
  NOR2_X1 U20869 ( .A1(n21868), .A2(n20954), .ZN(n18787) );
  INV_X1 U20870 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18800) );
  INV_X1 U20871 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18814) );
  NOR2_X1 U20872 ( .A1(n18800), .A2(n18814), .ZN(n18796) );
  NOR3_X1 U20873 ( .A1(n18824), .A2(n20922), .A3(n19549), .ZN(n18806) );
  AOI22_X1 U20874 ( .A1(n18796), .A2(n18806), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18881), .ZN(n18784) );
  NAND3_X1 U20875 ( .A1(n18795), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20940) );
  NOR2_X1 U20876 ( .A1(n18800), .A2(n20940), .ZN(n20962) );
  OAI21_X1 U20877 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n20962), .A(
        n18783), .ZN(n20957) );
  OAI22_X1 U20878 ( .A1(n18785), .A2(n18784), .B1(n18885), .B2(n20957), .ZN(
        n18786) );
  AOI211_X1 U20879 ( .C1(n18802), .C2(n21884), .A(n18787), .B(n18786), .ZN(
        n18788) );
  OAI221_X1 U20880 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18790), .C1(
        n21889), .C2(n18789), .A(n18788), .ZN(P3_U2821) );
  OAI21_X1 U20881 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18792), .A(
        n18791), .ZN(n21604) );
  AOI22_X1 U20882 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18793), .B1(
        n21762), .B2(n21600), .ZN(n18794) );
  XNOR2_X1 U20883 ( .A(n11224), .B(n18794), .ZN(n21606) );
  INV_X1 U20884 ( .A(n21606), .ZN(n21607) );
  INV_X1 U20885 ( .A(n18795), .ZN(n18805) );
  AOI21_X1 U20886 ( .B1(n18841), .B2(n18805), .A(n18840), .ZN(n18813) );
  AOI21_X1 U20887 ( .B1(n18800), .B2(n20940), .A(n20962), .ZN(n20942) );
  NAND2_X1 U20888 ( .A1(n18795), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18797) );
  AOI211_X1 U20889 ( .C1(n18800), .C2(n18797), .A(n18796), .B(n19549), .ZN(
        n18798) );
  AOI21_X1 U20890 ( .B1(n20942), .B2(n18873), .A(n18798), .ZN(n18799) );
  NAND2_X1 U20891 ( .A1(n21886), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n21608) );
  OAI211_X1 U20892 ( .C1(n18800), .C2(n18813), .A(n18799), .B(n21608), .ZN(
        n18801) );
  AOI221_X1 U20893 ( .B1(n18803), .B2(n21606), .C1(n18802), .C2(n21607), .A(
        n18801), .ZN(n18804) );
  OAI21_X1 U20894 ( .B1(n18892), .B2(n21604), .A(n18804), .ZN(P3_U2822) );
  NOR2_X1 U20895 ( .A1(n18805), .A2(n20857), .ZN(n20917) );
  OAI21_X1 U20896 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20917), .A(
        n20940), .ZN(n20927) );
  AOI22_X1 U20897 ( .A1(n21886), .A2(P3_REIP_REG_7__SCAN_IN), .B1(n18806), 
        .B2(n18814), .ZN(n18817) );
  INV_X1 U20898 ( .A(n18891), .ZN(n18882) );
  AOI21_X1 U20899 ( .B1(n21589), .B2(n18808), .A(n18807), .ZN(n21592) );
  OAI21_X1 U20900 ( .B1(n18811), .B2(n18810), .A(n18809), .ZN(n18812) );
  XNOR2_X1 U20901 ( .A(n18812), .B(n21589), .ZN(n21587) );
  OAI22_X1 U20902 ( .A1(n18892), .A2(n21587), .B1(n18814), .B2(n18813), .ZN(
        n18815) );
  AOI21_X1 U20903 ( .B1(n18882), .B2(n21592), .A(n18815), .ZN(n18816) );
  OAI211_X1 U20904 ( .C1(n18885), .C2(n20927), .A(n18817), .B(n18816), .ZN(
        P3_U2823) );
  INV_X1 U20905 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20929) );
  AOI21_X1 U20906 ( .B1(n18820), .B2(n18819), .A(n18818), .ZN(n21582) );
  NOR2_X1 U20907 ( .A1(n18824), .A2(n19549), .ZN(n18821) );
  AOI22_X1 U20908 ( .A1(n18882), .A2(n21582), .B1(n18821), .B2(n20922), .ZN(
        n18827) );
  OR2_X1 U20909 ( .A1(n18824), .A2(n20857), .ZN(n18834) );
  AOI21_X1 U20910 ( .B1(n20922), .B2(n18834), .A(n20917), .ZN(n20921) );
  OAI21_X1 U20911 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18823), .A(
        n18822), .ZN(n21585) );
  OAI21_X1 U20912 ( .B1(n19549), .B2(n18824), .A(n18881), .ZN(n18836) );
  OAI22_X1 U20913 ( .A1(n18892), .A2(n21585), .B1(n20922), .B2(n18836), .ZN(
        n18825) );
  AOI21_X1 U20914 ( .B1(n20921), .B2(n18873), .A(n18825), .ZN(n18826) );
  OAI211_X1 U20915 ( .C1(n21868), .C2(n20929), .A(n18827), .B(n18826), .ZN(
        P3_U2824) );
  OAI21_X1 U20916 ( .B1(n18830), .B2(n18829), .A(n18828), .ZN(n21577) );
  AOI21_X1 U20917 ( .B1(n18833), .B2(n18832), .A(n18831), .ZN(n21574) );
  AND2_X1 U20918 ( .A1(n18835), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20905) );
  OAI21_X1 U20919 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20905), .A(
        n18834), .ZN(n20906) );
  AOI21_X1 U20920 ( .B1(n18835), .B2(n18887), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18837) );
  OAI22_X1 U20921 ( .A1(n18885), .A2(n20906), .B1(n18837), .B2(n18836), .ZN(
        n18838) );
  AOI21_X1 U20922 ( .B1(n18882), .B2(n21574), .A(n18838), .ZN(n18839) );
  NAND2_X1 U20923 ( .A1(n21886), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n21575) );
  OAI211_X1 U20924 ( .C1(n18892), .C2(n21577), .A(n18839), .B(n21575), .ZN(
        P3_U2825) );
  AOI21_X1 U20925 ( .B1(n18841), .B2(n18851), .A(n18840), .ZN(n18863) );
  NOR3_X1 U20926 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18851), .A3(
        n19549), .ZN(n18842) );
  AOI21_X1 U20927 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n21886), .A(n18842), .ZN(
        n18853) );
  AOI21_X1 U20928 ( .B1(n18844), .B2(n11293), .A(n18843), .ZN(n18845) );
  NAND2_X1 U20929 ( .A1(n21895), .A2(n18845), .ZN(n18850) );
  OAI211_X1 U20930 ( .C1(n18848), .C2(n18847), .A(n21898), .B(n18846), .ZN(
        n18849) );
  NAND2_X1 U20931 ( .A1(n18850), .A2(n18849), .ZN(n21567) );
  OR2_X1 U20932 ( .A1(n18851), .A2(n20857), .ZN(n18857) );
  AOI21_X1 U20933 ( .B1(n20890), .B2(n18857), .A(n20905), .ZN(n20889) );
  AOI22_X1 U20934 ( .A1(n18871), .A2(n21567), .B1(n20889), .B2(n18873), .ZN(
        n18852) );
  OAI211_X1 U20935 ( .C1(n20890), .C2(n18863), .A(n18853), .B(n18852), .ZN(
        P3_U2826) );
  INV_X1 U20936 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20886) );
  NAND2_X1 U20937 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18887), .ZN(
        n18874) );
  AOI21_X1 U20938 ( .B1(n18856), .B2(n18855), .A(n18854), .ZN(n21556) );
  INV_X1 U20939 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20876) );
  NOR2_X1 U20940 ( .A1(n21868), .A2(n20876), .ZN(n21561) );
  INV_X1 U20941 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20862) );
  NOR2_X1 U20942 ( .A1(n20862), .A2(n20857), .ZN(n18872) );
  OAI21_X1 U20943 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18872), .A(
        n18857), .ZN(n20874) );
  OAI21_X1 U20944 ( .B1(n18860), .B2(n18859), .A(n18858), .ZN(n21557) );
  OAI22_X1 U20945 ( .A1(n18885), .A2(n20874), .B1(n18892), .B2(n21557), .ZN(
        n18861) );
  AOI211_X1 U20946 ( .C1(n18882), .C2(n21556), .A(n21561), .B(n18861), .ZN(
        n18862) );
  OAI221_X1 U20947 ( .B1(n18863), .B2(n20886), .C1(n18863), .C2(n18874), .A(
        n18862), .ZN(P3_U2827) );
  AOI21_X1 U20948 ( .B1(n18866), .B2(n18865), .A(n18864), .ZN(n18870) );
  XOR2_X1 U20949 ( .A(n18868), .B(n18867), .Z(n18869) );
  AOI22_X1 U20950 ( .A1(n21895), .A2(n18870), .B1(n21898), .B2(n18869), .ZN(
        n21544) );
  AOI21_X1 U20951 ( .B1(n20862), .B2(n20857), .A(n18872), .ZN(n20869) );
  AOI22_X1 U20952 ( .A1(n21886), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n20869), 
        .B2(n18873), .ZN(n18876) );
  OAI21_X1 U20953 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19715), .A(
        n18874), .ZN(n18875) );
  OAI211_X1 U20954 ( .C1(n21544), .C2(n11548), .A(n18876), .B(n18875), .ZN(
        P3_U2828) );
  NOR2_X1 U20955 ( .A1(n11152), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18877) );
  XNOR2_X1 U20956 ( .A(n18877), .B(n18880), .ZN(n21537) );
  AOI22_X1 U20957 ( .A1(n21886), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18878), 
        .B2(n21537), .ZN(n18884) );
  AOI21_X1 U20958 ( .B1(n18880), .B2(n18886), .A(n18879), .ZN(n21538) );
  AOI22_X1 U20959 ( .A1(n18882), .A2(n21538), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18881), .ZN(n18883) );
  OAI211_X1 U20960 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n18885), .A(
        n18884), .B(n18883), .ZN(P3_U2829) );
  OAI21_X1 U20961 ( .B1(n11152), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18886), .ZN(n21531) );
  INV_X1 U20962 ( .A(n21531), .ZN(n21530) );
  NAND3_X1 U20963 ( .A1(n21481), .A2(n18888), .A3(n18887), .ZN(n18889) );
  AOI22_X1 U20964 ( .A1(n21886), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18889), .ZN(n18890) );
  OAI221_X1 U20965 ( .B1(n21530), .B2(n18892), .C1(n21531), .C2(n18891), .A(
        n18890), .ZN(P3_U2830) );
  INV_X1 U20966 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21916) );
  NOR2_X1 U20967 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n21916), .ZN(
        n19414) );
  NOR2_X1 U20968 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19383), .ZN(
        n19433) );
  NOR2_X1 U20969 ( .A1(n19414), .A2(n19433), .ZN(n18894) );
  OAI22_X1 U20970 ( .A1(n18895), .A2(n21916), .B1(n18894), .B2(n18893), .ZN(
        P3_U2866) );
  NOR2_X1 U20971 ( .A1(n19380), .A2(n18896), .ZN(n18901) );
  INV_X1 U20972 ( .A(n18897), .ZN(n19428) );
  NAND3_X1 U20973 ( .A1(n19403), .A2(n18899), .A3(n18898), .ZN(n18900) );
  OAI221_X1 U20974 ( .B1(n19403), .B2(n18901), .C1(n19403), .C2(n19428), .A(
        n18900), .ZN(P3_U2864) );
  NOR4_X1 U20975 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18905) );
  NOR4_X1 U20976 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18904) );
  NOR4_X1 U20977 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18903) );
  NOR4_X1 U20978 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18902) );
  NAND4_X1 U20979 ( .A1(n18905), .A2(n18904), .A3(n18903), .A4(n18902), .ZN(
        n18911) );
  NOR4_X1 U20980 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18909) );
  AOI211_X1 U20981 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18908) );
  NOR4_X1 U20982 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18907) );
  NOR4_X1 U20983 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18906) );
  NAND4_X1 U20984 ( .A1(n18909), .A2(n18908), .A3(n18907), .A4(n18906), .ZN(
        n18910) );
  NOR2_X1 U20985 ( .A1(n18911), .A2(n18910), .ZN(n18919) );
  INV_X1 U20986 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18998) );
  OAI21_X1 U20987 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18919), .ZN(n18912) );
  OAI21_X1 U20988 ( .B1(n18919), .B2(n18998), .A(n18912), .ZN(P3_U3293) );
  INV_X1 U20989 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19002) );
  AOI21_X1 U20990 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18913) );
  INV_X1 U20991 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18963) );
  OAI221_X1 U20992 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18913), .C1(n18963), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18919), .ZN(n18914) );
  OAI21_X1 U20993 ( .B1(n18919), .B2(n19002), .A(n18914), .ZN(P3_U3292) );
  INV_X1 U20994 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19000) );
  NOR3_X1 U20995 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18916) );
  OAI21_X1 U20996 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18916), .A(n18919), .ZN(
        n18915) );
  OAI21_X1 U20997 ( .B1(n18919), .B2(n19000), .A(n18915), .ZN(P3_U2638) );
  INV_X1 U20998 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22280) );
  AOI21_X1 U20999 ( .B1(n18963), .B2(n22280), .A(n18916), .ZN(n18918) );
  INV_X1 U21000 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19004) );
  INV_X1 U21001 ( .A(n18919), .ZN(n18917) );
  AOI22_X1 U21002 ( .A1(n18919), .A2(n18918), .B1(n19004), .B2(n18917), .ZN(
        P3_U2639) );
  INV_X1 U21003 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19005) );
  AOI22_X1 U21004 ( .A1(n22288), .A2(n18920), .B1(n19005), .B2(n22333), .ZN(
        P3_U3297) );
  INV_X1 U21005 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18921) );
  AOI22_X1 U21006 ( .A1(n22288), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18921), 
        .B2(n22333), .ZN(P3_U3294) );
  AOI21_X1 U21007 ( .B1(n22335), .B2(n22284), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18922) );
  AOI22_X1 U21008 ( .A1(n22288), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18922), 
        .B2(n22333), .ZN(P3_U2635) );
  INV_X1 U21009 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21457) );
  AOI22_X1 U21010 ( .A1(n18957), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18923) );
  OAI21_X1 U21011 ( .B1(n21457), .B2(n18939), .A(n18923), .ZN(P3_U2767) );
  INV_X1 U21012 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n21446) );
  AOI22_X1 U21013 ( .A1(n18957), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18924) );
  OAI21_X1 U21014 ( .B1(n21446), .B2(n18939), .A(n18924), .ZN(P3_U2766) );
  INV_X1 U21015 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20819) );
  AOI22_X1 U21016 ( .A1(n18957), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18925) );
  OAI21_X1 U21017 ( .B1(n20819), .B2(n18939), .A(n18925), .ZN(P3_U2765) );
  INV_X1 U21018 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20821) );
  AOI22_X1 U21019 ( .A1(n18957), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18949), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18926) );
  OAI21_X1 U21020 ( .B1(n20821), .B2(n18939), .A(n18926), .ZN(P3_U2764) );
  INV_X1 U21021 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21308) );
  AOI22_X1 U21022 ( .A1(n18957), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18949), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18927) );
  OAI21_X1 U21023 ( .B1(n21308), .B2(n18939), .A(n18927), .ZN(P3_U2763) );
  INV_X1 U21024 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20824) );
  AOI22_X1 U21025 ( .A1(n18957), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18949), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18928) );
  OAI21_X1 U21026 ( .B1(n20824), .B2(n18939), .A(n18928), .ZN(P3_U2762) );
  INV_X1 U21027 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n21309) );
  AOI22_X1 U21028 ( .A1(n18957), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18949), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18929) );
  OAI21_X1 U21029 ( .B1(n21309), .B2(n18939), .A(n18929), .ZN(P3_U2761) );
  INV_X1 U21030 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20828) );
  INV_X2 U21031 ( .A(n21891), .ZN(n18957) );
  AOI22_X1 U21032 ( .A1(n18957), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18930) );
  OAI21_X1 U21033 ( .B1(n20828), .B2(n18939), .A(n18930), .ZN(P3_U2760) );
  INV_X1 U21034 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20830) );
  AOI22_X1 U21035 ( .A1(n18957), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18931) );
  OAI21_X1 U21036 ( .B1(n20830), .B2(n18939), .A(n18931), .ZN(P3_U2759) );
  INV_X1 U21037 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n21283) );
  AOI22_X1 U21038 ( .A1(n18957), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18932) );
  OAI21_X1 U21039 ( .B1(n21283), .B2(n18939), .A(n18932), .ZN(P3_U2758) );
  INV_X1 U21040 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20833) );
  AOI22_X1 U21041 ( .A1(n18957), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18933) );
  OAI21_X1 U21042 ( .B1(n20833), .B2(n18939), .A(n18933), .ZN(P3_U2757) );
  INV_X1 U21043 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n21295) );
  AOI22_X1 U21044 ( .A1(n18957), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18934) );
  OAI21_X1 U21045 ( .B1(n21295), .B2(n18939), .A(n18934), .ZN(P3_U2756) );
  INV_X1 U21046 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20836) );
  AOI22_X1 U21047 ( .A1(n18957), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18935) );
  OAI21_X1 U21048 ( .B1(n20836), .B2(n18939), .A(n18935), .ZN(P3_U2755) );
  INV_X1 U21049 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20838) );
  AOI22_X1 U21050 ( .A1(n18957), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18936) );
  OAI21_X1 U21051 ( .B1(n20838), .B2(n18939), .A(n18936), .ZN(P3_U2754) );
  INV_X1 U21052 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20840) );
  AOI22_X1 U21053 ( .A1(n18957), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18937) );
  OAI21_X1 U21054 ( .B1(n20840), .B2(n18939), .A(n18937), .ZN(P3_U2753) );
  INV_X1 U21055 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n21430) );
  AOI22_X1 U21056 ( .A1(n18957), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18938) );
  OAI21_X1 U21057 ( .B1(n21430), .B2(n18939), .A(n18938), .ZN(P3_U2752) );
  INV_X1 U21058 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20792) );
  NAND2_X1 U21059 ( .A1(n18940), .A2(n11381), .ZN(n18959) );
  AOI22_X1 U21060 ( .A1(n18957), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18941) );
  OAI21_X1 U21061 ( .B1(n20792), .B2(n18959), .A(n18941), .ZN(P3_U2751) );
  INV_X1 U21062 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n21357) );
  AOI22_X1 U21063 ( .A1(n18957), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18942) );
  OAI21_X1 U21064 ( .B1(n21357), .B2(n18959), .A(n18942), .ZN(P3_U2750) );
  INV_X1 U21065 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n21359) );
  AOI22_X1 U21066 ( .A1(n18957), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18943) );
  OAI21_X1 U21067 ( .B1(n21359), .B2(n18959), .A(n18943), .ZN(P3_U2749) );
  INV_X1 U21068 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20796) );
  AOI22_X1 U21069 ( .A1(n18957), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18949), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18944) );
  OAI21_X1 U21070 ( .B1(n20796), .B2(n18959), .A(n18944), .ZN(P3_U2748) );
  INV_X1 U21071 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n20798) );
  AOI22_X1 U21072 ( .A1(n18957), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18949), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18945) );
  OAI21_X1 U21073 ( .B1(n20798), .B2(n18959), .A(n18945), .ZN(P3_U2747) );
  INV_X1 U21074 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n21346) );
  AOI22_X1 U21075 ( .A1(n18957), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18949), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18946) );
  OAI21_X1 U21076 ( .B1(n21346), .B2(n18959), .A(n18946), .ZN(P3_U2746) );
  INV_X1 U21077 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20801) );
  AOI22_X1 U21078 ( .A1(n18957), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18949), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18947) );
  OAI21_X1 U21079 ( .B1(n20801), .B2(n18959), .A(n18947), .ZN(P3_U2745) );
  INV_X1 U21080 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20803) );
  AOI22_X1 U21081 ( .A1(n18957), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18949), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18948) );
  OAI21_X1 U21082 ( .B1(n20803), .B2(n18959), .A(n18948), .ZN(P3_U2744) );
  INV_X1 U21083 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20805) );
  AOI22_X1 U21084 ( .A1(n18957), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18949), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18950) );
  OAI21_X1 U21085 ( .B1(n20805), .B2(n18959), .A(n18950), .ZN(P3_U2743) );
  INV_X1 U21086 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20807) );
  AOI22_X1 U21087 ( .A1(n18957), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18951) );
  OAI21_X1 U21088 ( .B1(n20807), .B2(n18959), .A(n18951), .ZN(P3_U2742) );
  INV_X1 U21089 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n21377) );
  AOI22_X1 U21090 ( .A1(n18957), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18952) );
  OAI21_X1 U21091 ( .B1(n21377), .B2(n18959), .A(n18952), .ZN(P3_U2741) );
  INV_X1 U21092 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20811) );
  AOI22_X1 U21093 ( .A1(n18957), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18953) );
  OAI21_X1 U21094 ( .B1(n20811), .B2(n18959), .A(n18953), .ZN(P3_U2740) );
  INV_X1 U21095 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20813) );
  AOI22_X1 U21096 ( .A1(n18957), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18954) );
  OAI21_X1 U21097 ( .B1(n20813), .B2(n18959), .A(n18954), .ZN(P3_U2739) );
  INV_X1 U21098 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n21391) );
  AOI22_X1 U21099 ( .A1(n18957), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18955) );
  OAI21_X1 U21100 ( .B1(n21391), .B2(n18959), .A(n18955), .ZN(P3_U2738) );
  INV_X1 U21101 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n21387) );
  AOI22_X1 U21102 ( .A1(n18957), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18956), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18958) );
  OAI21_X1 U21103 ( .B1(n21387), .B2(n18959), .A(n18958), .ZN(P3_U2737) );
  NOR2_X1 U21104 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n18960), .ZN(n18961) );
  NOR2_X1 U21105 ( .A1(n22288), .A2(n18961), .ZN(P3_U2633) );
  OR2_X1 U21106 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22333), .ZN(n18992) );
  INV_X1 U21107 ( .A(n18992), .ZN(n18994) );
  AOI22_X1 U21108 ( .A1(n18994), .A2(P3_REIP_REG_2__SCAN_IN), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n22333), .ZN(n18962) );
  OAI21_X1 U21109 ( .B1(n18996), .B2(n18963), .A(n18962), .ZN(P3_U3032) );
  AOI22_X1 U21110 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18990), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n22333), .ZN(n18964) );
  OAI21_X1 U21111 ( .B1(n20876), .B2(n18992), .A(n18964), .ZN(P3_U3033) );
  AOI22_X1 U21112 ( .A1(n18994), .A2(P3_REIP_REG_4__SCAN_IN), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n22333), .ZN(n18965) );
  OAI21_X1 U21113 ( .B1(n18996), .B2(n20876), .A(n18965), .ZN(P3_U3034) );
  INV_X1 U21114 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20902) );
  AOI22_X1 U21115 ( .A1(n18994), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n22333), .ZN(n18966) );
  OAI21_X1 U21116 ( .B1(n18996), .B2(n20902), .A(n18966), .ZN(P3_U3035) );
  AOI22_X1 U21117 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n18990), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n22333), .ZN(n18967) );
  OAI21_X1 U21118 ( .B1(n20929), .B2(n18992), .A(n18967), .ZN(P3_U3036) );
  AOI22_X1 U21119 ( .A1(n18994), .A2(P3_REIP_REG_7__SCAN_IN), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n22333), .ZN(n18968) );
  OAI21_X1 U21120 ( .B1(n18996), .B2(n20929), .A(n18968), .ZN(P3_U3037) );
  INV_X1 U21121 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20947) );
  AOI22_X1 U21122 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n18990), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n22333), .ZN(n18969) );
  OAI21_X1 U21123 ( .B1(n20947), .B2(n18992), .A(n18969), .ZN(P3_U3038) );
  AOI22_X1 U21124 ( .A1(n18994), .A2(P3_REIP_REG_9__SCAN_IN), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n22333), .ZN(n18970) );
  OAI21_X1 U21125 ( .B1(n18996), .B2(n20947), .A(n18970), .ZN(P3_U3039) );
  AOI22_X1 U21126 ( .A1(n18994), .A2(P3_REIP_REG_10__SCAN_IN), .B1(
        P3_ADDRESS_REG_8__SCAN_IN), .B2(n22333), .ZN(n18971) );
  OAI21_X1 U21127 ( .B1(n18996), .B2(n20954), .A(n18971), .ZN(P3_U3040) );
  INV_X1 U21128 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20984) );
  AOI22_X1 U21129 ( .A1(n18994), .A2(P3_REIP_REG_11__SCAN_IN), .B1(
        P3_ADDRESS_REG_9__SCAN_IN), .B2(n22333), .ZN(n18972) );
  OAI21_X1 U21130 ( .B1(n18996), .B2(n20984), .A(n18972), .ZN(P3_U3041) );
  INV_X1 U21131 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20997) );
  AOI22_X1 U21132 ( .A1(n18994), .A2(P3_REIP_REG_12__SCAN_IN), .B1(
        P3_ADDRESS_REG_10__SCAN_IN), .B2(n22333), .ZN(n18973) );
  OAI21_X1 U21133 ( .B1(n18996), .B2(n20997), .A(n18973), .ZN(P3_U3042) );
  AOI22_X1 U21134 ( .A1(n18994), .A2(P3_REIP_REG_13__SCAN_IN), .B1(
        P3_ADDRESS_REG_11__SCAN_IN), .B2(n22333), .ZN(n18974) );
  OAI21_X1 U21135 ( .B1(n18996), .B2(n21005), .A(n18974), .ZN(P3_U3043) );
  INV_X1 U21136 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n21025) );
  AOI22_X1 U21137 ( .A1(n18994), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_ADDRESS_REG_12__SCAN_IN), .B2(n22333), .ZN(n18975) );
  OAI21_X1 U21138 ( .B1(n18996), .B2(n21025), .A(n18975), .ZN(P3_U3044) );
  INV_X1 U21139 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n21030) );
  AOI22_X1 U21140 ( .A1(n18994), .A2(P3_REIP_REG_15__SCAN_IN), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n22333), .ZN(n18976) );
  OAI21_X1 U21141 ( .B1(n18996), .B2(n21030), .A(n18976), .ZN(P3_U3045) );
  AOI22_X1 U21142 ( .A1(n18994), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_ADDRESS_REG_14__SCAN_IN), .B2(n22333), .ZN(n18977) );
  OAI21_X1 U21143 ( .B1(n18996), .B2(n21054), .A(n18977), .ZN(P3_U3046) );
  INV_X1 U21144 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n21075) );
  AOI22_X1 U21145 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18990), .B1(
        P3_ADDRESS_REG_15__SCAN_IN), .B2(n22333), .ZN(n18978) );
  OAI21_X1 U21146 ( .B1(n21075), .B2(n18992), .A(n18978), .ZN(P3_U3047) );
  AOI22_X1 U21147 ( .A1(n18994), .A2(P3_REIP_REG_18__SCAN_IN), .B1(
        P3_ADDRESS_REG_16__SCAN_IN), .B2(n22333), .ZN(n18979) );
  OAI21_X1 U21148 ( .B1(n18996), .B2(n21075), .A(n18979), .ZN(P3_U3048) );
  AOI22_X1 U21149 ( .A1(n18994), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_ADDRESS_REG_17__SCAN_IN), .B2(n22333), .ZN(n18980) );
  OAI21_X1 U21150 ( .B1(n18996), .B2(n21833), .A(n18980), .ZN(P3_U3049) );
  INV_X1 U21151 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n21104) );
  AOI22_X1 U21152 ( .A1(n18994), .A2(P3_REIP_REG_20__SCAN_IN), .B1(
        P3_ADDRESS_REG_18__SCAN_IN), .B2(n22333), .ZN(n18981) );
  OAI21_X1 U21153 ( .B1(n18996), .B2(n21104), .A(n18981), .ZN(P3_U3050) );
  AOI22_X1 U21154 ( .A1(n18994), .A2(P3_REIP_REG_21__SCAN_IN), .B1(
        P3_ADDRESS_REG_19__SCAN_IN), .B2(n22333), .ZN(n18982) );
  OAI21_X1 U21155 ( .B1(n18996), .B2(n21120), .A(n18982), .ZN(P3_U3051) );
  AOI22_X1 U21156 ( .A1(n18994), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_ADDRESS_REG_20__SCAN_IN), .B2(n22333), .ZN(n18983) );
  OAI21_X1 U21157 ( .B1(n18996), .B2(n21140), .A(n18983), .ZN(P3_U3052) );
  INV_X1 U21158 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n21141) );
  AOI22_X1 U21159 ( .A1(n18994), .A2(P3_REIP_REG_23__SCAN_IN), .B1(
        P3_ADDRESS_REG_21__SCAN_IN), .B2(n22333), .ZN(n18984) );
  OAI21_X1 U21160 ( .B1(n18996), .B2(n21141), .A(n18984), .ZN(P3_U3053) );
  INV_X1 U21161 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n21159) );
  AOI22_X1 U21162 ( .A1(n18994), .A2(P3_REIP_REG_24__SCAN_IN), .B1(
        P3_ADDRESS_REG_22__SCAN_IN), .B2(n22333), .ZN(n18985) );
  OAI21_X1 U21163 ( .B1(n18996), .B2(n21159), .A(n18985), .ZN(P3_U3054) );
  INV_X1 U21164 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n21177) );
  AOI22_X1 U21165 ( .A1(n18994), .A2(P3_REIP_REG_25__SCAN_IN), .B1(
        P3_ADDRESS_REG_23__SCAN_IN), .B2(n22333), .ZN(n18986) );
  OAI21_X1 U21166 ( .B1(n18996), .B2(n21177), .A(n18986), .ZN(P3_U3055) );
  AOI22_X1 U21167 ( .A1(n18994), .A2(P3_REIP_REG_26__SCAN_IN), .B1(
        P3_ADDRESS_REG_24__SCAN_IN), .B2(n22333), .ZN(n18987) );
  OAI21_X1 U21168 ( .B1(n18996), .B2(n21192), .A(n18987), .ZN(P3_U3056) );
  AOI22_X1 U21169 ( .A1(n18994), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_ADDRESS_REG_25__SCAN_IN), .B2(n22333), .ZN(n18988) );
  OAI21_X1 U21170 ( .B1(n18996), .B2(n21716), .A(n18988), .ZN(P3_U3057) );
  INV_X1 U21171 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n21216) );
  AOI22_X1 U21172 ( .A1(n18994), .A2(P3_REIP_REG_28__SCAN_IN), .B1(
        P3_ADDRESS_REG_26__SCAN_IN), .B2(n22333), .ZN(n18989) );
  OAI21_X1 U21173 ( .B1(n18996), .B2(n21216), .A(n18989), .ZN(P3_U3058) );
  AOI22_X1 U21174 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18990), .B1(
        P3_ADDRESS_REG_27__SCAN_IN), .B2(n22333), .ZN(n18991) );
  OAI21_X1 U21175 ( .B1(n21230), .B2(n18992), .A(n18991), .ZN(P3_U3059) );
  AOI22_X1 U21176 ( .A1(n18994), .A2(P3_REIP_REG_30__SCAN_IN), .B1(
        P3_ADDRESS_REG_28__SCAN_IN), .B2(n22333), .ZN(n18993) );
  OAI21_X1 U21177 ( .B1(n18996), .B2(n21230), .A(n18993), .ZN(P3_U3060) );
  AOI22_X1 U21178 ( .A1(n18994), .A2(P3_REIP_REG_31__SCAN_IN), .B1(
        P3_ADDRESS_REG_29__SCAN_IN), .B2(n22333), .ZN(n18995) );
  OAI21_X1 U21179 ( .B1(n18996), .B2(n21261), .A(n18995), .ZN(P3_U3061) );
  INV_X1 U21180 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18997) );
  AOI22_X1 U21181 ( .A1(n22288), .A2(n18998), .B1(n18997), .B2(n22333), .ZN(
        P3_U3277) );
  INV_X1 U21182 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18999) );
  AOI22_X1 U21183 ( .A1(n22288), .A2(n19000), .B1(n18999), .B2(n22333), .ZN(
        P3_U3276) );
  INV_X1 U21184 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19001) );
  AOI22_X1 U21185 ( .A1(n22288), .A2(n19002), .B1(n19001), .B2(n22333), .ZN(
        P3_U3275) );
  INV_X1 U21186 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19003) );
  AOI22_X1 U21187 ( .A1(n22288), .A2(n19004), .B1(n19003), .B2(n22333), .ZN(
        P3_U3274) );
  NOR4_X1 U21188 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n19007)
         );
  NOR4_X1 U21189 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n19005), .ZN(n19006) );
  INV_X2 U21190 ( .A(n19671), .ZN(U215) );
  NAND3_X1 U21191 ( .A1(n19007), .A2(n19006), .A3(U215), .ZN(U213) );
  OAI21_X1 U21192 ( .B1(n11354), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n22312), 
        .ZN(n19008) );
  NAND3_X1 U21193 ( .A1(n19009), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19008), 
        .ZN(n19012) );
  OAI21_X1 U21194 ( .B1(n22317), .B2(n19916), .A(n19010), .ZN(n19011) );
  NAND2_X1 U21195 ( .A1(n19012), .A2(n19011), .ZN(n19018) );
  OAI21_X1 U21196 ( .B1(n19341), .B2(n19014), .A(n19013), .ZN(n19015) );
  AOI21_X1 U21197 ( .B1(n19016), .B2(n19342), .A(n19015), .ZN(n19017) );
  MUX2_X1 U21198 ( .A(n19018), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n19017), 
        .Z(P2_U3610) );
  AOI22_X1 U21199 ( .A1(n19218), .A2(n19019), .B1(P2_EBX_REG_0__SCAN_IN), .B2(
        n19207), .ZN(n19022) );
  AOI22_X1 U21200 ( .A1(n19163), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19140), 
        .B2(n19020), .ZN(n19021) );
  OAI211_X1 U21201 ( .C1(n19023), .C2(n19165), .A(n19022), .B(n19021), .ZN(
        n19026) );
  OAI21_X1 U21202 ( .B1(n19124), .B2(n19092), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19024) );
  INV_X1 U21203 ( .A(n19024), .ZN(n19025) );
  AOI211_X1 U21204 ( .C1(n19040), .C2(n19027), .A(n19026), .B(n19025), .ZN(
        n19028) );
  OAI21_X1 U21205 ( .B1(n19030), .B2(n19029), .A(n19028), .ZN(P2_U2855) );
  NOR2_X1 U21206 ( .A1(n19193), .A2(n19031), .ZN(n19033) );
  XOR2_X1 U21207 ( .A(n19033), .B(n19032), .Z(n19043) );
  NOR2_X1 U21208 ( .A1(n19034), .A2(n19147), .ZN(n19037) );
  AOI22_X1 U21209 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19207), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19163), .ZN(n19035) );
  OAI211_X1 U21210 ( .C1(n19222), .C2(n19312), .A(n19035), .B(n19325), .ZN(
        n19036) );
  AOI211_X1 U21211 ( .C1(n19124), .C2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19037), .B(n19036), .ZN(n19042) );
  INV_X1 U21212 ( .A(n19038), .ZN(n20065) );
  INV_X1 U21213 ( .A(n19039), .ZN(n19316) );
  AOI22_X1 U21214 ( .A1(n20065), .A2(n19040), .B1(n19217), .B2(n19316), .ZN(
        n19041) );
  OAI211_X1 U21215 ( .C1(n19347), .C2(n19043), .A(n19042), .B(n19041), .ZN(
        P2_U2851) );
  OAI22_X1 U21216 ( .A1(n19045), .A2(n19147), .B1(n19182), .B2(n19044), .ZN(
        n19046) );
  INV_X1 U21217 ( .A(n19046), .ZN(n19047) );
  OAI21_X1 U21218 ( .B1(n19302), .B2(n19210), .A(n19047), .ZN(n19048) );
  AOI211_X1 U21219 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19207), .A(n19282), .B(
        n19048), .ZN(n19054) );
  NOR2_X1 U21220 ( .A1(n19193), .A2(n19049), .ZN(n19051) );
  XNOR2_X1 U21221 ( .A(n19051), .B(n19050), .ZN(n19052) );
  AOI22_X1 U21222 ( .A1(n19052), .A2(n19194), .B1(n19298), .B2(n19217), .ZN(
        n19053) );
  OAI211_X1 U21223 ( .C1(n19222), .C2(n19303), .A(n19054), .B(n19053), .ZN(
        P2_U2849) );
  AOI22_X1 U21224 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19208), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19163), .ZN(n19055) );
  OAI21_X1 U21225 ( .B1(n19056), .B2(n19147), .A(n19055), .ZN(n19057) );
  AOI211_X1 U21226 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n19207), .A(n19282), .B(
        n19057), .ZN(n19064) );
  NOR2_X1 U21227 ( .A1(n19193), .A2(n19058), .ZN(n19060) );
  XNOR2_X1 U21228 ( .A(n19060), .B(n19059), .ZN(n19062) );
  AOI22_X1 U21229 ( .A1(n19062), .A2(n19194), .B1(n19061), .B2(n19217), .ZN(
        n19063) );
  OAI211_X1 U21230 ( .C1(n19222), .C2(n19065), .A(n19064), .B(n19063), .ZN(
        P2_U2847) );
  AOI22_X1 U21231 ( .A1(n19066), .A2(n19218), .B1(n19208), .B2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n19067) );
  OAI21_X1 U21232 ( .B1(n19068), .B2(n19210), .A(n19067), .ZN(n19069) );
  AOI211_X1 U21233 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n19207), .A(n19282), .B(
        n19069), .ZN(n19076) );
  NOR2_X1 U21234 ( .A1(n19193), .A2(n19070), .ZN(n19072) );
  XNOR2_X1 U21235 ( .A(n19072), .B(n19071), .ZN(n19074) );
  AOI22_X1 U21236 ( .A1(n19074), .A2(n19194), .B1(n19073), .B2(n19217), .ZN(
        n19075) );
  OAI211_X1 U21237 ( .C1(n19077), .C2(n19222), .A(n19076), .B(n19075), .ZN(
        P2_U2845) );
  AOI22_X1 U21238 ( .A1(n19078), .A2(n19218), .B1(n19208), .B2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n19079) );
  OAI21_X1 U21239 ( .B1(n19080), .B2(n19210), .A(n19079), .ZN(n19081) );
  AOI211_X1 U21240 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n19207), .A(n19282), .B(
        n19081), .ZN(n19088) );
  NOR2_X1 U21241 ( .A1(n19193), .A2(n19082), .ZN(n19084) );
  XNOR2_X1 U21242 ( .A(n19084), .B(n19083), .ZN(n19086) );
  AOI22_X1 U21243 ( .A1(n19086), .A2(n19194), .B1(n19085), .B2(n19217), .ZN(
        n19087) );
  OAI211_X1 U21244 ( .C1(n19089), .C2(n19222), .A(n19088), .B(n19087), .ZN(
        P2_U2843) );
  OAI22_X1 U21245 ( .A1(n12110), .A2(n19199), .B1(n19090), .B2(n19210), .ZN(
        n19091) );
  AOI211_X1 U21246 ( .C1(n19095), .C2(n19092), .A(n19282), .B(n19091), .ZN(
        n19101) );
  AOI22_X1 U21247 ( .A1(n19093), .A2(n19218), .B1(n19124), .B2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19100) );
  AOI22_X1 U21248 ( .A1(n11273), .A2(n19217), .B1(n19823), .B2(n19140), .ZN(
        n19099) );
  OR2_X1 U21249 ( .A1(n19193), .A2(n19094), .ZN(n19106) );
  AOI211_X1 U21250 ( .C1(n19096), .C2(n19095), .A(n19347), .B(n19106), .ZN(
        n19097) );
  INV_X1 U21251 ( .A(n19097), .ZN(n19098) );
  NAND4_X1 U21252 ( .A1(n19101), .A2(n19100), .A3(n19099), .A4(n19098), .ZN(
        P2_U2842) );
  AOI22_X1 U21253 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19208), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19163), .ZN(n19102) );
  OAI21_X1 U21254 ( .B1(n19103), .B2(n19147), .A(n19102), .ZN(n19104) );
  AOI211_X1 U21255 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n19207), .A(n19282), .B(
        n19104), .ZN(n19109) );
  XOR2_X1 U21256 ( .A(n19106), .B(n19105), .Z(n19107) );
  AOI22_X1 U21257 ( .A1(n19107), .A2(n19194), .B1(n19260), .B2(n19217), .ZN(
        n19108) );
  OAI211_X1 U21258 ( .C1(n19256), .C2(n19222), .A(n19109), .B(n19108), .ZN(
        P2_U2841) );
  NOR2_X1 U21259 ( .A1(n19193), .A2(n19110), .ZN(n19111) );
  XNOR2_X1 U21260 ( .A(n19112), .B(n19111), .ZN(n19119) );
  OAI21_X1 U21261 ( .B1(n12124), .B2(n19199), .A(n19325), .ZN(n19115) );
  OAI22_X1 U21262 ( .A1(n19113), .A2(n19147), .B1(n12123), .B2(n19182), .ZN(
        n19114) );
  AOI211_X1 U21263 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19163), .A(n19115), 
        .B(n19114), .ZN(n19118) );
  XOR2_X1 U21264 ( .A(n16208), .B(n19116), .Z(n20318) );
  AOI22_X1 U21265 ( .A1(n19265), .A2(n19217), .B1(n19140), .B2(n20318), .ZN(
        n19117) );
  OAI211_X1 U21266 ( .C1(n19347), .C2(n19119), .A(n19118), .B(n19117), .ZN(
        P2_U2839) );
  OAI21_X1 U21267 ( .B1(n12132), .B2(n19199), .A(n19325), .ZN(n19123) );
  OAI22_X1 U21268 ( .A1(n19121), .A2(n19147), .B1(n19120), .B2(n19210), .ZN(
        n19122) );
  AOI211_X1 U21269 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19124), .A(
        n19123), .B(n19122), .ZN(n19131) );
  NOR2_X1 U21270 ( .A1(n19193), .A2(n19125), .ZN(n19127) );
  XNOR2_X1 U21271 ( .A(n19127), .B(n19126), .ZN(n19129) );
  AOI22_X1 U21272 ( .A1(n19129), .A2(n19194), .B1(n19128), .B2(n19217), .ZN(
        n19130) );
  OAI211_X1 U21273 ( .C1(n19132), .C2(n19222), .A(n19131), .B(n19130), .ZN(
        P2_U2837) );
  NAND2_X1 U21274 ( .A1(n11173), .A2(n19133), .ZN(n19134) );
  XOR2_X1 U21275 ( .A(n19135), .B(n19134), .Z(n19145) );
  AOI22_X1 U21276 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19208), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n19163), .ZN(n19136) );
  OAI21_X1 U21277 ( .B1(n19137), .B2(n19147), .A(n19136), .ZN(n19138) );
  AOI211_X1 U21278 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19207), .A(n19282), .B(
        n19138), .ZN(n19144) );
  INV_X1 U21279 ( .A(n19139), .ZN(n19142) );
  AOI22_X1 U21280 ( .A1(n19142), .A2(n19217), .B1(n19141), .B2(n19140), .ZN(
        n19143) );
  OAI211_X1 U21281 ( .C1(n19347), .C2(n19145), .A(n19144), .B(n19143), .ZN(
        P2_U2836) );
  INV_X1 U21282 ( .A(n19146), .ZN(n19148) );
  OAI222_X1 U21283 ( .A1(n19210), .A2(n19150), .B1(n19199), .B2(n19149), .C1(
        n19148), .C2(n19147), .ZN(n19154) );
  OAI22_X1 U21284 ( .A1(n19152), .A2(n19165), .B1(n19151), .B2(n19222), .ZN(
        n19153) );
  AOI211_X1 U21285 ( .C1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n19208), .A(
        n19154), .B(n19153), .ZN(n19158) );
  OAI211_X1 U21286 ( .C1(n19156), .C2(n19159), .A(n19194), .B(n19155), .ZN(
        n19157) );
  OAI211_X1 U21287 ( .C1(n19160), .C2(n19159), .A(n19158), .B(n19157), .ZN(
        P2_U2835) );
  INV_X1 U21288 ( .A(n19161), .ZN(n19168) );
  OAI22_X1 U21289 ( .A1(n19199), .A2(n12148), .B1(n12418), .B2(n19182), .ZN(
        n19162) );
  AOI21_X1 U21290 ( .B1(n19163), .B2(P2_REIP_REG_22__SCAN_IN), .A(n19162), 
        .ZN(n19164) );
  OAI21_X1 U21291 ( .B1(n19166), .B2(n19165), .A(n19164), .ZN(n19167) );
  AOI21_X1 U21292 ( .B1(n19168), .B2(n19218), .A(n19167), .ZN(n19175) );
  INV_X1 U21293 ( .A(n19169), .ZN(n19173) );
  NOR2_X1 U21294 ( .A1(n19193), .A2(n19170), .ZN(n19172) );
  AOI21_X1 U21295 ( .B1(n19173), .B2(n19172), .A(n19347), .ZN(n19171) );
  OAI21_X1 U21296 ( .B1(n19173), .B2(n19172), .A(n19171), .ZN(n19174) );
  OAI211_X1 U21297 ( .C1(n19222), .C2(n19176), .A(n19175), .B(n19174), .ZN(
        P2_U2833) );
  AND2_X1 U21298 ( .A1(n11173), .A2(n19177), .ZN(n19180) );
  OAI21_X1 U21299 ( .B1(n11751), .B2(n19180), .A(n19194), .ZN(n19179) );
  AOI21_X1 U21300 ( .B1(n11751), .B2(n19180), .A(n19179), .ZN(n19185) );
  OAI22_X1 U21301 ( .A1(n19183), .A2(n19182), .B1(n19181), .B2(n19210), .ZN(
        n19184) );
  AOI211_X1 U21302 ( .C1(n19207), .C2(P2_EBX_REG_25__SCAN_IN), .A(n19185), .B(
        n19184), .ZN(n19189) );
  AOI22_X1 U21303 ( .A1(n19187), .A2(n19218), .B1(n19217), .B2(n19186), .ZN(
        n19188) );
  OAI211_X1 U21304 ( .C1(n19190), .C2(n19222), .A(n19189), .B(n19188), .ZN(
        P2_U2830) );
  INV_X1 U21305 ( .A(n19191), .ZN(n19197) );
  NOR2_X1 U21306 ( .A1(n19193), .A2(n19192), .ZN(n19196) );
  OAI21_X1 U21307 ( .B1(n19197), .B2(n19196), .A(n19194), .ZN(n19195) );
  AOI21_X1 U21308 ( .B1(n19197), .B2(n19196), .A(n19195), .ZN(n19201) );
  OAI22_X1 U21309 ( .A1(n12164), .A2(n19199), .B1(n19198), .B2(n19210), .ZN(
        n19200) );
  AOI211_X1 U21310 ( .C1(n19208), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n19201), .B(n19200), .ZN(n19205) );
  AOI22_X1 U21311 ( .A1(n19203), .A2(n19218), .B1(n19217), .B2(n19202), .ZN(
        n19204) );
  OAI211_X1 U21312 ( .C1(n19206), .C2(n19222), .A(n19205), .B(n19204), .ZN(
        P2_U2829) );
  AOI22_X1 U21313 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19208), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19207), .ZN(n19209) );
  OAI21_X1 U21314 ( .B1(n19211), .B2(n19210), .A(n19209), .ZN(n19212) );
  AOI221_X1 U21315 ( .B1(n19215), .B2(n19214), .C1(n19213), .C2(n19214), .A(
        n19212), .ZN(n19221) );
  AOI22_X1 U21316 ( .A1(n19219), .A2(n19218), .B1(n19217), .B2(n19216), .ZN(
        n19220) );
  OAI211_X1 U21317 ( .C1(n19223), .C2(n19222), .A(n19221), .B(n19220), .ZN(
        P2_U2826) );
  OAI22_X1 U21318 ( .A1(n19327), .A2(n19226), .B1(n19225), .B2(n19224), .ZN(
        n19227) );
  INV_X1 U21319 ( .A(n19227), .ZN(n19236) );
  NAND2_X1 U21320 ( .A1(n19271), .A2(n19228), .ZN(n19232) );
  AOI21_X1 U21321 ( .B1(n19329), .B2(n19230), .A(n19229), .ZN(n19231) );
  OAI211_X1 U21322 ( .C1(n19304), .C2(n19233), .A(n19232), .B(n19231), .ZN(
        n19234) );
  INV_X1 U21323 ( .A(n19234), .ZN(n19235) );
  OAI211_X1 U21324 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19237), .A(
        n19236), .B(n19235), .ZN(P2_U3046) );
  AOI22_X1 U21325 ( .A1(n19281), .A2(n19238), .B1(P2_REIP_REG_11__SCAN_IN), 
        .B2(n19282), .ZN(n19250) );
  INV_X1 U21326 ( .A(n19239), .ZN(n19241) );
  OAI22_X1 U21327 ( .A1(n19241), .A2(n19304), .B1(n19285), .B2(n19240), .ZN(
        n19242) );
  AOI21_X1 U21328 ( .B1(n19271), .B2(n19243), .A(n19242), .ZN(n19249) );
  OAI21_X1 U21329 ( .B1(n19245), .B2(n19244), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n19248) );
  NAND4_X1 U21330 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n19253), .A4(n19246), .ZN(
        n19247) );
  NAND4_X1 U21331 ( .A1(n19250), .A2(n19249), .A3(n19248), .A4(n19247), .ZN(
        P2_U3035) );
  AOI21_X1 U21332 ( .B1(n19252), .B2(n19251), .A(n14033), .ZN(n19258) );
  NAND2_X1 U21333 ( .A1(n19254), .A2(n19253), .ZN(n19255) );
  OAI22_X1 U21334 ( .A1(n19327), .A2(n19256), .B1(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n19255), .ZN(n19257) );
  AOI211_X1 U21335 ( .C1(n19282), .C2(P2_REIP_REG_14__SCAN_IN), .A(n19258), 
        .B(n19257), .ZN(n19263) );
  INV_X1 U21336 ( .A(n19259), .ZN(n19261) );
  AOI22_X1 U21337 ( .A1(n19261), .A2(n19335), .B1(n19329), .B2(n19260), .ZN(
        n19262) );
  OAI211_X1 U21338 ( .C1(n19332), .C2(n19264), .A(n19263), .B(n19262), .ZN(
        P2_U3032) );
  AOI22_X1 U21339 ( .A1(n19265), .A2(n19329), .B1(n19281), .B2(n20318), .ZN(
        n19279) );
  INV_X1 U21340 ( .A(n19266), .ZN(n19267) );
  AOI22_X1 U21341 ( .A1(n19269), .A2(n19268), .B1(n19335), .B2(n19267), .ZN(
        n19278) );
  NOR2_X1 U21342 ( .A1(n19271), .A2(n19270), .ZN(n19273) );
  OAI21_X1 U21343 ( .B1(n19274), .B2(n19273), .A(n19272), .ZN(n19275) );
  NAND2_X1 U21344 ( .A1(n19275), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n19276) );
  NAND4_X1 U21345 ( .A1(n19279), .A2(n19278), .A3(n19277), .A4(n19276), .ZN(
        P2_U3030) );
  INV_X1 U21346 ( .A(n19280), .ZN(n19293) );
  NAND2_X1 U21347 ( .A1(n19281), .A2(n19829), .ZN(n19284) );
  NAND2_X1 U21348 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19282), .ZN(n19283) );
  OAI211_X1 U21349 ( .C1(n19286), .C2(n19285), .A(n19284), .B(n19283), .ZN(
        n19287) );
  AOI21_X1 U21350 ( .B1(n19288), .B2(n19335), .A(n19287), .ZN(n19289) );
  OAI21_X1 U21351 ( .B1(n19290), .B2(n19332), .A(n19289), .ZN(n19291) );
  INV_X1 U21352 ( .A(n19291), .ZN(n19292) );
  OAI221_X1 U21353 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n19295), .C1(
        n19294), .C2(n19293), .A(n19292), .ZN(P2_U3039) );
  INV_X1 U21354 ( .A(n19296), .ZN(n19297) );
  NOR2_X1 U21355 ( .A1(n19297), .A2(n19338), .ZN(n19300) );
  AOI22_X1 U21356 ( .A1(n19300), .A2(n19299), .B1(n19298), .B2(n19329), .ZN(
        n19310) );
  INV_X1 U21357 ( .A(n19301), .ZN(n19308) );
  OAI22_X1 U21358 ( .A1(n19327), .A2(n19303), .B1(n19302), .B2(n19325), .ZN(
        n19307) );
  NOR2_X1 U21359 ( .A1(n19305), .A2(n19304), .ZN(n19306) );
  AOI211_X1 U21360 ( .C1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n19308), .A(
        n19307), .B(n19306), .ZN(n19309) );
  OAI211_X1 U21361 ( .C1(n19332), .C2(n19311), .A(n19310), .B(n19309), .ZN(
        P2_U3040) );
  NOR2_X1 U21362 ( .A1(n19327), .A2(n19312), .ZN(n19315) );
  OAI22_X1 U21363 ( .A1(n19325), .A2(n12076), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19313), .ZN(n19314) );
  AOI211_X1 U21364 ( .C1(n19316), .C2(n19329), .A(n19315), .B(n19314), .ZN(
        n19322) );
  NOR2_X1 U21365 ( .A1(n19318), .A2(n19317), .ZN(n19319) );
  AOI21_X1 U21366 ( .B1(n19320), .B2(n19335), .A(n19319), .ZN(n19321) );
  OAI211_X1 U21367 ( .C1(n19323), .C2(n19332), .A(n19322), .B(n19321), .ZN(
        P2_U3042) );
  INV_X1 U21368 ( .A(n19324), .ZN(n19333) );
  OAI22_X1 U21369 ( .A1(n20155), .A2(n19327), .B1(n19326), .B2(n19325), .ZN(
        n19328) );
  AOI21_X1 U21370 ( .B1(n19330), .B2(n19329), .A(n19328), .ZN(n19331) );
  OAI21_X1 U21371 ( .B1(n19333), .B2(n19332), .A(n19331), .ZN(n19334) );
  AOI21_X1 U21372 ( .B1(n19336), .B2(n19335), .A(n19334), .ZN(n19337) );
  OAI221_X1 U21373 ( .B1(n19340), .B2(n19339), .C1(n19340), .C2(n19338), .A(
        n19337), .ZN(P2_U3043) );
  AOI21_X1 U21374 ( .B1(n19343), .B2(n19342), .A(n19341), .ZN(n19348) );
  OAI211_X1 U21375 ( .C1(n19345), .C2(n19344), .A(n22317), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19346) );
  OAI211_X1 U21376 ( .C1(n19349), .C2(n19348), .A(n19347), .B(n19346), .ZN(
        P2_U3177) );
  NOR2_X1 U21377 ( .A1(n19351), .A2(n19350), .ZN(n19354) );
  MUX2_X1 U21378 ( .A(P2_MORE_REG_SCAN_IN), .B(n19352), .S(n19354), .Z(
        P2_U3609) );
  OAI21_X1 U21379 ( .B1(n19354), .B2(n14073), .A(n19353), .ZN(P2_U2819) );
  INV_X1 U21380 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20778) );
  INV_X1 U21381 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19379) );
  AOI22_X1 U21382 ( .A1(n19671), .A2(n20778), .B1(n19379), .B2(U215), .ZN(U282) );
  OAI22_X1 U21383 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19671), .ZN(n19355) );
  INV_X1 U21384 ( .A(n19355), .ZN(U281) );
  OAI22_X1 U21385 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19671), .ZN(n19356) );
  INV_X1 U21386 ( .A(n19356), .ZN(U280) );
  INV_X1 U21387 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n19357) );
  INV_X1 U21388 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n21401) );
  AOI22_X1 U21389 ( .A1(n19671), .A2(n19357), .B1(n21401), .B2(U215), .ZN(U279) );
  OAI22_X1 U21390 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19671), .ZN(n19358) );
  INV_X1 U21391 ( .A(n19358), .ZN(U278) );
  OAI22_X1 U21392 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19671), .ZN(n19359) );
  INV_X1 U21393 ( .A(n19359), .ZN(U277) );
  OAI22_X1 U21394 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19713), .ZN(n19360) );
  INV_X1 U21395 ( .A(n19360), .ZN(U276) );
  OAI22_X1 U21396 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19713), .ZN(n19361) );
  INV_X1 U21397 ( .A(n19361), .ZN(U275) );
  OAI22_X1 U21398 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19713), .ZN(n19362) );
  INV_X1 U21399 ( .A(n19362), .ZN(U274) );
  OAI22_X1 U21400 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19713), .ZN(n19363) );
  INV_X1 U21401 ( .A(n19363), .ZN(U273) );
  INV_X1 U21402 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n19364) );
  INV_X1 U21403 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n21337) );
  AOI22_X1 U21404 ( .A1(n19671), .A2(n19364), .B1(n21337), .B2(U215), .ZN(U272) );
  OAI22_X1 U21405 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19671), .ZN(n19365) );
  INV_X1 U21406 ( .A(n19365), .ZN(U271) );
  OAI22_X1 U21407 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19713), .ZN(n19366) );
  INV_X1 U21408 ( .A(n19366), .ZN(U270) );
  OAI22_X1 U21409 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19671), .ZN(n19367) );
  INV_X1 U21410 ( .A(n19367), .ZN(U269) );
  OAI22_X1 U21411 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19671), .ZN(n19368) );
  INV_X1 U21412 ( .A(n19368), .ZN(U268) );
  OAI22_X1 U21413 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19671), .ZN(n19369) );
  INV_X1 U21414 ( .A(n19369), .ZN(U267) );
  OAI22_X1 U21415 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19671), .ZN(n19370) );
  INV_X1 U21416 ( .A(n19370), .ZN(U266) );
  OAI22_X1 U21417 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19671), .ZN(n19371) );
  INV_X1 U21418 ( .A(n19371), .ZN(U265) );
  OAI22_X1 U21419 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19671), .ZN(n19372) );
  INV_X1 U21420 ( .A(n19372), .ZN(U264) );
  INV_X1 U21421 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n19373) );
  INV_X1 U21422 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n21292) );
  AOI22_X1 U21423 ( .A1(n19671), .A2(n19373), .B1(n21292), .B2(U215), .ZN(U263) );
  OAI22_X1 U21424 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19671), .ZN(n19374) );
  INV_X1 U21425 ( .A(n19374), .ZN(U262) );
  INV_X1 U21426 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n19375) );
  INV_X1 U21427 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n21300) );
  AOI22_X1 U21428 ( .A1(n19671), .A2(n19375), .B1(n21300), .B2(U215), .ZN(U261) );
  INV_X1 U21429 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n19376) );
  INV_X1 U21430 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n21306) );
  AOI22_X1 U21431 ( .A1(n19713), .A2(n19376), .B1(n21306), .B2(U215), .ZN(U260) );
  INV_X1 U21432 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n19377) );
  INV_X1 U21433 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n21442) );
  AOI22_X1 U21434 ( .A1(n19713), .A2(n19377), .B1(n21442), .B2(U215), .ZN(U259) );
  INV_X1 U21435 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n19378) );
  INV_X1 U21436 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n21311) );
  AOI22_X1 U21437 ( .A1(n19671), .A2(n19378), .B1(n21311), .B2(U215), .ZN(U258) );
  NOR3_X1 U21438 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19383), .A3(
        n21916), .ZN(n19381) );
  NAND2_X1 U21439 ( .A1(n19381), .A2(n19392), .ZN(n19675) );
  NOR2_X1 U21440 ( .A1(n19379), .A2(n19549), .ZN(n19452) );
  INV_X1 U21441 ( .A(n19381), .ZN(n19394) );
  NOR2_X2 U21442 ( .A1(n19392), .A2(n19394), .ZN(n19810) );
  NAND2_X1 U21443 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19715), .ZN(n19458) );
  NOR2_X2 U21444 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21937), .ZN(n21930) );
  NAND2_X1 U21445 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19411), .ZN(
        n19388) );
  NOR2_X1 U21446 ( .A1(n21930), .A2(n19388), .ZN(n19717) );
  NOR2_X2 U21447 ( .A1(n21311), .A2(n19591), .ZN(n19460) );
  AOI22_X1 U21448 ( .A1(n19810), .A2(n19461), .B1(n19717), .B2(n19460), .ZN(
        n19387) );
  INV_X1 U21449 ( .A(n19388), .ZN(n19455) );
  NOR2_X1 U21450 ( .A1(n19380), .A2(n19591), .ZN(n19393) );
  AOI22_X1 U21451 ( .A1(n19715), .A2(n19381), .B1(n19455), .B2(n19393), .ZN(
        n19719) );
  NOR2_X1 U21452 ( .A1(n19392), .A2(n19403), .ZN(n21904) );
  INV_X1 U21453 ( .A(n21904), .ZN(n19382) );
  NOR3_X2 U21454 ( .A1(n19383), .A2(n21916), .A3(n19382), .ZN(n19794) );
  NAND2_X1 U21455 ( .A1(n19385), .A2(n19384), .ZN(n19718) );
  NOR2_X2 U21456 ( .A1(n21438), .A2(n19718), .ZN(n19465) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19719), .B1(
        n19794), .B2(n19465), .ZN(n19386) );
  OAI211_X1 U21458 ( .C1(n19675), .C2(n19468), .A(n19387), .B(n19386), .ZN(
        P3_U2995) );
  NAND2_X1 U21459 ( .A1(n21904), .A2(n19414), .ZN(n19727) );
  INV_X1 U21460 ( .A(n19675), .ZN(n19734) );
  NOR2_X2 U21461 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19388), .ZN(
        n19801) );
  NOR2_X1 U21462 ( .A1(n19810), .A2(n19801), .ZN(n19389) );
  NOR2_X1 U21463 ( .A1(n21930), .A2(n19389), .ZN(n19723) );
  AOI22_X1 U21464 ( .A1(n19734), .A2(n19461), .B1(n19460), .B2(n19723), .ZN(
        n19391) );
  NAND2_X1 U21465 ( .A1(n19675), .A2(n19727), .ZN(n19399) );
  AOI21_X1 U21466 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19591), .ZN(n19463) );
  INV_X1 U21467 ( .A(n19389), .ZN(n19464) );
  AOI22_X1 U21468 ( .A1(n19715), .A2(n19399), .B1(n19463), .B2(n19464), .ZN(
        n19724) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19724), .B1(
        n19465), .B2(n19801), .ZN(n19390) );
  OAI211_X1 U21470 ( .C1(n19468), .C2(n19727), .A(n19391), .B(n19390), .ZN(
        P3_U2987) );
  NAND3_X1 U21471 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19414), .A3(
        n19392), .ZN(n19732) );
  INV_X1 U21472 ( .A(n19727), .ZN(n19739) );
  NOR2_X1 U21473 ( .A1(n21930), .A2(n19394), .ZN(n19728) );
  AOI22_X1 U21474 ( .A1(n19461), .A2(n19739), .B1(n19460), .B2(n19728), .ZN(
        n19397) );
  NAND2_X1 U21475 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19414), .ZN(
        n19402) );
  INV_X1 U21476 ( .A(n19393), .ZN(n19413) );
  OAI22_X1 U21477 ( .A1(n19549), .A2(n19402), .B1(n19394), .B2(n19413), .ZN(
        n19395) );
  INV_X1 U21478 ( .A(n19395), .ZN(n19729) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19729), .B1(
        n19465), .B2(n19810), .ZN(n19396) );
  OAI211_X1 U21480 ( .C1(n19468), .C2(n19732), .A(n19397), .B(n19396), .ZN(
        P3_U2979) );
  INV_X1 U21481 ( .A(n19414), .ZN(n19412) );
  NAND2_X1 U21482 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19403), .ZN(
        n19418) );
  NOR2_X2 U21483 ( .A1(n19412), .A2(n19418), .ZN(n19752) );
  INV_X1 U21484 ( .A(n19399), .ZN(n19398) );
  NOR2_X1 U21485 ( .A1(n21930), .A2(n19398), .ZN(n19733) );
  AOI22_X1 U21486 ( .A1(n19452), .A2(n19752), .B1(n19460), .B2(n19733), .ZN(
        n19401) );
  INV_X1 U21487 ( .A(n19752), .ZN(n19743) );
  NAND2_X1 U21488 ( .A1(n19732), .A2(n19743), .ZN(n19406) );
  AOI22_X1 U21489 ( .A1(n19715), .A2(n19406), .B1(n19463), .B2(n19399), .ZN(
        n19735) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19465), .ZN(n19400) );
  OAI211_X1 U21491 ( .C1(n19458), .C2(n19732), .A(n19401), .B(n19400), .ZN(
        P3_U2971) );
  NOR2_X1 U21492 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21907) );
  INV_X1 U21493 ( .A(n21907), .ZN(n19442) );
  NOR2_X2 U21494 ( .A1(n19442), .A2(n19412), .ZN(n19758) );
  NOR2_X1 U21495 ( .A1(n21930), .A2(n19402), .ZN(n19738) );
  AOI22_X1 U21496 ( .A1(n19452), .A2(n19758), .B1(n19460), .B2(n19738), .ZN(
        n19405) );
  AOI21_X1 U21497 ( .B1(n19403), .B2(n19428), .A(n19413), .ZN(n19444) );
  NAND2_X1 U21498 ( .A1(n19414), .A2(n19444), .ZN(n19740) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19740), .B1(
        n19465), .B2(n19739), .ZN(n19404) );
  OAI211_X1 U21500 ( .C1(n19458), .C2(n19743), .A(n19405), .B(n19404), .ZN(
        P3_U2963) );
  NAND2_X1 U21501 ( .A1(n21904), .A2(n19433), .ZN(n19688) );
  INV_X1 U21502 ( .A(n19406), .ZN(n19407) );
  NOR2_X1 U21503 ( .A1(n21930), .A2(n19407), .ZN(n19744) );
  AOI22_X1 U21504 ( .A1(n19461), .A2(n19758), .B1(n19460), .B2(n19744), .ZN(
        n19410) );
  INV_X1 U21505 ( .A(n19688), .ZN(n19764) );
  NOR2_X1 U21506 ( .A1(n19758), .A2(n19764), .ZN(n19419) );
  OAI21_X1 U21507 ( .B1(n19419), .B2(n19428), .A(n19407), .ZN(n19408) );
  OAI211_X1 U21508 ( .C1(n19745), .C2(n21937), .A(n19716), .B(n19408), .ZN(
        n19746) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19746), .B1(
        n19465), .B2(n19745), .ZN(n19409) );
  OAI211_X1 U21510 ( .C1(n19468), .C2(n19688), .A(n19410), .B(n19409), .ZN(
        P3_U2955) );
  NAND2_X1 U21511 ( .A1(n19411), .A2(n21916), .ZN(n19423) );
  NOR2_X2 U21512 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19423), .ZN(
        n19771) );
  AOI22_X1 U21513 ( .A1(n19452), .A2(n19771), .B1(n19460), .B2(n19750), .ZN(
        n19417) );
  INV_X1 U21514 ( .A(n19423), .ZN(n19415) );
  NOR2_X1 U21515 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19413), .ZN(
        n19454) );
  AOI22_X1 U21516 ( .A1(n19715), .A2(n19415), .B1(n19414), .B2(n19454), .ZN(
        n19753) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19753), .B1(
        n19465), .B2(n19752), .ZN(n19416) );
  OAI211_X1 U21518 ( .C1(n19458), .C2(n19688), .A(n19417), .B(n19416), .ZN(
        P3_U2947) );
  INV_X1 U21519 ( .A(n19418), .ZN(n19437) );
  NAND2_X1 U21520 ( .A1(n19437), .A2(n19433), .ZN(n19768) );
  NOR2_X1 U21521 ( .A1(n21930), .A2(n19419), .ZN(n19757) );
  AOI22_X1 U21522 ( .A1(n19461), .A2(n19771), .B1(n19460), .B2(n19757), .ZN(
        n19422) );
  NAND2_X1 U21523 ( .A1(n19762), .A2(n19768), .ZN(n19426) );
  INV_X1 U21524 ( .A(n19419), .ZN(n19420) );
  AOI22_X1 U21525 ( .A1(n19715), .A2(n19426), .B1(n19463), .B2(n19420), .ZN(
        n19759) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19759), .B1(
        n19465), .B2(n19758), .ZN(n19421) );
  OAI211_X1 U21527 ( .C1(n19468), .C2(n19768), .A(n19422), .B(n19421), .ZN(
        P3_U2939) );
  NAND2_X1 U21528 ( .A1(n21907), .A2(n19433), .ZN(n19774) );
  INV_X1 U21529 ( .A(n19768), .ZN(n19776) );
  NOR2_X1 U21530 ( .A1(n21930), .A2(n19423), .ZN(n19763) );
  AOI22_X1 U21531 ( .A1(n19461), .A2(n19776), .B1(n19460), .B2(n19763), .ZN(
        n19425) );
  NAND2_X1 U21532 ( .A1(n19444), .A2(n19433), .ZN(n19765) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19765), .B1(
        n19465), .B2(n19764), .ZN(n19424) );
  OAI211_X1 U21534 ( .C1(n19468), .C2(n19774), .A(n19425), .B(n19424), .ZN(
        P3_U2931) );
  NOR2_X1 U21535 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19453) );
  NAND2_X1 U21536 ( .A1(n21904), .A2(n19453), .ZN(n19780) );
  INV_X1 U21537 ( .A(n19426), .ZN(n19427) );
  NOR2_X1 U21538 ( .A1(n21930), .A2(n19427), .ZN(n19769) );
  AOI22_X1 U21539 ( .A1(n19461), .A2(n19782), .B1(n19460), .B2(n19769), .ZN(
        n19431) );
  INV_X1 U21540 ( .A(n19780), .ZN(n19788) );
  NOR2_X1 U21541 ( .A1(n19782), .A2(n19788), .ZN(n19438) );
  OAI21_X1 U21542 ( .B1(n19438), .B2(n19428), .A(n19427), .ZN(n19429) );
  OAI211_X1 U21543 ( .C1(n19771), .C2(n21937), .A(n19716), .B(n19429), .ZN(
        n19770) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19770), .B1(
        n19465), .B2(n19771), .ZN(n19430) );
  OAI211_X1 U21545 ( .C1(n19468), .C2(n19780), .A(n19431), .B(n19430), .ZN(
        P3_U2923) );
  NAND2_X1 U21546 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19453), .ZN(
        n19443) );
  NOR2_X2 U21547 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19443), .ZN(
        n19795) );
  INV_X1 U21548 ( .A(n19433), .ZN(n19432) );
  AOI22_X1 U21549 ( .A1(n19452), .A2(n19795), .B1(n19460), .B2(n19775), .ZN(
        n19436) );
  INV_X1 U21550 ( .A(n19443), .ZN(n19434) );
  AOI22_X1 U21551 ( .A1(n19715), .A2(n19434), .B1(n19433), .B2(n19454), .ZN(
        n19777) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19777), .B1(
        n19465), .B2(n19776), .ZN(n19435) );
  OAI211_X1 U21553 ( .C1(n19458), .C2(n19780), .A(n19436), .B(n19435), .ZN(
        P3_U2915) );
  NAND2_X1 U21554 ( .A1(n19437), .A2(n19453), .ZN(n19792) );
  NOR2_X1 U21555 ( .A1(n21930), .A2(n19438), .ZN(n19781) );
  AOI22_X1 U21556 ( .A1(n19461), .A2(n19795), .B1(n19460), .B2(n19781), .ZN(
        n19441) );
  INV_X1 U21557 ( .A(n19795), .ZN(n19786) );
  NAND2_X1 U21558 ( .A1(n19786), .A2(n19792), .ZN(n19448) );
  INV_X1 U21559 ( .A(n19438), .ZN(n19439) );
  AOI22_X1 U21560 ( .A1(n19715), .A2(n19448), .B1(n19463), .B2(n19439), .ZN(
        n19783) );
  AOI22_X1 U21561 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19783), .B1(
        n19465), .B2(n19782), .ZN(n19440) );
  OAI211_X1 U21562 ( .C1(n19468), .C2(n19792), .A(n19441), .B(n19440), .ZN(
        P3_U2907) );
  INV_X1 U21563 ( .A(n19453), .ZN(n19451) );
  NOR2_X2 U21564 ( .A1(n19442), .A2(n19451), .ZN(n19812) );
  NOR2_X1 U21565 ( .A1(n21930), .A2(n19443), .ZN(n19787) );
  AOI22_X1 U21566 ( .A1(n19452), .A2(n19812), .B1(n19460), .B2(n19787), .ZN(
        n19446) );
  NAND2_X1 U21567 ( .A1(n19444), .A2(n19453), .ZN(n19789) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19789), .B1(
        n19465), .B2(n19788), .ZN(n19445) );
  OAI211_X1 U21569 ( .C1(n19458), .C2(n19792), .A(n19446), .B(n19445), .ZN(
        P3_U2899) );
  INV_X1 U21570 ( .A(n19448), .ZN(n19447) );
  NOR2_X1 U21571 ( .A1(n21930), .A2(n19447), .ZN(n19793) );
  AOI22_X1 U21572 ( .A1(n19461), .A2(n19812), .B1(n19460), .B2(n19793), .ZN(
        n19450) );
  INV_X1 U21573 ( .A(n19812), .ZN(n19799) );
  NAND2_X1 U21574 ( .A1(n19806), .A2(n19799), .ZN(n19462) );
  AOI22_X1 U21575 ( .A1(n19715), .A2(n19462), .B1(n19463), .B2(n19448), .ZN(
        n19796) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19796), .B1(
        n19465), .B2(n19795), .ZN(n19449) );
  OAI211_X1 U21577 ( .C1(n19468), .C2(n19806), .A(n19450), .B(n19449), .ZN(
        P3_U2891) );
  AOI22_X1 U21578 ( .A1(n19452), .A2(n19801), .B1(n19460), .B2(n19800), .ZN(
        n19457) );
  AOI22_X1 U21579 ( .A1(n19715), .A2(n19455), .B1(n19454), .B2(n19453), .ZN(
        n19803) );
  INV_X1 U21580 ( .A(n19792), .ZN(n19802) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19803), .B1(
        n19465), .B2(n19802), .ZN(n19456) );
  OAI211_X1 U21582 ( .C1(n19806), .C2(n19458), .A(n19457), .B(n19456), .ZN(
        P3_U2883) );
  INV_X1 U21583 ( .A(n19810), .ZN(n19722) );
  INV_X1 U21584 ( .A(n19462), .ZN(n19459) );
  NOR2_X1 U21585 ( .A1(n21930), .A2(n19459), .ZN(n19808) );
  AOI22_X1 U21586 ( .A1(n19461), .A2(n19801), .B1(n19460), .B2(n19808), .ZN(
        n19467) );
  AOI22_X1 U21587 ( .A1(n19715), .A2(n19464), .B1(n19463), .B2(n19462), .ZN(
        n19813) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19813), .B1(
        n19465), .B2(n19812), .ZN(n19466) );
  OAI211_X1 U21589 ( .C1(n19468), .C2(n19722), .A(n19467), .B(n19466), .ZN(
        P3_U2875) );
  INV_X1 U21590 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n19469) );
  INV_X1 U21591 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21316) );
  AOI22_X1 U21592 ( .A1(n19713), .A2(n19469), .B1(n21316), .B2(U215), .ZN(U257) );
  NAND2_X1 U21593 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19715), .ZN(n19500) );
  NAND2_X1 U21594 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19715), .ZN(n19508) );
  INV_X1 U21595 ( .A(n19508), .ZN(n19497) );
  NOR2_X2 U21596 ( .A1(n21316), .A2(n19591), .ZN(n19503) );
  AOI22_X1 U21597 ( .A1(n19810), .A2(n19497), .B1(n19717), .B2(n19503), .ZN(
        n19472) );
  NOR2_X2 U21598 ( .A1(n19470), .A2(n19718), .ZN(n19505) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19719), .B1(
        n19794), .B2(n19505), .ZN(n19471) );
  OAI211_X1 U21600 ( .C1(n19675), .C2(n19500), .A(n19472), .B(n19471), .ZN(
        P3_U2994) );
  INV_X1 U21601 ( .A(n19500), .ZN(n19504) );
  AOI22_X1 U21602 ( .A1(n19739), .A2(n19504), .B1(n19723), .B2(n19503), .ZN(
        n19474) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19724), .B1(
        n19801), .B2(n19505), .ZN(n19473) );
  OAI211_X1 U21604 ( .C1(n19675), .C2(n19508), .A(n19474), .B(n19473), .ZN(
        P3_U2986) );
  AOI22_X1 U21605 ( .A1(n19739), .A2(n19497), .B1(n19728), .B2(n19503), .ZN(
        n19476) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19729), .B1(
        n19810), .B2(n19505), .ZN(n19475) );
  OAI211_X1 U21607 ( .C1(n19732), .C2(n19500), .A(n19476), .B(n19475), .ZN(
        P3_U2978) );
  AOI22_X1 U21608 ( .A1(n19752), .A2(n19504), .B1(n19733), .B2(n19503), .ZN(
        n19478) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19505), .ZN(n19477) );
  OAI211_X1 U21610 ( .C1(n19732), .C2(n19508), .A(n19478), .B(n19477), .ZN(
        P3_U2970) );
  AOI22_X1 U21611 ( .A1(n19738), .A2(n19503), .B1(n19758), .B2(n19504), .ZN(
        n19480) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n19505), .ZN(n19479) );
  OAI211_X1 U21613 ( .C1(n19743), .C2(n19508), .A(n19480), .B(n19479), .ZN(
        P3_U2962) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19746), .B1(
        n19744), .B2(n19503), .ZN(n19482) );
  AOI22_X1 U21615 ( .A1(n19745), .A2(n19505), .B1(n19758), .B2(n19497), .ZN(
        n19481) );
  OAI211_X1 U21616 ( .C1(n19688), .C2(n19500), .A(n19482), .B(n19481), .ZN(
        P3_U2954) );
  AOI22_X1 U21617 ( .A1(n19764), .A2(n19497), .B1(n19750), .B2(n19503), .ZN(
        n19484) );
  AOI22_X1 U21618 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n19505), .ZN(n19483) );
  OAI211_X1 U21619 ( .C1(n19762), .C2(n19500), .A(n19484), .B(n19483), .ZN(
        P3_U2946) );
  AOI22_X1 U21620 ( .A1(n19776), .A2(n19504), .B1(n19757), .B2(n19503), .ZN(
        n19486) );
  AOI22_X1 U21621 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19759), .B1(
        n19758), .B2(n19505), .ZN(n19485) );
  OAI211_X1 U21622 ( .C1(n19762), .C2(n19508), .A(n19486), .B(n19485), .ZN(
        P3_U2938) );
  AOI22_X1 U21623 ( .A1(n19776), .A2(n19497), .B1(n19763), .B2(n19503), .ZN(
        n19488) );
  AOI22_X1 U21624 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19765), .B1(
        n19764), .B2(n19505), .ZN(n19487) );
  OAI211_X1 U21625 ( .C1(n19774), .C2(n19500), .A(n19488), .B(n19487), .ZN(
        P3_U2930) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19503), .ZN(n19490) );
  AOI22_X1 U21627 ( .A1(n19771), .A2(n19505), .B1(n19788), .B2(n19504), .ZN(
        n19489) );
  OAI211_X1 U21628 ( .C1(n19774), .C2(n19508), .A(n19490), .B(n19489), .ZN(
        P3_U2922) );
  AOI22_X1 U21629 ( .A1(n19795), .A2(n19504), .B1(n19775), .B2(n19503), .ZN(
        n19492) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19505), .ZN(n19491) );
  OAI211_X1 U21631 ( .C1(n19780), .C2(n19508), .A(n19492), .B(n19491), .ZN(
        P3_U2914) );
  AOI22_X1 U21632 ( .A1(n19802), .A2(n19504), .B1(n19781), .B2(n19503), .ZN(
        n19494) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19505), .ZN(n19493) );
  OAI211_X1 U21634 ( .C1(n19786), .C2(n19508), .A(n19494), .B(n19493), .ZN(
        P3_U2906) );
  AOI22_X1 U21635 ( .A1(n19802), .A2(n19497), .B1(n19787), .B2(n19503), .ZN(
        n19496) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19789), .B1(
        n19788), .B2(n19505), .ZN(n19495) );
  OAI211_X1 U21637 ( .C1(n19799), .C2(n19500), .A(n19496), .B(n19495), .ZN(
        P3_U2898) );
  AOI22_X1 U21638 ( .A1(n19812), .A2(n19497), .B1(n19793), .B2(n19503), .ZN(
        n19499) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19796), .B1(
        n19795), .B2(n19505), .ZN(n19498) );
  OAI211_X1 U21640 ( .C1(n19806), .C2(n19500), .A(n19499), .B(n19498), .ZN(
        P3_U2890) );
  AOI22_X1 U21641 ( .A1(n19801), .A2(n19504), .B1(n19800), .B2(n19503), .ZN(
        n19502) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19803), .B1(
        n19802), .B2(n19505), .ZN(n19501) );
  OAI211_X1 U21643 ( .C1(n19806), .C2(n19508), .A(n19502), .B(n19501), .ZN(
        P3_U2882) );
  INV_X1 U21644 ( .A(n19801), .ZN(n19817) );
  AOI22_X1 U21645 ( .A1(n19810), .A2(n19504), .B1(n19808), .B2(n19503), .ZN(
        n19507) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n19505), .ZN(n19506) );
  OAI211_X1 U21647 ( .C1(n19817), .C2(n19508), .A(n19507), .B(n19506), .ZN(
        P3_U2874) );
  INV_X1 U21648 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n19509) );
  INV_X1 U21649 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21320) );
  AOI22_X1 U21650 ( .A1(n19671), .A2(n19509), .B1(n21320), .B2(U215), .ZN(U256) );
  NAND2_X1 U21651 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19715), .ZN(n19541) );
  NOR2_X1 U21652 ( .A1(n19549), .A2(n21337), .ZN(n19538) );
  NOR2_X2 U21653 ( .A1(n19591), .A2(n21320), .ZN(n19542) );
  AOI22_X1 U21654 ( .A1(n19810), .A2(n19538), .B1(n19717), .B2(n19542), .ZN(
        n19511) );
  NOR2_X2 U21655 ( .A1(n21335), .A2(n19718), .ZN(n19544) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19719), .B1(
        n19794), .B2(n19544), .ZN(n19510) );
  OAI211_X1 U21657 ( .C1(n19675), .C2(n19541), .A(n19511), .B(n19510), .ZN(
        P3_U2993) );
  INV_X1 U21658 ( .A(n19538), .ZN(n19547) );
  INV_X1 U21659 ( .A(n19541), .ZN(n19543) );
  AOI22_X1 U21660 ( .A1(n19739), .A2(n19543), .B1(n19723), .B2(n19542), .ZN(
        n19513) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19724), .B1(
        n19801), .B2(n19544), .ZN(n19512) );
  OAI211_X1 U21662 ( .C1(n19675), .C2(n19547), .A(n19513), .B(n19512), .ZN(
        P3_U2985) );
  AOI22_X1 U21663 ( .A1(n19745), .A2(n19543), .B1(n19728), .B2(n19542), .ZN(
        n19515) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19729), .B1(
        n19810), .B2(n19544), .ZN(n19514) );
  OAI211_X1 U21665 ( .C1(n19727), .C2(n19547), .A(n19515), .B(n19514), .ZN(
        P3_U2977) );
  AOI22_X1 U21666 ( .A1(n19752), .A2(n19543), .B1(n19733), .B2(n19542), .ZN(
        n19517) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19544), .ZN(n19516) );
  OAI211_X1 U21668 ( .C1(n19732), .C2(n19547), .A(n19517), .B(n19516), .ZN(
        P3_U2969) );
  INV_X1 U21669 ( .A(n19758), .ZN(n19749) );
  AOI22_X1 U21670 ( .A1(n19752), .A2(n19538), .B1(n19738), .B2(n19542), .ZN(
        n19519) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n19544), .ZN(n19518) );
  OAI211_X1 U21672 ( .C1(n19749), .C2(n19541), .A(n19519), .B(n19518), .ZN(
        P3_U2961) );
  AOI22_X1 U21673 ( .A1(n19764), .A2(n19543), .B1(n19744), .B2(n19542), .ZN(
        n19521) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n19544), .ZN(n19520) );
  OAI211_X1 U21675 ( .C1(n19749), .C2(n19547), .A(n19521), .B(n19520), .ZN(
        P3_U2953) );
  AOI22_X1 U21676 ( .A1(n19771), .A2(n19543), .B1(n19750), .B2(n19542), .ZN(
        n19523) );
  AOI22_X1 U21677 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n19544), .ZN(n19522) );
  OAI211_X1 U21678 ( .C1(n19688), .C2(n19547), .A(n19523), .B(n19522), .ZN(
        P3_U2945) );
  AOI22_X1 U21679 ( .A1(n19776), .A2(n19543), .B1(n19757), .B2(n19542), .ZN(
        n19525) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19759), .B1(
        n19758), .B2(n19544), .ZN(n19524) );
  OAI211_X1 U21681 ( .C1(n19762), .C2(n19547), .A(n19525), .B(n19524), .ZN(
        P3_U2937) );
  AOI22_X1 U21682 ( .A1(n19776), .A2(n19538), .B1(n19763), .B2(n19542), .ZN(
        n19527) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19765), .B1(
        n19764), .B2(n19544), .ZN(n19526) );
  OAI211_X1 U21684 ( .C1(n19774), .C2(n19541), .A(n19527), .B(n19526), .ZN(
        P3_U2929) );
  AOI22_X1 U21685 ( .A1(n19782), .A2(n19538), .B1(n19769), .B2(n19542), .ZN(
        n19529) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19770), .B1(
        n19771), .B2(n19544), .ZN(n19528) );
  OAI211_X1 U21687 ( .C1(n19780), .C2(n19541), .A(n19529), .B(n19528), .ZN(
        P3_U2921) );
  AOI22_X1 U21688 ( .A1(n19795), .A2(n19543), .B1(n19775), .B2(n19542), .ZN(
        n19531) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19544), .ZN(n19530) );
  OAI211_X1 U21690 ( .C1(n19780), .C2(n19547), .A(n19531), .B(n19530), .ZN(
        P3_U2913) );
  AOI22_X1 U21691 ( .A1(n19795), .A2(n19538), .B1(n19781), .B2(n19542), .ZN(
        n19533) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19544), .ZN(n19532) );
  OAI211_X1 U21693 ( .C1(n19792), .C2(n19541), .A(n19533), .B(n19532), .ZN(
        P3_U2905) );
  AOI22_X1 U21694 ( .A1(n19812), .A2(n19543), .B1(n19787), .B2(n19542), .ZN(
        n19535) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19789), .B1(
        n19788), .B2(n19544), .ZN(n19534) );
  OAI211_X1 U21696 ( .C1(n19792), .C2(n19547), .A(n19535), .B(n19534), .ZN(
        P3_U2897) );
  AOI22_X1 U21697 ( .A1(n19812), .A2(n19538), .B1(n19793), .B2(n19542), .ZN(
        n19537) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19796), .B1(
        n19795), .B2(n19544), .ZN(n19536) );
  OAI211_X1 U21699 ( .C1(n19806), .C2(n19541), .A(n19537), .B(n19536), .ZN(
        P3_U2889) );
  AOI22_X1 U21700 ( .A1(n19794), .A2(n19538), .B1(n19800), .B2(n19542), .ZN(
        n19540) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19803), .B1(
        n19802), .B2(n19544), .ZN(n19539) );
  OAI211_X1 U21702 ( .C1(n19817), .C2(n19541), .A(n19540), .B(n19539), .ZN(
        P3_U2881) );
  AOI22_X1 U21703 ( .A1(n19810), .A2(n19543), .B1(n19808), .B2(n19542), .ZN(
        n19546) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n19544), .ZN(n19545) );
  OAI211_X1 U21705 ( .C1(n19817), .C2(n19547), .A(n19546), .B(n19545), .ZN(
        P3_U2873) );
  INV_X1 U21706 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n19548) );
  AOI22_X1 U21707 ( .A1(n19671), .A2(n19548), .B1(n21325), .B2(U215), .ZN(U255) );
  NAND2_X1 U21708 ( .A1(n19715), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19582) );
  NOR2_X1 U21709 ( .A1(n21401), .A2(n19549), .ZN(n19579) );
  NOR2_X2 U21710 ( .A1(n19591), .A2(n21325), .ZN(n19583) );
  AOI22_X1 U21711 ( .A1(n19734), .A2(n19579), .B1(n19717), .B2(n19583), .ZN(
        n19552) );
  NOR2_X2 U21712 ( .A1(n19550), .A2(n19718), .ZN(n19585) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19719), .B1(
        n19794), .B2(n19585), .ZN(n19551) );
  OAI211_X1 U21714 ( .C1(n19722), .C2(n19582), .A(n19552), .B(n19551), .ZN(
        P3_U2992) );
  AOI22_X1 U21715 ( .A1(n19739), .A2(n19579), .B1(n19723), .B2(n19583), .ZN(
        n19554) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19724), .B1(
        n19801), .B2(n19585), .ZN(n19553) );
  OAI211_X1 U21717 ( .C1(n19675), .C2(n19582), .A(n19554), .B(n19553), .ZN(
        P3_U2984) );
  AOI22_X1 U21718 ( .A1(n19745), .A2(n19579), .B1(n19728), .B2(n19583), .ZN(
        n19556) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19729), .B1(
        n19810), .B2(n19585), .ZN(n19555) );
  OAI211_X1 U21720 ( .C1(n19727), .C2(n19582), .A(n19556), .B(n19555), .ZN(
        P3_U2976) );
  INV_X1 U21721 ( .A(n19579), .ZN(n19588) );
  INV_X1 U21722 ( .A(n19582), .ZN(n19584) );
  AOI22_X1 U21723 ( .A1(n19745), .A2(n19584), .B1(n19733), .B2(n19583), .ZN(
        n19558) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19585), .ZN(n19557) );
  OAI211_X1 U21725 ( .C1(n19743), .C2(n19588), .A(n19558), .B(n19557), .ZN(
        P3_U2968) );
  AOI22_X1 U21726 ( .A1(n19752), .A2(n19584), .B1(n19738), .B2(n19583), .ZN(
        n19560) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n19585), .ZN(n19559) );
  OAI211_X1 U21728 ( .C1(n19749), .C2(n19588), .A(n19560), .B(n19559), .ZN(
        P3_U2960) );
  AOI22_X1 U21729 ( .A1(n19764), .A2(n19579), .B1(n19744), .B2(n19583), .ZN(
        n19562) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n19585), .ZN(n19561) );
  OAI211_X1 U21731 ( .C1(n19749), .C2(n19582), .A(n19562), .B(n19561), .ZN(
        P3_U2952) );
  AOI22_X1 U21732 ( .A1(n19764), .A2(n19584), .B1(n19750), .B2(n19583), .ZN(
        n19564) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n19585), .ZN(n19563) );
  OAI211_X1 U21734 ( .C1(n19762), .C2(n19588), .A(n19564), .B(n19563), .ZN(
        P3_U2944) );
  AOI22_X1 U21735 ( .A1(n19776), .A2(n19579), .B1(n19757), .B2(n19583), .ZN(
        n19566) );
  AOI22_X1 U21736 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19759), .B1(
        n19758), .B2(n19585), .ZN(n19565) );
  OAI211_X1 U21737 ( .C1(n19762), .C2(n19582), .A(n19566), .B(n19565), .ZN(
        P3_U2936) );
  AOI22_X1 U21738 ( .A1(n19782), .A2(n19579), .B1(n19763), .B2(n19583), .ZN(
        n19568) );
  AOI22_X1 U21739 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19765), .B1(
        n19764), .B2(n19585), .ZN(n19567) );
  OAI211_X1 U21740 ( .C1(n19768), .C2(n19582), .A(n19568), .B(n19567), .ZN(
        P3_U2928) );
  AOI22_X1 U21741 ( .A1(n19782), .A2(n19584), .B1(n19769), .B2(n19583), .ZN(
        n19570) );
  AOI22_X1 U21742 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19770), .B1(
        n19771), .B2(n19585), .ZN(n19569) );
  OAI211_X1 U21743 ( .C1(n19780), .C2(n19588), .A(n19570), .B(n19569), .ZN(
        P3_U2920) );
  AOI22_X1 U21744 ( .A1(n19795), .A2(n19579), .B1(n19775), .B2(n19583), .ZN(
        n19572) );
  AOI22_X1 U21745 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19585), .ZN(n19571) );
  OAI211_X1 U21746 ( .C1(n19780), .C2(n19582), .A(n19572), .B(n19571), .ZN(
        P3_U2912) );
  AOI22_X1 U21747 ( .A1(n19802), .A2(n19579), .B1(n19781), .B2(n19583), .ZN(
        n19574) );
  AOI22_X1 U21748 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19585), .ZN(n19573) );
  OAI211_X1 U21749 ( .C1(n19786), .C2(n19582), .A(n19574), .B(n19573), .ZN(
        P3_U2904) );
  AOI22_X1 U21750 ( .A1(n19802), .A2(n19584), .B1(n19787), .B2(n19583), .ZN(
        n19576) );
  AOI22_X1 U21751 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19789), .B1(
        n19788), .B2(n19585), .ZN(n19575) );
  OAI211_X1 U21752 ( .C1(n19799), .C2(n19588), .A(n19576), .B(n19575), .ZN(
        P3_U2896) );
  AOI22_X1 U21753 ( .A1(n19794), .A2(n19579), .B1(n19793), .B2(n19583), .ZN(
        n19578) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19796), .B1(
        n19795), .B2(n19585), .ZN(n19577) );
  OAI211_X1 U21755 ( .C1(n19799), .C2(n19582), .A(n19578), .B(n19577), .ZN(
        P3_U2888) );
  AOI22_X1 U21756 ( .A1(n19801), .A2(n19579), .B1(n19800), .B2(n19583), .ZN(
        n19581) );
  AOI22_X1 U21757 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19803), .B1(
        n19802), .B2(n19585), .ZN(n19580) );
  OAI211_X1 U21758 ( .C1(n19806), .C2(n19582), .A(n19581), .B(n19580), .ZN(
        P3_U2880) );
  AOI22_X1 U21759 ( .A1(n19801), .A2(n19584), .B1(n19808), .B2(n19583), .ZN(
        n19587) );
  AOI22_X1 U21760 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n19585), .ZN(n19586) );
  OAI211_X1 U21761 ( .C1(n19722), .C2(n19588), .A(n19587), .B(n19586), .ZN(
        P3_U2872) );
  INV_X1 U21762 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n19590) );
  INV_X1 U21763 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n21329) );
  AOI22_X1 U21764 ( .A1(n19713), .A2(n19590), .B1(n21329), .B2(U215), .ZN(U254) );
  NAND2_X1 U21765 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19715), .ZN(n19630) );
  NAND2_X1 U21766 ( .A1(n19715), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19624) );
  INV_X1 U21767 ( .A(n19624), .ZN(n19626) );
  NOR2_X2 U21768 ( .A1(n19591), .A2(n21329), .ZN(n19625) );
  AOI22_X1 U21769 ( .A1(n19810), .A2(n19626), .B1(n19717), .B2(n19625), .ZN(
        n19594) );
  NOR2_X2 U21770 ( .A1(n19592), .A2(n19718), .ZN(n19627) );
  AOI22_X1 U21771 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19719), .B1(
        n19794), .B2(n19627), .ZN(n19593) );
  OAI211_X1 U21772 ( .C1(n19675), .C2(n19630), .A(n19594), .B(n19593), .ZN(
        P3_U2991) );
  INV_X1 U21773 ( .A(n19630), .ZN(n19621) );
  AOI22_X1 U21774 ( .A1(n19739), .A2(n19621), .B1(n19723), .B2(n19625), .ZN(
        n19596) );
  AOI22_X1 U21775 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19724), .B1(
        n19801), .B2(n19627), .ZN(n19595) );
  OAI211_X1 U21776 ( .C1(n19675), .C2(n19624), .A(n19596), .B(n19595), .ZN(
        P3_U2983) );
  AOI22_X1 U21777 ( .A1(n19739), .A2(n19626), .B1(n19728), .B2(n19625), .ZN(
        n19598) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19729), .B1(
        n19810), .B2(n19627), .ZN(n19597) );
  OAI211_X1 U21779 ( .C1(n19732), .C2(n19630), .A(n19598), .B(n19597), .ZN(
        P3_U2975) );
  AOI22_X1 U21780 ( .A1(n19745), .A2(n19626), .B1(n19733), .B2(n19625), .ZN(
        n19600) );
  AOI22_X1 U21781 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19627), .ZN(n19599) );
  OAI211_X1 U21782 ( .C1(n19743), .C2(n19630), .A(n19600), .B(n19599), .ZN(
        P3_U2967) );
  AOI22_X1 U21783 ( .A1(n19752), .A2(n19626), .B1(n19738), .B2(n19625), .ZN(
        n19602) );
  AOI22_X1 U21784 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n19627), .ZN(n19601) );
  OAI211_X1 U21785 ( .C1(n19749), .C2(n19630), .A(n19602), .B(n19601), .ZN(
        P3_U2959) );
  AOI22_X1 U21786 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19746), .B1(
        n19744), .B2(n19625), .ZN(n19604) );
  AOI22_X1 U21787 ( .A1(n19745), .A2(n19627), .B1(n19764), .B2(n19621), .ZN(
        n19603) );
  OAI211_X1 U21788 ( .C1(n19749), .C2(n19624), .A(n19604), .B(n19603), .ZN(
        P3_U2951) );
  AOI22_X1 U21789 ( .A1(n19771), .A2(n19621), .B1(n19750), .B2(n19625), .ZN(
        n19606) );
  AOI22_X1 U21790 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n19627), .ZN(n19605) );
  OAI211_X1 U21791 ( .C1(n19688), .C2(n19624), .A(n19606), .B(n19605), .ZN(
        P3_U2943) );
  AOI22_X1 U21792 ( .A1(n19771), .A2(n19626), .B1(n19757), .B2(n19625), .ZN(
        n19608) );
  AOI22_X1 U21793 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19759), .B1(
        n19758), .B2(n19627), .ZN(n19607) );
  OAI211_X1 U21794 ( .C1(n19768), .C2(n19630), .A(n19608), .B(n19607), .ZN(
        P3_U2935) );
  AOI22_X1 U21795 ( .A1(n19776), .A2(n19626), .B1(n19763), .B2(n19625), .ZN(
        n19610) );
  AOI22_X1 U21796 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19765), .B1(
        n19764), .B2(n19627), .ZN(n19609) );
  OAI211_X1 U21797 ( .C1(n19774), .C2(n19630), .A(n19610), .B(n19609), .ZN(
        P3_U2927) );
  AOI22_X1 U21798 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19625), .ZN(n19612) );
  AOI22_X1 U21799 ( .A1(n19771), .A2(n19627), .B1(n19788), .B2(n19621), .ZN(
        n19611) );
  OAI211_X1 U21800 ( .C1(n19774), .C2(n19624), .A(n19612), .B(n19611), .ZN(
        P3_U2919) );
  AOI22_X1 U21801 ( .A1(n19795), .A2(n19621), .B1(n19775), .B2(n19625), .ZN(
        n19614) );
  AOI22_X1 U21802 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19627), .ZN(n19613) );
  OAI211_X1 U21803 ( .C1(n19780), .C2(n19624), .A(n19614), .B(n19613), .ZN(
        P3_U2911) );
  AOI22_X1 U21804 ( .A1(n19795), .A2(n19626), .B1(n19781), .B2(n19625), .ZN(
        n19616) );
  AOI22_X1 U21805 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19627), .ZN(n19615) );
  OAI211_X1 U21806 ( .C1(n19792), .C2(n19630), .A(n19616), .B(n19615), .ZN(
        P3_U2903) );
  AOI22_X1 U21807 ( .A1(n19812), .A2(n19621), .B1(n19787), .B2(n19625), .ZN(
        n19618) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19789), .B1(
        n19788), .B2(n19627), .ZN(n19617) );
  OAI211_X1 U21809 ( .C1(n19792), .C2(n19624), .A(n19618), .B(n19617), .ZN(
        P3_U2895) );
  AOI22_X1 U21810 ( .A1(n19812), .A2(n19626), .B1(n19793), .B2(n19625), .ZN(
        n19620) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19796), .B1(
        n19795), .B2(n19627), .ZN(n19619) );
  OAI211_X1 U21812 ( .C1(n19806), .C2(n19630), .A(n19620), .B(n19619), .ZN(
        P3_U2887) );
  AOI22_X1 U21813 ( .A1(n19801), .A2(n19621), .B1(n19800), .B2(n19625), .ZN(
        n19623) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19803), .B1(
        n19802), .B2(n19627), .ZN(n19622) );
  OAI211_X1 U21815 ( .C1(n19806), .C2(n19624), .A(n19623), .B(n19622), .ZN(
        P3_U2879) );
  AOI22_X1 U21816 ( .A1(n19801), .A2(n19626), .B1(n19808), .B2(n19625), .ZN(
        n19629) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n19627), .ZN(n19628) );
  OAI211_X1 U21818 ( .C1(n19722), .C2(n19630), .A(n19629), .B(n19628), .ZN(
        P3_U2871) );
  OAI22_X1 U21819 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19671), .ZN(n19631) );
  INV_X1 U21820 ( .A(n19631), .ZN(U253) );
  NAND2_X1 U21821 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19715), .ZN(n19670) );
  NAND2_X1 U21822 ( .A1(n19715), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19664) );
  INV_X1 U21823 ( .A(n19664), .ZN(n19666) );
  AND2_X1 U21824 ( .A1(n19716), .A2(BUF2_REG_2__SCAN_IN), .ZN(n19665) );
  AOI22_X1 U21825 ( .A1(n19810), .A2(n19666), .B1(n19717), .B2(n19665), .ZN(
        n19634) );
  NOR2_X2 U21826 ( .A1(n19632), .A2(n19718), .ZN(n19667) );
  AOI22_X1 U21827 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19719), .B1(
        n19794), .B2(n19667), .ZN(n19633) );
  OAI211_X1 U21828 ( .C1(n19675), .C2(n19670), .A(n19634), .B(n19633), .ZN(
        P3_U2990) );
  AOI22_X1 U21829 ( .A1(n19734), .A2(n19666), .B1(n19723), .B2(n19665), .ZN(
        n19636) );
  AOI22_X1 U21830 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19724), .B1(
        n19801), .B2(n19667), .ZN(n19635) );
  OAI211_X1 U21831 ( .C1(n19727), .C2(n19670), .A(n19636), .B(n19635), .ZN(
        P3_U2982) );
  INV_X1 U21832 ( .A(n19670), .ZN(n19661) );
  AOI22_X1 U21833 ( .A1(n19745), .A2(n19661), .B1(n19728), .B2(n19665), .ZN(
        n19638) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19729), .B1(
        n19810), .B2(n19667), .ZN(n19637) );
  OAI211_X1 U21835 ( .C1(n19727), .C2(n19664), .A(n19638), .B(n19637), .ZN(
        P3_U2974) );
  AOI22_X1 U21836 ( .A1(n19752), .A2(n19661), .B1(n19733), .B2(n19665), .ZN(
        n19640) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19667), .ZN(n19639) );
  OAI211_X1 U21838 ( .C1(n19732), .C2(n19664), .A(n19640), .B(n19639), .ZN(
        P3_U2966) );
  AOI22_X1 U21839 ( .A1(n19752), .A2(n19666), .B1(n19738), .B2(n19665), .ZN(
        n19642) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n19667), .ZN(n19641) );
  OAI211_X1 U21841 ( .C1(n19749), .C2(n19670), .A(n19642), .B(n19641), .ZN(
        P3_U2958) );
  AOI22_X1 U21842 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19746), .B1(
        n19744), .B2(n19665), .ZN(n19644) );
  AOI22_X1 U21843 ( .A1(n19745), .A2(n19667), .B1(n19764), .B2(n19661), .ZN(
        n19643) );
  OAI211_X1 U21844 ( .C1(n19749), .C2(n19664), .A(n19644), .B(n19643), .ZN(
        P3_U2950) );
  AOI22_X1 U21845 ( .A1(n19764), .A2(n19666), .B1(n19750), .B2(n19665), .ZN(
        n19646) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n19667), .ZN(n19645) );
  OAI211_X1 U21847 ( .C1(n19762), .C2(n19670), .A(n19646), .B(n19645), .ZN(
        P3_U2942) );
  AOI22_X1 U21848 ( .A1(n19776), .A2(n19661), .B1(n19757), .B2(n19665), .ZN(
        n19648) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19759), .B1(
        n19758), .B2(n19667), .ZN(n19647) );
  OAI211_X1 U21850 ( .C1(n19762), .C2(n19664), .A(n19648), .B(n19647), .ZN(
        P3_U2934) );
  AOI22_X1 U21851 ( .A1(n19782), .A2(n19661), .B1(n19763), .B2(n19665), .ZN(
        n19650) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19765), .B1(
        n19764), .B2(n19667), .ZN(n19649) );
  OAI211_X1 U21853 ( .C1(n19768), .C2(n19664), .A(n19650), .B(n19649), .ZN(
        P3_U2926) );
  AOI22_X1 U21854 ( .A1(n19788), .A2(n19661), .B1(n19769), .B2(n19665), .ZN(
        n19652) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19770), .B1(
        n19771), .B2(n19667), .ZN(n19651) );
  OAI211_X1 U21856 ( .C1(n19774), .C2(n19664), .A(n19652), .B(n19651), .ZN(
        P3_U2918) );
  AOI22_X1 U21857 ( .A1(n19788), .A2(n19666), .B1(n19775), .B2(n19665), .ZN(
        n19654) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19667), .ZN(n19653) );
  OAI211_X1 U21859 ( .C1(n19786), .C2(n19670), .A(n19654), .B(n19653), .ZN(
        P3_U2910) );
  AOI22_X1 U21860 ( .A1(n19802), .A2(n19661), .B1(n19781), .B2(n19665), .ZN(
        n19656) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19667), .ZN(n19655) );
  OAI211_X1 U21862 ( .C1(n19786), .C2(n19664), .A(n19656), .B(n19655), .ZN(
        P3_U2902) );
  AOI22_X1 U21863 ( .A1(n19812), .A2(n19661), .B1(n19787), .B2(n19665), .ZN(
        n19658) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19789), .B1(
        n19788), .B2(n19667), .ZN(n19657) );
  OAI211_X1 U21865 ( .C1(n19792), .C2(n19664), .A(n19658), .B(n19657), .ZN(
        P3_U2894) );
  AOI22_X1 U21866 ( .A1(n19812), .A2(n19666), .B1(n19793), .B2(n19665), .ZN(
        n19660) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19796), .B1(
        n19795), .B2(n19667), .ZN(n19659) );
  OAI211_X1 U21868 ( .C1(n19806), .C2(n19670), .A(n19660), .B(n19659), .ZN(
        P3_U2886) );
  AOI22_X1 U21869 ( .A1(n19801), .A2(n19661), .B1(n19800), .B2(n19665), .ZN(
        n19663) );
  AOI22_X1 U21870 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19803), .B1(
        n19802), .B2(n19667), .ZN(n19662) );
  OAI211_X1 U21871 ( .C1(n19806), .C2(n19664), .A(n19663), .B(n19662), .ZN(
        P3_U2878) );
  AOI22_X1 U21872 ( .A1(n19801), .A2(n19666), .B1(n19808), .B2(n19665), .ZN(
        n19669) );
  AOI22_X1 U21873 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n19667), .ZN(n19668) );
  OAI211_X1 U21874 ( .C1(n19722), .C2(n19670), .A(n19669), .B(n19668), .ZN(
        P3_U2870) );
  OAI22_X1 U21875 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19671), .ZN(n19672) );
  INV_X1 U21876 ( .A(n19672), .ZN(U252) );
  NAND2_X1 U21877 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19715), .ZN(n19706) );
  NAND2_X1 U21878 ( .A1(n19715), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19712) );
  AND2_X1 U21879 ( .A1(n19716), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19707) );
  AOI22_X1 U21880 ( .A1(n19810), .A2(n19703), .B1(n19717), .B2(n19707), .ZN(
        n19674) );
  NOR2_X2 U21881 ( .A1(n21279), .A2(n19718), .ZN(n19709) );
  AOI22_X1 U21882 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19719), .B1(
        n19794), .B2(n19709), .ZN(n19673) );
  OAI211_X1 U21883 ( .C1(n19675), .C2(n19706), .A(n19674), .B(n19673), .ZN(
        P3_U2989) );
  AOI22_X1 U21884 ( .A1(n19734), .A2(n19703), .B1(n19723), .B2(n19707), .ZN(
        n19677) );
  AOI22_X1 U21885 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19724), .B1(
        n19801), .B2(n19709), .ZN(n19676) );
  OAI211_X1 U21886 ( .C1(n19727), .C2(n19706), .A(n19677), .B(n19676), .ZN(
        P3_U2981) );
  AOI22_X1 U21887 ( .A1(n19739), .A2(n19703), .B1(n19728), .B2(n19707), .ZN(
        n19679) );
  AOI22_X1 U21888 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19729), .B1(
        n19810), .B2(n19709), .ZN(n19678) );
  OAI211_X1 U21889 ( .C1(n19732), .C2(n19706), .A(n19679), .B(n19678), .ZN(
        P3_U2973) );
  AOI22_X1 U21890 ( .A1(n19745), .A2(n19703), .B1(n19733), .B2(n19707), .ZN(
        n19681) );
  AOI22_X1 U21891 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19709), .ZN(n19680) );
  OAI211_X1 U21892 ( .C1(n19743), .C2(n19706), .A(n19681), .B(n19680), .ZN(
        P3_U2965) );
  INV_X1 U21893 ( .A(n19706), .ZN(n19708) );
  AOI22_X1 U21894 ( .A1(n19738), .A2(n19707), .B1(n19758), .B2(n19708), .ZN(
        n19683) );
  AOI22_X1 U21895 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n19709), .ZN(n19682) );
  OAI211_X1 U21896 ( .C1(n19743), .C2(n19712), .A(n19683), .B(n19682), .ZN(
        P3_U2957) );
  AOI22_X1 U21897 ( .A1(n19758), .A2(n19703), .B1(n19744), .B2(n19707), .ZN(
        n19685) );
  AOI22_X1 U21898 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n19709), .ZN(n19684) );
  OAI211_X1 U21899 ( .C1(n19688), .C2(n19706), .A(n19685), .B(n19684), .ZN(
        P3_U2949) );
  AOI22_X1 U21900 ( .A1(n19771), .A2(n19708), .B1(n19750), .B2(n19707), .ZN(
        n19687) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n19709), .ZN(n19686) );
  OAI211_X1 U21902 ( .C1(n19688), .C2(n19712), .A(n19687), .B(n19686), .ZN(
        P3_U2941) );
  AOI22_X1 U21903 ( .A1(n19771), .A2(n19703), .B1(n19757), .B2(n19707), .ZN(
        n19690) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19759), .B1(
        n19758), .B2(n19709), .ZN(n19689) );
  OAI211_X1 U21905 ( .C1(n19768), .C2(n19706), .A(n19690), .B(n19689), .ZN(
        P3_U2933) );
  AOI22_X1 U21906 ( .A1(n19782), .A2(n19708), .B1(n19763), .B2(n19707), .ZN(
        n19692) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19765), .B1(
        n19764), .B2(n19709), .ZN(n19691) );
  OAI211_X1 U21908 ( .C1(n19768), .C2(n19712), .A(n19692), .B(n19691), .ZN(
        P3_U2925) );
  AOI22_X1 U21909 ( .A1(n19788), .A2(n19708), .B1(n19769), .B2(n19707), .ZN(
        n19694) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19770), .B1(
        n19771), .B2(n19709), .ZN(n19693) );
  OAI211_X1 U21911 ( .C1(n19774), .C2(n19712), .A(n19694), .B(n19693), .ZN(
        P3_U2917) );
  AOI22_X1 U21912 ( .A1(n19795), .A2(n19708), .B1(n19775), .B2(n19707), .ZN(
        n19696) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19709), .ZN(n19695) );
  OAI211_X1 U21914 ( .C1(n19780), .C2(n19712), .A(n19696), .B(n19695), .ZN(
        P3_U2909) );
  AOI22_X1 U21915 ( .A1(n19795), .A2(n19703), .B1(n19781), .B2(n19707), .ZN(
        n19698) );
  AOI22_X1 U21916 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19709), .ZN(n19697) );
  OAI211_X1 U21917 ( .C1(n19792), .C2(n19706), .A(n19698), .B(n19697), .ZN(
        P3_U2901) );
  AOI22_X1 U21918 ( .A1(n19812), .A2(n19708), .B1(n19787), .B2(n19707), .ZN(
        n19700) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19789), .B1(
        n19788), .B2(n19709), .ZN(n19699) );
  OAI211_X1 U21920 ( .C1(n19792), .C2(n19712), .A(n19700), .B(n19699), .ZN(
        P3_U2893) );
  AOI22_X1 U21921 ( .A1(n19812), .A2(n19703), .B1(n19793), .B2(n19707), .ZN(
        n19702) );
  AOI22_X1 U21922 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19796), .B1(
        n19795), .B2(n19709), .ZN(n19701) );
  OAI211_X1 U21923 ( .C1(n19806), .C2(n19706), .A(n19702), .B(n19701), .ZN(
        P3_U2885) );
  AOI22_X1 U21924 ( .A1(n19794), .A2(n19703), .B1(n19800), .B2(n19707), .ZN(
        n19705) );
  AOI22_X1 U21925 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19803), .B1(
        n19802), .B2(n19709), .ZN(n19704) );
  OAI211_X1 U21926 ( .C1(n19817), .C2(n19706), .A(n19705), .B(n19704), .ZN(
        P3_U2877) );
  AOI22_X1 U21927 ( .A1(n19810), .A2(n19708), .B1(n19808), .B2(n19707), .ZN(
        n19711) );
  AOI22_X1 U21928 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n19709), .ZN(n19710) );
  OAI211_X1 U21929 ( .C1(n19817), .C2(n19712), .A(n19711), .B(n19710), .ZN(
        P3_U2869) );
  OAI22_X1 U21930 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19713), .ZN(n19714) );
  INV_X1 U21931 ( .A(n19714), .ZN(U251) );
  NAND2_X1 U21932 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n19715), .ZN(n19816) );
  NAND2_X1 U21933 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19715), .ZN(n19756) );
  INV_X1 U21934 ( .A(n19756), .ZN(n19809) );
  AND2_X1 U21935 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n19716), .ZN(n19807) );
  AOI22_X1 U21936 ( .A1(n19734), .A2(n19809), .B1(n19717), .B2(n19807), .ZN(
        n19721) );
  NOR2_X2 U21937 ( .A1(n21278), .A2(n19718), .ZN(n19811) );
  AOI22_X1 U21938 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19719), .B1(
        n19794), .B2(n19811), .ZN(n19720) );
  OAI211_X1 U21939 ( .C1(n19722), .C2(n19816), .A(n19721), .B(n19720), .ZN(
        P3_U2988) );
  INV_X1 U21940 ( .A(n19816), .ZN(n19751) );
  AOI22_X1 U21941 ( .A1(n19734), .A2(n19751), .B1(n19723), .B2(n19807), .ZN(
        n19726) );
  AOI22_X1 U21942 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19724), .B1(
        n19801), .B2(n19811), .ZN(n19725) );
  OAI211_X1 U21943 ( .C1(n19727), .C2(n19756), .A(n19726), .B(n19725), .ZN(
        P3_U2980) );
  AOI22_X1 U21944 ( .A1(n19739), .A2(n19751), .B1(n19728), .B2(n19807), .ZN(
        n19731) );
  AOI22_X1 U21945 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19729), .B1(
        n19810), .B2(n19811), .ZN(n19730) );
  OAI211_X1 U21946 ( .C1(n19732), .C2(n19756), .A(n19731), .B(n19730), .ZN(
        P3_U2972) );
  AOI22_X1 U21947 ( .A1(n19745), .A2(n19751), .B1(n19733), .B2(n19807), .ZN(
        n19737) );
  AOI22_X1 U21948 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19811), .ZN(n19736) );
  OAI211_X1 U21949 ( .C1(n19743), .C2(n19756), .A(n19737), .B(n19736), .ZN(
        P3_U2964) );
  AOI22_X1 U21950 ( .A1(n19738), .A2(n19807), .B1(n19758), .B2(n19809), .ZN(
        n19742) );
  AOI22_X1 U21951 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19740), .B1(
        n19739), .B2(n19811), .ZN(n19741) );
  OAI211_X1 U21952 ( .C1(n19743), .C2(n19816), .A(n19742), .B(n19741), .ZN(
        P3_U2956) );
  AOI22_X1 U21953 ( .A1(n19764), .A2(n19809), .B1(n19744), .B2(n19807), .ZN(
        n19748) );
  AOI22_X1 U21954 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n19811), .ZN(n19747) );
  OAI211_X1 U21955 ( .C1(n19749), .C2(n19816), .A(n19748), .B(n19747), .ZN(
        P3_U2948) );
  AOI22_X1 U21956 ( .A1(n19764), .A2(n19751), .B1(n19750), .B2(n19807), .ZN(
        n19755) );
  AOI22_X1 U21957 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n19811), .ZN(n19754) );
  OAI211_X1 U21958 ( .C1(n19762), .C2(n19756), .A(n19755), .B(n19754), .ZN(
        P3_U2940) );
  AOI22_X1 U21959 ( .A1(n19776), .A2(n19809), .B1(n19757), .B2(n19807), .ZN(
        n19761) );
  AOI22_X1 U21960 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19759), .B1(
        n19758), .B2(n19811), .ZN(n19760) );
  OAI211_X1 U21961 ( .C1(n19762), .C2(n19816), .A(n19761), .B(n19760), .ZN(
        P3_U2932) );
  AOI22_X1 U21962 ( .A1(n19782), .A2(n19809), .B1(n19763), .B2(n19807), .ZN(
        n19767) );
  AOI22_X1 U21963 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19765), .B1(
        n19764), .B2(n19811), .ZN(n19766) );
  OAI211_X1 U21964 ( .C1(n19768), .C2(n19816), .A(n19767), .B(n19766), .ZN(
        P3_U2924) );
  AOI22_X1 U21965 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19807), .ZN(n19773) );
  AOI22_X1 U21966 ( .A1(n19771), .A2(n19811), .B1(n19788), .B2(n19809), .ZN(
        n19772) );
  OAI211_X1 U21967 ( .C1(n19774), .C2(n19816), .A(n19773), .B(n19772), .ZN(
        P3_U2916) );
  AOI22_X1 U21968 ( .A1(n19795), .A2(n19809), .B1(n19775), .B2(n19807), .ZN(
        n19779) );
  AOI22_X1 U21969 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19777), .B1(
        n19776), .B2(n19811), .ZN(n19778) );
  OAI211_X1 U21970 ( .C1(n19780), .C2(n19816), .A(n19779), .B(n19778), .ZN(
        P3_U2908) );
  AOI22_X1 U21971 ( .A1(n19802), .A2(n19809), .B1(n19781), .B2(n19807), .ZN(
        n19785) );
  AOI22_X1 U21972 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19811), .ZN(n19784) );
  OAI211_X1 U21973 ( .C1(n19786), .C2(n19816), .A(n19785), .B(n19784), .ZN(
        P3_U2900) );
  AOI22_X1 U21974 ( .A1(n19812), .A2(n19809), .B1(n19787), .B2(n19807), .ZN(
        n19791) );
  AOI22_X1 U21975 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19789), .B1(
        n19788), .B2(n19811), .ZN(n19790) );
  OAI211_X1 U21976 ( .C1(n19792), .C2(n19816), .A(n19791), .B(n19790), .ZN(
        P3_U2892) );
  AOI22_X1 U21977 ( .A1(n19794), .A2(n19809), .B1(n19793), .B2(n19807), .ZN(
        n19798) );
  AOI22_X1 U21978 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19796), .B1(
        n19795), .B2(n19811), .ZN(n19797) );
  OAI211_X1 U21979 ( .C1(n19799), .C2(n19816), .A(n19798), .B(n19797), .ZN(
        P3_U2884) );
  AOI22_X1 U21980 ( .A1(n19801), .A2(n19809), .B1(n19800), .B2(n19807), .ZN(
        n19805) );
  AOI22_X1 U21981 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19803), .B1(
        n19802), .B2(n19811), .ZN(n19804) );
  OAI211_X1 U21982 ( .C1(n19806), .C2(n19816), .A(n19805), .B(n19804), .ZN(
        P3_U2876) );
  AOI22_X1 U21983 ( .A1(n19810), .A2(n19809), .B1(n19808), .B2(n19807), .ZN(
        n19815) );
  AOI22_X1 U21984 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19813), .B1(
        n19812), .B2(n19811), .ZN(n19814) );
  OAI211_X1 U21985 ( .C1(n19817), .C2(n19816), .A(n19815), .B(n19814), .ZN(
        P3_U2868) );
  AOI22_X1 U21986 ( .A1(n17542), .A2(n20319), .B1(n20316), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19819) );
  AOI22_X1 U21987 ( .A1(n20317), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n20313), .ZN(n19818) );
  NAND2_X1 U21988 ( .A1(n19819), .A2(n19818), .ZN(P2_U2888) );
  AOI22_X1 U21989 ( .A1(n20064), .A2(n19820), .B1(P2_EAX_REG_15__SCAN_IN), 
        .B2(n20313), .ZN(n19821) );
  OAI21_X1 U21990 ( .B1(n20257), .B2(n19822), .A(n19821), .ZN(P2_U2904) );
  AOI22_X1 U21991 ( .A1(n20064), .A2(n19823), .B1(P2_EAX_REG_13__SCAN_IN), 
        .B2(n20313), .ZN(n19824) );
  OAI21_X1 U21992 ( .B1(n19825), .B2(n20257), .A(n19824), .ZN(P2_U2906) );
  AOI22_X1 U21993 ( .A1(n20064), .A2(n19826), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n20313), .ZN(n19827) );
  OAI21_X1 U21994 ( .B1(n19828), .B2(n20257), .A(n19827), .ZN(P2_U2910) );
  AOI22_X1 U21995 ( .A1(n20064), .A2(n19829), .B1(P2_EAX_REG_7__SCAN_IN), .B2(
        n20313), .ZN(n19830) );
  OAI21_X1 U21996 ( .B1(n19833), .B2(n20257), .A(n19830), .ZN(P2_U2912) );
  OAI21_X1 U21997 ( .B1(n19831), .B2(n20325), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19832) );
  OAI21_X1 U21998 ( .B1(n19845), .B2(n20002), .A(n19832), .ZN(n20326) );
  NOR2_X2 U21999 ( .A1(n19835), .A2(n20261), .ZN(n20016) );
  AOI22_X1 U22000 ( .A1(n20326), .A2(n19834), .B1(n20016), .B2(n20325), .ZN(
        n19842) );
  INV_X1 U22001 ( .A(n19844), .ZN(n19862) );
  INV_X1 U22002 ( .A(n19836), .ZN(n19928) );
  NOR2_X1 U22003 ( .A1(n19862), .A2(n19928), .ZN(n19840) );
  OAI21_X1 U22004 ( .B1(n19846), .B2(n20325), .A(n19932), .ZN(n19837) );
  OAI21_X1 U22005 ( .B1(n13931), .B2(n19941), .A(n19837), .ZN(n19838) );
  OAI21_X1 U22006 ( .B1(n19840), .B2(n19839), .A(n19838), .ZN(n20327) );
  AOI22_X1 U22007 ( .A1(n20264), .A2(BUF2_REG_23__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n20015) );
  AOI22_X1 U22008 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20327), .B1(
        n20430), .B2(n20018), .ZN(n19841) );
  OAI211_X1 U22009 ( .C1(n19979), .C2(n20336), .A(n19842), .B(n19841), .ZN(
        P2_U3175) );
  NOR2_X1 U22010 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19845), .ZN(
        n20330) );
  AOI22_X1 U22011 ( .A1(n20018), .A2(n20210), .B1(n20016), .B2(n20330), .ZN(
        n19857) );
  NAND2_X1 U22012 ( .A1(n20336), .A2(n19846), .ZN(n19848) );
  INV_X1 U22013 ( .A(n19847), .ZN(n19912) );
  OAI21_X1 U22014 ( .B1(n19848), .B2(n20331), .A(n19912), .ZN(n19853) );
  NOR2_X1 U22015 ( .A1(n20000), .A2(n19861), .ZN(n20337) );
  INV_X1 U22016 ( .A(n20337), .ZN(n19863) );
  OR2_X1 U22017 ( .A1(n19851), .A2(n19941), .ZN(n19849) );
  AOI22_X1 U22018 ( .A1(n19853), .A2(n19863), .B1(n19985), .B2(n19849), .ZN(
        n19850) );
  INV_X1 U22019 ( .A(n19853), .ZN(n19855) );
  INV_X1 U22020 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19916) );
  NOR2_X1 U22021 ( .A1(n19851), .A2(n19916), .ZN(n19852) );
  OAI22_X1 U22022 ( .A1(n19853), .A2(P2_STATE2_REG_2__SCAN_IN), .B1(n20330), 
        .B2(n19852), .ZN(n19854) );
  AOI22_X1 U22023 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20333), .B1(
        n19834), .B2(n20332), .ZN(n19856) );
  OAI211_X1 U22024 ( .C1(n19979), .C2(n20343), .A(n19857), .B(n19856), .ZN(
        P2_U3167) );
  OAI21_X1 U22025 ( .B1(n19858), .B2(n20337), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19859) );
  OAI21_X1 U22026 ( .B1(n19861), .B2(n20002), .A(n19859), .ZN(n20338) );
  AOI22_X1 U22027 ( .A1(n20338), .A2(n19834), .B1(n20016), .B2(n20337), .ZN(
        n19868) );
  OR2_X1 U22028 ( .A1(n19860), .A2(n22273), .ZN(n20005) );
  OAI21_X1 U22029 ( .B1(n19862), .B2(n20005), .A(n19861), .ZN(n19866) );
  OAI211_X1 U22030 ( .C1(n19864), .C2(n19941), .A(n19863), .B(n20002), .ZN(
        n19865) );
  NAND3_X1 U22031 ( .A1(n19866), .A2(n19932), .A3(n19865), .ZN(n20340) );
  AOI22_X1 U22032 ( .A1(n20340), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n20331), .B2(n20018), .ZN(n19867) );
  OAI211_X1 U22033 ( .C1(n19979), .C2(n20215), .A(n19868), .B(n19867), .ZN(
        P2_U3159) );
  AOI22_X1 U22034 ( .A1(n20272), .A2(n19834), .B1(n20271), .B2(n20016), .ZN(
        n19871) );
  AOI22_X1 U22035 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20273), .B1(
        n20339), .B2(n20018), .ZN(n19870) );
  OAI211_X1 U22036 ( .C1(n19979), .C2(n20349), .A(n19871), .B(n19870), .ZN(
        P2_U3151) );
  NAND3_X1 U22037 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19884), .ZN(n19885) );
  AND2_X1 U22038 ( .A1(n19884), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19873) );
  NAND2_X1 U22039 ( .A1(n19873), .A2(n19872), .ZN(n19877) );
  INV_X1 U22040 ( .A(n19877), .ZN(n20344) );
  OAI21_X1 U22041 ( .B1(n19874), .B2(n20344), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19875) );
  OAI21_X1 U22042 ( .B1(n19885), .B2(n20002), .A(n19875), .ZN(n20345) );
  AOI22_X1 U22043 ( .A1(n20345), .A2(n19834), .B1(n20344), .B2(n20016), .ZN(
        n19881) );
  OAI21_X1 U22044 ( .B1(n19876), .B2(n19981), .A(n19885), .ZN(n19879) );
  OAI211_X1 U22045 ( .C1(n13924), .C2(n19941), .A(n20002), .B(n19877), .ZN(
        n19878) );
  NAND3_X1 U22046 ( .A1(n19879), .A2(n19932), .A3(n19878), .ZN(n20346) );
  AOI22_X1 U22047 ( .A1(n20172), .A2(n20018), .B1(n20346), .B2(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n19880) );
  OAI211_X1 U22048 ( .C1(n19979), .C2(n20280), .A(n19881), .B(n19880), .ZN(
        P2_U3143) );
  NAND3_X1 U22049 ( .A1(n20356), .A2(n20280), .A3(n14357), .ZN(n19883) );
  NAND2_X1 U22050 ( .A1(n19883), .A2(n19912), .ZN(n19891) );
  NAND3_X1 U22051 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12216), .A3(
        n19884), .ZN(n19911) );
  NOR2_X1 U22052 ( .A1(n20000), .A2(n19911), .ZN(n20357) );
  NOR2_X1 U22053 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19885), .ZN(
        n20350) );
  NOR2_X1 U22054 ( .A1(n20357), .A2(n20350), .ZN(n19894) );
  NAND2_X1 U22055 ( .A1(n19891), .A2(n19894), .ZN(n19890) );
  OR2_X1 U22056 ( .A1(n19886), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19888) );
  NOR2_X1 U22057 ( .A1(n19846), .A2(n20350), .ZN(n19887) );
  AOI21_X1 U22058 ( .B1(n19888), .B2(n19887), .A(n20259), .ZN(n19889) );
  INV_X1 U22059 ( .A(n19979), .ZN(n20017) );
  AOI22_X1 U22060 ( .A1(n20017), .A2(n20358), .B1(n20016), .B2(n20350), .ZN(
        n19897) );
  INV_X1 U22061 ( .A(n19891), .ZN(n19895) );
  OAI21_X1 U22062 ( .B1(n19892), .B2(n20350), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19893) );
  AOI22_X1 U22063 ( .A1(n19834), .A2(n20352), .B1(n20351), .B2(n20018), .ZN(
        n19896) );
  OAI211_X1 U22064 ( .C1(n20175), .C2(n19898), .A(n19897), .B(n19896), .ZN(
        P2_U3135) );
  AOI22_X1 U22065 ( .A1(n20018), .A2(n20358), .B1(n20016), .B2(n20357), .ZN(
        n19909) );
  OAI21_X1 U22066 ( .B1(n19900), .B2(n20005), .A(n19846), .ZN(n19907) );
  INV_X1 U22067 ( .A(n19911), .ZN(n19903) );
  OAI21_X1 U22068 ( .B1(n19846), .B2(n20357), .A(n19932), .ZN(n19901) );
  OAI21_X1 U22069 ( .B1(n19904), .B2(n19941), .A(n19901), .ZN(n19902) );
  OAI21_X1 U22070 ( .B1(n19907), .B2(n19903), .A(n19902), .ZN(n20360) );
  INV_X1 U22071 ( .A(n19904), .ZN(n19905) );
  OAI21_X1 U22072 ( .B1(n19905), .B2(n20357), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19906) );
  AOI22_X1 U22073 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20360), .B1(
        n19834), .B2(n20359), .ZN(n19908) );
  OAI211_X1 U22074 ( .C1(n19979), .C2(n20363), .A(n19909), .B(n19908), .ZN(
        P2_U3127) );
  INV_X1 U22075 ( .A(n19962), .ZN(n19910) );
  NOR2_X1 U22076 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19911), .ZN(
        n20364) );
  AOI22_X1 U22077 ( .A1(n20365), .A2(n20018), .B1(n20016), .B2(n20364), .ZN(
        n19923) );
  NAND2_X1 U22078 ( .A1(n20363), .A2(n19846), .ZN(n19913) );
  OAI21_X1 U22079 ( .B1(n19913), .B2(n20373), .A(n19912), .ZN(n19919) );
  INV_X1 U22080 ( .A(n19919), .ZN(n19921) );
  INV_X1 U22081 ( .A(n19929), .ZN(n20371) );
  NOR2_X1 U22082 ( .A1(n19921), .A2(n20371), .ZN(n19914) );
  AOI211_X1 U22083 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19917), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19914), .ZN(n19915) );
  NOR2_X1 U22084 ( .A1(n19917), .A2(n19916), .ZN(n19918) );
  OAI22_X1 U22085 ( .A1(n19919), .A2(P2_STATE2_REG_2__SCAN_IN), .B1(n20364), 
        .B2(n19918), .ZN(n19920) );
  AOI22_X1 U22086 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n19834), .ZN(n19922) );
  OAI211_X1 U22087 ( .C1(n19979), .C2(n20370), .A(n19923), .B(n19922), .ZN(
        P2_U3119) );
  NAND2_X1 U22088 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n14348), .ZN(
        n19927) );
  OAI21_X1 U22089 ( .B1(n19925), .B2(n20371), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19926) );
  OAI21_X1 U22090 ( .B1(n19927), .B2(n20002), .A(n19926), .ZN(n20372) );
  AOI22_X1 U22091 ( .A1(n20372), .A2(n19834), .B1(n20371), .B2(n20016), .ZN(
        n19935) );
  OAI22_X1 U22092 ( .A1(n19952), .A2(n19928), .B1(n19964), .B2(n12216), .ZN(
        n19933) );
  OAI211_X1 U22093 ( .C1(n19930), .C2(n19941), .A(n20002), .B(n19929), .ZN(
        n19931) );
  NAND3_X1 U22094 ( .A1(n19933), .A2(n19932), .A3(n19931), .ZN(n20374) );
  AOI22_X1 U22095 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20374), .B1(
        n20018), .B2(n20373), .ZN(n19934) );
  OAI211_X1 U22096 ( .C1(n19979), .C2(n20382), .A(n19935), .B(n19934), .ZN(
        P2_U3111) );
  INV_X1 U22097 ( .A(n19942), .ZN(n19937) );
  AND3_X1 U22098 ( .A1(n20000), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        n14348), .ZN(n20377) );
  OAI21_X1 U22099 ( .B1(n19937), .B2(n20377), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19938) );
  OAI21_X1 U22100 ( .B1(n19939), .B2(n19964), .A(n19938), .ZN(n20378) );
  AOI22_X1 U22101 ( .A1(n20378), .A2(n19834), .B1(n20016), .B2(n20377), .ZN(
        n19949) );
  NOR2_X1 U22102 ( .A1(n19846), .A2(n20377), .ZN(n19940) );
  OAI21_X1 U22103 ( .B1(n19942), .B2(n19941), .A(n19940), .ZN(n19947) );
  NAND3_X1 U22104 ( .A1(n19965), .A2(n14348), .A3(n19980), .ZN(n19943) );
  OAI221_X1 U22105 ( .B1(n22273), .B2(n20382), .C1(n22273), .C2(n20393), .A(
        n19943), .ZN(n19944) );
  INV_X1 U22106 ( .A(n19944), .ZN(n19945) );
  NOR2_X1 U22107 ( .A1(n20259), .A2(n19945), .ZN(n19946) );
  NAND2_X1 U22108 ( .A1(n19947), .A2(n19946), .ZN(n20379) );
  AOI22_X1 U22109 ( .A1(n20287), .A2(n20018), .B1(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n20379), .ZN(n19948) );
  OAI211_X1 U22110 ( .C1(n19979), .C2(n20393), .A(n19949), .B(n19948), .ZN(
        P2_U3103) );
  INV_X1 U22111 ( .A(n20393), .ZN(n20290) );
  NAND2_X1 U22112 ( .A1(n14348), .A2(n12216), .ZN(n19958) );
  NOR2_X1 U22113 ( .A1(n20000), .A2(n19958), .ZN(n20386) );
  AOI22_X1 U22114 ( .A1(n20290), .A2(n20018), .B1(n20016), .B2(n20386), .ZN(
        n19961) );
  OAI21_X1 U22115 ( .B1(n19952), .B2(n20005), .A(n19846), .ZN(n19959) );
  INV_X1 U22116 ( .A(n19958), .ZN(n19955) );
  INV_X1 U22117 ( .A(n19985), .ZN(n20007) );
  AOI211_X1 U22118 ( .C1(n19956), .C2(n20008), .A(n20007), .B(n20386), .ZN(
        n19953) );
  NOR2_X1 U22119 ( .A1(n20259), .A2(n19953), .ZN(n19954) );
  OAI21_X1 U22120 ( .B1(n19959), .B2(n19955), .A(n19954), .ZN(n20390) );
  OAI21_X1 U22121 ( .B1(n19956), .B2(n20386), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19957) );
  OAI21_X1 U22122 ( .B1(n19959), .B2(n19958), .A(n19957), .ZN(n20389) );
  AOI22_X1 U22123 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20390), .B1(
        n19834), .B2(n20389), .ZN(n19960) );
  OAI211_X1 U22124 ( .C1(n19979), .C2(n20396), .A(n19961), .B(n19960), .ZN(
        P2_U3095) );
  INV_X1 U22125 ( .A(n20006), .ZN(n19963) );
  NOR2_X1 U22126 ( .A1(n19965), .A2(n19964), .ZN(n20394) );
  AOI22_X1 U22127 ( .A1(n20293), .A2(n20018), .B1(n20016), .B2(n20394), .ZN(
        n19978) );
  OAI21_X1 U22128 ( .B1(n20297), .B2(n20293), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19966) );
  NAND2_X1 U22129 ( .A1(n19966), .A2(n19846), .ZN(n19976) );
  INV_X1 U22130 ( .A(n19967), .ZN(n19968) );
  NAND2_X1 U22131 ( .A1(n19969), .A2(n19968), .ZN(n19975) );
  INV_X1 U22132 ( .A(n19975), .ZN(n19973) );
  AOI211_X1 U22133 ( .C1(n13857), .C2(n20008), .A(n20007), .B(n20394), .ZN(
        n19971) );
  NOR2_X1 U22134 ( .A1(n20259), .A2(n19971), .ZN(n19972) );
  OAI21_X1 U22135 ( .B1(n13857), .B2(n20394), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19974) );
  AOI22_X1 U22136 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20399), .B1(
        n19834), .B2(n20398), .ZN(n19977) );
  OAI211_X1 U22137 ( .C1(n19979), .C2(n20404), .A(n19978), .B(n19977), .ZN(
        P2_U3087) );
  NOR2_X1 U22138 ( .A1(n19980), .A2(n20004), .ZN(n20296) );
  AOI22_X1 U22139 ( .A1(n20017), .A2(n20415), .B1(n20296), .B2(n20016), .ZN(
        n19994) );
  OAI21_X1 U22140 ( .B1(n19982), .B2(n19981), .A(n19846), .ZN(n19992) );
  NOR2_X1 U22141 ( .A1(n12216), .A2(n20004), .ZN(n19988) );
  INV_X1 U22142 ( .A(n20296), .ZN(n20402) );
  NAND2_X1 U22143 ( .A1(n19983), .A2(n20402), .ZN(n19984) );
  OAI21_X1 U22144 ( .B1(n20008), .B2(n20296), .A(n19984), .ZN(n19986) );
  AOI21_X1 U22145 ( .B1(n19986), .B2(n19985), .A(n20259), .ZN(n19987) );
  OAI21_X1 U22146 ( .B1(n19992), .B2(n19988), .A(n19987), .ZN(n20407) );
  INV_X1 U22147 ( .A(n19988), .ZN(n19991) );
  OAI21_X1 U22148 ( .B1(n19989), .B2(n20296), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19990) );
  OAI21_X1 U22149 ( .B1(n19992), .B2(n19991), .A(n19990), .ZN(n20406) );
  AOI22_X1 U22150 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20407), .B1(
        n19834), .B2(n20406), .ZN(n19993) );
  OAI211_X1 U22151 ( .C1(n20015), .C2(n20404), .A(n19994), .B(n19993), .ZN(
        P2_U3079) );
  INV_X1 U22152 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n19997) );
  AOI22_X1 U22153 ( .A1(n20413), .A2(n19834), .B1(n20016), .B2(n20412), .ZN(
        n19996) );
  AOI22_X1 U22154 ( .A1(n20415), .A2(n20018), .B1(n20414), .B2(n20017), .ZN(
        n19995) );
  OAI211_X1 U22155 ( .C1(n20419), .C2(n19997), .A(n19996), .B(n19995), .ZN(
        P2_U3071) );
  INV_X1 U22156 ( .A(n20004), .ZN(n19998) );
  NAND2_X1 U22157 ( .A1(n19998), .A2(n12216), .ZN(n20003) );
  INV_X1 U22158 ( .A(n19999), .ZN(n20009) );
  NOR3_X2 U22159 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20000), .A3(
        n20004), .ZN(n20420) );
  OAI21_X1 U22160 ( .B1(n20009), .B2(n20420), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20001) );
  OAI21_X1 U22161 ( .B1(n20003), .B2(n20002), .A(n20001), .ZN(n20421) );
  AOI22_X1 U22162 ( .A1(n20421), .A2(n19834), .B1(n20016), .B2(n20420), .ZN(
        n20014) );
  OAI22_X1 U22163 ( .A1(n20006), .A2(n20005), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n20004), .ZN(n20012) );
  AOI211_X1 U22164 ( .C1(n20009), .C2(n20008), .A(n20007), .B(n20420), .ZN(
        n20010) );
  NOR2_X1 U22165 ( .A1(n20259), .A2(n20010), .ZN(n20011) );
  NAND2_X1 U22166 ( .A1(n20012), .A2(n20011), .ZN(n20422) );
  AOI22_X1 U22167 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20422), .B1(
        n20432), .B2(n20017), .ZN(n20013) );
  OAI211_X1 U22168 ( .C1(n20015), .C2(n20425), .A(n20014), .B(n20013), .ZN(
        P2_U3063) );
  INV_X1 U22169 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20021) );
  AOI22_X1 U22170 ( .A1(n20017), .A2(n20430), .B1(n20427), .B2(n20016), .ZN(
        n20020) );
  AOI22_X1 U22171 ( .A1(n19834), .A2(n20433), .B1(n20432), .B2(n20018), .ZN(
        n20019) );
  OAI211_X1 U22172 ( .C1(n20438), .C2(n20021), .A(n20020), .B(n20019), .ZN(
        P2_U3055) );
  AOI22_X1 U22173 ( .A1(n20264), .A2(BUF2_REG_30__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n20051) );
  NOR2_X2 U22174 ( .A1(n14353), .A2(n20261), .ZN(n20057) );
  AOI22_X1 U22175 ( .A1(n20326), .A2(n20023), .B1(n20057), .B2(n20325), .ZN(
        n20025) );
  AOI22_X1 U22176 ( .A1(n20264), .A2(BUF2_REG_22__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n20056) );
  AOI22_X1 U22177 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20327), .B1(
        n20430), .B2(n20059), .ZN(n20024) );
  OAI211_X1 U22178 ( .C1(n20051), .C2(n20336), .A(n20025), .B(n20024), .ZN(
        P2_U3174) );
  INV_X1 U22179 ( .A(n20051), .ZN(n20058) );
  AOI22_X1 U22180 ( .A1(n20058), .A2(n20331), .B1(n20057), .B2(n20330), .ZN(
        n20027) );
  AOI22_X1 U22181 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20333), .B1(
        n20023), .B2(n20332), .ZN(n20026) );
  OAI211_X1 U22182 ( .C1(n20056), .C2(n20336), .A(n20027), .B(n20026), .ZN(
        P2_U3166) );
  AOI22_X1 U22183 ( .A1(n20338), .A2(n20023), .B1(n20057), .B2(n20337), .ZN(
        n20029) );
  AOI22_X1 U22184 ( .A1(n20340), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n20059), .B2(n20331), .ZN(n20028) );
  OAI211_X1 U22185 ( .C1(n20051), .C2(n20215), .A(n20029), .B(n20028), .ZN(
        P2_U3158) );
  AOI22_X1 U22186 ( .A1(n20272), .A2(n20023), .B1(n20271), .B2(n20057), .ZN(
        n20031) );
  AOI22_X1 U22187 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20273), .B1(
        n20339), .B2(n20059), .ZN(n20030) );
  OAI211_X1 U22188 ( .C1(n20051), .C2(n20349), .A(n20031), .B(n20030), .ZN(
        P2_U3150) );
  AOI22_X1 U22189 ( .A1(n20345), .A2(n20023), .B1(n20344), .B2(n20057), .ZN(
        n20033) );
  AOI22_X1 U22190 ( .A1(n20058), .A2(n20351), .B1(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n20346), .ZN(n20032) );
  OAI211_X1 U22191 ( .C1(n20056), .C2(n20349), .A(n20033), .B(n20032), .ZN(
        P2_U3142) );
  AOI22_X1 U22192 ( .A1(n20058), .A2(n20358), .B1(n20057), .B2(n20350), .ZN(
        n20035) );
  AOI22_X1 U22193 ( .A1(n20023), .A2(n20352), .B1(n20351), .B2(n20059), .ZN(
        n20034) );
  OAI211_X1 U22194 ( .C1(n20175), .C2(n20036), .A(n20035), .B(n20034), .ZN(
        P2_U3134) );
  AOI22_X1 U22195 ( .A1(n20059), .A2(n20358), .B1(n20057), .B2(n20357), .ZN(
        n20038) );
  AOI22_X1 U22196 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20360), .B1(
        n20023), .B2(n20359), .ZN(n20037) );
  OAI211_X1 U22197 ( .C1(n20051), .C2(n20363), .A(n20038), .B(n20037), .ZN(
        P2_U3126) );
  AOI22_X1 U22198 ( .A1(n20365), .A2(n20059), .B1(n20057), .B2(n20364), .ZN(
        n20040) );
  AOI22_X1 U22199 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20023), .ZN(n20039) );
  OAI211_X1 U22200 ( .C1(n20051), .C2(n20370), .A(n20040), .B(n20039), .ZN(
        P2_U3118) );
  AOI22_X1 U22201 ( .A1(n20372), .A2(n20023), .B1(n20371), .B2(n20057), .ZN(
        n20042) );
  AOI22_X1 U22202 ( .A1(n20058), .A2(n20287), .B1(
        P2_INSTQUEUE_REG_7__6__SCAN_IN), .B2(n20374), .ZN(n20041) );
  OAI211_X1 U22203 ( .C1(n20056), .C2(n20370), .A(n20042), .B(n20041), .ZN(
        P2_U3110) );
  AOI22_X1 U22204 ( .A1(n20378), .A2(n20023), .B1(n20057), .B2(n20377), .ZN(
        n20044) );
  AOI22_X1 U22205 ( .A1(n20059), .A2(n20287), .B1(
        P2_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n20379), .ZN(n20043) );
  OAI211_X1 U22206 ( .C1(n20051), .C2(n20393), .A(n20044), .B(n20043), .ZN(
        P2_U3102) );
  AOI22_X1 U22207 ( .A1(n20058), .A2(n20293), .B1(n20057), .B2(n20386), .ZN(
        n20046) );
  AOI22_X1 U22208 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20390), .B1(
        n20023), .B2(n20389), .ZN(n20045) );
  OAI211_X1 U22209 ( .C1(n20056), .C2(n20393), .A(n20046), .B(n20045), .ZN(
        P2_U3094) );
  AOI22_X1 U22210 ( .A1(n20059), .A2(n20293), .B1(n20057), .B2(n20394), .ZN(
        n20048) );
  AOI22_X1 U22211 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20399), .B1(
        n20023), .B2(n20398), .ZN(n20047) );
  OAI211_X1 U22212 ( .C1(n20051), .C2(n20404), .A(n20048), .B(n20047), .ZN(
        P2_U3086) );
  INV_X1 U22213 ( .A(n20415), .ZN(n20410) );
  AOI22_X1 U22214 ( .A1(n20059), .A2(n20297), .B1(n20296), .B2(n20057), .ZN(
        n20050) );
  AOI22_X1 U22215 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20407), .B1(
        n20023), .B2(n20406), .ZN(n20049) );
  OAI211_X1 U22216 ( .C1(n20051), .C2(n20410), .A(n20050), .B(n20049), .ZN(
        P2_U3078) );
  AOI22_X1 U22217 ( .A1(n20413), .A2(n20023), .B1(n20057), .B2(n20412), .ZN(
        n20053) );
  AOI22_X1 U22218 ( .A1(n20415), .A2(n20059), .B1(n20414), .B2(n20058), .ZN(
        n20052) );
  OAI211_X1 U22219 ( .C1(n20419), .C2(n14462), .A(n20053), .B(n20052), .ZN(
        P2_U3070) );
  AOI22_X1 U22220 ( .A1(n20421), .A2(n20023), .B1(n20057), .B2(n20420), .ZN(
        n20055) );
  AOI22_X1 U22221 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20422), .B1(
        n20432), .B2(n20058), .ZN(n20054) );
  OAI211_X1 U22222 ( .C1(n20056), .C2(n20425), .A(n20055), .B(n20054), .ZN(
        P2_U3062) );
  AOI22_X1 U22223 ( .A1(n20058), .A2(n20430), .B1(n20427), .B2(n20057), .ZN(
        n20061) );
  AOI22_X1 U22224 ( .A1(n20023), .A2(n20433), .B1(n20432), .B2(n20059), .ZN(
        n20060) );
  OAI211_X1 U22225 ( .C1(n20438), .C2(n20062), .A(n20061), .B(n20060), .ZN(
        P2_U3054) );
  AOI22_X1 U22226 ( .A1(n20064), .A2(n20063), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n20313), .ZN(n20068) );
  NAND3_X1 U22227 ( .A1(n20066), .A2(n20065), .A3(n20320), .ZN(n20067) );
  OAI211_X1 U22228 ( .C1(n20069), .C2(n20257), .A(n20068), .B(n20067), .ZN(
        P2_U2914) );
  AOI22_X1 U22229 ( .A1(n20264), .A2(BUF2_REG_29__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n20095) );
  NOR2_X2 U22230 ( .A1(n11843), .A2(n20261), .ZN(n20103) );
  AOI22_X1 U22231 ( .A1(n20326), .A2(n20070), .B1(n20103), .B2(n20325), .ZN(
        n20072) );
  AOI22_X1 U22232 ( .A1(n20264), .A2(BUF2_REG_21__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n20102) );
  AOI22_X1 U22233 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20327), .B1(
        n20430), .B2(n20105), .ZN(n20071) );
  OAI211_X1 U22234 ( .C1(n20095), .C2(n20336), .A(n20072), .B(n20071), .ZN(
        P2_U3173) );
  INV_X1 U22235 ( .A(n20095), .ZN(n20104) );
  AOI22_X1 U22236 ( .A1(n20104), .A2(n20331), .B1(n20103), .B2(n20330), .ZN(
        n20074) );
  AOI22_X1 U22237 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20333), .B1(
        n20070), .B2(n20332), .ZN(n20073) );
  OAI211_X1 U22238 ( .C1(n20102), .C2(n20336), .A(n20074), .B(n20073), .ZN(
        P2_U3165) );
  AOI22_X1 U22239 ( .A1(n20338), .A2(n20070), .B1(n20103), .B2(n20337), .ZN(
        n20076) );
  AOI22_X1 U22240 ( .A1(n20340), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n20105), .B2(n20331), .ZN(n20075) );
  OAI211_X1 U22241 ( .C1(n20095), .C2(n20215), .A(n20076), .B(n20075), .ZN(
        P2_U3157) );
  AOI22_X1 U22242 ( .A1(n20272), .A2(n20070), .B1(n20271), .B2(n20103), .ZN(
        n20078) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20273), .B1(
        n20339), .B2(n20105), .ZN(n20077) );
  OAI211_X1 U22244 ( .C1(n20095), .C2(n20349), .A(n20078), .B(n20077), .ZN(
        P2_U3149) );
  AOI22_X1 U22245 ( .A1(n20345), .A2(n20070), .B1(n20344), .B2(n20103), .ZN(
        n20080) );
  AOI22_X1 U22246 ( .A1(n20105), .A2(n20172), .B1(n20346), .B2(
        P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n20079) );
  OAI211_X1 U22247 ( .C1(n20095), .C2(n20280), .A(n20080), .B(n20079), .ZN(
        P2_U3141) );
  AOI22_X1 U22248 ( .A1(n20105), .A2(n20351), .B1(n20103), .B2(n20350), .ZN(
        n20082) );
  AOI22_X1 U22249 ( .A1(n20070), .A2(n20352), .B1(n20358), .B2(n20104), .ZN(
        n20081) );
  OAI211_X1 U22250 ( .C1(n20175), .C2(n13933), .A(n20082), .B(n20081), .ZN(
        P2_U3133) );
  AOI22_X1 U22251 ( .A1(n20104), .A2(n20365), .B1(n20103), .B2(n20357), .ZN(
        n20084) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20360), .B1(
        n20070), .B2(n20359), .ZN(n20083) );
  OAI211_X1 U22253 ( .C1(n20102), .C2(n20356), .A(n20084), .B(n20083), .ZN(
        P2_U3125) );
  AOI22_X1 U22254 ( .A1(n20105), .A2(n20365), .B1(n20103), .B2(n20364), .ZN(
        n20086) );
  AOI22_X1 U22255 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20070), .ZN(n20085) );
  OAI211_X1 U22256 ( .C1(n20095), .C2(n20370), .A(n20086), .B(n20085), .ZN(
        P2_U3117) );
  AOI22_X1 U22257 ( .A1(n20372), .A2(n20070), .B1(n20371), .B2(n20103), .ZN(
        n20088) );
  AOI22_X1 U22258 ( .A1(n20104), .A2(n20287), .B1(n20374), .B2(
        P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n20087) );
  OAI211_X1 U22259 ( .C1(n20102), .C2(n20370), .A(n20088), .B(n20087), .ZN(
        P2_U3109) );
  AOI22_X1 U22260 ( .A1(n20378), .A2(n20070), .B1(n20103), .B2(n20377), .ZN(
        n20090) );
  AOI22_X1 U22261 ( .A1(n20105), .A2(n20287), .B1(
        P2_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n20379), .ZN(n20089) );
  OAI211_X1 U22262 ( .C1(n20095), .C2(n20393), .A(n20090), .B(n20089), .ZN(
        P2_U3101) );
  AOI22_X1 U22263 ( .A1(n20104), .A2(n20293), .B1(n20103), .B2(n20386), .ZN(
        n20092) );
  AOI22_X1 U22264 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20390), .B1(
        n20070), .B2(n20389), .ZN(n20091) );
  OAI211_X1 U22265 ( .C1(n20102), .C2(n20393), .A(n20092), .B(n20091), .ZN(
        P2_U3093) );
  AOI22_X1 U22266 ( .A1(n20105), .A2(n20293), .B1(n20103), .B2(n20394), .ZN(
        n20094) );
  AOI22_X1 U22267 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20399), .B1(
        n20070), .B2(n20398), .ZN(n20093) );
  OAI211_X1 U22268 ( .C1(n20095), .C2(n20404), .A(n20094), .B(n20093), .ZN(
        P2_U3085) );
  AOI22_X1 U22269 ( .A1(n20104), .A2(n20415), .B1(n20296), .B2(n20103), .ZN(
        n20097) );
  AOI22_X1 U22270 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20407), .B1(
        n20070), .B2(n20406), .ZN(n20096) );
  OAI211_X1 U22271 ( .C1(n20102), .C2(n20404), .A(n20097), .B(n20096), .ZN(
        P2_U3077) );
  AOI22_X1 U22272 ( .A1(n20413), .A2(n20070), .B1(n20103), .B2(n20412), .ZN(
        n20099) );
  AOI22_X1 U22273 ( .A1(n20415), .A2(n20105), .B1(n20414), .B2(n20104), .ZN(
        n20098) );
  OAI211_X1 U22274 ( .C1(n20419), .C2(n13948), .A(n20099), .B(n20098), .ZN(
        P2_U3069) );
  AOI22_X1 U22275 ( .A1(n20421), .A2(n20070), .B1(n20103), .B2(n20420), .ZN(
        n20101) );
  AOI22_X1 U22276 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20422), .B1(
        n20432), .B2(n20104), .ZN(n20100) );
  OAI211_X1 U22277 ( .C1(n20102), .C2(n20425), .A(n20101), .B(n20100), .ZN(
        P2_U3061) );
  AOI22_X1 U22278 ( .A1(n20104), .A2(n20430), .B1(n20427), .B2(n20103), .ZN(
        n20107) );
  AOI22_X1 U22279 ( .A1(n20070), .A2(n20433), .B1(n20432), .B2(n20105), .ZN(
        n20106) );
  OAI211_X1 U22280 ( .C1(n20438), .C2(n20108), .A(n20107), .B(n20106), .ZN(
        P2_U3053) );
  AOI22_X1 U22281 ( .A1(n20264), .A2(BUF2_REG_28__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n20138) );
  INV_X1 U22282 ( .A(n20109), .ZN(n20110) );
  NOR2_X2 U22283 ( .A1(n20112), .A2(n20261), .ZN(n20147) );
  AOI22_X1 U22284 ( .A1(n20326), .A2(n20111), .B1(n20147), .B2(n20325), .ZN(
        n20114) );
  AOI22_X1 U22285 ( .A1(n20264), .A2(BUF2_REG_20__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n20146) );
  AOI22_X1 U22286 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20327), .B1(
        n20430), .B2(n20149), .ZN(n20113) );
  OAI211_X1 U22287 ( .C1(n20138), .C2(n20336), .A(n20114), .B(n20113), .ZN(
        P2_U3172) );
  INV_X1 U22288 ( .A(n20138), .ZN(n20148) );
  AOI22_X1 U22289 ( .A1(n20148), .A2(n20331), .B1(n20147), .B2(n20330), .ZN(
        n20116) );
  AOI22_X1 U22290 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20333), .B1(
        n20111), .B2(n20332), .ZN(n20115) );
  OAI211_X1 U22291 ( .C1(n20146), .C2(n20336), .A(n20116), .B(n20115), .ZN(
        P2_U3164) );
  AOI22_X1 U22292 ( .A1(n20338), .A2(n20111), .B1(n20147), .B2(n20337), .ZN(
        n20118) );
  AOI22_X1 U22293 ( .A1(n20340), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n20149), .B2(n20331), .ZN(n20117) );
  OAI211_X1 U22294 ( .C1(n20138), .C2(n20215), .A(n20118), .B(n20117), .ZN(
        P2_U3156) );
  AOI22_X1 U22295 ( .A1(n20272), .A2(n20111), .B1(n20271), .B2(n20147), .ZN(
        n20120) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20273), .B1(
        n20339), .B2(n20149), .ZN(n20119) );
  OAI211_X1 U22297 ( .C1(n20138), .C2(n20349), .A(n20120), .B(n20119), .ZN(
        P2_U3148) );
  AOI22_X1 U22298 ( .A1(n20345), .A2(n20111), .B1(n20344), .B2(n20147), .ZN(
        n20122) );
  AOI22_X1 U22299 ( .A1(n20148), .A2(n20351), .B1(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n20346), .ZN(n20121) );
  OAI211_X1 U22300 ( .C1(n20146), .C2(n20349), .A(n20122), .B(n20121), .ZN(
        P2_U3140) );
  INV_X1 U22301 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n20125) );
  AOI22_X1 U22302 ( .A1(n20149), .A2(n20351), .B1(n20147), .B2(n20350), .ZN(
        n20124) );
  AOI22_X1 U22303 ( .A1(n20111), .A2(n20352), .B1(n20358), .B2(n20148), .ZN(
        n20123) );
  OAI211_X1 U22304 ( .C1(n20175), .C2(n20125), .A(n20124), .B(n20123), .ZN(
        P2_U3132) );
  AOI22_X1 U22305 ( .A1(n20149), .A2(n20358), .B1(n20147), .B2(n20357), .ZN(
        n20127) );
  AOI22_X1 U22306 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20360), .B1(
        n20111), .B2(n20359), .ZN(n20126) );
  OAI211_X1 U22307 ( .C1(n20138), .C2(n20363), .A(n20127), .B(n20126), .ZN(
        P2_U3124) );
  AOI22_X1 U22308 ( .A1(n20148), .A2(n20373), .B1(n20147), .B2(n20364), .ZN(
        n20129) );
  AOI22_X1 U22309 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20111), .ZN(n20128) );
  OAI211_X1 U22310 ( .C1(n20146), .C2(n20363), .A(n20129), .B(n20128), .ZN(
        P2_U3116) );
  AOI22_X1 U22311 ( .A1(n20372), .A2(n20111), .B1(n20371), .B2(n20147), .ZN(
        n20131) );
  AOI22_X1 U22312 ( .A1(n20149), .A2(n20373), .B1(n20374), .B2(
        P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n20130) );
  OAI211_X1 U22313 ( .C1(n20138), .C2(n20382), .A(n20131), .B(n20130), .ZN(
        P2_U3108) );
  AOI22_X1 U22314 ( .A1(n20378), .A2(n20111), .B1(n20147), .B2(n20377), .ZN(
        n20133) );
  AOI22_X1 U22315 ( .A1(n20149), .A2(n20287), .B1(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n20379), .ZN(n20132) );
  OAI211_X1 U22316 ( .C1(n20138), .C2(n20393), .A(n20133), .B(n20132), .ZN(
        P2_U3100) );
  AOI22_X1 U22317 ( .A1(n20148), .A2(n20293), .B1(n20147), .B2(n20386), .ZN(
        n20135) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20390), .B1(
        n20111), .B2(n20389), .ZN(n20134) );
  OAI211_X1 U22319 ( .C1(n20146), .C2(n20393), .A(n20135), .B(n20134), .ZN(
        P2_U3092) );
  AOI22_X1 U22320 ( .A1(n20149), .A2(n20293), .B1(n20147), .B2(n20394), .ZN(
        n20137) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20399), .B1(
        n20111), .B2(n20398), .ZN(n20136) );
  OAI211_X1 U22322 ( .C1(n20138), .C2(n20404), .A(n20137), .B(n20136), .ZN(
        P2_U3084) );
  AOI22_X1 U22323 ( .A1(n20148), .A2(n20415), .B1(n20296), .B2(n20147), .ZN(
        n20140) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20407), .B1(
        n20111), .B2(n20406), .ZN(n20139) );
  OAI211_X1 U22325 ( .C1(n20146), .C2(n20404), .A(n20140), .B(n20139), .ZN(
        P2_U3076) );
  INV_X1 U22326 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n20143) );
  AOI22_X1 U22327 ( .A1(n20413), .A2(n20111), .B1(n20147), .B2(n20412), .ZN(
        n20142) );
  AOI22_X1 U22328 ( .A1(n20414), .A2(n20148), .B1(n20415), .B2(n20149), .ZN(
        n20141) );
  OAI211_X1 U22329 ( .C1(n20419), .C2(n20143), .A(n20142), .B(n20141), .ZN(
        P2_U3068) );
  AOI22_X1 U22330 ( .A1(n20421), .A2(n20111), .B1(n20147), .B2(n20420), .ZN(
        n20145) );
  AOI22_X1 U22331 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20422), .B1(
        n20432), .B2(n20148), .ZN(n20144) );
  OAI211_X1 U22332 ( .C1(n20146), .C2(n20425), .A(n20145), .B(n20144), .ZN(
        P2_U3060) );
  INV_X1 U22333 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20152) );
  AOI22_X1 U22334 ( .A1(n20148), .A2(n20430), .B1(n20427), .B2(n20147), .ZN(
        n20151) );
  AOI22_X1 U22335 ( .A1(n20111), .A2(n20433), .B1(n20432), .B2(n20149), .ZN(
        n20150) );
  OAI211_X1 U22336 ( .C1(n20438), .C2(n20152), .A(n20151), .B(n20150), .ZN(
        P2_U3052) );
  OAI22_X1 U22337 ( .A1(n20155), .A2(n20154), .B1(n20153), .B2(n18056), .ZN(
        n20156) );
  INV_X1 U22338 ( .A(n20156), .ZN(n20162) );
  AOI21_X1 U22339 ( .B1(n20159), .B2(n20158), .A(n20157), .ZN(n20160) );
  OR2_X1 U22340 ( .A1(n20160), .A2(n20253), .ZN(n20161) );
  OAI211_X1 U22341 ( .C1(n20163), .C2(n20257), .A(n20162), .B(n20161), .ZN(
        P2_U2916) );
  AOI22_X1 U22342 ( .A1(n20326), .A2(n16029), .B1(n20194), .B2(n20325), .ZN(
        n20165) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20327), .B1(
        n20430), .B2(n20188), .ZN(n20164) );
  OAI211_X1 U22344 ( .C1(n20191), .C2(n20336), .A(n20165), .B(n20164), .ZN(
        P2_U3171) );
  AOI22_X1 U22345 ( .A1(n20195), .A2(n20331), .B1(n20194), .B2(n20330), .ZN(
        n20167) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20333), .B1(
        n16029), .B2(n20332), .ZN(n20166) );
  OAI211_X1 U22347 ( .C1(n20198), .C2(n20336), .A(n20167), .B(n20166), .ZN(
        P2_U3163) );
  AOI22_X1 U22348 ( .A1(n20338), .A2(n16029), .B1(n20194), .B2(n20337), .ZN(
        n20169) );
  AOI22_X1 U22349 ( .A1(n20340), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n20188), .B2(n20331), .ZN(n20168) );
  OAI211_X1 U22350 ( .C1(n20191), .C2(n20215), .A(n20169), .B(n20168), .ZN(
        P2_U3155) );
  AOI22_X1 U22351 ( .A1(n20272), .A2(n16029), .B1(n20271), .B2(n20194), .ZN(
        n20171) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20273), .B1(
        n20339), .B2(n20188), .ZN(n20170) );
  OAI211_X1 U22353 ( .C1(n20191), .C2(n20349), .A(n20171), .B(n20170), .ZN(
        P2_U3147) );
  AOI22_X1 U22354 ( .A1(n20345), .A2(n16029), .B1(n20194), .B2(n20344), .ZN(
        n20174) );
  AOI22_X1 U22355 ( .A1(n20188), .A2(n20172), .B1(n20346), .B2(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n20173) );
  OAI211_X1 U22356 ( .C1(n20191), .C2(n20280), .A(n20174), .B(n20173), .ZN(
        P2_U3139) );
  AOI22_X1 U22357 ( .A1(n20195), .A2(n20358), .B1(n20194), .B2(n20350), .ZN(
        n20177) );
  AOI22_X1 U22358 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20353), .B1(
        n16029), .B2(n20352), .ZN(n20176) );
  OAI211_X1 U22359 ( .C1(n20198), .C2(n20280), .A(n20177), .B(n20176), .ZN(
        P2_U3131) );
  AOI22_X1 U22360 ( .A1(n20188), .A2(n20358), .B1(n20194), .B2(n20357), .ZN(
        n20179) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20360), .B1(
        n16029), .B2(n20359), .ZN(n20178) );
  OAI211_X1 U22362 ( .C1(n20191), .C2(n20363), .A(n20179), .B(n20178), .ZN(
        P2_U3123) );
  AOI22_X1 U22363 ( .A1(n20195), .A2(n20373), .B1(n20194), .B2(n20364), .ZN(
        n20181) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n16029), .ZN(n20180) );
  OAI211_X1 U22365 ( .C1(n20198), .C2(n20363), .A(n20181), .B(n20180), .ZN(
        P2_U3115) );
  AOI22_X1 U22366 ( .A1(n20372), .A2(n16029), .B1(n20371), .B2(n20194), .ZN(
        n20183) );
  AOI22_X1 U22367 ( .A1(n20195), .A2(n20287), .B1(
        P2_INSTQUEUE_REG_7__3__SCAN_IN), .B2(n20374), .ZN(n20182) );
  OAI211_X1 U22368 ( .C1(n20198), .C2(n20370), .A(n20183), .B(n20182), .ZN(
        P2_U3107) );
  AOI22_X1 U22369 ( .A1(n20378), .A2(n16029), .B1(n20194), .B2(n20377), .ZN(
        n20185) );
  AOI22_X1 U22370 ( .A1(n20188), .A2(n20287), .B1(
        P2_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n20379), .ZN(n20184) );
  OAI211_X1 U22371 ( .C1(n20191), .C2(n20393), .A(n20185), .B(n20184), .ZN(
        P2_U3099) );
  AOI22_X1 U22372 ( .A1(n20188), .A2(n20290), .B1(n20194), .B2(n20386), .ZN(
        n20187) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20390), .B1(
        n16029), .B2(n20389), .ZN(n20186) );
  OAI211_X1 U22374 ( .C1(n20191), .C2(n20396), .A(n20187), .B(n20186), .ZN(
        P2_U3091) );
  AOI22_X1 U22375 ( .A1(n20188), .A2(n20293), .B1(n20194), .B2(n20394), .ZN(
        n20190) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20399), .B1(
        n16029), .B2(n20398), .ZN(n20189) );
  OAI211_X1 U22377 ( .C1(n20191), .C2(n20404), .A(n20190), .B(n20189), .ZN(
        P2_U3083) );
  AOI22_X1 U22378 ( .A1(n20195), .A2(n20415), .B1(n20194), .B2(n20296), .ZN(
        n20193) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20407), .B1(
        n16029), .B2(n20406), .ZN(n20192) );
  OAI211_X1 U22380 ( .C1(n20198), .C2(n20404), .A(n20193), .B(n20192), .ZN(
        P2_U3075) );
  AOI22_X1 U22381 ( .A1(n20421), .A2(n16029), .B1(n20194), .B2(n20420), .ZN(
        n20197) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20422), .B1(
        n20432), .B2(n20195), .ZN(n20196) );
  OAI211_X1 U22383 ( .C1(n20198), .C2(n20425), .A(n20197), .B(n20196), .ZN(
        P2_U3059) );
  AOI22_X1 U22384 ( .A1(n20199), .A2(n20319), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n20313), .ZN(n20204) );
  XNOR2_X1 U22385 ( .A(n20201), .B(n20200), .ZN(n20202) );
  NAND2_X1 U22386 ( .A1(n20202), .A2(n20320), .ZN(n20203) );
  OAI211_X1 U22387 ( .C1(n20205), .C2(n20257), .A(n20204), .B(n20203), .ZN(
        P2_U2917) );
  NOR2_X2 U22388 ( .A1(n20207), .A2(n20261), .ZN(n20243) );
  AOI22_X1 U22389 ( .A1(n20326), .A2(n20206), .B1(n20243), .B2(n20325), .ZN(
        n20209) );
  AOI22_X1 U22390 ( .A1(n20264), .A2(BUF2_REG_18__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n20242) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20327), .B1(
        n20430), .B2(n20245), .ZN(n20208) );
  OAI211_X1 U22392 ( .C1(n20236), .C2(n20336), .A(n20209), .B(n20208), .ZN(
        P2_U3170) );
  AOI22_X1 U22393 ( .A1(n20245), .A2(n20210), .B1(n20243), .B2(n20330), .ZN(
        n20212) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20333), .B1(
        n20206), .B2(n20332), .ZN(n20211) );
  OAI211_X1 U22395 ( .C1(n20236), .C2(n20343), .A(n20212), .B(n20211), .ZN(
        P2_U3162) );
  AOI22_X1 U22396 ( .A1(n20338), .A2(n20206), .B1(n20243), .B2(n20337), .ZN(
        n20214) );
  AOI22_X1 U22397 ( .A1(n20340), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n20331), .B2(n20245), .ZN(n20213) );
  OAI211_X1 U22398 ( .C1(n20236), .C2(n20215), .A(n20214), .B(n20213), .ZN(
        P2_U3154) );
  AOI22_X1 U22399 ( .A1(n20272), .A2(n20206), .B1(n20271), .B2(n20243), .ZN(
        n20217) );
  AOI22_X1 U22400 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20273), .B1(
        n20339), .B2(n20245), .ZN(n20216) );
  OAI211_X1 U22401 ( .C1(n20236), .C2(n20349), .A(n20217), .B(n20216), .ZN(
        P2_U3146) );
  AOI22_X1 U22402 ( .A1(n20345), .A2(n20206), .B1(n20344), .B2(n20243), .ZN(
        n20219) );
  INV_X1 U22403 ( .A(n20236), .ZN(n20244) );
  AOI22_X1 U22404 ( .A1(n20244), .A2(n20351), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n20346), .ZN(n20218) );
  OAI211_X1 U22405 ( .C1(n20242), .C2(n20349), .A(n20219), .B(n20218), .ZN(
        P2_U3138) );
  AOI22_X1 U22406 ( .A1(n20245), .A2(n20351), .B1(n20243), .B2(n20350), .ZN(
        n20221) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20353), .B1(
        n20206), .B2(n20352), .ZN(n20220) );
  OAI211_X1 U22408 ( .C1(n20236), .C2(n20356), .A(n20221), .B(n20220), .ZN(
        P2_U3130) );
  AOI22_X1 U22409 ( .A1(n20245), .A2(n20358), .B1(n20243), .B2(n20357), .ZN(
        n20223) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20360), .B1(
        n20206), .B2(n20359), .ZN(n20222) );
  OAI211_X1 U22411 ( .C1(n20236), .C2(n20363), .A(n20223), .B(n20222), .ZN(
        P2_U3122) );
  AOI22_X1 U22412 ( .A1(n20365), .A2(n20245), .B1(n20243), .B2(n20364), .ZN(
        n20225) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20206), .ZN(n20224) );
  OAI211_X1 U22414 ( .C1(n20236), .C2(n20370), .A(n20225), .B(n20224), .ZN(
        P2_U3114) );
  AOI22_X1 U22415 ( .A1(n20372), .A2(n20206), .B1(n20371), .B2(n20243), .ZN(
        n20227) );
  AOI22_X1 U22416 ( .A1(n20373), .A2(n20245), .B1(n20374), .B2(
        P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n20226) );
  OAI211_X1 U22417 ( .C1(n20236), .C2(n20382), .A(n20227), .B(n20226), .ZN(
        P2_U3106) );
  AOI22_X1 U22418 ( .A1(n20378), .A2(n20206), .B1(n20243), .B2(n20377), .ZN(
        n20229) );
  AOI22_X1 U22419 ( .A1(n20245), .A2(n20287), .B1(
        P2_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n20379), .ZN(n20228) );
  OAI211_X1 U22420 ( .C1(n20236), .C2(n20393), .A(n20229), .B(n20228), .ZN(
        P2_U3098) );
  AOI22_X1 U22421 ( .A1(n20244), .A2(n20293), .B1(n20243), .B2(n20386), .ZN(
        n20231) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20390), .B1(
        n20206), .B2(n20389), .ZN(n20230) );
  OAI211_X1 U22423 ( .C1(n20242), .C2(n20393), .A(n20231), .B(n20230), .ZN(
        P2_U3090) );
  AOI22_X1 U22424 ( .A1(n20245), .A2(n20293), .B1(n20243), .B2(n20394), .ZN(
        n20233) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20399), .B1(
        n20206), .B2(n20398), .ZN(n20232) );
  OAI211_X1 U22426 ( .C1(n20236), .C2(n20404), .A(n20233), .B(n20232), .ZN(
        P2_U3082) );
  AOI22_X1 U22427 ( .A1(n20297), .A2(n20245), .B1(n20296), .B2(n20243), .ZN(
        n20235) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20407), .B1(
        n20206), .B2(n20406), .ZN(n20234) );
  OAI211_X1 U22429 ( .C1(n20236), .C2(n20410), .A(n20235), .B(n20234), .ZN(
        P2_U3074) );
  INV_X1 U22430 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n20239) );
  AOI22_X1 U22431 ( .A1(n20413), .A2(n20206), .B1(n20243), .B2(n20412), .ZN(
        n20238) );
  AOI22_X1 U22432 ( .A1(n20415), .A2(n20245), .B1(n20414), .B2(n20244), .ZN(
        n20237) );
  OAI211_X1 U22433 ( .C1(n20419), .C2(n20239), .A(n20238), .B(n20237), .ZN(
        P2_U3066) );
  AOI22_X1 U22434 ( .A1(n20421), .A2(n20206), .B1(n20243), .B2(n20420), .ZN(
        n20241) );
  AOI22_X1 U22435 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20422), .B1(
        n20432), .B2(n20244), .ZN(n20240) );
  OAI211_X1 U22436 ( .C1(n20242), .C2(n20425), .A(n20241), .B(n20240), .ZN(
        P2_U3058) );
  AOI22_X1 U22437 ( .A1(n20244), .A2(n20430), .B1(n20427), .B2(n20243), .ZN(
        n20247) );
  AOI22_X1 U22438 ( .A1(n20206), .A2(n20433), .B1(n20432), .B2(n20245), .ZN(
        n20246) );
  OAI211_X1 U22439 ( .C1(n20438), .C2(n20248), .A(n20247), .B(n20246), .ZN(
        P2_U3050) );
  AOI22_X1 U22440 ( .A1(n20319), .A2(n20249), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n20313), .ZN(n20256) );
  AOI21_X1 U22441 ( .B1(n20252), .B2(n20251), .A(n20250), .ZN(n20254) );
  OR2_X1 U22442 ( .A1(n20254), .A2(n20253), .ZN(n20255) );
  OAI211_X1 U22443 ( .C1(n20258), .C2(n20257), .A(n20256), .B(n20255), .ZN(
        P2_U2918) );
  AOI22_X1 U22444 ( .A1(n20264), .A2(BUF2_REG_25__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n20300) );
  NOR2_X2 U22445 ( .A1(n14120), .A2(n20261), .ZN(n20307) );
  AOI22_X1 U22446 ( .A1(n20326), .A2(n20260), .B1(n20307), .B2(n20325), .ZN(
        n20266) );
  AOI22_X1 U22447 ( .A1(n20264), .A2(BUF2_REG_17__SCAN_IN), .B1(n20263), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n20306) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20327), .B1(
        n20430), .B2(n20309), .ZN(n20265) );
  OAI211_X1 U22449 ( .C1(n20300), .C2(n20336), .A(n20266), .B(n20265), .ZN(
        P2_U3169) );
  INV_X1 U22450 ( .A(n20300), .ZN(n20308) );
  AOI22_X1 U22451 ( .A1(n20308), .A2(n20331), .B1(n20307), .B2(n20330), .ZN(
        n20268) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20333), .B1(
        n20260), .B2(n20332), .ZN(n20267) );
  OAI211_X1 U22453 ( .C1(n20306), .C2(n20336), .A(n20268), .B(n20267), .ZN(
        P2_U3161) );
  AOI22_X1 U22454 ( .A1(n20338), .A2(n20260), .B1(n20307), .B2(n20337), .ZN(
        n20270) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20340), .B1(
        n20308), .B2(n20339), .ZN(n20269) );
  OAI211_X1 U22456 ( .C1(n20306), .C2(n20343), .A(n20270), .B(n20269), .ZN(
        P2_U3153) );
  AOI22_X1 U22457 ( .A1(n20272), .A2(n20260), .B1(n20271), .B2(n20307), .ZN(
        n20275) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20273), .B1(
        n20339), .B2(n20309), .ZN(n20274) );
  OAI211_X1 U22459 ( .C1(n20300), .C2(n20349), .A(n20275), .B(n20274), .ZN(
        P2_U3145) );
  AOI22_X1 U22460 ( .A1(n20345), .A2(n20260), .B1(n20344), .B2(n20307), .ZN(
        n20277) );
  AOI22_X1 U22461 ( .A1(n20308), .A2(n20351), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n20346), .ZN(n20276) );
  OAI211_X1 U22462 ( .C1(n20306), .C2(n20349), .A(n20277), .B(n20276), .ZN(
        P2_U3137) );
  AOI22_X1 U22463 ( .A1(n20308), .A2(n20358), .B1(n20307), .B2(n20350), .ZN(
        n20279) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20353), .B1(
        n20260), .B2(n20352), .ZN(n20278) );
  OAI211_X1 U22465 ( .C1(n20306), .C2(n20280), .A(n20279), .B(n20278), .ZN(
        P2_U3129) );
  AOI22_X1 U22466 ( .A1(n20309), .A2(n20358), .B1(n20307), .B2(n20357), .ZN(
        n20282) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20360), .B1(
        n20260), .B2(n20359), .ZN(n20281) );
  OAI211_X1 U22468 ( .C1(n20300), .C2(n20363), .A(n20282), .B(n20281), .ZN(
        P2_U3121) );
  AOI22_X1 U22469 ( .A1(n20308), .A2(n20373), .B1(n20307), .B2(n20364), .ZN(
        n20284) );
  AOI22_X1 U22470 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20260), .ZN(n20283) );
  OAI211_X1 U22471 ( .C1(n20306), .C2(n20363), .A(n20284), .B(n20283), .ZN(
        P2_U3113) );
  AOI22_X1 U22472 ( .A1(n20372), .A2(n20260), .B1(n20371), .B2(n20307), .ZN(
        n20286) );
  AOI22_X1 U22473 ( .A1(n20309), .A2(n20373), .B1(n20374), .B2(
        P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n20285) );
  OAI211_X1 U22474 ( .C1(n20300), .C2(n20382), .A(n20286), .B(n20285), .ZN(
        P2_U3105) );
  AOI22_X1 U22475 ( .A1(n20378), .A2(n20260), .B1(n20307), .B2(n20377), .ZN(
        n20289) );
  AOI22_X1 U22476 ( .A1(n20309), .A2(n20287), .B1(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n20379), .ZN(n20288) );
  OAI211_X1 U22477 ( .C1(n20300), .C2(n20393), .A(n20289), .B(n20288), .ZN(
        P2_U3097) );
  AOI22_X1 U22478 ( .A1(n20309), .A2(n20290), .B1(n20307), .B2(n20386), .ZN(
        n20292) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20390), .B1(
        n20260), .B2(n20389), .ZN(n20291) );
  OAI211_X1 U22480 ( .C1(n20300), .C2(n20396), .A(n20292), .B(n20291), .ZN(
        P2_U3089) );
  AOI22_X1 U22481 ( .A1(n20309), .A2(n20293), .B1(n20307), .B2(n20394), .ZN(
        n20295) );
  AOI22_X1 U22482 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20399), .B1(
        n20260), .B2(n20398), .ZN(n20294) );
  OAI211_X1 U22483 ( .C1(n20300), .C2(n20404), .A(n20295), .B(n20294), .ZN(
        P2_U3081) );
  AOI22_X1 U22484 ( .A1(n20309), .A2(n20297), .B1(n20296), .B2(n20307), .ZN(
        n20299) );
  AOI22_X1 U22485 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20407), .B1(
        n20260), .B2(n20406), .ZN(n20298) );
  OAI211_X1 U22486 ( .C1(n20300), .C2(n20410), .A(n20299), .B(n20298), .ZN(
        P2_U3073) );
  AOI22_X1 U22487 ( .A1(n20413), .A2(n20260), .B1(n20307), .B2(n20412), .ZN(
        n20302) );
  AOI22_X1 U22488 ( .A1(n20414), .A2(n20308), .B1(n20415), .B2(n20309), .ZN(
        n20301) );
  OAI211_X1 U22489 ( .C1(n20419), .C2(n20303), .A(n20302), .B(n20301), .ZN(
        P2_U3065) );
  AOI22_X1 U22490 ( .A1(n20421), .A2(n20260), .B1(n20307), .B2(n20420), .ZN(
        n20305) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20422), .B1(
        n20432), .B2(n20308), .ZN(n20304) );
  OAI211_X1 U22492 ( .C1(n20306), .C2(n20425), .A(n20305), .B(n20304), .ZN(
        P2_U3057) );
  AOI22_X1 U22493 ( .A1(n20308), .A2(n20430), .B1(n20427), .B2(n20307), .ZN(
        n20311) );
  AOI22_X1 U22494 ( .A1(n20260), .A2(n20433), .B1(n20432), .B2(n20309), .ZN(
        n20310) );
  OAI211_X1 U22495 ( .C1(n20438), .C2(n20312), .A(n20311), .B(n20310), .ZN(
        P2_U3049) );
  AOI22_X1 U22496 ( .A1(n20315), .A2(n20314), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n20313), .ZN(n20324) );
  AOI22_X1 U22497 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20317), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20316), .ZN(n20323) );
  AOI22_X1 U22498 ( .A1(n20321), .A2(n20320), .B1(n20319), .B2(n20318), .ZN(
        n20322) );
  NAND3_X1 U22499 ( .A1(n20324), .A2(n20323), .A3(n20322), .ZN(P2_U2903) );
  AOI22_X1 U22500 ( .A1(n20326), .A2(n20434), .B1(n20428), .B2(n20325), .ZN(
        n20329) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20327), .B1(
        n20430), .B2(n20431), .ZN(n20328) );
  OAI211_X1 U22502 ( .C1(n20411), .C2(n20336), .A(n20329), .B(n20328), .ZN(
        P2_U3168) );
  INV_X1 U22503 ( .A(n20411), .ZN(n20429) );
  AOI22_X1 U22504 ( .A1(n20331), .A2(n20429), .B1(n20428), .B2(n20330), .ZN(
        n20335) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20333), .B1(
        n20434), .B2(n20332), .ZN(n20334) );
  OAI211_X1 U22506 ( .C1(n20426), .C2(n20336), .A(n20335), .B(n20334), .ZN(
        P2_U3160) );
  AOI22_X1 U22507 ( .A1(n20338), .A2(n20434), .B1(n20428), .B2(n20337), .ZN(
        n20342) );
  AOI22_X1 U22508 ( .A1(n20340), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n20339), .B2(n20429), .ZN(n20341) );
  OAI211_X1 U22509 ( .C1(n20426), .C2(n20343), .A(n20342), .B(n20341), .ZN(
        P2_U3152) );
  AOI22_X1 U22510 ( .A1(n20345), .A2(n20434), .B1(n20428), .B2(n20344), .ZN(
        n20348) );
  AOI22_X1 U22511 ( .A1(n20346), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n20351), .B2(n20429), .ZN(n20347) );
  OAI211_X1 U22512 ( .C1(n20426), .C2(n20349), .A(n20348), .B(n20347), .ZN(
        P2_U3136) );
  AOI22_X1 U22513 ( .A1(n20351), .A2(n20431), .B1(n20428), .B2(n20350), .ZN(
        n20355) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20353), .B1(
        n20434), .B2(n20352), .ZN(n20354) );
  OAI211_X1 U22515 ( .C1(n20411), .C2(n20356), .A(n20355), .B(n20354), .ZN(
        P2_U3128) );
  AOI22_X1 U22516 ( .A1(n20358), .A2(n20431), .B1(n20428), .B2(n20357), .ZN(
        n20362) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20360), .B1(
        n20434), .B2(n20359), .ZN(n20361) );
  OAI211_X1 U22518 ( .C1(n20411), .C2(n20363), .A(n20362), .B(n20361), .ZN(
        P2_U3120) );
  AOI22_X1 U22519 ( .A1(n20365), .A2(n20431), .B1(n20428), .B2(n20364), .ZN(
        n20369) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20367), .B1(
        n20434), .B2(n20366), .ZN(n20368) );
  OAI211_X1 U22521 ( .C1(n20411), .C2(n20370), .A(n20369), .B(n20368), .ZN(
        P2_U3112) );
  AOI22_X1 U22522 ( .A1(n20372), .A2(n20434), .B1(n20371), .B2(n20428), .ZN(
        n20376) );
  AOI22_X1 U22523 ( .A1(n20374), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n20373), .B2(n20431), .ZN(n20375) );
  OAI211_X1 U22524 ( .C1(n20411), .C2(n20382), .A(n20376), .B(n20375), .ZN(
        P2_U3104) );
  AOI22_X1 U22525 ( .A1(n20378), .A2(n20434), .B1(n20428), .B2(n20377), .ZN(
        n20385) );
  INV_X1 U22526 ( .A(n20379), .ZN(n20381) );
  INV_X1 U22527 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n20380) );
  OAI22_X1 U22528 ( .A1(n20382), .A2(n20426), .B1(n20381), .B2(n20380), .ZN(
        n20383) );
  INV_X1 U22529 ( .A(n20383), .ZN(n20384) );
  OAI211_X1 U22530 ( .C1(n20411), .C2(n20393), .A(n20385), .B(n20384), .ZN(
        P2_U3096) );
  INV_X1 U22531 ( .A(n20386), .ZN(n20387) );
  OAI22_X1 U22532 ( .A1(n20396), .A2(n20411), .B1(n20403), .B2(n20387), .ZN(
        n20388) );
  INV_X1 U22533 ( .A(n20388), .ZN(n20392) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20390), .B1(
        n20434), .B2(n20389), .ZN(n20391) );
  OAI211_X1 U22535 ( .C1(n20426), .C2(n20393), .A(n20392), .B(n20391), .ZN(
        P2_U3088) );
  INV_X1 U22536 ( .A(n20394), .ZN(n20395) );
  OAI22_X1 U22537 ( .A1(n20396), .A2(n20426), .B1(n20403), .B2(n20395), .ZN(
        n20397) );
  INV_X1 U22538 ( .A(n20397), .ZN(n20401) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20399), .B1(
        n20434), .B2(n20398), .ZN(n20400) );
  OAI211_X1 U22540 ( .C1(n20411), .C2(n20404), .A(n20401), .B(n20400), .ZN(
        P2_U3080) );
  OAI22_X1 U22541 ( .A1(n20404), .A2(n20426), .B1(n20403), .B2(n20402), .ZN(
        n20405) );
  INV_X1 U22542 ( .A(n20405), .ZN(n20409) );
  AOI22_X1 U22543 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20407), .B1(
        n20434), .B2(n20406), .ZN(n20408) );
  OAI211_X1 U22544 ( .C1(n20411), .C2(n20410), .A(n20409), .B(n20408), .ZN(
        P2_U3072) );
  INV_X1 U22545 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n20418) );
  AOI22_X1 U22546 ( .A1(n20413), .A2(n20434), .B1(n20428), .B2(n20412), .ZN(
        n20417) );
  AOI22_X1 U22547 ( .A1(n20415), .A2(n20431), .B1(n20414), .B2(n20429), .ZN(
        n20416) );
  OAI211_X1 U22548 ( .C1(n20419), .C2(n20418), .A(n20417), .B(n20416), .ZN(
        P2_U3064) );
  AOI22_X1 U22549 ( .A1(n20421), .A2(n20434), .B1(n20428), .B2(n20420), .ZN(
        n20424) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20422), .B1(
        n20432), .B2(n20429), .ZN(n20423) );
  OAI211_X1 U22551 ( .C1(n20426), .C2(n20425), .A(n20424), .B(n20423), .ZN(
        P2_U3056) );
  AOI22_X1 U22552 ( .A1(n20430), .A2(n20429), .B1(n20428), .B2(n20427), .ZN(
        n20436) );
  AOI22_X1 U22553 ( .A1(n20434), .A2(n20433), .B1(n20432), .B2(n20431), .ZN(
        n20435) );
  OAI211_X1 U22554 ( .C1(n20438), .C2(n20437), .A(n20436), .B(n20435), .ZN(
        P2_U3048) );
  INV_X1 U22555 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20775) );
  INV_X1 U22556 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20439) );
  AOI222_X1 U22557 ( .A1(n20775), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20778), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n20439), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n20440) );
  INV_X2 U22558 ( .A(n20440), .ZN(n20500) );
  INV_X1 U22559 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20442) );
  AOI22_X1 U22560 ( .A1(n20489), .A2(n20442), .B1(n20441), .B2(n20500), .ZN(
        U376) );
  INV_X1 U22561 ( .A(n20500), .ZN(n20503) );
  INV_X1 U22562 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n20444) );
  AOI22_X1 U22563 ( .A1(n20503), .A2(n20444), .B1(n20443), .B2(n20500), .ZN(
        U365) );
  INV_X1 U22564 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n20446) );
  AOI22_X1 U22565 ( .A1(n20489), .A2(n20446), .B1(n20445), .B2(n20500), .ZN(
        U354) );
  INV_X1 U22566 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n20448) );
  AOI22_X1 U22567 ( .A1(n20489), .A2(n20448), .B1(n20447), .B2(n20500), .ZN(
        U353) );
  INV_X1 U22568 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n20450) );
  AOI22_X1 U22569 ( .A1(n20489), .A2(n20450), .B1(n20449), .B2(n20500), .ZN(
        U352) );
  INV_X1 U22570 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n20452) );
  AOI22_X1 U22571 ( .A1(n20489), .A2(n20452), .B1(n20451), .B2(n20500), .ZN(
        U351) );
  INV_X1 U22572 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n20454) );
  AOI22_X1 U22573 ( .A1(n20503), .A2(n20454), .B1(n20453), .B2(n20500), .ZN(
        U350) );
  INV_X1 U22574 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n20456) );
  AOI22_X1 U22575 ( .A1(n20489), .A2(n20456), .B1(n20455), .B2(n20500), .ZN(
        U349) );
  INV_X1 U22576 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20458) );
  AOI22_X1 U22577 ( .A1(n20489), .A2(n20458), .B1(n20457), .B2(n20500), .ZN(
        U348) );
  INV_X1 U22578 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n20460) );
  AOI22_X1 U22579 ( .A1(n20489), .A2(n20460), .B1(n20459), .B2(n20500), .ZN(
        U347) );
  INV_X1 U22580 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20462) );
  AOI22_X1 U22581 ( .A1(n20489), .A2(n20462), .B1(n20461), .B2(n20500), .ZN(
        U375) );
  INV_X1 U22582 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20464) );
  AOI22_X1 U22583 ( .A1(n20489), .A2(n20464), .B1(n20463), .B2(n20500), .ZN(
        U374) );
  INV_X1 U22584 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20466) );
  AOI22_X1 U22585 ( .A1(n20489), .A2(n20466), .B1(n20465), .B2(n20500), .ZN(
        U373) );
  INV_X1 U22586 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20468) );
  AOI22_X1 U22587 ( .A1(n20489), .A2(n20468), .B1(n20467), .B2(n20500), .ZN(
        U372) );
  INV_X1 U22588 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20470) );
  AOI22_X1 U22589 ( .A1(n20489), .A2(n20470), .B1(n20469), .B2(n20500), .ZN(
        U371) );
  INV_X1 U22590 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20472) );
  AOI22_X1 U22591 ( .A1(n20489), .A2(n20472), .B1(n20471), .B2(n20500), .ZN(
        U370) );
  INV_X1 U22592 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20474) );
  AOI22_X1 U22593 ( .A1(n20489), .A2(n20474), .B1(n20473), .B2(n20500), .ZN(
        U369) );
  INV_X1 U22594 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20476) );
  AOI22_X1 U22595 ( .A1(n20489), .A2(n20476), .B1(n20475), .B2(n20500), .ZN(
        U368) );
  INV_X1 U22596 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20478) );
  AOI22_X1 U22597 ( .A1(n20489), .A2(n20478), .B1(n20477), .B2(n20500), .ZN(
        U367) );
  INV_X1 U22598 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20480) );
  AOI22_X1 U22599 ( .A1(n20489), .A2(n20480), .B1(n20479), .B2(n20500), .ZN(
        U366) );
  INV_X1 U22600 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20482) );
  AOI22_X1 U22601 ( .A1(n20489), .A2(n20482), .B1(n20481), .B2(n20500), .ZN(
        U364) );
  INV_X1 U22602 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n20484) );
  AOI22_X1 U22603 ( .A1(n20489), .A2(n20484), .B1(n20483), .B2(n20500), .ZN(
        U363) );
  INV_X1 U22604 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20486) );
  AOI22_X1 U22605 ( .A1(n20489), .A2(n20486), .B1(n20485), .B2(n20500), .ZN(
        U362) );
  INV_X1 U22606 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20488) );
  AOI22_X1 U22607 ( .A1(n20489), .A2(n20488), .B1(n20487), .B2(n20500), .ZN(
        U361) );
  INV_X1 U22608 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20491) );
  AOI22_X1 U22609 ( .A1(n20503), .A2(n20491), .B1(n20490), .B2(n20500), .ZN(
        U360) );
  INV_X1 U22610 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20493) );
  AOI22_X1 U22611 ( .A1(n20503), .A2(n20493), .B1(n20492), .B2(n20500), .ZN(
        U359) );
  INV_X1 U22612 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20495) );
  AOI22_X1 U22613 ( .A1(n20503), .A2(n20495), .B1(n20494), .B2(n20500), .ZN(
        U358) );
  INV_X1 U22614 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20497) );
  AOI22_X1 U22615 ( .A1(n20503), .A2(n20497), .B1(n20496), .B2(n20500), .ZN(
        U357) );
  INV_X1 U22616 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20499) );
  AOI22_X1 U22617 ( .A1(n20503), .A2(n20499), .B1(n20498), .B2(n20500), .ZN(
        U356) );
  INV_X1 U22618 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20502) );
  AOI22_X1 U22619 ( .A1(n20503), .A2(n20502), .B1(n20501), .B2(n20500), .ZN(
        U355) );
  AOI22_X1 U22620 ( .A1(n21955), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20505) );
  OAI21_X1 U22621 ( .B1(n20506), .B2(n20526), .A(n20505), .ZN(P1_U2936) );
  AOI22_X1 U22622 ( .A1(n21955), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20507) );
  OAI21_X1 U22623 ( .B1(n13076), .B2(n20526), .A(n20507), .ZN(P1_U2935) );
  AOI22_X1 U22624 ( .A1(n21955), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20508) );
  OAI21_X1 U22625 ( .B1(n13067), .B2(n20526), .A(n20508), .ZN(P1_U2934) );
  AOI22_X1 U22626 ( .A1(n20521), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20509) );
  OAI21_X1 U22627 ( .B1(n13098), .B2(n20526), .A(n20509), .ZN(P1_U2933) );
  AOI22_X1 U22628 ( .A1(n20521), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20510) );
  OAI21_X1 U22629 ( .B1(n20511), .B2(n20526), .A(n20510), .ZN(P1_U2932) );
  AOI22_X1 U22630 ( .A1(n20521), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20512) );
  OAI21_X1 U22631 ( .B1(n20513), .B2(n20526), .A(n20512), .ZN(P1_U2931) );
  AOI22_X1 U22632 ( .A1(n20521), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20515) );
  OAI21_X1 U22633 ( .B1(n13127), .B2(n20526), .A(n20515), .ZN(P1_U2930) );
  AOI22_X1 U22634 ( .A1(n20521), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20516) );
  OAI21_X1 U22635 ( .B1(n13140), .B2(n20526), .A(n20516), .ZN(P1_U2929) );
  AOI22_X1 U22636 ( .A1(n20521), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20517) );
  OAI21_X1 U22637 ( .B1(n16199), .B2(n20526), .A(n20517), .ZN(P1_U2928) );
  INV_X1 U22638 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n22352) );
  AOI22_X1 U22639 ( .A1(n20521), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20518) );
  OAI21_X1 U22640 ( .B1(n22352), .B2(n20526), .A(n20518), .ZN(P1_U2927) );
  AOI22_X1 U22641 ( .A1(n20521), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20519) );
  OAI21_X1 U22642 ( .B1(n16271), .B2(n20526), .A(n20519), .ZN(P1_U2926) );
  AOI22_X1 U22643 ( .A1(n20521), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20520) );
  OAI21_X1 U22644 ( .B1(n16279), .B2(n20526), .A(n20520), .ZN(P1_U2925) );
  INV_X1 U22645 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n22366) );
  AOI22_X1 U22646 ( .A1(n20521), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20522) );
  OAI21_X1 U22647 ( .B1(n22366), .B2(n20526), .A(n20522), .ZN(P1_U2924) );
  AOI22_X1 U22648 ( .A1(n21955), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20523) );
  OAI21_X1 U22649 ( .B1(n16790), .B2(n20526), .A(n20523), .ZN(P1_U2923) );
  AOI22_X1 U22650 ( .A1(n21955), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20524) );
  OAI21_X1 U22651 ( .B1(n16786), .B2(n20526), .A(n20524), .ZN(P1_U2922) );
  AOI22_X1 U22652 ( .A1(n21955), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20514), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20525) );
  OAI21_X1 U22653 ( .B1(n20527), .B2(n20526), .A(n20525), .ZN(P1_U2921) );
  INV_X1 U22654 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n22295) );
  AND2_X1 U22655 ( .A1(n20780), .A2(n22295), .ZN(n20544) );
  AND2_X1 U22656 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20780), .ZN(n20546) );
  INV_X2 U22657 ( .A(n20546), .ZN(n20577) );
  OAI222_X1 U22658 ( .A1(n11157), .A2(n20529), .B1(n20528), .B2(n20780), .C1(
        n20592), .C2(n20577), .ZN(P1_U3197) );
  INV_X1 U22659 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20530) );
  OAI222_X1 U22660 ( .A1(n11157), .A2(n15820), .B1(n20530), .B2(n20780), .C1(
        n20529), .C2(n20577), .ZN(P1_U3198) );
  INV_X1 U22661 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20531) );
  OAI222_X1 U22662 ( .A1(n11157), .A2(n20532), .B1(n20531), .B2(n20780), .C1(
        n15820), .C2(n20577), .ZN(P1_U3199) );
  INV_X1 U22663 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20533) );
  OAI222_X1 U22664 ( .A1(n11157), .A2(n20535), .B1(n20533), .B2(n20780), .C1(
        n20532), .C2(n20577), .ZN(P1_U3200) );
  INV_X1 U22665 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20534) );
  OAI222_X1 U22666 ( .A1(n20577), .A2(n20535), .B1(n20534), .B2(n20780), .C1(
        n20536), .C2(n11157), .ZN(P1_U3201) );
  INV_X1 U22667 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20537) );
  OAI222_X1 U22668 ( .A1(n11157), .A2(n22158), .B1(n20537), .B2(n20780), .C1(
        n20536), .C2(n20577), .ZN(P1_U3202) );
  INV_X1 U22669 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20538) );
  OAI222_X1 U22670 ( .A1(n20577), .A2(n22158), .B1(n20538), .B2(n20780), .C1(
        n22164), .C2(n11157), .ZN(P1_U3203) );
  INV_X1 U22671 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20539) );
  OAI222_X1 U22672 ( .A1(n20577), .A2(n22164), .B1(n20539), .B2(n20780), .C1(
        n22183), .C2(n11157), .ZN(P1_U3204) );
  INV_X1 U22673 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20540) );
  OAI222_X1 U22674 ( .A1(n20577), .A2(n22183), .B1(n20540), .B2(n20780), .C1(
        n14777), .C2(n11157), .ZN(P1_U3205) );
  INV_X1 U22675 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20541) );
  OAI222_X1 U22676 ( .A1(n20577), .A2(n14777), .B1(n20541), .B2(n20780), .C1(
        n20653), .C2(n11157), .ZN(P1_U3206) );
  INV_X1 U22677 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n22220) );
  INV_X1 U22678 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20542) );
  OAI222_X1 U22679 ( .A1(n11157), .A2(n22220), .B1(n20542), .B2(n20780), .C1(
        n20653), .C2(n20577), .ZN(P1_U3207) );
  INV_X1 U22680 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20543) );
  OAI222_X1 U22681 ( .A1(n11157), .A2(n21966), .B1(n20543), .B2(n20780), .C1(
        n22220), .C2(n20577), .ZN(P1_U3208) );
  AOI22_X1 U22682 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n20544), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n22778), .ZN(n20545) );
  OAI21_X1 U22683 ( .B1(n21966), .B2(n20577), .A(n20545), .ZN(P1_U3209) );
  AOI22_X1 U22684 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n20546), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n22778), .ZN(n20547) );
  OAI21_X1 U22685 ( .B1(n20549), .B2(n11157), .A(n20547), .ZN(P1_U3210) );
  INV_X1 U22686 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20548) );
  OAI222_X1 U22687 ( .A1(n20577), .A2(n20549), .B1(n20548), .B2(n20780), .C1(
        n22227), .C2(n11157), .ZN(P1_U3211) );
  INV_X1 U22688 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20550) );
  OAI222_X1 U22689 ( .A1(n20577), .A2(n22227), .B1(n20550), .B2(n20780), .C1(
        n20551), .C2(n11157), .ZN(P1_U3212) );
  INV_X1 U22690 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20552) );
  OAI222_X1 U22691 ( .A1(n11157), .A2(n20554), .B1(n20552), .B2(n20780), .C1(
        n20551), .C2(n20577), .ZN(P1_U3213) );
  INV_X1 U22692 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20553) );
  OAI222_X1 U22693 ( .A1(n20577), .A2(n20554), .B1(n20553), .B2(n20780), .C1(
        n22067), .C2(n11157), .ZN(P1_U3214) );
  INV_X1 U22694 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20555) );
  OAI222_X1 U22695 ( .A1(n11157), .A2(n20557), .B1(n20555), .B2(n20780), .C1(
        n22067), .C2(n20577), .ZN(P1_U3215) );
  INV_X1 U22696 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20556) );
  OAI222_X1 U22697 ( .A1(n20577), .A2(n20557), .B1(n20556), .B2(n20780), .C1(
        n20559), .C2(n11157), .ZN(P1_U3216) );
  INV_X1 U22698 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20558) );
  OAI222_X1 U22699 ( .A1(n20577), .A2(n20559), .B1(n20558), .B2(n20780), .C1(
        n20561), .C2(n11157), .ZN(P1_U3217) );
  INV_X1 U22700 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20560) );
  OAI222_X1 U22701 ( .A1(n20577), .A2(n20561), .B1(n20560), .B2(n20780), .C1(
        n20563), .C2(n11157), .ZN(P1_U3218) );
  INV_X1 U22702 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20562) );
  OAI222_X1 U22703 ( .A1(n20577), .A2(n20563), .B1(n20562), .B2(n20780), .C1(
        n20565), .C2(n11157), .ZN(P1_U3219) );
  INV_X1 U22704 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20564) );
  INV_X1 U22705 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n22092) );
  OAI222_X1 U22706 ( .A1(n20577), .A2(n20565), .B1(n20564), .B2(n20780), .C1(
        n22092), .C2(n11157), .ZN(P1_U3220) );
  INV_X1 U22707 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20566) );
  OAI222_X1 U22708 ( .A1(n11157), .A2(n20568), .B1(n20566), .B2(n20780), .C1(
        n22092), .C2(n20577), .ZN(P1_U3221) );
  INV_X1 U22709 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20567) );
  OAI222_X1 U22710 ( .A1(n20577), .A2(n20568), .B1(n20567), .B2(n20780), .C1(
        n22085), .C2(n11157), .ZN(P1_U3222) );
  INV_X1 U22711 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20569) );
  OAI222_X1 U22712 ( .A1(n20577), .A2(n22085), .B1(n20569), .B2(n20780), .C1(
        n20570), .C2(n11157), .ZN(P1_U3223) );
  INV_X1 U22713 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20571) );
  OAI222_X1 U22714 ( .A1(n11157), .A2(n20573), .B1(n20571), .B2(n20780), .C1(
        n20570), .C2(n20577), .ZN(P1_U3224) );
  INV_X1 U22715 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20572) );
  OAI222_X1 U22716 ( .A1(n20577), .A2(n20573), .B1(n20572), .B2(n20780), .C1(
        n20576), .C2(n11157), .ZN(P1_U3225) );
  INV_X1 U22717 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20575) );
  OAI222_X1 U22718 ( .A1(n20577), .A2(n20576), .B1(n20575), .B2(n20780), .C1(
        n20574), .C2(n11157), .ZN(P1_U3226) );
  INV_X1 U22719 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20578) );
  AOI22_X1 U22720 ( .A1(n20780), .A2(n20579), .B1(n20578), .B2(n22778), .ZN(
        P1_U3458) );
  AOI221_X1 U22721 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20590) );
  NOR4_X1 U22722 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20583) );
  NOR4_X1 U22723 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20582) );
  NOR4_X1 U22724 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20581) );
  NOR4_X1 U22725 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20580) );
  NAND4_X1 U22726 ( .A1(n20583), .A2(n20582), .A3(n20581), .A4(n20580), .ZN(
        n20589) );
  NOR4_X1 U22727 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20587) );
  AOI211_X1 U22728 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20586) );
  NOR4_X1 U22729 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20585) );
  NOR4_X1 U22730 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20584) );
  NAND4_X1 U22731 ( .A1(n20587), .A2(n20586), .A3(n20585), .A4(n20584), .ZN(
        n20588) );
  NOR2_X1 U22732 ( .A1(n20589), .A2(n20588), .ZN(n20603) );
  MUX2_X1 U22733 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(n20590), .S(n20603), 
        .Z(P1_U2808) );
  INV_X1 U22734 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20595) );
  INV_X1 U22735 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20591) );
  AOI22_X1 U22736 ( .A1(n20780), .A2(n20595), .B1(n20591), .B2(n22778), .ZN(
        P1_U3459) );
  AOI21_X1 U22737 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20593) );
  OAI221_X1 U22738 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20593), .C1(n20592), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20603), .ZN(n20594) );
  OAI21_X1 U22739 ( .B1(n20603), .B2(n20595), .A(n20594), .ZN(P1_U3481) );
  INV_X1 U22740 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20596) );
  AOI22_X1 U22741 ( .A1(n20780), .A2(n20599), .B1(n20596), .B2(n22778), .ZN(
        P1_U3460) );
  NOR3_X1 U22742 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20597) );
  OAI21_X1 U22743 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20597), .A(n20603), .ZN(
        n20598) );
  OAI21_X1 U22744 ( .B1(n20603), .B2(n20599), .A(n20598), .ZN(P1_U2807) );
  INV_X1 U22745 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20600) );
  AOI22_X1 U22746 ( .A1(n20780), .A2(n20602), .B1(n20600), .B2(n22778), .ZN(
        P1_U3461) );
  OAI21_X1 U22747 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .A(n20603), .ZN(n20601) );
  OAI21_X1 U22748 ( .B1(n20603), .B2(n20602), .A(n20601), .ZN(P1_U3482) );
  INV_X1 U22749 ( .A(n20604), .ZN(n20605) );
  AOI22_X1 U22750 ( .A1(n20605), .A2(n20618), .B1(n20617), .B2(n21995), .ZN(
        n20606) );
  OAI21_X1 U22751 ( .B1(n20621), .B2(n20607), .A(n20606), .ZN(P1_U2869) );
  XNOR2_X1 U22752 ( .A(n20609), .B(n20608), .ZN(n22189) );
  AOI22_X1 U22753 ( .A1(n22192), .A2(n20618), .B1(n20617), .B2(n22189), .ZN(
        n20610) );
  OAI21_X1 U22754 ( .B1(n20621), .B2(n20611), .A(n20610), .ZN(P1_U2862) );
  NOR2_X1 U22755 ( .A1(n20612), .A2(n16724), .ZN(n20613) );
  AOI21_X1 U22756 ( .B1(n20614), .B2(n20618), .A(n20613), .ZN(n20615) );
  OAI21_X1 U22757 ( .B1(n20621), .B2(n20616), .A(n20615), .ZN(P1_U2857) );
  AOI22_X1 U22758 ( .A1(n20677), .A2(n20618), .B1(n20617), .B2(n21976), .ZN(
        n20619) );
  OAI21_X1 U22759 ( .B1(n20621), .B2(n20620), .A(n20619), .ZN(P1_U2858) );
  INV_X1 U22760 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20626) );
  INV_X1 U22761 ( .A(n22173), .ZN(n20622) );
  OAI22_X1 U22762 ( .A1(n22179), .A2(n20623), .B1(n16724), .B2(n20622), .ZN(
        n20624) );
  INV_X1 U22763 ( .A(n20624), .ZN(n20625) );
  OAI21_X1 U22764 ( .B1(n20621), .B2(n20626), .A(n20625), .ZN(P1_U2863) );
  INV_X1 U22765 ( .A(n20627), .ZN(n20630) );
  INV_X1 U22766 ( .A(n20628), .ZN(n20629) );
  AOI21_X1 U22767 ( .B1(n20630), .B2(n22123), .A(n20629), .ZN(n22119) );
  OR2_X1 U22768 ( .A1(n20694), .A2(n20631), .ZN(n20632) );
  AOI22_X1 U22769 ( .A1(n22119), .A2(n13804), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20632), .ZN(n20633) );
  NAND2_X1 U22770 ( .A1(n22102), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n22113) );
  OAI211_X1 U22771 ( .C1(n20634), .C2(n20697), .A(n20633), .B(n22113), .ZN(
        P1_U2999) );
  AOI222_X1 U22772 ( .A1(n20637), .A2(n13804), .B1(n20636), .B2(n20689), .C1(
        n20635), .C2(n20676), .ZN(n20639) );
  OAI211_X1 U22773 ( .C1(n20646), .C2(n20640), .A(n20639), .B(n20638), .ZN(
        P1_U2994) );
  INV_X1 U22774 ( .A(n22148), .ZN(n20641) );
  AOI222_X1 U22775 ( .A1(n20642), .A2(n13804), .B1(n20689), .B2(n22155), .C1(
        n20641), .C2(n20676), .ZN(n20644) );
  OAI211_X1 U22776 ( .C1(n20646), .C2(n20645), .A(n20644), .B(n20643), .ZN(
        P1_U2992) );
  MUX2_X1 U22777 ( .A(n20647), .B(n20669), .S(n11670), .Z(n20648) );
  INV_X1 U22778 ( .A(n20648), .ZN(n20649) );
  OAI21_X1 U22779 ( .B1(n20649), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n20656), .ZN(n22015) );
  AOI22_X1 U22780 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20694), .B1(
        n22102), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n20652) );
  INV_X1 U22781 ( .A(n20650), .ZN(n22191) );
  AOI22_X1 U22782 ( .A1(n22192), .A2(n20689), .B1(n22191), .B2(n20676), .ZN(
        n20651) );
  OAI211_X1 U22783 ( .C1(n20696), .C2(n22015), .A(n20652), .B(n20651), .ZN(
        P1_U2989) );
  NOR2_X1 U22784 ( .A1(n22093), .A2(n20653), .ZN(n22031) );
  NAND2_X1 U22785 ( .A1(n20656), .A2(n20654), .ZN(n20655) );
  MUX2_X1 U22786 ( .A(n20656), .B(n20655), .S(n11670), .Z(n20658) );
  INV_X1 U22787 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20657) );
  OAI22_X1 U22788 ( .A1(n22029), .A2(n20696), .B1(n20703), .B2(n22209), .ZN(
        n20659) );
  OAI21_X1 U22789 ( .B1(n20697), .B2(n20661), .A(n20660), .ZN(P1_U2988) );
  AOI21_X1 U22790 ( .B1(n20664), .B2(n20663), .A(n20662), .ZN(n22028) );
  AOI22_X1 U22791 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20694), .B1(
        n22102), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n20667) );
  INV_X1 U22792 ( .A(n20665), .ZN(n22214) );
  AOI22_X1 U22793 ( .A1(n20676), .A2(n22217), .B1(n20689), .B2(n22214), .ZN(
        n20666) );
  OAI211_X1 U22794 ( .C1(n22028), .C2(n20696), .A(n20667), .B(n20666), .ZN(
        P1_U2987) );
  NOR2_X1 U22795 ( .A1(n20669), .A2(n20668), .ZN(n20672) );
  OAI21_X1 U22796 ( .B1(n20672), .B2(n20671), .A(n20670), .ZN(n20674) );
  XNOR2_X1 U22797 ( .A(n11667), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n20673) );
  XNOR2_X1 U22798 ( .A(n20674), .B(n20673), .ZN(n21979) );
  AOI22_X1 U22799 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20694), .B1(
        n22102), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n20679) );
  AOI22_X1 U22800 ( .A1(n20677), .A2(n20689), .B1(n20676), .B2(n20675), .ZN(
        n20678) );
  OAI211_X1 U22801 ( .C1(n21979), .C2(n20696), .A(n20679), .B(n20678), .ZN(
        P1_U2985) );
  AOI22_X1 U22802 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n20694), .B1(
        n22102), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n20687) );
  OAI21_X1 U22803 ( .B1(n11670), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n20680), .ZN(n20684) );
  OAI21_X1 U22804 ( .B1(n11670), .B2(n20682), .A(n20681), .ZN(n20683) );
  XNOR2_X1 U22805 ( .A(n20684), .B(n20683), .ZN(n22059) );
  AOI22_X1 U22806 ( .A1(n20685), .A2(n20689), .B1(n13804), .B2(n22059), .ZN(
        n20686) );
  OAI211_X1 U22807 ( .C1(n20703), .C2(n22245), .A(n20687), .B(n20686), .ZN(
        P1_U2983) );
  AOI22_X1 U22808 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20694), .B1(
        n22102), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n20692) );
  AOI22_X1 U22809 ( .A1(n20690), .A2(n20689), .B1(n13804), .B2(n20688), .ZN(
        n20691) );
  OAI211_X1 U22810 ( .C1(n20703), .C2(n20693), .A(n20692), .B(n20691), .ZN(
        P1_U2979) );
  AOI22_X1 U22811 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20694), .B1(
        n22102), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n20701) );
  OAI22_X1 U22812 ( .A1(n20698), .A2(n20697), .B1(n20696), .B2(n20695), .ZN(
        n20699) );
  INV_X1 U22813 ( .A(n20699), .ZN(n20700) );
  OAI211_X1 U22814 ( .C1(n20703), .C2(n20702), .A(n20701), .B(n20700), .ZN(
        P1_U2977) );
  AND2_X1 U22815 ( .A1(n20705), .A2(n20704), .ZN(n20708) );
  OAI22_X1 U22816 ( .A1(n20708), .A2(n20707), .B1(n22256), .B2(n20706), .ZN(
        P1_U2803) );
  OAI21_X1 U22817 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n22295), .A(n22302), 
        .ZN(n20709) );
  AOI22_X1 U22818 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n20780), .B1(n20710), 
        .B2(n20709), .ZN(P1_U2804) );
  INV_X1 U22819 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20713) );
  AOI22_X1 U22820 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n11155), .ZN(n20712) );
  OAI21_X1 U22821 ( .B1(n20713), .B2(n20777), .A(n20712), .ZN(U247) );
  AOI22_X1 U22822 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n11155), .ZN(n20714) );
  OAI21_X1 U22823 ( .B1(n20715), .B2(n20777), .A(n20714), .ZN(U246) );
  INV_X1 U22824 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20717) );
  AOI22_X1 U22825 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n11155), .ZN(n20716) );
  OAI21_X1 U22826 ( .B1(n20717), .B2(n20777), .A(n20716), .ZN(U245) );
  AOI22_X1 U22827 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n11155), .ZN(n20718) );
  OAI21_X1 U22828 ( .B1(n20719), .B2(n20777), .A(n20718), .ZN(U244) );
  AOI22_X1 U22829 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n11155), .ZN(n20720) );
  OAI21_X1 U22830 ( .B1(n20721), .B2(n20777), .A(n20720), .ZN(U243) );
  INV_X1 U22831 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20723) );
  AOI22_X1 U22832 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n11155), .ZN(n20722) );
  OAI21_X1 U22833 ( .B1(n20723), .B2(n20777), .A(n20722), .ZN(U242) );
  INV_X1 U22834 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20725) );
  AOI22_X1 U22835 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n11155), .ZN(n20724) );
  OAI21_X1 U22836 ( .B1(n20725), .B2(n20777), .A(n20724), .ZN(U241) );
  AOI22_X1 U22837 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n11155), .ZN(n20726) );
  OAI21_X1 U22838 ( .B1(n20727), .B2(n20777), .A(n20726), .ZN(U240) );
  AOI22_X1 U22839 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n11155), .ZN(n20728) );
  OAI21_X1 U22840 ( .B1(n20729), .B2(n20777), .A(n20728), .ZN(U239) );
  AOI22_X1 U22841 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n11155), .ZN(n20730) );
  OAI21_X1 U22842 ( .B1(n20731), .B2(n20777), .A(n20730), .ZN(U238) );
  INV_X1 U22843 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20733) );
  AOI22_X1 U22844 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n11155), .ZN(n20732) );
  OAI21_X1 U22845 ( .B1(n20733), .B2(n20777), .A(n20732), .ZN(U237) );
  AOI22_X1 U22846 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n11155), .ZN(n20734) );
  OAI21_X1 U22847 ( .B1(n20735), .B2(n20777), .A(n20734), .ZN(U236) );
  AOI22_X1 U22848 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n11155), .ZN(n20736) );
  OAI21_X1 U22849 ( .B1(n20737), .B2(n20777), .A(n20736), .ZN(U235) );
  AOI22_X1 U22850 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n11155), .ZN(n20738) );
  OAI21_X1 U22851 ( .B1(n20739), .B2(n20777), .A(n20738), .ZN(U234) );
  INV_X1 U22852 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20741) );
  AOI22_X1 U22853 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n11155), .ZN(n20740) );
  OAI21_X1 U22854 ( .B1(n20741), .B2(n20777), .A(n20740), .ZN(U233) );
  INV_X1 U22855 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n20743) );
  AOI22_X1 U22856 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n11155), .ZN(n20742) );
  OAI21_X1 U22857 ( .B1(n20743), .B2(n20777), .A(n20742), .ZN(U232) );
  AOI22_X1 U22858 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n11155), .ZN(n20744) );
  OAI21_X1 U22859 ( .B1(n20745), .B2(n20777), .A(n20744), .ZN(U231) );
  AOI22_X1 U22860 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n11155), .ZN(n20746) );
  OAI21_X1 U22861 ( .B1(n20747), .B2(n20777), .A(n20746), .ZN(U230) );
  AOI22_X1 U22862 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n11155), .ZN(n20748) );
  OAI21_X1 U22863 ( .B1(n20749), .B2(n20777), .A(n20748), .ZN(U229) );
  AOI22_X1 U22864 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n11155), .ZN(n20750) );
  OAI21_X1 U22865 ( .B1(n20751), .B2(n20777), .A(n20750), .ZN(U228) );
  AOI22_X1 U22866 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n11155), .ZN(n20752) );
  OAI21_X1 U22867 ( .B1(n20753), .B2(n20777), .A(n20752), .ZN(U227) );
  AOI22_X1 U22868 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n11155), .ZN(n20754) );
  OAI21_X1 U22869 ( .B1(n20755), .B2(n20777), .A(n20754), .ZN(U226) );
  AOI22_X1 U22870 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n11155), .ZN(n20756) );
  OAI21_X1 U22871 ( .B1(n20757), .B2(n20777), .A(n20756), .ZN(U225) );
  AOI22_X1 U22872 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n11155), .ZN(n20758) );
  OAI21_X1 U22873 ( .B1(n20759), .B2(n20777), .A(n20758), .ZN(U224) );
  AOI22_X1 U22874 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n11155), .ZN(n20760) );
  OAI21_X1 U22875 ( .B1(n20761), .B2(n20777), .A(n20760), .ZN(U223) );
  AOI22_X1 U22876 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n11155), .ZN(n20762) );
  OAI21_X1 U22877 ( .B1(n20763), .B2(n20777), .A(n20762), .ZN(U222) );
  AOI22_X1 U22878 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n11155), .ZN(n20765) );
  OAI21_X1 U22879 ( .B1(n20766), .B2(n20777), .A(n20765), .ZN(U221) );
  AOI22_X1 U22880 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n11155), .ZN(n20767) );
  OAI21_X1 U22881 ( .B1(n20768), .B2(n20777), .A(n20767), .ZN(U220) );
  AOI22_X1 U22882 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n11155), .ZN(n20769) );
  OAI21_X1 U22883 ( .B1(n20770), .B2(n20777), .A(n20769), .ZN(U219) );
  AOI22_X1 U22884 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n11155), .ZN(n20771) );
  OAI21_X1 U22885 ( .B1(n20772), .B2(n20777), .A(n20771), .ZN(U218) );
  AOI22_X1 U22886 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20764), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n11155), .ZN(n20773) );
  OAI21_X1 U22887 ( .B1(n20774), .B2(n20777), .A(n20773), .ZN(U217) );
  OAI222_X1 U22888 ( .A1(U212), .A2(n20778), .B1(n20777), .B2(n20776), .C1(
        U214), .C2(n20775), .ZN(U216) );
  AOI22_X1 U22889 ( .A1(n20780), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20779), 
        .B2(n22778), .ZN(P1_U3483) );
  OAI21_X1 U22890 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20850), .A(n20851), 
        .ZN(n20781) );
  AOI211_X1 U22891 ( .C1(n20782), .C2(n20781), .A(n22285), .B(n21808), .ZN(
        n20784) );
  INV_X1 U22892 ( .A(n21939), .ZN(n20783) );
  OAI21_X1 U22893 ( .B1(n20784), .B2(n20846), .A(n20783), .ZN(n20788) );
  OAI21_X1 U22894 ( .B1(n22285), .B2(n21891), .A(n20848), .ZN(n20785) );
  AOI21_X1 U22895 ( .B1(n20786), .B2(n21948), .A(n20785), .ZN(n20787) );
  MUX2_X1 U22896 ( .A(n20788), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n20787), 
        .Z(P3_U3296) );
  NAND3_X1 U22897 ( .A1(n21921), .A2(n21926), .A3(n22332), .ZN(n21281) );
  AOI22_X1 U22898 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20808), .ZN(n20791) );
  OAI21_X1 U22899 ( .B1(n20792), .B2(n20844), .A(n20791), .ZN(P3_U2768) );
  AOI22_X1 U22900 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20808), .ZN(n20793) );
  OAI21_X1 U22901 ( .B1(n21357), .B2(n20844), .A(n20793), .ZN(P3_U2769) );
  AOI22_X1 U22902 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20808), .ZN(n20794) );
  OAI21_X1 U22903 ( .B1(n21359), .B2(n20844), .A(n20794), .ZN(P3_U2770) );
  AOI22_X1 U22904 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20808), .ZN(n20795) );
  OAI21_X1 U22905 ( .B1(n20796), .B2(n20844), .A(n20795), .ZN(P3_U2771) );
  AOI22_X1 U22906 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20808), .ZN(n20797) );
  OAI21_X1 U22907 ( .B1(n20798), .B2(n20844), .A(n20797), .ZN(P3_U2772) );
  AOI22_X1 U22908 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20808), .ZN(n20799) );
  OAI21_X1 U22909 ( .B1(n21346), .B2(n20844), .A(n20799), .ZN(P3_U2773) );
  AOI22_X1 U22910 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20808), .ZN(n20800) );
  OAI21_X1 U22911 ( .B1(n20801), .B2(n20844), .A(n20800), .ZN(P3_U2774) );
  AOI22_X1 U22912 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20808), .ZN(n20802) );
  OAI21_X1 U22913 ( .B1(n20803), .B2(n20844), .A(n20802), .ZN(P3_U2775) );
  AOI22_X1 U22914 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20808), .ZN(n20804) );
  OAI21_X1 U22915 ( .B1(n20805), .B2(n20844), .A(n20804), .ZN(P3_U2776) );
  AOI22_X1 U22916 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20808), .ZN(n20806) );
  OAI21_X1 U22917 ( .B1(n20807), .B2(n20844), .A(n20806), .ZN(P3_U2777) );
  AOI22_X1 U22918 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20841), .ZN(n20809) );
  OAI21_X1 U22919 ( .B1(n21377), .B2(n20844), .A(n20809), .ZN(P3_U2778) );
  AOI22_X1 U22920 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20841), .ZN(n20810) );
  OAI21_X1 U22921 ( .B1(n20811), .B2(n20844), .A(n20810), .ZN(P3_U2779) );
  AOI22_X1 U22922 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20842), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20841), .ZN(n20812) );
  OAI21_X1 U22923 ( .B1(n20813), .B2(n20844), .A(n20812), .ZN(P3_U2780) );
  AOI22_X1 U22924 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20826), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20841), .ZN(n20814) );
  OAI21_X1 U22925 ( .B1(n21391), .B2(n20844), .A(n20814), .ZN(P3_U2781) );
  AOI22_X1 U22926 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20826), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20841), .ZN(n20815) );
  OAI21_X1 U22927 ( .B1(n21387), .B2(n20844), .A(n20815), .ZN(P3_U2782) );
  AOI22_X1 U22928 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20826), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20841), .ZN(n20816) );
  OAI21_X1 U22929 ( .B1(n21457), .B2(n20844), .A(n20816), .ZN(P3_U2783) );
  AOI22_X1 U22930 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20826), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20841), .ZN(n20817) );
  OAI21_X1 U22931 ( .B1(n21446), .B2(n20844), .A(n20817), .ZN(P3_U2784) );
  AOI22_X1 U22932 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20826), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20841), .ZN(n20818) );
  OAI21_X1 U22933 ( .B1(n20819), .B2(n20844), .A(n20818), .ZN(P3_U2785) );
  AOI22_X1 U22934 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20826), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20841), .ZN(n20820) );
  OAI21_X1 U22935 ( .B1(n20821), .B2(n20844), .A(n20820), .ZN(P3_U2786) );
  AOI22_X1 U22936 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20826), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20841), .ZN(n20822) );
  OAI21_X1 U22937 ( .B1(n21308), .B2(n20844), .A(n20822), .ZN(P3_U2787) );
  AOI22_X1 U22938 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20826), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20841), .ZN(n20823) );
  OAI21_X1 U22939 ( .B1(n20824), .B2(n20844), .A(n20823), .ZN(P3_U2788) );
  AOI22_X1 U22940 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20826), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20841), .ZN(n20825) );
  OAI21_X1 U22941 ( .B1(n21309), .B2(n20844), .A(n20825), .ZN(P3_U2789) );
  AOI22_X1 U22942 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20826), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20841), .ZN(n20827) );
  OAI21_X1 U22943 ( .B1(n20828), .B2(n20844), .A(n20827), .ZN(P3_U2790) );
  AOI22_X1 U22944 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20842), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20841), .ZN(n20829) );
  OAI21_X1 U22945 ( .B1(n20830), .B2(n20844), .A(n20829), .ZN(P3_U2791) );
  AOI22_X1 U22946 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20842), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20841), .ZN(n20831) );
  OAI21_X1 U22947 ( .B1(n21283), .B2(n20844), .A(n20831), .ZN(P3_U2792) );
  AOI22_X1 U22948 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20842), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20841), .ZN(n20832) );
  OAI21_X1 U22949 ( .B1(n20833), .B2(n20844), .A(n20832), .ZN(P3_U2793) );
  AOI22_X1 U22950 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20842), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20841), .ZN(n20834) );
  OAI21_X1 U22951 ( .B1(n21295), .B2(n20844), .A(n20834), .ZN(P3_U2794) );
  AOI22_X1 U22952 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20842), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20841), .ZN(n20835) );
  OAI21_X1 U22953 ( .B1(n20836), .B2(n20844), .A(n20835), .ZN(P3_U2795) );
  AOI22_X1 U22954 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20842), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20841), .ZN(n20837) );
  OAI21_X1 U22955 ( .B1(n20838), .B2(n20844), .A(n20837), .ZN(P3_U2796) );
  AOI22_X1 U22956 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20842), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20841), .ZN(n20839) );
  OAI21_X1 U22957 ( .B1(n20840), .B2(n20844), .A(n20839), .ZN(P3_U2797) );
  AOI22_X1 U22958 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20842), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20841), .ZN(n20843) );
  OAI21_X1 U22959 ( .B1(n21430), .B2(n20844), .A(n20843), .ZN(P3_U2798) );
  NAND2_X1 U22960 ( .A1(n22332), .A2(n22278), .ZN(n20845) );
  NAND4_X1 U22961 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n20846), .A3(n21808), 
        .A4(n22278), .ZN(n21248) );
  INV_X1 U22962 ( .A(n21248), .ZN(n21934) );
  INV_X1 U22963 ( .A(n21929), .ZN(n20847) );
  NAND2_X1 U22964 ( .A1(n20847), .A2(n21930), .ZN(n21945) );
  AND2_X1 U22965 ( .A1(n20849), .A2(n21485), .ZN(n21466) );
  AOI22_X1 U22966 ( .A1(n21193), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n21466), 
        .B2(n20891), .ZN(n20860) );
  INV_X1 U22967 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21009) );
  NOR2_X1 U22968 ( .A1(n21114), .A2(n21248), .ZN(n21053) );
  INV_X1 U22969 ( .A(n21053), .ZN(n20887) );
  OAI21_X1 U22970 ( .B1(n21009), .B2(n20887), .A(n21228), .ZN(n20858) );
  AOI21_X1 U22971 ( .B1(n11463), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n21248), .ZN(n21059) );
  OAI211_X1 U22972 ( .C1(n20851), .C2(n20850), .A(n22332), .B(n22278), .ZN(
        n21928) );
  INV_X1 U22973 ( .A(n21928), .ZN(n20852) );
  OAI22_X1 U22974 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n21269), .B1(n21268), 
        .B2(n20855), .ZN(n20856) );
  AOI221_X1 U22975 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20858), .C1(
        n20857), .C2(n21059), .A(n20856), .ZN(n20859) );
  OAI211_X1 U22976 ( .C1(n21267), .C2(n20861), .A(n20860), .B(n20859), .ZN(
        P3_U2670) );
  INV_X1 U22977 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20872) );
  NOR2_X1 U22978 ( .A1(n11463), .A2(n21179), .ZN(n21092) );
  NAND2_X1 U22979 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n21009), .ZN(
        n21066) );
  OAI21_X1 U22980 ( .B1(n20862), .B2(n21066), .A(n11463), .ZN(n20873) );
  AOI211_X1 U22981 ( .C1(n20869), .C2(n21066), .A(n21248), .B(n20873), .ZN(
        n20868) );
  INV_X1 U22982 ( .A(n20891), .ZN(n21275) );
  NAND2_X1 U22983 ( .A1(n21491), .A2(n21485), .ZN(n21489) );
  INV_X1 U22984 ( .A(n21489), .ZN(n21488) );
  OR2_X1 U22985 ( .A1(n20878), .A2(n21488), .ZN(n21476) );
  AOI22_X1 U22986 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n21254), .B1(
        n21193), .B2(P3_REIP_REG_2__SCAN_IN), .ZN(n20866) );
  NOR2_X1 U22987 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n20864) );
  NOR3_X1 U22988 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20883) );
  INV_X1 U22989 ( .A(n20883), .ZN(n20863) );
  OAI211_X1 U22990 ( .C1(n20864), .C2(n20872), .A(n21235), .B(n20863), .ZN(
        n20865) );
  OAI211_X1 U22991 ( .C1(n21275), .C2(n21476), .A(n20866), .B(n20865), .ZN(
        n20867) );
  AOI211_X1 U22992 ( .C1(n20869), .C2(n21092), .A(n20868), .B(n20867), .ZN(
        n20871) );
  NAND2_X1 U22993 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n20875) );
  OAI211_X1 U22994 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n21232), .B(n20875), .ZN(n20870) );
  OAI211_X1 U22995 ( .C1(n20872), .C2(n21268), .A(n20871), .B(n20870), .ZN(
        P3_U2669) );
  XOR2_X1 U22996 ( .A(n20874), .B(n20873), .Z(n20881) );
  NAND3_X1 U22997 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n20901) );
  AOI21_X1 U22998 ( .B1(n21232), .B2(n20901), .A(n21193), .ZN(n20900) );
  AOI221_X1 U22999 ( .B1(n21269), .B2(n20876), .C1(n20875), .C2(n20876), .A(
        n20900), .ZN(n20880) );
  NOR2_X1 U23000 ( .A1(n20878), .A2(n20877), .ZN(n21497) );
  NOR2_X1 U23001 ( .A1(n18468), .A2(n21497), .ZN(n21506) );
  OAI22_X1 U23002 ( .A1(n21506), .A2(n21275), .B1(n21268), .B2(n20882), .ZN(
        n20879) );
  AOI211_X1 U23003 ( .C1(n21934), .C2(n20881), .A(n20880), .B(n20879), .ZN(
        n20885) );
  NAND2_X1 U23004 ( .A1(n20883), .A2(n20882), .ZN(n20888) );
  OAI211_X1 U23005 ( .C1(n20883), .C2(n20882), .A(n21235), .B(n20888), .ZN(
        n20884) );
  OAI211_X1 U23006 ( .C1(n21228), .C2(n20886), .A(n20885), .B(n20884), .ZN(
        P3_U2668) );
  AOI211_X1 U23007 ( .C1(n20905), .C2(n21009), .A(n20889), .B(n20887), .ZN(
        n20898) );
  NOR2_X1 U23008 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20888), .ZN(n20911) );
  AOI211_X1 U23009 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20888), .A(n20911), .B(
        n21267), .ZN(n20897) );
  NOR3_X1 U23010 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n21269), .A3(n20901), .ZN(
        n20896) );
  AOI22_X1 U23011 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n21254), .B1(
        n21253), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n20894) );
  OAI211_X1 U23012 ( .C1(n21114), .C2(n20890), .A(n20889), .B(n21059), .ZN(
        n20893) );
  OAI21_X1 U23013 ( .B1(n12577), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n20891), .ZN(n20892) );
  NAND4_X1 U23014 ( .A1(n20894), .A2(n21868), .A3(n20893), .A4(n20892), .ZN(
        n20895) );
  NOR4_X1 U23015 ( .A1(n20898), .A2(n20897), .A3(n20896), .A4(n20895), .ZN(
        n20899) );
  OAI21_X1 U23016 ( .B1(n20902), .B2(n20900), .A(n20899), .ZN(P3_U2667) );
  AOI22_X1 U23017 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n21254), .B1(
        n21253), .B2(P3_EBX_REG_5__SCAN_IN), .ZN(n20915) );
  NOR2_X1 U23018 ( .A1(n20902), .A2(n20901), .ZN(n20904) );
  NAND2_X1 U23019 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n20904), .ZN(n20928) );
  NAND2_X1 U23020 ( .A1(n20928), .A2(n21232), .ZN(n20908) );
  INV_X1 U23021 ( .A(n20908), .ZN(n20903) );
  AOI21_X1 U23022 ( .B1(n20904), .B2(n20903), .A(n21801), .ZN(n20914) );
  AOI21_X1 U23023 ( .B1(n20905), .B2(n21009), .A(n21114), .ZN(n20907) );
  XNOR2_X1 U23024 ( .A(n20907), .B(n20906), .ZN(n20909) );
  NAND2_X1 U23025 ( .A1(n21272), .A2(n20908), .ZN(n20934) );
  AOI22_X1 U23026 ( .A1(n21934), .A2(n20909), .B1(P3_REIP_REG_5__SCAN_IN), 
        .B2(n20934), .ZN(n20913) );
  NAND2_X1 U23027 ( .A1(n20911), .A2(n20910), .ZN(n20916) );
  OAI211_X1 U23028 ( .C1(n20911), .C2(n20910), .A(n21235), .B(n20916), .ZN(
        n20912) );
  NAND4_X1 U23029 ( .A1(n20915), .A2(n20914), .A3(n20913), .A4(n20912), .ZN(
        P3_U2666) );
  NOR3_X1 U23030 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n21269), .A3(n20928), .ZN(
        n20935) );
  AOI211_X1 U23031 ( .C1(n21253), .C2(P3_EBX_REG_6__SCAN_IN), .A(n21886), .B(
        n20935), .ZN(n20925) );
  AOI211_X1 U23032 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20916), .A(n20936), .B(
        n21267), .ZN(n20920) );
  NAND2_X1 U23033 ( .A1(n20917), .A2(n21009), .ZN(n20958) );
  NAND3_X1 U23034 ( .A1(n21934), .A2(n11463), .A3(n20958), .ZN(n20918) );
  OAI22_X1 U23035 ( .A1(n20921), .A2(n20918), .B1(n20922), .B2(n21228), .ZN(
        n20919) );
  AOI211_X1 U23036 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n20934), .A(n20920), .B(
        n20919), .ZN(n20924) );
  OAI211_X1 U23037 ( .C1(n21092), .C2(n20922), .A(n20921), .B(n21059), .ZN(
        n20923) );
  NAND3_X1 U23038 ( .A1(n20925), .A2(n20924), .A3(n20923), .ZN(P3_U2665) );
  NAND2_X1 U23039 ( .A1(n11463), .A2(n20958), .ZN(n20926) );
  XNOR2_X1 U23040 ( .A(n20927), .B(n20926), .ZN(n20932) );
  NOR2_X1 U23041 ( .A1(n20929), .A2(n20928), .ZN(n20945) );
  NOR2_X1 U23042 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n21269), .ZN(n20930) );
  AOI22_X1 U23043 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n21254), .B1(
        n20945), .B2(n20930), .ZN(n20931) );
  OAI211_X1 U23044 ( .C1(n21179), .C2(n20932), .A(n20931), .B(n21868), .ZN(
        n20933) );
  AOI221_X1 U23045 ( .B1(n20935), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n20934), 
        .C2(P3_REIP_REG_7__SCAN_IN), .A(n20933), .ZN(n20938) );
  NAND2_X1 U23046 ( .A1(n20936), .A2(n20939), .ZN(n20943) );
  OAI211_X1 U23047 ( .C1(n20936), .C2(n20939), .A(n21235), .B(n20943), .ZN(
        n20937) );
  OAI211_X1 U23048 ( .C1(n20939), .C2(n21268), .A(n20938), .B(n20937), .ZN(
        P3_U2664) );
  OAI21_X1 U23049 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20940), .A(
        n11463), .ZN(n20941) );
  XOR2_X1 U23050 ( .A(n20942), .B(n20941), .Z(n20951) );
  NOR2_X1 U23051 ( .A1(n20970), .A2(n21267), .ZN(n20952) );
  NAND2_X1 U23052 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20943), .ZN(n20944) );
  AOI22_X1 U23053 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n21254), .B1(
        n20952), .B2(n20944), .ZN(n20950) );
  NAND2_X1 U23054 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20945), .ZN(n20946) );
  NOR2_X1 U23055 ( .A1(n20947), .A2(n20946), .ZN(n20972) );
  OAI21_X1 U23056 ( .B1(n20972), .B2(n21269), .A(n21272), .ZN(n20978) );
  INV_X1 U23057 ( .A(n20978), .ZN(n20953) );
  AOI221_X1 U23058 ( .B1(n21269), .B2(n20947), .C1(n20946), .C2(n20947), .A(
        n20953), .ZN(n20948) );
  AOI211_X1 U23059 ( .C1(n21253), .C2(P3_EBX_REG_8__SCAN_IN), .A(n21886), .B(
        n20948), .ZN(n20949) );
  OAI211_X1 U23060 ( .C1(n21179), .C2(n20951), .A(n20950), .B(n20949), .ZN(
        P3_U2663) );
  NOR2_X1 U23061 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n21269), .ZN(n20979) );
  AOI22_X1 U23062 ( .A1(n20979), .A2(n20972), .B1(n20952), .B2(n20969), .ZN(
        n20966) );
  AOI21_X1 U23063 ( .B1(n21235), .B2(n20970), .A(n21253), .ZN(n20955) );
  OAI22_X1 U23064 ( .A1(n20969), .A2(n20955), .B1(n20954), .B2(n20953), .ZN(
        n20956) );
  INV_X1 U23065 ( .A(n20956), .ZN(n20965) );
  INV_X1 U23066 ( .A(n20957), .ZN(n20961) );
  OAI21_X1 U23067 ( .B1(n20959), .B2(n20958), .A(n11463), .ZN(n20967) );
  NOR3_X1 U23068 ( .A1(n20961), .A2(n21248), .A3(n20967), .ZN(n20960) );
  AOI211_X1 U23069 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n21254), .A(
        n21801), .B(n20960), .ZN(n20964) );
  OAI211_X1 U23070 ( .C1(n20962), .C2(n21092), .A(n20961), .B(n21059), .ZN(
        n20963) );
  NAND4_X1 U23071 ( .A1(n20966), .A2(n20965), .A3(n20964), .A4(n20963), .ZN(
        P3_U2662) );
  XOR2_X1 U23072 ( .A(n20968), .B(n20967), .Z(n20982) );
  NAND2_X1 U23073 ( .A1(n20970), .A2(n20969), .ZN(n20971) );
  AOI211_X1 U23074 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20971), .A(n20991), .B(
        n21267), .ZN(n20977) );
  NAND2_X1 U23075 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20972), .ZN(n20983) );
  NOR3_X1 U23076 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n21269), .A3(n20983), 
        .ZN(n20976) );
  OAI22_X1 U23077 ( .A1(n20974), .A2(n21228), .B1(n21268), .B2(n20973), .ZN(
        n20975) );
  NOR4_X1 U23078 ( .A1(n21801), .A2(n20977), .A3(n20976), .A4(n20975), .ZN(
        n20981) );
  OAI21_X1 U23079 ( .B1(n20979), .B2(n20978), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n20980) );
  OAI211_X1 U23080 ( .C1(n21179), .C2(n20982), .A(n20981), .B(n20980), .ZN(
        P3_U2661) );
  NOR2_X1 U23081 ( .A1(n20984), .A2(n20983), .ZN(n21000) );
  NAND2_X1 U23082 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n21000), .ZN(n21154) );
  AOI21_X1 U23083 ( .B1(n21154), .B2(n21232), .A(n21193), .ZN(n21028) );
  NAND2_X1 U23084 ( .A1(n21232), .A2(n21000), .ZN(n20996) );
  OAI21_X1 U23085 ( .B1(n18549), .B2(n21066), .A(n11463), .ZN(n21002) );
  INV_X1 U23086 ( .A(n21002), .ZN(n20988) );
  INV_X1 U23087 ( .A(n20985), .ZN(n20986) );
  AOI221_X1 U23088 ( .B1(n20986), .B2(n20989), .C1(n21066), .C2(n20989), .A(
        n21248), .ZN(n20987) );
  OAI22_X1 U23089 ( .A1(n20989), .A2(n20988), .B1(n21092), .B2(n20987), .ZN(
        n20993) );
  INV_X1 U23090 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20990) );
  NAND2_X1 U23091 ( .A1(n20991), .A2(n20990), .ZN(n20998) );
  OAI211_X1 U23092 ( .C1(n20991), .C2(n20990), .A(n21235), .B(n20998), .ZN(
        n20992) );
  OAI211_X1 U23093 ( .C1(n21228), .C2(n11470), .A(n20993), .B(n20992), .ZN(
        n20994) );
  AOI211_X1 U23094 ( .C1(n21253), .C2(P3_EBX_REG_11__SCAN_IN), .A(n21801), .B(
        n20994), .ZN(n20995) );
  OAI221_X1 U23095 ( .B1(n21028), .B2(n20997), .C1(n21028), .C2(n20996), .A(
        n20995), .ZN(P3_U2660) );
  AOI211_X1 U23096 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20998), .A(n21014), .B(
        n21267), .ZN(n20999) );
  AOI211_X1 U23097 ( .C1(n21253), .C2(P3_EBX_REG_12__SCAN_IN), .A(n21886), .B(
        n20999), .ZN(n21007) );
  NAND3_X1 U23098 ( .A1(n21232), .A2(P3_REIP_REG_11__SCAN_IN), .A3(n21000), 
        .ZN(n21152) );
  INV_X1 U23099 ( .A(n21028), .ZN(n21076) );
  OAI21_X1 U23100 ( .B1(n21003), .B2(n21002), .A(n21934), .ZN(n21001) );
  AOI21_X1 U23101 ( .B1(n21003), .B2(n21002), .A(n21001), .ZN(n21004) );
  AOI221_X1 U23102 ( .B1(n21087), .B2(n21005), .C1(n21076), .C2(
        P3_REIP_REG_12__SCAN_IN), .A(n21004), .ZN(n21006) );
  OAI211_X1 U23103 ( .C1(n21008), .C2(n21228), .A(n21007), .B(n21006), .ZN(
        P3_U2659) );
  NAND2_X1 U23104 ( .A1(n21934), .A2(n21009), .ZN(n21011) );
  INV_X1 U23105 ( .A(n21092), .ZN(n21010) );
  OAI21_X1 U23106 ( .B1(n21012), .B2(n21011), .A(n21010), .ZN(n21019) );
  AOI22_X1 U23107 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n21254), .B1(
        n21253), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n21017) );
  NAND2_X1 U23108 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_12__SCAN_IN), 
        .ZN(n21031) );
  OAI211_X1 U23109 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(P3_REIP_REG_12__SCAN_IN), .A(n21087), .B(n21031), .ZN(n21016) );
  NAND2_X1 U23110 ( .A1(n21014), .A2(n21013), .ZN(n21032) );
  OAI211_X1 U23111 ( .C1(n21014), .C2(n21013), .A(n21235), .B(n21032), .ZN(
        n21015) );
  NAND4_X1 U23112 ( .A1(n21017), .A2(n21868), .A3(n21016), .A4(n21015), .ZN(
        n21018) );
  AOI21_X1 U23113 ( .B1(n21021), .B2(n21019), .A(n21018), .ZN(n21024) );
  NOR3_X1 U23114 ( .A1(n18549), .A2(n21020), .A3(n21066), .ZN(n21038) );
  NOR2_X1 U23115 ( .A1(n21038), .A2(n21114), .ZN(n21027) );
  INV_X1 U23116 ( .A(n21021), .ZN(n21022) );
  NAND3_X1 U23117 ( .A1(n21934), .A2(n21027), .A3(n21022), .ZN(n21023) );
  OAI211_X1 U23118 ( .C1(n21028), .C2(n21025), .A(n21024), .B(n21023), .ZN(
        P3_U2658) );
  XOR2_X1 U23119 ( .A(n21027), .B(n21026), .Z(n21037) );
  AOI21_X1 U23120 ( .B1(n21253), .B2(P3_EBX_REG_14__SCAN_IN), .A(n21801), .ZN(
        n21036) );
  NOR2_X1 U23121 ( .A1(n21030), .A2(n21031), .ZN(n21073) );
  OAI21_X1 U23122 ( .B1(n21073), .B2(n21269), .A(n21028), .ZN(n21057) );
  INV_X1 U23123 ( .A(n21057), .ZN(n21029) );
  AOI221_X1 U23124 ( .B1(n21031), .B2(n21030), .C1(n21152), .C2(n21030), .A(
        n21029), .ZN(n21034) );
  AOI211_X1 U23125 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n21032), .A(n21044), .B(
        n21267), .ZN(n21033) );
  AOI211_X1 U23126 ( .C1(n21254), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n21034), .B(n21033), .ZN(n21035) );
  OAI211_X1 U23127 ( .C1(n21248), .C2(n21037), .A(n21036), .B(n21035), .ZN(
        P3_U2657) );
  AOI22_X1 U23128 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n21254), .B1(
        n21253), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n21047) );
  AND2_X1 U23129 ( .A1(n21073), .A2(n21087), .ZN(n21056) );
  NAND2_X1 U23130 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n21038), .ZN(
        n21050) );
  NAND2_X1 U23131 ( .A1(n11463), .A2(n21050), .ZN(n21040) );
  OAI21_X1 U23132 ( .B1(n21041), .B2(n21040), .A(n21934), .ZN(n21039) );
  AOI21_X1 U23133 ( .B1(n21041), .B2(n21040), .A(n21039), .ZN(n21042) );
  AOI221_X1 U23134 ( .B1(n21056), .B2(n21054), .C1(n21057), .C2(
        P3_REIP_REG_15__SCAN_IN), .A(n21042), .ZN(n21046) );
  NAND2_X1 U23135 ( .A1(n21044), .A2(n21043), .ZN(n21048) );
  OAI211_X1 U23136 ( .C1(n21044), .C2(n21043), .A(n21235), .B(n21048), .ZN(
        n21045) );
  NAND4_X1 U23137 ( .A1(n21047), .A2(n21046), .A3(n21868), .A4(n21045), .ZN(
        P3_U2656) );
  AOI211_X1 U23138 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n21048), .A(n21070), .B(
        n21267), .ZN(n21049) );
  AOI211_X1 U23139 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n21254), .A(
        n21886), .B(n21049), .ZN(n21065) );
  NOR2_X1 U23140 ( .A1(n21051), .A2(n21050), .ZN(n21115) );
  NOR2_X1 U23141 ( .A1(n21115), .A2(n21060), .ZN(n21052) );
  AOI22_X1 U23142 ( .A1(n21253), .A2(P3_EBX_REG_16__SCAN_IN), .B1(n21053), 
        .B2(n21052), .ZN(n21064) );
  XNOR2_X1 U23143 ( .A(P3_REIP_REG_16__SCAN_IN), .B(n21054), .ZN(n21055) );
  AOI22_X1 U23144 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n21057), .B1(n21056), 
        .B2(n21055), .ZN(n21063) );
  INV_X1 U23145 ( .A(n21058), .ZN(n21061) );
  OAI211_X1 U23146 ( .C1(n21061), .C2(n21114), .A(n21060), .B(n21059), .ZN(
        n21062) );
  NAND4_X1 U23147 ( .A1(n21065), .A2(n21064), .A3(n21063), .A4(n21062), .ZN(
        P3_U2655) );
  OAI21_X1 U23148 ( .B1(n21067), .B2(n21066), .A(n11463), .ZN(n21068) );
  XNOR2_X1 U23149 ( .A(n21069), .B(n21068), .ZN(n21083) );
  NAND2_X1 U23150 ( .A1(n21070), .A2(n21072), .ZN(n21084) );
  OAI211_X1 U23151 ( .C1(n21070), .C2(n21072), .A(n21235), .B(n21084), .ZN(
        n21071) );
  OAI211_X1 U23152 ( .C1(n21268), .C2(n21072), .A(n21868), .B(n21071), .ZN(
        n21081) );
  NAND3_X1 U23153 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n21073), .ZN(n21074) );
  NOR2_X1 U23154 ( .A1(n21074), .A2(n21152), .ZN(n21079) );
  NOR2_X1 U23155 ( .A1(n21075), .A2(n21074), .ZN(n21151) );
  INV_X1 U23156 ( .A(n21151), .ZN(n21077) );
  AOI21_X1 U23157 ( .B1(n21232), .B2(n21077), .A(n21076), .ZN(n21113) );
  INV_X1 U23158 ( .A(n21113), .ZN(n21078) );
  MUX2_X1 U23159 ( .A(n21079), .B(n21078), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n21080) );
  AOI211_X1 U23160 ( .C1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n21254), .A(
        n21081), .B(n21080), .ZN(n21082) );
  OAI21_X1 U23161 ( .B1(n21179), .B2(n21083), .A(n21082), .ZN(P3_U2654) );
  AOI211_X1 U23162 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n21084), .A(n21100), .B(
        n21267), .ZN(n21097) );
  INV_X1 U23163 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n21085) );
  OAI22_X1 U23164 ( .A1(n21086), .A2(n21228), .B1(n21268), .B2(n21085), .ZN(
        n21096) );
  NAND2_X1 U23165 ( .A1(n21151), .A2(n21087), .ZN(n21111) );
  AOI21_X1 U23166 ( .B1(n21115), .B2(n21088), .A(n21114), .ZN(n21098) );
  INV_X1 U23167 ( .A(n21115), .ZN(n21090) );
  AOI221_X1 U23168 ( .B1(n21090), .B2(n21093), .C1(n21089), .C2(n21093), .A(
        n21179), .ZN(n21091) );
  OAI22_X1 U23169 ( .A1(n21093), .A2(n21098), .B1(n21092), .B2(n21091), .ZN(
        n21094) );
  OAI221_X1 U23170 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n21111), .C1(n21833), 
        .C2(n21113), .A(n21094), .ZN(n21095) );
  OR4_X1 U23171 ( .A1(n21886), .A2(n21097), .A3(n21096), .A4(n21095), .ZN(
        P3_U2653) );
  XOR2_X1 U23172 ( .A(n21099), .B(n21098), .Z(n21108) );
  NAND2_X1 U23173 ( .A1(n21100), .A2(n21102), .ZN(n21109) );
  OAI211_X1 U23174 ( .C1(n21100), .C2(n21102), .A(n21235), .B(n21109), .ZN(
        n21101) );
  OAI211_X1 U23175 ( .C1(n21268), .C2(n21102), .A(n21868), .B(n21101), .ZN(
        n21106) );
  NAND2_X1 U23176 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n21112) );
  OAI21_X1 U23177 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(P3_REIP_REG_19__SCAN_IN), 
        .A(n21112), .ZN(n21103) );
  OAI22_X1 U23178 ( .A1(n21113), .A2(n21104), .B1(n21111), .B2(n21103), .ZN(
        n21105) );
  AOI211_X1 U23179 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n21254), .A(
        n21106), .B(n21105), .ZN(n21107) );
  OAI21_X1 U23180 ( .B1(n21179), .B2(n21108), .A(n21107), .ZN(P3_U2652) );
  AOI211_X1 U23181 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n21109), .A(n21130), .B(
        n21267), .ZN(n21110) );
  AOI21_X1 U23182 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n21253), .A(n21110), .ZN(
        n21122) );
  NOR2_X1 U23183 ( .A1(n21112), .A2(n21111), .ZN(n21124) );
  NOR2_X1 U23184 ( .A1(n21120), .A2(n21112), .ZN(n21150) );
  OAI21_X1 U23185 ( .B1(n21150), .B2(n21269), .A(n21113), .ZN(n21146) );
  NOR2_X1 U23186 ( .A1(n21118), .A2(n21117), .ZN(n21126) );
  AOI211_X1 U23187 ( .C1(n21118), .C2(n21117), .A(n21126), .B(n21179), .ZN(
        n21119) );
  AOI221_X1 U23188 ( .B1(n21124), .B2(n21120), .C1(n21146), .C2(
        P3_REIP_REG_20__SCAN_IN), .A(n21119), .ZN(n21121) );
  OAI211_X1 U23189 ( .C1(n21123), .C2(n21228), .A(n21122), .B(n21121), .ZN(
        P3_U2651) );
  NAND2_X1 U23190 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n21124), .ZN(n21139) );
  INV_X1 U23191 ( .A(n21146), .ZN(n21136) );
  INV_X1 U23192 ( .A(n21125), .ZN(n21128) );
  AOI211_X1 U23193 ( .C1(n21128), .C2(n21127), .A(n21142), .B(n21179), .ZN(
        n21134) );
  NAND2_X1 U23194 ( .A1(n21130), .A2(n21129), .ZN(n21137) );
  OAI211_X1 U23195 ( .C1(n21130), .C2(n21129), .A(n21235), .B(n21137), .ZN(
        n21131) );
  OAI21_X1 U23196 ( .B1(n21228), .B2(n21132), .A(n21131), .ZN(n21133) );
  AOI211_X1 U23197 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n21253), .A(n21134), .B(
        n21133), .ZN(n21135) );
  OAI221_X1 U23198 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n21139), .C1(n21140), 
        .C2(n21136), .A(n21135), .ZN(P3_U2650) );
  AOI211_X1 U23199 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n21137), .A(n21162), .B(
        n21267), .ZN(n21138) );
  AOI21_X1 U23200 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n21253), .A(n21138), .ZN(
        n21148) );
  AOI221_X1 U23201 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n21141), .C2(n21140), .A(n21139), .ZN(n21145) );
  AOI211_X1 U23202 ( .C1(n21143), .C2(n11282), .A(n21155), .B(n21179), .ZN(
        n21144) );
  AOI211_X1 U23203 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n21146), .A(n21145), 
        .B(n21144), .ZN(n21147) );
  OAI211_X1 U23204 ( .C1(n21149), .C2(n21228), .A(n21148), .B(n21147), .ZN(
        P3_U2649) );
  AOI22_X1 U23205 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n21254), .B1(
        n21253), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n21165) );
  NAND4_X1 U23206 ( .A1(n21151), .A2(n21150), .A3(P3_REIP_REG_22__SCAN_IN), 
        .A4(P3_REIP_REG_21__SCAN_IN), .ZN(n21153) );
  NOR2_X1 U23207 ( .A1(n21153), .A2(n21152), .ZN(n21160) );
  NOR3_X1 U23208 ( .A1(n21159), .A2(n21154), .A3(n21153), .ZN(n21181) );
  OAI21_X1 U23209 ( .B1(n21181), .B2(n21269), .A(n21272), .ZN(n21176) );
  NOR2_X1 U23210 ( .A1(n21155), .A2(n21114), .ZN(n21156) );
  AOI211_X1 U23211 ( .C1(n21157), .C2(n21156), .A(n21166), .B(n21179), .ZN(
        n21158) );
  AOI221_X1 U23212 ( .B1(n21160), .B2(n21159), .C1(n21176), .C2(
        P3_REIP_REG_23__SCAN_IN), .A(n21158), .ZN(n21164) );
  NAND2_X1 U23213 ( .A1(n21162), .A2(n21161), .ZN(n21169) );
  OAI211_X1 U23214 ( .C1(n21162), .C2(n21161), .A(n21235), .B(n21169), .ZN(
        n21163) );
  NAND3_X1 U23215 ( .A1(n21165), .A2(n21164), .A3(n21163), .ZN(P3_U2648) );
  INV_X1 U23216 ( .A(n21176), .ZN(n21175) );
  AOI22_X1 U23217 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n21254), .B1(
        n21253), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n21174) );
  NOR2_X1 U23218 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21269), .ZN(n21172) );
  NOR2_X1 U23219 ( .A1(n21166), .A2(n21114), .ZN(n21167) );
  AOI211_X1 U23220 ( .C1(n21168), .C2(n21167), .A(n21178), .B(n21179), .ZN(
        n21171) );
  NOR2_X1 U23221 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n21169), .ZN(n21187) );
  AOI211_X1 U23222 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n21169), .A(n21187), .B(
        n21267), .ZN(n21170) );
  AOI211_X1 U23223 ( .C1(n21172), .C2(n21181), .A(n21171), .B(n21170), .ZN(
        n21173) );
  OAI211_X1 U23224 ( .C1(n21175), .C2(n21177), .A(n21174), .B(n21173), .ZN(
        P3_U2647) );
  AOI21_X1 U23225 ( .B1(n21232), .B2(n21177), .A(n21176), .ZN(n21190) );
  AOI211_X1 U23226 ( .C1(n21180), .C2(n11290), .A(n21196), .B(n21179), .ZN(
        n21185) );
  NAND2_X1 U23227 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21181), .ZN(n21191) );
  NAND2_X1 U23228 ( .A1(n21232), .A2(n21192), .ZN(n21182) );
  OAI22_X1 U23229 ( .A1(n21183), .A2(n21228), .B1(n21191), .B2(n21182), .ZN(
        n21184) );
  AOI211_X1 U23230 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n21253), .A(n21185), .B(
        n21184), .ZN(n21189) );
  NAND2_X1 U23231 ( .A1(n21187), .A2(n21186), .ZN(n21195) );
  OAI211_X1 U23232 ( .C1(n21187), .C2(n21186), .A(n21235), .B(n21195), .ZN(
        n21188) );
  OAI211_X1 U23233 ( .C1(n21190), .C2(n21192), .A(n21189), .B(n21188), .ZN(
        P3_U2646) );
  OR2_X1 U23234 ( .A1(n21192), .A2(n21191), .ZN(n21194) );
  NOR2_X1 U23235 ( .A1(n21269), .A2(n21194), .ZN(n21208) );
  AOI22_X1 U23236 ( .A1(n21253), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n21208), 
        .B2(n21716), .ZN(n21202) );
  AOI221_X1 U23237 ( .B1(n21232), .B2(n21716), .C1(n21232), .C2(n21194), .A(
        n21193), .ZN(n21218) );
  INV_X1 U23238 ( .A(n21218), .ZN(n21231) );
  NOR2_X1 U23239 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n21195), .ZN(n21213) );
  AOI211_X1 U23240 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n21195), .A(n21213), .B(
        n21267), .ZN(n21200) );
  AOI211_X1 U23241 ( .C1(n21198), .C2(n21197), .A(n21205), .B(n21248), .ZN(
        n21199) );
  AOI211_X1 U23242 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n21231), .A(n21200), 
        .B(n21199), .ZN(n21201) );
  OAI211_X1 U23243 ( .C1(n21203), .C2(n21228), .A(n21202), .B(n21201), .ZN(
        P3_U2645) );
  INV_X1 U23244 ( .A(n21204), .ZN(n21207) );
  NOR2_X1 U23245 ( .A1(n21205), .A2(n21114), .ZN(n21206) );
  NOR2_X1 U23246 ( .A1(n21207), .A2(n21206), .ZN(n21220) );
  AOI211_X1 U23247 ( .C1(n21207), .C2(n21206), .A(n21220), .B(n21248), .ZN(
        n21211) );
  NAND2_X1 U23248 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n21208), .ZN(n21245) );
  OAI22_X1 U23249 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n21245), .B1(n21209), 
        .B2(n21228), .ZN(n21210) );
  AOI211_X1 U23250 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n21253), .A(n21211), .B(
        n21210), .ZN(n21215) );
  INV_X1 U23251 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n21212) );
  NAND2_X1 U23252 ( .A1(n21213), .A2(n21212), .ZN(n21219) );
  OAI211_X1 U23253 ( .C1(n21213), .C2(n21212), .A(n21235), .B(n21219), .ZN(
        n21214) );
  OAI211_X1 U23254 ( .C1(n21218), .C2(n21216), .A(n21215), .B(n21214), .ZN(
        P3_U2644) );
  NOR2_X1 U23255 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n21245), .ZN(n21217) );
  AOI22_X1 U23256 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n21217), .B1(n21253), 
        .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n21227) );
  OAI21_X1 U23257 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n21245), .A(n21218), 
        .ZN(n21225) );
  NOR2_X1 U23258 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n21219), .ZN(n21234) );
  AOI211_X1 U23259 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n21219), .A(n21234), .B(
        n21267), .ZN(n21224) );
  NOR2_X1 U23260 ( .A1(n21220), .A2(n21114), .ZN(n21221) );
  AOI211_X1 U23261 ( .C1(n21222), .C2(n21221), .A(n21237), .B(n21248), .ZN(
        n21223) );
  AOI211_X1 U23262 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n21225), .A(n21224), 
        .B(n21223), .ZN(n21226) );
  OAI211_X1 U23263 ( .C1(n21229), .C2(n21228), .A(n21227), .B(n21226), .ZN(
        P3_U2643) );
  NAND3_X1 U23264 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n21230), .ZN(n21244) );
  AOI22_X1 U23265 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n21254), .B1(
        n21253), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n21243) );
  NAND3_X1 U23266 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n21246) );
  AOI21_X1 U23267 ( .B1(n21232), .B2(n21246), .A(n21231), .ZN(n21252) );
  INV_X1 U23268 ( .A(n21252), .ZN(n21257) );
  INV_X1 U23269 ( .A(n21234), .ZN(n21236) );
  NAND2_X1 U23270 ( .A1(n21234), .A2(n21233), .ZN(n21247) );
  NAND2_X1 U23271 ( .A1(n21235), .A2(n21247), .ZN(n21249) );
  AOI21_X1 U23272 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n21236), .A(n21249), .ZN(
        n21241) );
  AOI211_X1 U23273 ( .C1(n21239), .C2(n21238), .A(n21259), .B(n21248), .ZN(
        n21240) );
  AOI211_X1 U23274 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n21257), .A(n21241), 
        .B(n21240), .ZN(n21242) );
  OAI211_X1 U23275 ( .C1(n21245), .C2(n21244), .A(n21243), .B(n21242), .ZN(
        P3_U2642) );
  NOR2_X1 U23276 ( .A1(n21246), .A2(n21245), .ZN(n21260) );
  AOI22_X1 U23277 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n21254), .B1(
        n21260), .B2(n21261), .ZN(n21251) );
  NOR2_X1 U23278 ( .A1(n21267), .A2(n21247), .ZN(n21256) );
  OAI211_X1 U23279 ( .C1(n21252), .C2(n21261), .A(n21251), .B(n21250), .ZN(
        P3_U2641) );
  AOI22_X1 U23280 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n21254), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n21253), .ZN(n21266) );
  INV_X1 U23281 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n21255) );
  AOI22_X1 U23282 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n21257), .B1(n21256), 
        .B2(n21255), .ZN(n21265) );
  NAND4_X1 U23283 ( .A1(n11463), .A2(n21934), .A3(n21259), .A4(n21258), .ZN(
        n21264) );
  OAI221_X1 U23284 ( .B1(P3_REIP_REG_31__SCAN_IN), .B2(P3_REIP_REG_30__SCAN_IN), .C1(n21262), .C2(n21261), .A(n21260), .ZN(n21263) );
  NAND4_X1 U23285 ( .A1(n21266), .A2(n21265), .A3(n21264), .A4(n21263), .ZN(
        P3_U2640) );
  NAND2_X1 U23286 ( .A1(n21268), .A2(n21267), .ZN(n21271) );
  NAND2_X1 U23287 ( .A1(n21272), .A2(n21269), .ZN(n21270) );
  AOI22_X1 U23288 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n21271), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n21270), .ZN(n21274) );
  NAND3_X1 U23289 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21272), .A3(
        n21507), .ZN(n21273) );
  OAI211_X1 U23290 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n21275), .A(
        n21274), .B(n21273), .ZN(P3_U2671) );
  NAND3_X1 U23291 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .ZN(n21307) );
  NAND4_X1 U23292 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n21276) );
  NOR3_X1 U23293 ( .A1(n21307), .A2(n21309), .A3(n21276), .ZN(n21334) );
  INV_X1 U23294 ( .A(n21334), .ZN(n21437) );
  NAND3_X1 U23295 ( .A1(n21279), .A2(n21278), .A3(n21277), .ZN(n21280) );
  NAND2_X1 U23296 ( .A1(n21438), .A2(n21456), .ZN(n21458) );
  NAND2_X1 U23297 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21435), .ZN(n21301) );
  NAND2_X1 U23298 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n21305), .ZN(n21296) );
  NOR2_X1 U23299 ( .A1(n21295), .A2(n21296), .ZN(n21289) );
  NAND2_X1 U23300 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n21289), .ZN(n21288) );
  NAND3_X1 U23301 ( .A1(n21447), .A2(P3_EAX_REG_13__SCAN_IN), .A3(n21288), 
        .ZN(n21287) );
  NAND2_X1 U23302 ( .A1(n21284), .A2(n21456), .ZN(n21443) );
  AOI22_X1 U23303 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21454), .B1(n21453), .B2(
        n21285), .ZN(n21286) );
  OAI211_X1 U23304 ( .C1(P3_EAX_REG_13__SCAN_IN), .C2(n21288), .A(n21287), .B(
        n21286), .ZN(P3_U2722) );
  INV_X1 U23305 ( .A(n21288), .ZN(n21424) );
  AOI21_X1 U23306 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n21447), .A(n21289), .ZN(
        n21291) );
  OAI222_X1 U23307 ( .A1(n21443), .A2(n21292), .B1(n21424), .B2(n21291), .C1(
        n21450), .C2(n21290), .ZN(P3_U2723) );
  NAND2_X1 U23308 ( .A1(n21447), .A2(n21296), .ZN(n21299) );
  AOI22_X1 U23309 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21454), .B1(n21453), .B2(
        n21293), .ZN(n21294) );
  OAI221_X1 U23310 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n21296), .C1(n21295), 
        .C2(n21299), .A(n21294), .ZN(P3_U2724) );
  NOR2_X1 U23311 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n21305), .ZN(n21298) );
  OAI222_X1 U23312 ( .A1(n21443), .A2(n21300), .B1(n21299), .B2(n21298), .C1(
        n21450), .C2(n21297), .ZN(P3_U2725) );
  INV_X1 U23313 ( .A(n21301), .ZN(n21302) );
  AOI21_X1 U23314 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n21447), .A(n21302), .ZN(
        n21304) );
  OAI222_X1 U23315 ( .A1(n21443), .A2(n21306), .B1(n21305), .B2(n21304), .C1(
        n21450), .C2(n21303), .ZN(P3_U2726) );
  NOR2_X1 U23316 ( .A1(n21307), .A2(n21458), .ZN(n21333) );
  NAND2_X1 U23317 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n21333), .ZN(n21321) );
  NOR2_X1 U23318 ( .A1(n21308), .A2(n21321), .ZN(n21324) );
  NAND2_X1 U23319 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n21324), .ZN(n21312) );
  NOR2_X1 U23320 ( .A1(n21309), .A2(n21312), .ZN(n21315) );
  AOI21_X1 U23321 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n21447), .A(n21315), .ZN(
        n21310) );
  OAI222_X1 U23322 ( .A1(n21311), .A2(n21443), .B1(n21435), .B2(n21310), .C1(
        n21450), .C2(n21751), .ZN(P3_U2728) );
  INV_X1 U23323 ( .A(n21312), .ZN(n21319) );
  AOI21_X1 U23324 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n21447), .A(n21319), .ZN(
        n21314) );
  OAI222_X1 U23325 ( .A1(n21316), .A2(n21443), .B1(n21315), .B2(n21314), .C1(
        n21450), .C2(n21313), .ZN(P3_U2729) );
  AOI21_X1 U23326 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n21447), .A(n21324), .ZN(
        n21318) );
  OAI222_X1 U23327 ( .A1(n21320), .A2(n21443), .B1(n21319), .B2(n21318), .C1(
        n21450), .C2(n21317), .ZN(P3_U2730) );
  INV_X1 U23328 ( .A(n21321), .ZN(n21328) );
  AOI21_X1 U23329 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n21447), .A(n21328), .ZN(
        n21323) );
  OAI222_X1 U23330 ( .A1(n21325), .A2(n21443), .B1(n21324), .B2(n21323), .C1(
        n21450), .C2(n21322), .ZN(P3_U2731) );
  AOI21_X1 U23331 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n21447), .A(n21333), .ZN(
        n21327) );
  OAI222_X1 U23332 ( .A1(n21329), .A2(n21443), .B1(n21328), .B2(n21327), .C1(
        n21450), .C2(n21326), .ZN(P3_U2732) );
  NAND2_X1 U23333 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n21456), .ZN(n21445) );
  NOR2_X1 U23334 ( .A1(n21446), .A2(n21445), .ZN(n21444) );
  OAI21_X1 U23335 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n21444), .A(n21447), .ZN(
        n21332) );
  AOI22_X1 U23336 ( .A1(n21454), .A2(BUF2_REG_2__SCAN_IN), .B1(n21453), .B2(
        n21330), .ZN(n21331) );
  OAI21_X1 U23337 ( .B1(n21333), .B2(n21332), .A(n21331), .ZN(P3_U2733) );
  NAND2_X1 U23338 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n21370) );
  NOR3_X1 U23339 ( .A1(n21371), .A2(n21420), .A3(n21370), .ZN(n21358) );
  NAND2_X1 U23340 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n21358), .ZN(n21353) );
  INV_X1 U23341 ( .A(n21353), .ZN(n21341) );
  NAND2_X1 U23342 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n21341), .ZN(n21345) );
  NAND2_X1 U23343 ( .A1(n21447), .A2(n21345), .ZN(n21348) );
  NAND2_X1 U23344 ( .A1(n21336), .A2(n21389), .ZN(n21402) );
  OAI22_X1 U23345 ( .A1(n21338), .A2(n21450), .B1(n21337), .B2(n21402), .ZN(
        n21339) );
  AOI21_X1 U23346 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n21418), .A(n21339), .ZN(
        n21340) );
  OAI221_X1 U23347 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21345), .C1(n21346), 
        .C2(n21348), .A(n21340), .ZN(P3_U2714) );
  AOI22_X1 U23348 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n21418), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n21419), .ZN(n21343) );
  OAI211_X1 U23349 ( .C1(n21341), .C2(P3_EAX_REG_20__SCAN_IN), .A(n21447), .B(
        n21345), .ZN(n21342) );
  OAI211_X1 U23350 ( .C1(n21344), .C2(n21450), .A(n21343), .B(n21342), .ZN(
        P3_U2715) );
  OR2_X1 U23351 ( .A1(n21346), .A2(n21345), .ZN(n21352) );
  AOI22_X1 U23352 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n21419), .B1(n21453), .B2(
        n21347), .ZN(n21351) );
  OAI21_X1 U23353 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21458), .A(n21348), .ZN(
        n21349) );
  AOI22_X1 U23354 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n21418), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n21349), .ZN(n21350) );
  OAI211_X1 U23355 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n21352), .A(n21351), .B(
        n21350), .ZN(P3_U2713) );
  AOI22_X1 U23356 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n21418), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n21419), .ZN(n21355) );
  OAI211_X1 U23357 ( .C1(n21358), .C2(P3_EAX_REG_19__SCAN_IN), .A(n21447), .B(
        n21353), .ZN(n21354) );
  OAI211_X1 U23358 ( .C1(n21356), .C2(n21450), .A(n21355), .B(n21354), .ZN(
        P3_U2716) );
  AOI22_X1 U23359 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n21418), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n21419), .ZN(n21362) );
  OR2_X1 U23360 ( .A1(n21357), .A2(n21420), .ZN(n21364) );
  AOI211_X1 U23361 ( .C1(n21359), .C2(n21364), .A(n21358), .B(n21389), .ZN(
        n21360) );
  INV_X1 U23362 ( .A(n21360), .ZN(n21361) );
  OAI211_X1 U23363 ( .C1(n21363), .C2(n21450), .A(n21362), .B(n21361), .ZN(
        P3_U2717) );
  AOI22_X1 U23364 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21418), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n21419), .ZN(n21367) );
  INV_X1 U23365 ( .A(n21420), .ZN(n21365) );
  OAI211_X1 U23366 ( .C1(n21365), .C2(P3_EAX_REG_17__SCAN_IN), .A(n21447), .B(
        n21364), .ZN(n21366) );
  OAI211_X1 U23367 ( .C1(n21368), .C2(n21450), .A(n21367), .B(n21366), .ZN(
        P3_U2718) );
  AOI22_X1 U23368 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n21418), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n21419), .ZN(n21374) );
  NAND4_X1 U23369 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(P3_EAX_REG_20__SCAN_IN), .ZN(n21369)
         );
  NAND2_X1 U23370 ( .A1(n21414), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n21413) );
  NOR2_X1 U23371 ( .A1(n21371), .A2(n21413), .ZN(n21409) );
  NAND2_X1 U23372 ( .A1(n21409), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n21408) );
  OAI211_X1 U23373 ( .C1(n21372), .C2(P3_EAX_REG_25__SCAN_IN), .A(n21447), .B(
        n21376), .ZN(n21373) );
  OAI211_X1 U23374 ( .C1(n21375), .C2(n21450), .A(n21374), .B(n21373), .ZN(
        P3_U2710) );
  AOI22_X1 U23375 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21418), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n21419), .ZN(n21380) );
  AOI211_X1 U23376 ( .C1(n21377), .C2(n21376), .A(n21404), .B(n21389), .ZN(
        n21378) );
  INV_X1 U23377 ( .A(n21378), .ZN(n21379) );
  OAI211_X1 U23378 ( .C1(n21381), .C2(n21450), .A(n21380), .B(n21379), .ZN(
        P3_U2709) );
  NAND2_X1 U23379 ( .A1(n21390), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n21382) );
  INV_X1 U23380 ( .A(n21383), .ZN(n21384) );
  AOI22_X1 U23381 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n21419), .B1(n21453), .B2(
        n21384), .ZN(n21386) );
  AOI22_X1 U23382 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21418), .B1(n21390), .B2(
        n21387), .ZN(n21385) );
  OAI211_X1 U23383 ( .C1(n21388), .C2(n21387), .A(n21386), .B(n21385), .ZN(
        P3_U2705) );
  AOI22_X1 U23384 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21418), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n21419), .ZN(n21394) );
  AOI211_X1 U23385 ( .C1(n21391), .C2(n21397), .A(n21390), .B(n21389), .ZN(
        n21392) );
  INV_X1 U23386 ( .A(n21392), .ZN(n21393) );
  OAI211_X1 U23387 ( .C1(n21450), .C2(n21395), .A(n21394), .B(n21393), .ZN(
        P3_U2706) );
  AOI22_X1 U23388 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n21418), .B1(n21453), .B2(
        n21396), .ZN(n21400) );
  OAI211_X1 U23389 ( .C1(n21398), .C2(P3_EAX_REG_28__SCAN_IN), .A(n21447), .B(
        n21397), .ZN(n21399) );
  OAI211_X1 U23390 ( .C1(n21402), .C2(n21401), .A(n21400), .B(n21399), .ZN(
        P3_U2707) );
  AOI22_X1 U23391 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21418), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n21419), .ZN(n21406) );
  OAI211_X1 U23392 ( .C1(n21404), .C2(P3_EAX_REG_27__SCAN_IN), .A(n21447), .B(
        n21403), .ZN(n21405) );
  OAI211_X1 U23393 ( .C1(n21407), .C2(n21450), .A(n21406), .B(n21405), .ZN(
        P3_U2708) );
  AOI22_X1 U23394 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n21419), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n21418), .ZN(n21411) );
  OAI211_X1 U23395 ( .C1(n21409), .C2(P3_EAX_REG_24__SCAN_IN), .A(n21447), .B(
        n21408), .ZN(n21410) );
  OAI211_X1 U23396 ( .C1(n21412), .C2(n21450), .A(n21411), .B(n21410), .ZN(
        P3_U2711) );
  AOI22_X1 U23397 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n21418), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n21419), .ZN(n21416) );
  OAI211_X1 U23398 ( .C1(n21414), .C2(P3_EAX_REG_23__SCAN_IN), .A(n21447), .B(
        n21413), .ZN(n21415) );
  OAI211_X1 U23399 ( .C1(n21417), .C2(n21450), .A(n21416), .B(n21415), .ZN(
        P3_U2712) );
  AOI22_X1 U23400 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n21419), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n21418), .ZN(n21422) );
  OAI211_X1 U23401 ( .C1(n21429), .C2(P3_EAX_REG_16__SCAN_IN), .A(n21447), .B(
        n21420), .ZN(n21421) );
  OAI211_X1 U23402 ( .C1(n21423), .C2(n21450), .A(n21422), .B(n21421), .ZN(
        P3_U2719) );
  NAND2_X1 U23403 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n21424), .ZN(n21428) );
  AOI22_X1 U23404 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21454), .B1(n21453), .B2(
        n21425), .ZN(n21427) );
  NAND3_X1 U23405 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n21447), .A3(n21431), 
        .ZN(n21426) );
  OAI211_X1 U23406 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n21428), .A(n21427), .B(
        n21426), .ZN(P3_U2721) );
  AOI21_X1 U23407 ( .B1(n21431), .B2(n21430), .A(n21429), .ZN(n21432) );
  AOI22_X1 U23408 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n21454), .B1(n21432), .B2(
        n21447), .ZN(n21433) );
  OAI21_X1 U23409 ( .B1(n21434), .B2(n21450), .A(n21433), .ZN(P3_U2720) );
  NOR2_X1 U23410 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21435), .ZN(n21441) );
  AOI21_X1 U23411 ( .B1(n21438), .B2(n21437), .A(n21436), .ZN(n21440) );
  OAI222_X1 U23412 ( .A1(n21443), .A2(n21442), .B1(n21441), .B2(n21440), .C1(
        n21450), .C2(n21439), .ZN(P3_U2727) );
  AOI21_X1 U23413 ( .B1(n21446), .B2(n21445), .A(n21444), .ZN(n21448) );
  AOI22_X1 U23414 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21454), .B1(n21448), .B2(
        n21447), .ZN(n21449) );
  OAI21_X1 U23415 ( .B1(n21451), .B2(n21450), .A(n21449), .ZN(P3_U2734) );
  AOI22_X1 U23416 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n21454), .B1(n21453), .B2(
        n11152), .ZN(n21455) );
  OAI221_X1 U23417 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n21458), .C1(n21457), 
        .C2(n21456), .A(n21455), .ZN(P3_U2735) );
  INV_X1 U23418 ( .A(n21508), .ZN(n21468) );
  OR2_X1 U23419 ( .A1(n21528), .A2(n21459), .ZN(n21464) );
  AOI22_X1 U23420 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21865), .B1(
        n21464), .B2(n21460), .ZN(n21905) );
  OAI222_X1 U23421 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21481), .B1(
        n21905), .B2(n21507), .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(
        n21505), .ZN(n21461) );
  OAI22_X1 U23422 ( .A1(n21468), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n21461), .B2(n21508), .ZN(n21462) );
  INV_X1 U23423 ( .A(n21462), .ZN(P3_U3290) );
  INV_X1 U23424 ( .A(n21479), .ZN(n21463) );
  AOI22_X1 U23425 ( .A1(n21466), .A2(n21464), .B1(n21492), .B2(n21463), .ZN(
        n21906) );
  INV_X1 U23426 ( .A(n21906), .ZN(n21467) );
  INV_X1 U23427 ( .A(n21507), .ZN(n21484) );
  AOI22_X1 U23428 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12574), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21543), .ZN(n21480) );
  NOR2_X1 U23429 ( .A1(n21481), .A2(n21615), .ZN(n21465) );
  AOI222_X1 U23430 ( .A1(n21467), .A2(n21484), .B1(n21466), .B2(n21938), .C1(
        n21480), .C2(n21465), .ZN(n21469) );
  AOI22_X1 U23431 ( .A1(n21508), .A2(n21492), .B1(n21469), .B2(n21468), .ZN(
        P3_U3289) );
  NAND2_X1 U23432 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21491), .ZN(
        n21478) );
  INV_X1 U23433 ( .A(n21826), .ZN(n21899) );
  AOI22_X1 U23434 ( .A1(n21473), .A2(n21472), .B1(n21471), .B2(n21470), .ZN(
        n21490) );
  OAI21_X1 U23435 ( .B1(n21503), .B2(n21492), .A(n21495), .ZN(n21474) );
  AOI21_X1 U23436 ( .B1(n21490), .B2(n21474), .A(n21491), .ZN(n21475) );
  AOI22_X1 U23437 ( .A1(n21899), .A2(n21476), .B1(n21475), .B2(n21485), .ZN(
        n21477) );
  OAI21_X1 U23438 ( .B1(n21479), .B2(n21478), .A(n21477), .ZN(n21909) );
  NOR3_X1 U23439 ( .A1(n21481), .A2(n21615), .A3(n21480), .ZN(n21483) );
  NOR3_X1 U23440 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21485), .A3(
        n21505), .ZN(n21482) );
  AOI211_X1 U23441 ( .C1(n21484), .C2(n21909), .A(n21483), .B(n21482), .ZN(
        n21487) );
  AOI21_X1 U23442 ( .B1(n21938), .B2(n21485), .A(n21508), .ZN(n21486) );
  OAI22_X1 U23443 ( .A1(n21508), .A2(n21487), .B1(n21486), .B2(n21491), .ZN(
        P3_U3288) );
  NOR2_X1 U23444 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20877), .ZN(
        n21504) );
  AOI221_X1 U23445 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n21489), 
        .C1(n20877), .C2(n21488), .A(n21826), .ZN(n21502) );
  INV_X1 U23446 ( .A(n21490), .ZN(n21496) );
  NOR2_X1 U23447 ( .A1(n21492), .A2(n21491), .ZN(n21493) );
  OAI22_X1 U23448 ( .A1(n21493), .A2(n20877), .B1(n21500), .B2(n11547), .ZN(
        n21494) );
  AOI22_X1 U23449 ( .A1(n21497), .A2(n21496), .B1(n21495), .B2(n21494), .ZN(
        n21498) );
  OAI221_X1 U23450 ( .B1(n21500), .B2(n21499), .C1(n21500), .C2(n21460), .A(
        n21498), .ZN(n21501) );
  AOI211_X1 U23451 ( .C1(n21504), .C2(n21503), .A(n21502), .B(n21501), .ZN(
        n21913) );
  OAI22_X1 U23452 ( .A1(n21913), .A2(n21507), .B1(n21506), .B2(n21505), .ZN(
        n21509) );
  MUX2_X1 U23453 ( .A(n21509), .B(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n21508), .Z(P3_U3285) );
  NOR2_X1 U23454 ( .A1(n21829), .A2(n21510), .ZN(n21512) );
  OAI22_X1 U23455 ( .A1(n21511), .A2(n21792), .B1(n21794), .B2(n21616), .ZN(
        n21613) );
  AOI21_X1 U23456 ( .B1(n21512), .B2(n21613), .A(n21687), .ZN(n21677) );
  NOR2_X1 U23457 ( .A1(n21677), .A2(n21821), .ZN(n21806) );
  AOI21_X1 U23458 ( .B1(n21514), .B2(n21806), .A(n21513), .ZN(n21526) );
  INV_X1 U23459 ( .A(n21515), .ZN(n21521) );
  INV_X1 U23460 ( .A(n21516), .ZN(n21518) );
  OAI21_X1 U23461 ( .B1(n21522), .B2(n21800), .A(n21865), .ZN(n21517) );
  OAI21_X1 U23462 ( .B1(n21518), .B2(n21826), .A(n21517), .ZN(n21797) );
  NOR2_X1 U23463 ( .A1(n21899), .A2(n21865), .ZN(n21866) );
  OAI22_X1 U23464 ( .A1(n21523), .A2(n21866), .B1(n21519), .B2(n21792), .ZN(
        n21520) );
  AOI211_X1 U23465 ( .C1(n21819), .C2(n21521), .A(n21797), .B(n21520), .ZN(
        n21679) );
  AOI221_X1 U23466 ( .B1(n21522), .B2(n21528), .C1(n21615), .C2(n21528), .A(
        n21821), .ZN(n21799) );
  OAI211_X1 U23467 ( .C1(n21523), .C2(n21875), .A(n21679), .B(n21799), .ZN(
        n21524) );
  NAND3_X1 U23468 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21868), .A3(
        n21524), .ZN(n21525) );
  OAI211_X1 U23469 ( .C1(n21527), .C2(n21849), .A(n21526), .B(n21525), .ZN(
        P3_U2841) );
  NOR2_X1 U23470 ( .A1(n21821), .A2(n21792), .ZN(n21708) );
  INV_X1 U23471 ( .A(n21559), .ZN(n21593) );
  NOR2_X1 U23472 ( .A1(n21899), .A2(n21528), .ZN(n21809) );
  AOI221_X1 U23473 ( .B1(n21876), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n21809), .C2(n21615), .A(n21821), .ZN(n21529) );
  AOI221_X1 U23474 ( .B1(n21708), .B2(n21531), .C1(n21593), .C2(n21530), .A(
        n21529), .ZN(n21533) );
  NAND2_X1 U23475 ( .A1(n21886), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n21532) );
  OAI211_X1 U23476 ( .C1(n21773), .C2(n21615), .A(n21533), .B(n21532), .ZN(
        P3_U2862) );
  NOR2_X1 U23477 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21809), .ZN(
        n21536) );
  NOR2_X1 U23478 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21843), .ZN(
        n21534) );
  AOI22_X1 U23479 ( .A1(n21536), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n21535), .B2(n21534), .ZN(n21541) );
  AOI22_X1 U23480 ( .A1(n21886), .A2(P3_REIP_REG_1__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21881), .ZN(n21540) );
  AOI22_X1 U23481 ( .A1(n21593), .A2(n21538), .B1(n21708), .B2(n21537), .ZN(
        n21539) );
  OAI211_X1 U23482 ( .C1(n21821), .C2(n21541), .A(n21540), .B(n21539), .ZN(
        P3_U2861) );
  NAND2_X1 U23483 ( .A1(n21886), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n21549) );
  NOR3_X1 U23484 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21543), .A3(
        n21554), .ZN(n21547) );
  NOR3_X1 U23485 ( .A1(n21826), .A2(n21543), .A3(n21615), .ZN(n21542) );
  NOR2_X1 U23486 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21875), .ZN(
        n21822) );
  AOI211_X1 U23487 ( .C1(n21828), .C2(n21543), .A(n21542), .B(n21822), .ZN(
        n21545) );
  NAND2_X1 U23488 ( .A1(n21899), .A2(n21555), .ZN(n21551) );
  OAI211_X1 U23489 ( .C1(n21545), .C2(n12536), .A(n21544), .B(n21551), .ZN(
        n21546) );
  OAI21_X1 U23490 ( .B1(n21547), .B2(n21546), .A(n21856), .ZN(n21548) );
  OAI211_X1 U23491 ( .C1(n21773), .C2(n12536), .A(n21549), .B(n21548), .ZN(
        P3_U2860) );
  INV_X1 U23492 ( .A(n21822), .ZN(n21550) );
  OAI211_X1 U23493 ( .C1(n11246), .C2(n21552), .A(n21551), .B(n21550), .ZN(
        n21571) );
  OAI21_X1 U23494 ( .B1(n21564), .B2(n21571), .A(n21856), .ZN(n21563) );
  OAI22_X1 U23495 ( .A1(n21555), .A2(n21826), .B1(n21554), .B2(n21553), .ZN(
        n21599) );
  INV_X1 U23496 ( .A(n21599), .ZN(n21612) );
  INV_X1 U23497 ( .A(n21556), .ZN(n21558) );
  INV_X1 U23498 ( .A(n21708), .ZN(n21588) );
  OAI22_X1 U23499 ( .A1(n21559), .A2(n21558), .B1(n21588), .B2(n21557), .ZN(
        n21560) );
  AOI211_X1 U23500 ( .C1(n21881), .C2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n21561), .B(n21560), .ZN(n21562) );
  OAI221_X1 U23501 ( .B1(n21563), .B2(n21612), .C1(n21563), .C2(n21564), .A(
        n21562), .ZN(P3_U2859) );
  NOR3_X1 U23502 ( .A1(n21843), .A2(n11585), .A3(n21563), .ZN(n21566) );
  NAND2_X1 U23503 ( .A1(n21856), .A2(n21599), .ZN(n21579) );
  NOR3_X1 U23504 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21564), .A3(
        n21579), .ZN(n21565) );
  AOI211_X1 U23505 ( .C1(n21856), .C2(n21567), .A(n21566), .B(n21565), .ZN(
        n21569) );
  NAND2_X1 U23506 ( .A1(n21886), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n21568) );
  OAI211_X1 U23507 ( .C1(n21773), .C2(n11585), .A(n21569), .B(n21568), .ZN(
        P3_U2858) );
  NAND2_X1 U23508 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21570) );
  NOR2_X1 U23509 ( .A1(n21570), .A2(n21579), .ZN(n21572) );
  AOI21_X1 U23510 ( .B1(n21788), .B2(n21580), .A(n21571), .ZN(n21586) );
  AOI21_X1 U23511 ( .B1(n21856), .B2(n21586), .A(n21801), .ZN(n21578) );
  MUX2_X1 U23512 ( .A(n21572), .B(n21578), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n21573) );
  AOI21_X1 U23513 ( .B1(n21593), .B2(n21574), .A(n21573), .ZN(n21576) );
  OAI211_X1 U23514 ( .C1(n21588), .C2(n21577), .A(n21576), .B(n21575), .ZN(
        P3_U2857) );
  AOI22_X1 U23515 ( .A1(n21886), .A2(P3_REIP_REG_6__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n21578), .ZN(n21584) );
  NOR3_X1 U23516 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21580), .A3(
        n21579), .ZN(n21581) );
  AOI21_X1 U23517 ( .B1(n21582), .B2(n21593), .A(n21581), .ZN(n21583) );
  OAI211_X1 U23518 ( .C1(n21588), .C2(n21585), .A(n21584), .B(n21583), .ZN(
        P3_U2856) );
  NAND2_X1 U23519 ( .A1(n21601), .A2(n21599), .ZN(n21597) );
  OAI211_X1 U23520 ( .C1(n21843), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n21586), .ZN(n21598) );
  NAND2_X1 U23521 ( .A1(n21856), .A2(n21598), .ZN(n21596) );
  AOI21_X1 U23522 ( .B1(n21856), .B2(n21598), .A(n21881), .ZN(n21590) );
  OAI22_X1 U23523 ( .A1(n21590), .A2(n21589), .B1(n21588), .B2(n21587), .ZN(
        n21591) );
  AOI21_X1 U23524 ( .B1(n21593), .B2(n21592), .A(n21591), .ZN(n21595) );
  NAND2_X1 U23525 ( .A1(n21886), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n21594) );
  OAI211_X1 U23526 ( .C1(n21597), .C2(n21596), .A(n21595), .B(n21594), .ZN(
        P3_U2855) );
  NAND3_X1 U23527 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21788), .A3(
        n21598), .ZN(n21603) );
  NAND4_X1 U23528 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21601), .A3(
        n21600), .A4(n21599), .ZN(n21602) );
  OAI211_X1 U23529 ( .C1(n21604), .C2(n21792), .A(n21603), .B(n21602), .ZN(
        n21605) );
  AOI21_X1 U23530 ( .B1(n21819), .B2(n21606), .A(n21605), .ZN(n21610) );
  AOI22_X1 U23531 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21881), .B1(
        n21885), .B2(n21607), .ZN(n21609) );
  OAI211_X1 U23532 ( .C1(n21610), .C2(n21821), .A(n21609), .B(n21608), .ZN(
        P3_U2854) );
  NOR3_X1 U23533 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21622), .A3(
        n21890), .ZN(n21614) );
  AOI21_X1 U23534 ( .B1(P3_REIP_REG_11__SCAN_IN), .B2(n21886), .A(n21614), 
        .ZN(n21626) );
  NOR2_X1 U23535 ( .A1(n21819), .A2(n21898), .ZN(n21620) );
  NOR2_X1 U23536 ( .A1(n21615), .A2(n21864), .ZN(n21874) );
  AOI21_X1 U23537 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21874), .A(
        n21875), .ZN(n21618) );
  NOR2_X1 U23538 ( .A1(n21663), .A2(n21826), .ZN(n21880) );
  NAND2_X1 U23539 ( .A1(n21819), .A2(n21616), .ZN(n21815) );
  OAI21_X1 U23540 ( .B1(n21617), .B2(n21792), .A(n21815), .ZN(n21883) );
  NOR4_X1 U23541 ( .A1(n21618), .A2(n21880), .A3(n21821), .A4(n21883), .ZN(
        n21619) );
  OAI21_X1 U23542 ( .B1(n21621), .B2(n21620), .A(n21619), .ZN(n21869) );
  NAND2_X1 U23543 ( .A1(n21899), .A2(n21635), .ZN(n21623) );
  OAI21_X1 U23544 ( .B1(n21622), .B2(n21864), .A(n21865), .ZN(n21631) );
  OAI211_X1 U23545 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n21875), .A(
        n21623), .B(n21631), .ZN(n21624) );
  OAI211_X1 U23546 ( .C1(n21869), .C2(n21624), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n21868), .ZN(n21625) );
  OAI211_X1 U23547 ( .C1(n21627), .C2(n21849), .A(n21626), .B(n21625), .ZN(
        P3_U2851) );
  AOI22_X1 U23548 ( .A1(n21886), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n21885), 
        .B2(n21628), .ZN(n21639) );
  AOI21_X1 U23549 ( .B1(n21629), .B2(n21874), .A(n21875), .ZN(n21640) );
  AOI21_X1 U23550 ( .B1(n21630), .B2(n21663), .A(n21826), .ZN(n21643) );
  OAI21_X1 U23551 ( .B1(n21632), .B2(n21792), .A(n21631), .ZN(n21633) );
  AOI211_X1 U23552 ( .C1(n21819), .C2(n21634), .A(n21643), .B(n21633), .ZN(
        n21857) );
  OAI211_X1 U23553 ( .C1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n21876), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n21857), .ZN(n21637) );
  OAI22_X1 U23554 ( .A1(n21821), .A2(n21853), .B1(n21635), .B2(n21890), .ZN(
        n21636) );
  OAI21_X1 U23555 ( .B1(n21640), .B2(n21637), .A(n21636), .ZN(n21638) );
  OAI211_X1 U23556 ( .C1(n21773), .C2(n21853), .A(n21639), .B(n21638), .ZN(
        P3_U2850) );
  AOI22_X1 U23557 ( .A1(n21886), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21881), .ZN(n21653) );
  AOI21_X1 U23558 ( .B1(n21899), .B2(n21853), .A(n21640), .ZN(n21855) );
  INV_X1 U23559 ( .A(n21809), .ZN(n21644) );
  INV_X1 U23560 ( .A(n21864), .ZN(n21641) );
  AOI21_X1 U23561 ( .B1(n21642), .B2(n21641), .A(n21876), .ZN(n21659) );
  AOI211_X1 U23562 ( .C1(n12552), .C2(n21644), .A(n21659), .B(n21643), .ZN(
        n21649) );
  NOR2_X1 U23563 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21645), .ZN(
        n21646) );
  AOI22_X1 U23564 ( .A1(n21819), .A2(n21647), .B1(n21665), .B2(n21646), .ZN(
        n21648) );
  OAI221_X1 U23565 ( .B1(n21661), .B2(n21855), .C1(n21661), .C2(n21649), .A(
        n21648), .ZN(n21651) );
  AOI22_X1 U23566 ( .A1(n21856), .A2(n21651), .B1(n21708), .B2(n21650), .ZN(
        n21652) );
  OAI211_X1 U23567 ( .C1(n21654), .C2(n21849), .A(n21653), .B(n21652), .ZN(
        P3_U2848) );
  NOR2_X1 U23568 ( .A1(n21655), .A2(n21794), .ZN(n21669) );
  NOR2_X1 U23569 ( .A1(n21667), .A2(n21792), .ZN(n21656) );
  AOI22_X1 U23570 ( .A1(n21658), .A2(n21669), .B1(n21657), .B2(n21656), .ZN(
        n21676) );
  AOI22_X1 U23571 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21820), .B1(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n21875), .ZN(n21660) );
  AOI211_X1 U23572 ( .C1(n21661), .C2(n21865), .A(n21660), .B(n21659), .ZN(
        n21662) );
  OAI221_X1 U23573 ( .B1(n21826), .B2(n21664), .C1(n21826), .C2(n21663), .A(
        n21662), .ZN(n21666) );
  NAND3_X1 U23574 ( .A1(n21665), .A2(n21664), .A3(n21666), .ZN(n21675) );
  INV_X1 U23575 ( .A(n21666), .ZN(n21841) );
  OAI21_X1 U23576 ( .B1(n21667), .B2(n21792), .A(n21856), .ZN(n21668) );
  NOR2_X1 U23577 ( .A1(n21669), .A2(n21668), .ZN(n21842) );
  INV_X1 U23578 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21670) );
  AOI211_X1 U23579 ( .C1(n21841), .C2(n21842), .A(n21801), .B(n21670), .ZN(
        n21672) );
  AOI211_X1 U23580 ( .C1(n21885), .C2(n21673), .A(n21672), .B(n21671), .ZN(
        n21674) );
  OAI221_X1 U23581 ( .B1(n21821), .B2(n21676), .C1(n21821), .C2(n21675), .A(
        n21674), .ZN(P3_U2847) );
  NAND2_X1 U23582 ( .A1(n21801), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n21685) );
  INV_X1 U23583 ( .A(n21677), .ZN(n21678) );
  NAND2_X1 U23584 ( .A1(n21678), .A2(n21688), .ZN(n21784) );
  INV_X1 U23585 ( .A(n21784), .ZN(n21723) );
  OAI211_X1 U23586 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n21866), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n21679), .ZN(n21680) );
  OAI21_X1 U23587 ( .B1(n21681), .B2(n21680), .A(n21856), .ZN(n21682) );
  OAI21_X1 U23588 ( .B1(n21773), .B2(n21770), .A(n21682), .ZN(n21683) );
  OAI21_X1 U23589 ( .B1(n21723), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n21683), .ZN(n21684) );
  OAI211_X1 U23590 ( .C1(n21686), .C2(n21849), .A(n21685), .B(n21684), .ZN(
        P3_U2840) );
  NAND2_X1 U23591 ( .A1(n21688), .A2(n21687), .ZN(n21689) );
  NOR4_X1 U23592 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21690), .A3(
        n21783), .A4(n21689), .ZN(n21697) );
  NAND2_X1 U23593 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21693) );
  NOR2_X1 U23594 ( .A1(n21691), .A2(n21826), .ZN(n21777) );
  INV_X1 U23595 ( .A(n21775), .ZN(n21692) );
  AOI211_X1 U23596 ( .C1(n21788), .C2(n21693), .A(n21777), .B(n21692), .ZN(
        n21704) );
  OAI22_X1 U23597 ( .A1(n21704), .A2(n21695), .B1(n21792), .B2(n21694), .ZN(
        n21696) );
  AOI211_X1 U23598 ( .C1(n21698), .C2(n21819), .A(n21697), .B(n21696), .ZN(
        n21702) );
  AOI22_X1 U23599 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21881), .B1(
        n21885), .B2(n21699), .ZN(n21701) );
  NAND2_X1 U23600 ( .A1(n21886), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21700) );
  OAI211_X1 U23601 ( .C1(n21702), .C2(n21821), .A(n21701), .B(n21700), .ZN(
        P3_U2837) );
  NAND2_X1 U23602 ( .A1(n21819), .A2(n21719), .ZN(n21703) );
  OAI211_X1 U23603 ( .C1(n21843), .C2(n21705), .A(n21704), .B(n21703), .ZN(
        n21706) );
  AOI22_X1 U23604 ( .A1(n21856), .A2(n21706), .B1(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n21881), .ZN(n21712) );
  NAND2_X1 U23605 ( .A1(n21708), .A2(n21707), .ZN(n21724) );
  NAND4_X1 U23606 ( .A1(n21723), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A4(n21709), .ZN(n21710) );
  AOI22_X1 U23607 ( .A1(n21712), .A2(n21724), .B1(n21711), .B2(n21710), .ZN(
        n21713) );
  AOI21_X1 U23608 ( .B1(n21714), .B2(n21885), .A(n21713), .ZN(n21715) );
  OAI21_X1 U23609 ( .B1(n21868), .B2(n21716), .A(n21715), .ZN(P3_U2836) );
  NOR2_X1 U23610 ( .A1(n21717), .A2(n21759), .ZN(n21732) );
  AOI22_X1 U23611 ( .A1(n21819), .A2(n21719), .B1(n21828), .B2(n21718), .ZN(
        n21720) );
  NAND3_X1 U23612 ( .A1(n21775), .A2(n21732), .A3(n21720), .ZN(n21721) );
  AOI22_X1 U23613 ( .A1(n21856), .A2(n21721), .B1(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21881), .ZN(n21725) );
  NAND2_X1 U23614 ( .A1(n21723), .A2(n21722), .ZN(n21760) );
  AOI22_X1 U23615 ( .A1(n21725), .A2(n21724), .B1(n21760), .B2(n21759), .ZN(
        n21726) );
  AOI21_X1 U23616 ( .B1(n21885), .B2(n21727), .A(n21726), .ZN(n21729) );
  NAND2_X1 U23617 ( .A1(n21729), .A2(n21728), .ZN(P3_U2835) );
  OAI22_X1 U23618 ( .A1(n21876), .A2(n21733), .B1(n21732), .B2(n21826), .ZN(
        n21734) );
  AOI221_X1 U23619 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21736), 
        .C1(n21809), .C2(n21736), .A(n12570), .ZN(n21740) );
  AND2_X1 U23620 ( .A1(n21898), .A2(n21753), .ZN(n21737) );
  AOI211_X1 U23621 ( .C1(n21754), .C2(n21819), .A(n21738), .B(n21737), .ZN(
        n21744) );
  NOR3_X1 U23622 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21744), .A3(
        n21821), .ZN(n21739) );
  OAI21_X1 U23623 ( .B1(n21742), .B2(n21849), .A(n21741), .ZN(P3_U2833) );
  AOI22_X1 U23624 ( .A1(n21886), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n21885), 
        .B2(n21743), .ZN(n21749) );
  OAI21_X1 U23625 ( .B1(n21744), .B2(n12570), .A(n12569), .ZN(n21745) );
  OAI211_X1 U23626 ( .C1(n21747), .C2(n21746), .A(n21856), .B(n21745), .ZN(
        n21748) );
  OAI211_X1 U23627 ( .C1(n12569), .C2(n21773), .A(n21749), .B(n21748), .ZN(
        P3_U2832) );
  NAND2_X1 U23628 ( .A1(n21895), .A2(n21750), .ZN(n21761) );
  OAI21_X1 U23629 ( .B1(n21751), .B2(n21761), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21757) );
  OAI211_X1 U23630 ( .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n21866), .A(
        n21752), .B(n21773), .ZN(n21756) );
  OAI22_X1 U23631 ( .A1(n21754), .A2(n21794), .B1(n21753), .B2(n21792), .ZN(
        n21755) );
  AOI211_X1 U23632 ( .C1(n21758), .C2(n21757), .A(n21756), .B(n21755), .ZN(
        n21769) );
  OAI22_X1 U23633 ( .A1(n21762), .A2(n21761), .B1(n21760), .B2(n21759), .ZN(
        n21763) );
  OAI221_X1 U23634 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21856), 
        .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n21763), .A(n21868), .ZN(
        n21768) );
  OR3_X1 U23635 ( .A1(n21765), .A2(n21849), .A3(n21764), .ZN(n21766) );
  OAI211_X1 U23636 ( .C1(n21769), .C2(n21768), .A(n21767), .B(n21766), .ZN(
        P3_U2834) );
  NOR3_X1 U23637 ( .A1(n21881), .A2(n21770), .A3(n21784), .ZN(n21779) );
  AOI22_X1 U23638 ( .A1(n21819), .A2(n21772), .B1(n21898), .B2(n21771), .ZN(
        n21774) );
  NAND3_X1 U23639 ( .A1(n21775), .A2(n21774), .A3(n21773), .ZN(n21787) );
  NOR3_X1 U23640 ( .A1(n21777), .A2(n21776), .A3(n21787), .ZN(n21778) );
  NOR2_X1 U23641 ( .A1(n21778), .A2(n21886), .ZN(n21786) );
  OAI21_X1 U23642 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n21779), .A(
        n21786), .ZN(n21780) );
  OAI211_X1 U23643 ( .C1(n21782), .C2(n21849), .A(n21781), .B(n21780), .ZN(
        P3_U2839) );
  NOR4_X1 U23644 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21784), .A3(
        n21821), .A4(n21783), .ZN(n21785) );
  AOI21_X1 U23645 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n21886), .A(n21785), 
        .ZN(n21790) );
  OAI211_X1 U23646 ( .C1(n21788), .C2(n21787), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n21786), .ZN(n21789) );
  OAI211_X1 U23647 ( .C1(n21791), .C2(n21849), .A(n21790), .B(n21789), .ZN(
        P3_U2838) );
  OAI22_X1 U23648 ( .A1(n21795), .A2(n21794), .B1(n21793), .B2(n21792), .ZN(
        n21796) );
  NOR2_X1 U23649 ( .A1(n21797), .A2(n21796), .ZN(n21798) );
  AOI21_X1 U23650 ( .B1(n21799), .B2(n21798), .A(n21801), .ZN(n21811) );
  AOI22_X1 U23651 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21811), .B1(
        n21806), .B2(n21800), .ZN(n21803) );
  NAND2_X1 U23652 ( .A1(n21801), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n21802) );
  OAI211_X1 U23653 ( .C1(n21804), .C2(n21849), .A(n21803), .B(n21802), .ZN(
        P3_U2843) );
  AOI21_X1 U23654 ( .B1(n21807), .B2(n21806), .A(n21805), .ZN(n21813) );
  NOR3_X1 U23655 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21809), .A3(
        n21808), .ZN(n21810) );
  OAI21_X1 U23656 ( .B1(n21811), .B2(n21810), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21812) );
  OAI211_X1 U23657 ( .C1(n21814), .C2(n21849), .A(n21813), .B(n21812), .ZN(
        P3_U2842) );
  NAND2_X1 U23658 ( .A1(n21816), .A2(n21815), .ZN(n21818) );
  OAI22_X1 U23659 ( .A1(n21819), .A2(n21898), .B1(n21818), .B2(n21817), .ZN(
        n21825) );
  NAND2_X1 U23660 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21820), .ZN(
        n21823) );
  AOI211_X1 U23661 ( .C1(n21828), .C2(n21823), .A(n21822), .B(n21821), .ZN(
        n21824) );
  OAI211_X1 U23662 ( .C1(n21827), .C2(n21826), .A(n21825), .B(n21824), .ZN(
        n21836) );
  OAI221_X1 U23663 ( .B1(n21836), .B2(n21828), .C1(n21836), .C2(n21837), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21834) );
  NOR2_X1 U23664 ( .A1(n21829), .A2(n21890), .ZN(n21845) );
  AOI22_X1 U23665 ( .A1(n21885), .A2(n21831), .B1(n21845), .B2(n21830), .ZN(
        n21832) );
  OAI221_X1 U23666 ( .B1(n21886), .B2(n21834), .C1(n21868), .C2(n21833), .A(
        n21832), .ZN(P3_U2844) );
  AOI22_X1 U23667 ( .A1(n21886), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n21885), 
        .B2(n21835), .ZN(n21840) );
  NAND3_X1 U23668 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21868), .A3(
        n21836), .ZN(n21839) );
  NAND3_X1 U23669 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21845), .A3(
        n21837), .ZN(n21838) );
  NAND3_X1 U23670 ( .A1(n21840), .A2(n21839), .A3(n21838), .ZN(P3_U2845) );
  AOI221_X1 U23671 ( .B1(n21843), .B2(n21842), .C1(n21841), .C2(n21842), .A(
        n21886), .ZN(n21846) );
  AOI22_X1 U23672 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21846), .B1(
        n21845), .B2(n21844), .ZN(n21848) );
  OAI211_X1 U23673 ( .C1(n21850), .C2(n21849), .A(n21848), .B(n21847), .ZN(
        P3_U2846) );
  AOI22_X1 U23674 ( .A1(n21886), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21885), 
        .B2(n21851), .ZN(n21860) );
  OAI21_X1 U23675 ( .B1(n21853), .B2(n21852), .A(n21865), .ZN(n21854) );
  NAND4_X1 U23676 ( .A1(n21857), .A2(n21856), .A3(n21855), .A4(n21854), .ZN(
        n21858) );
  NAND3_X1 U23677 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21868), .A3(
        n21858), .ZN(n21859) );
  OAI211_X1 U23678 ( .C1(n21890), .C2(n21861), .A(n21860), .B(n21859), .ZN(
        P3_U2849) );
  NAND2_X1 U23679 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21862), .ZN(
        n21873) );
  AOI22_X1 U23680 ( .A1(n21886), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21885), 
        .B2(n21863), .ZN(n21872) );
  NAND2_X1 U23681 ( .A1(n21865), .A2(n21864), .ZN(n21867) );
  AOI21_X1 U23682 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21867), .A(
        n21866), .ZN(n21870) );
  OAI211_X1 U23683 ( .C1(n21870), .C2(n21869), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n21868), .ZN(n21871) );
  OAI211_X1 U23684 ( .C1(n21873), .C2(n21890), .A(n21872), .B(n21871), .ZN(
        P3_U2852) );
  AOI211_X1 U23685 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n21875), .A(
        n11246), .B(n21874), .ZN(n21879) );
  AOI21_X1 U23686 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21877), .A(
        n21876), .ZN(n21878) );
  OR4_X1 U23687 ( .A1(n21881), .A2(n21880), .A3(n21879), .A4(n21878), .ZN(
        n21882) );
  OAI21_X1 U23688 ( .B1(n21883), .B2(n21882), .A(n21868), .ZN(n21888) );
  AOI22_X1 U23689 ( .A1(n21886), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n21885), 
        .B2(n21884), .ZN(n21887) );
  OAI221_X1 U23690 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21890), .C1(
        n21889), .C2(n21888), .A(n21887), .ZN(P3_U2853) );
  NOR2_X1 U23691 ( .A1(n22332), .A2(n21891), .ZN(n21933) );
  NAND3_X1 U23692 ( .A1(n21894), .A2(n21893), .A3(n21892), .ZN(n21896) );
  AOI21_X1 U23693 ( .B1(n21897), .B2(n21896), .A(n21895), .ZN(n21902) );
  NOR2_X1 U23694 ( .A1(n21899), .A2(n21898), .ZN(n21900) );
  OAI22_X1 U23695 ( .A1(n21903), .A2(n21902), .B1(n21901), .B2(n21900), .ZN(
        n21950) );
  AOI222_X1 U23696 ( .A1(n21906), .A2(n21905), .B1(n21906), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C1(n21905), .C2(n21904), .ZN(
        n21908) );
  AOI21_X1 U23697 ( .B1(n21908), .B2(n21912), .A(n21907), .ZN(n21911) );
  AOI22_X1 U23698 ( .A1(n21925), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21909), .B2(n21912), .ZN(n21914) );
  OR2_X1 U23699 ( .A1(n21914), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21910) );
  AOI221_X1 U23700 ( .B1(n21911), .B2(n21910), .C1(n21914), .C2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21918) );
  AOI22_X1 U23701 ( .A1(n21925), .A2(n20877), .B1(n21913), .B2(n21912), .ZN(
        n21917) );
  OAI21_X1 U23702 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n21914), .ZN(n21915) );
  AND3_X1 U23703 ( .A1(n21921), .A2(n21920), .A3(n21919), .ZN(n21949) );
  OAI21_X1 U23704 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n21949), .ZN(n21922) );
  OAI21_X1 U23705 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n22332), .A(n21936), 
        .ZN(n21941) );
  NOR3_X1 U23706 ( .A1(n21930), .A2(n21929), .A3(n21941), .ZN(n21931) );
  OR4_X1 U23707 ( .A1(n21934), .A2(n21933), .A3(n21932), .A4(n21931), .ZN(
        P3_U2997) );
  OAI221_X1 U23708 ( .B1(n21937), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21937), 
        .C2(n21936), .A(n21935), .ZN(P3_U3282) );
  AOI22_X1 U23709 ( .A1(n21939), .A2(n21938), .B1(n22285), .B2(n18957), .ZN(
        n21940) );
  INV_X1 U23710 ( .A(n21940), .ZN(n21944) );
  NOR2_X1 U23711 ( .A1(n21942), .A2(n21941), .ZN(n21943) );
  MUX2_X1 U23712 ( .A(n21944), .B(n21943), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n21946) );
  OAI211_X1 U23713 ( .C1(n21947), .C2(n21948), .A(n21946), .B(n21945), .ZN(
        P3_U2996) );
  NOR2_X1 U23714 ( .A1(n21949), .A2(n21948), .ZN(n21952) );
  MUX2_X1 U23715 ( .A(P3_MORE_REG_SCAN_IN), .B(n21950), .S(n21952), .Z(
        P3_U3295) );
  OAI21_X1 U23716 ( .B1(n21952), .B2(n21951), .A(n11548), .ZN(P3_U2637) );
  AOI211_X1 U23717 ( .C1(n22248), .C2(n21955), .A(n21954), .B(n21953), .ZN(
        n21962) );
  INV_X1 U23718 ( .A(n21956), .ZN(n21957) );
  OAI21_X1 U23719 ( .B1(n21957), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n21959) );
  OAI21_X1 U23720 ( .B1(n21959), .B2(n21958), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n21961) );
  NOR2_X1 U23721 ( .A1(n21962), .A2(n22260), .ZN(n21960) );
  AOI22_X1 U23722 ( .A1(n21963), .A2(n21962), .B1(n21961), .B2(n21960), .ZN(
        P1_U3485) );
  AOI22_X1 U23723 ( .A1(n21965), .A2(n22118), .B1(n22106), .B2(n21964), .ZN(
        n21970) );
  NOR2_X1 U23724 ( .A1(n22093), .A2(n21966), .ZN(n21967) );
  AOI221_X1 U23725 ( .B1(n21968), .B2(n13773), .C1(n22038), .C2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(n21967), .ZN(n21969) );
  NAND2_X1 U23726 ( .A1(n21970), .A2(n21969), .ZN(P1_U3018) );
  INV_X1 U23727 ( .A(n22038), .ZN(n21971) );
  OAI21_X1 U23728 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n21972), .A(
        n21971), .ZN(n21973) );
  AOI22_X1 U23729 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21973), .B1(
        n22102), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n21978) );
  NOR2_X1 U23730 ( .A1(n21974), .A2(n22007), .ZN(n22008) );
  NAND2_X1 U23731 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n22008), .ZN(
        n22033) );
  NOR4_X1 U23732 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n20657), .A3(
        n22025), .A4(n22033), .ZN(n21975) );
  AOI22_X1 U23733 ( .A1(n21976), .A2(n22106), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n21975), .ZN(n21977) );
  OAI211_X1 U23734 ( .C1(n21979), .C2(n22043), .A(n21978), .B(n21977), .ZN(
        P1_U3017) );
  OAI21_X1 U23735 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n21996), .ZN(n21992) );
  AOI211_X1 U23736 ( .C1(n21983), .C2(n21982), .A(n21981), .B(n21980), .ZN(
        n22000) );
  INV_X1 U23737 ( .A(n21984), .ZN(n21985) );
  OAI21_X1 U23738 ( .B1(n22000), .B2(n21986), .A(n21985), .ZN(n21989) );
  NOR2_X1 U23739 ( .A1(n21987), .A2(n22043), .ZN(n21988) );
  AOI211_X1 U23740 ( .C1(n22106), .C2(n21990), .A(n21989), .B(n21988), .ZN(
        n21991) );
  OAI21_X1 U23741 ( .B1(n21993), .B2(n21992), .A(n21991), .ZN(P1_U3027) );
  AOI21_X1 U23742 ( .B1(n22106), .B2(n21995), .A(n21994), .ZN(n21999) );
  AOI22_X1 U23743 ( .A1(n21997), .A2(n22118), .B1(n13719), .B2(n21996), .ZN(
        n21998) );
  OAI211_X1 U23744 ( .C1(n22000), .C2(n13719), .A(n21999), .B(n21998), .ZN(
        P1_U3028) );
  OAI22_X1 U23745 ( .A1(n22001), .A2(n22043), .B1(n22115), .B2(n22139), .ZN(
        n22002) );
  NOR2_X1 U23746 ( .A1(n22003), .A2(n22002), .ZN(n22004) );
  OAI221_X1 U23747 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n22007), .C1(
        n22006), .C2(n22005), .A(n22004), .ZN(P1_U3025) );
  AOI22_X1 U23748 ( .A1(n22189), .A2(n22106), .B1(n22102), .B2(
        P1_REIP_REG_10__SCAN_IN), .ZN(n22014) );
  INV_X1 U23749 ( .A(n22008), .ZN(n22012) );
  NOR2_X1 U23750 ( .A1(n22010), .A2(n22009), .ZN(n22011) );
  MUX2_X1 U23751 ( .A(n22012), .B(n22011), .S(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(n22013) );
  OAI211_X1 U23752 ( .C1(n22043), .C2(n22015), .A(n22014), .B(n22013), .ZN(
        P1_U3021) );
  NOR2_X1 U23753 ( .A1(n20657), .A2(n22033), .ZN(n22026) );
  OAI21_X1 U23754 ( .B1(n22018), .B2(n22017), .A(n22016), .ZN(n22019) );
  AOI21_X1 U23755 ( .B1(n22021), .B2(n22020), .A(n22019), .ZN(n22037) );
  OAI21_X1 U23756 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n22022), .A(
        n22037), .ZN(n22024) );
  OAI22_X1 U23757 ( .A1(n22211), .A2(n22115), .B1(n22093), .B2(n22220), .ZN(
        n22023) );
  AOI221_X1 U23758 ( .B1(n22026), .B2(n22025), .C1(n22024), .C2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n22023), .ZN(n22027) );
  OAI21_X1 U23759 ( .B1(n22028), .B2(n22043), .A(n22027), .ZN(P1_U3019) );
  INV_X1 U23760 ( .A(n22029), .ZN(n22035) );
  INV_X1 U23761 ( .A(n22030), .ZN(n22200) );
  AOI21_X1 U23762 ( .B1(n22200), .B2(n22106), .A(n22031), .ZN(n22032) );
  OAI21_X1 U23763 ( .B1(n22033), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n22032), .ZN(n22034) );
  AOI21_X1 U23764 ( .B1(n22035), .B2(n22118), .A(n22034), .ZN(n22036) );
  OAI21_X1 U23765 ( .B1(n22037), .B2(n20657), .A(n22036), .ZN(P1_U3020) );
  AOI21_X1 U23766 ( .B1(n22039), .B2(n22041), .A(n22038), .ZN(n22056) );
  NOR3_X1 U23767 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n22041), .A3(
        n22040), .ZN(n22046) );
  OAI22_X1 U23768 ( .A1(n22044), .A2(n22043), .B1(n22115), .B2(n22042), .ZN(
        n22045) );
  AOI211_X1 U23769 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n22102), .A(n22046), 
        .B(n22045), .ZN(n22047) );
  OAI21_X1 U23770 ( .B1(n22056), .B2(n22048), .A(n22047), .ZN(P1_U3013) );
  AOI21_X1 U23771 ( .B1(n22049), .B2(n22061), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n22055) );
  INV_X1 U23772 ( .A(n22050), .ZN(n22052) );
  AOI22_X1 U23773 ( .A1(n22052), .A2(n22118), .B1(n22106), .B2(n22051), .ZN(
        n22054) );
  NAND2_X1 U23774 ( .A1(n22102), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n22053) );
  OAI211_X1 U23775 ( .C1(n22056), .C2(n22055), .A(n22054), .B(n22053), .ZN(
        P1_U3014) );
  OAI22_X1 U23776 ( .A1(n22057), .A2(n20682), .B1(n22115), .B2(n22236), .ZN(
        n22058) );
  AOI21_X1 U23777 ( .B1(n22118), .B2(n22059), .A(n22058), .ZN(n22063) );
  OAI211_X1 U23778 ( .C1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n22061), .B(n22060), .ZN(
        n22062) );
  OAI211_X1 U23779 ( .C1(n22227), .C2(n22093), .A(n22063), .B(n22062), .ZN(
        P1_U3015) );
  INV_X1 U23780 ( .A(n22064), .ZN(n22066) );
  AOI22_X1 U23781 ( .A1(n22066), .A2(n22118), .B1(n22106), .B2(n22065), .ZN(
        n22072) );
  NOR2_X1 U23782 ( .A1(n22093), .A2(n22067), .ZN(n22068) );
  AOI211_X1 U23783 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n22070), .A(
        n22069), .B(n22068), .ZN(n22071) );
  NAND2_X1 U23784 ( .A1(n22072), .A2(n22071), .ZN(P1_U3012) );
  AOI21_X1 U23785 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n22102), .A(n22073), 
        .ZN(n22079) );
  INV_X1 U23786 ( .A(n22074), .ZN(n22077) );
  INV_X1 U23787 ( .A(n22075), .ZN(n22076) );
  AOI22_X1 U23788 ( .A1(n22077), .A2(n22118), .B1(n22106), .B2(n22076), .ZN(
        n22078) );
  OAI211_X1 U23789 ( .C1(n16859), .C2(n22080), .A(n22079), .B(n22078), .ZN(
        P1_U3010) );
  INV_X1 U23790 ( .A(n22081), .ZN(n22083) );
  AOI22_X1 U23791 ( .A1(n22083), .A2(n22118), .B1(n22106), .B2(n22082), .ZN(
        n22091) );
  INV_X1 U23792 ( .A(n22084), .ZN(n22088) );
  NOR2_X1 U23793 ( .A1(n22093), .A2(n22085), .ZN(n22086) );
  AOI221_X1 U23794 ( .B1(n22089), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), 
        .C1(n22088), .C2(n22087), .A(n22086), .ZN(n22090) );
  NAND2_X1 U23795 ( .A1(n22091), .A2(n22090), .ZN(P1_U3004) );
  NOR2_X1 U23796 ( .A1(n22093), .A2(n22092), .ZN(n22096) );
  NOR3_X1 U23797 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n22110), .A3(
        n22094), .ZN(n22095) );
  AOI22_X1 U23798 ( .A1(n22099), .A2(n22106), .B1(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n22098), .ZN(n22100) );
  NAND2_X1 U23799 ( .A1(n22101), .A2(n22100), .ZN(P1_U3006) );
  AOI22_X1 U23800 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n22103), .B1(
        n22102), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n22109) );
  INV_X1 U23801 ( .A(n22104), .ZN(n22107) );
  AOI22_X1 U23802 ( .A1(n22107), .A2(n22118), .B1(n22106), .B2(n22105), .ZN(
        n22108) );
  OAI211_X1 U23803 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n22110), .A(
        n22109), .B(n22108), .ZN(P1_U3008) );
  AOI21_X1 U23804 ( .B1(n22112), .B2(n22111), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n22117) );
  OAI21_X1 U23805 ( .B1(n22115), .B2(n22114), .A(n22113), .ZN(n22116) );
  AOI211_X1 U23806 ( .C1(n22119), .C2(n22118), .A(n22117), .B(n22116), .ZN(
        n22120) );
  OAI221_X1 U23807 ( .B1(n22123), .B2(n22122), .C1(n22123), .C2(n22121), .A(
        n22120), .ZN(P1_U3031) );
  INV_X1 U23808 ( .A(n22124), .ZN(n22134) );
  NAND2_X1 U23809 ( .A1(n22199), .A2(n22125), .ZN(n22126) );
  OAI21_X1 U23810 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n22197), .A(n22126), .ZN(
        n22132) );
  AND2_X1 U23811 ( .A1(n22501), .A2(n22127), .ZN(n22131) );
  AOI22_X1 U23812 ( .A1(n22242), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n22162), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n22128) );
  OAI21_X1 U23813 ( .B1(n22235), .B2(n22129), .A(n22128), .ZN(n22130) );
  OR3_X1 U23814 ( .A1(n22132), .A2(n22131), .A3(n22130), .ZN(n22133) );
  AOI21_X1 U23815 ( .B1(n22135), .B2(n22134), .A(n22133), .ZN(n22136) );
  OAI21_X1 U23816 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n22244), .A(
        n22136), .ZN(P1_U2839) );
  AOI21_X1 U23817 ( .B1(n22222), .B2(n22137), .A(P1_REIP_REG_6__SCAN_IN), .ZN(
        n22146) );
  AOI21_X1 U23818 ( .B1(n22222), .B2(n22147), .A(n22162), .ZN(n22157) );
  OAI22_X1 U23819 ( .A1(n22237), .A2(n22139), .B1(n22138), .B2(n22235), .ZN(
        n22140) );
  AOI211_X1 U23820 ( .C1(n22242), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n22213), .B(n22140), .ZN(n22145) );
  INV_X1 U23821 ( .A(n22141), .ZN(n22142) );
  AOI22_X1 U23822 ( .A1(n22143), .A2(n22215), .B1(n22142), .B2(n22216), .ZN(
        n22144) );
  OAI211_X1 U23823 ( .C1(n22146), .C2(n22157), .A(n22145), .B(n22144), .ZN(
        P1_U2834) );
  NOR3_X1 U23824 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n22197), .A3(n22147), .ZN(
        n22154) );
  OAI21_X1 U23825 ( .B1(n22244), .B2(n22148), .A(n22232), .ZN(n22149) );
  AOI21_X1 U23826 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n22242), .A(
        n22149), .ZN(n22152) );
  NAND2_X1 U23827 ( .A1(n22150), .A2(n22199), .ZN(n22151) );
  OAI211_X1 U23828 ( .C1(n22235), .C2(n16048), .A(n22152), .B(n22151), .ZN(
        n22153) );
  AOI211_X1 U23829 ( .C1(n22155), .C2(n22215), .A(n22154), .B(n22153), .ZN(
        n22156) );
  OAI21_X1 U23830 ( .B1(n22158), .B2(n22157), .A(n22156), .ZN(P1_U2833) );
  AND3_X1 U23831 ( .A1(n22222), .A2(n22172), .A3(n22159), .ZN(n22160) );
  AOI21_X1 U23832 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n22201), .A(n22160), .ZN(
        n22171) );
  OAI21_X1 U23833 ( .B1(n22162), .B2(n22172), .A(n22161), .ZN(n22184) );
  OAI22_X1 U23834 ( .A1(n22184), .A2(n22164), .B1(n22237), .B2(n22163), .ZN(
        n22165) );
  AOI211_X1 U23835 ( .C1(n22242), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n22213), .B(n22165), .ZN(n22170) );
  INV_X1 U23836 ( .A(n22166), .ZN(n22167) );
  AOI22_X1 U23837 ( .A1(n22168), .A2(n22215), .B1(n22167), .B2(n22216), .ZN(
        n22169) );
  NAND3_X1 U23838 ( .A1(n22171), .A2(n22170), .A3(n22169), .ZN(P1_U2832) );
  NOR2_X1 U23839 ( .A1(n22172), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n22177) );
  AOI22_X1 U23840 ( .A1(n22173), .A2(n22199), .B1(n22201), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n22174) );
  OAI211_X1 U23841 ( .C1(n22204), .C2(n22175), .A(n22174), .B(n22232), .ZN(
        n22176) );
  AOI21_X1 U23842 ( .B1(n22177), .B2(n22222), .A(n22176), .ZN(n22182) );
  OAI22_X1 U23843 ( .A1(n22179), .A2(n22238), .B1(n22244), .B2(n22178), .ZN(
        n22180) );
  INV_X1 U23844 ( .A(n22180), .ZN(n22181) );
  OAI211_X1 U23845 ( .C1(n22184), .C2(n22183), .A(n22182), .B(n22181), .ZN(
        P1_U2831) );
  INV_X1 U23846 ( .A(n22185), .ZN(n22198) );
  INV_X1 U23847 ( .A(n22186), .ZN(n22187) );
  NOR3_X1 U23848 ( .A1(n22197), .A2(n22198), .A3(n22187), .ZN(n22188) );
  AOI21_X1 U23849 ( .B1(n22189), .B2(n22199), .A(n22188), .ZN(n22196) );
  OAI21_X1 U23850 ( .B1(n22197), .B2(n22198), .A(n22190), .ZN(n22218) );
  AOI22_X1 U23851 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n22242), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n22218), .ZN(n22195) );
  AOI21_X1 U23852 ( .B1(n22201), .B2(P1_EBX_REG_10__SCAN_IN), .A(n22213), .ZN(
        n22194) );
  AOI22_X1 U23853 ( .A1(n22192), .A2(n22215), .B1(n22191), .B2(n22216), .ZN(
        n22193) );
  NAND4_X1 U23854 ( .A1(n22196), .A2(n22195), .A3(n22194), .A4(n22193), .ZN(
        P1_U2830) );
  NOR2_X1 U23855 ( .A1(n22197), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n22219) );
  AOI22_X1 U23856 ( .A1(n22200), .A2(n22199), .B1(n22198), .B2(n22219), .ZN(
        n22208) );
  INV_X1 U23857 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n22203) );
  AOI22_X1 U23858 ( .A1(n22218), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n22201), 
        .B2(P1_EBX_REG_11__SCAN_IN), .ZN(n22202) );
  OAI211_X1 U23859 ( .C1(n22204), .C2(n22203), .A(n22202), .B(n22232), .ZN(
        n22205) );
  AOI21_X1 U23860 ( .B1(n22215), .B2(n22206), .A(n22205), .ZN(n22207) );
  OAI211_X1 U23861 ( .C1(n22209), .C2(n22244), .A(n22208), .B(n22207), .ZN(
        P1_U2829) );
  OAI22_X1 U23862 ( .A1(n22211), .A2(n22237), .B1(n22235), .B2(n22210), .ZN(
        n22212) );
  AOI211_X1 U23863 ( .C1(n22242), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n22213), .B(n22212), .ZN(n22226) );
  AOI22_X1 U23864 ( .A1(n22217), .A2(n22216), .B1(n22215), .B2(n22214), .ZN(
        n22225) );
  OAI21_X1 U23865 ( .B1(n22219), .B2(n22218), .A(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n22224) );
  NAND3_X1 U23866 ( .A1(n22222), .A2(n22221), .A3(n22220), .ZN(n22223) );
  NAND4_X1 U23867 ( .A1(n22226), .A2(n22225), .A3(n22224), .A4(n22223), .ZN(
        P1_U2828) );
  NOR2_X1 U23868 ( .A1(n22228), .A2(n22227), .ZN(n22230) );
  OAI21_X1 U23869 ( .B1(n22231), .B2(n22230), .A(n22229), .ZN(n22233) );
  OAI211_X1 U23870 ( .C1(n22235), .C2(n22234), .A(n22233), .B(n22232), .ZN(
        n22241) );
  OAI22_X1 U23871 ( .A1(n22239), .A2(n22238), .B1(n22237), .B2(n22236), .ZN(
        n22240) );
  AOI211_X1 U23872 ( .C1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n22242), .A(
        n22241), .B(n22240), .ZN(n22243) );
  OAI21_X1 U23873 ( .B1(n22245), .B2(n22244), .A(n22243), .ZN(P1_U2824) );
  OAI21_X1 U23874 ( .B1(n22247), .B2(n22246), .A(n20696), .ZN(P1_U2806) );
  NAND2_X1 U23875 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22248), .ZN(n22254) );
  INV_X1 U23876 ( .A(n22257), .ZN(n22249) );
  OAI21_X1 U23877 ( .B1(n22250), .B2(n22249), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n22251) );
  OAI211_X1 U23878 ( .C1(n22254), .C2(n22253), .A(n22252), .B(n22251), .ZN(
        P1_U3163) );
  OAI22_X1 U23879 ( .A1(n22257), .A2(n22452), .B1(n22256), .B2(n22255), .ZN(
        P1_U3466) );
  AOI21_X1 U23880 ( .B1(n22260), .B2(n22259), .A(n22258), .ZN(n22261) );
  OAI22_X1 U23881 ( .A1(n22263), .A2(n22262), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n22261), .ZN(n22264) );
  OAI21_X1 U23882 ( .B1(n22266), .B2(n22265), .A(n22264), .ZN(P1_U3161) );
  INV_X1 U23883 ( .A(n22267), .ZN(n22269) );
  OAI21_X1 U23884 ( .B1(n22271), .B2(n22268), .A(n22269), .ZN(P1_U2805) );
  INV_X1 U23885 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22270) );
  OAI21_X1 U23886 ( .B1(n22271), .B2(n22270), .A(n22269), .ZN(P1_U3465) );
  INV_X1 U23887 ( .A(n22272), .ZN(n22274) );
  OAI21_X1 U23888 ( .B1(n22276), .B2(n22273), .A(n22274), .ZN(P2_U2818) );
  OAI21_X1 U23889 ( .B1(n22276), .B2(n22275), .A(n22274), .ZN(P2_U3592) );
  INV_X1 U23890 ( .A(n22277), .ZN(n22279) );
  OAI21_X1 U23891 ( .B1(n22281), .B2(n22278), .A(n22279), .ZN(P3_U2636) );
  OAI21_X1 U23892 ( .B1(n22281), .B2(n22280), .A(n22279), .ZN(P3_U3281) );
  INV_X1 U23893 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22282) );
  AOI21_X1 U23894 ( .B1(HOLD), .B2(n22283), .A(n22282), .ZN(n22287) );
  AOI21_X1 U23895 ( .B1(n22285), .B2(P3_STATE_REG_1__SCAN_IN), .A(n22284), 
        .ZN(n22340) );
  OAI21_X1 U23896 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n22336), .A(
        P3_STATE_REG_2__SCAN_IN), .ZN(n22339) );
  INV_X1 U23897 ( .A(n22339), .ZN(n22286) );
  OAI22_X1 U23898 ( .A1(n22288), .A2(n22287), .B1(n22340), .B2(n22286), .ZN(
        P3_U3029) );
  AOI21_X1 U23899 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n22295), .A(n22334), .ZN(n22291) );
  AOI21_X1 U23900 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(
        P1_STATE_REG_1__SCAN_IN), .A(n22291), .ZN(n22294) );
  INV_X1 U23901 ( .A(n22289), .ZN(n22290) );
  AOI22_X1 U23902 ( .A1(n22296), .A2(n22336), .B1(n22291), .B2(n22290), .ZN(
        n22293) );
  NOR2_X1 U23903 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n22336), .ZN(n22292) );
  AOI21_X1 U23904 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n22296), .A(n22302), 
        .ZN(n22304) );
  OAI33_X1 U23905 ( .A1(n22302), .A2(n22294), .A3(n22293), .B1(n22295), .B2(
        n22292), .B3(n22304), .ZN(P1_U3196) );
  OAI21_X1 U23906 ( .B1(n22295), .B2(n22334), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22300) );
  OAI221_X1 U23907 ( .B1(n22296), .B2(HOLD), .C1(n22296), .C2(n22295), .A(
        P1_STATE_REG_1__SCAN_IN), .ZN(n22298) );
  OAI211_X1 U23908 ( .C1(n22302), .C2(n22300), .A(n22298), .B(n22297), .ZN(
        P1_U3195) );
  NOR2_X1 U23909 ( .A1(n22299), .A2(n22334), .ZN(n22301) );
  AOI211_X1 U23910 ( .C1(NA), .C2(n22302), .A(n22301), .B(n22300), .ZN(n22303)
         );
  OAI22_X1 U23911 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22304), .B1(n20780), 
        .B2(n22303), .ZN(P1_U3194) );
  AOI21_X1 U23912 ( .B1(n22317), .B2(P2_STATE_REG_1__SCAN_IN), .A(n22323), 
        .ZN(n22319) );
  OAI21_X1 U23913 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n22319), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22309) );
  NOR2_X1 U23914 ( .A1(n22305), .A2(n22336), .ZN(n22318) );
  AOI211_X1 U23915 ( .C1(n22320), .C2(n22307), .A(n22334), .B(n22306), .ZN(
        n22308) );
  AOI211_X1 U23916 ( .C1(n18096), .C2(n22309), .A(n22318), .B(n22308), .ZN(
        n22310) );
  INV_X1 U23917 ( .A(n22310), .ZN(P2_U3209) );
  AOI21_X1 U23918 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n22320), .A(n22334), .ZN(n22316) );
  AOI21_X1 U23919 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(
        P2_STATE_REG_1__SCAN_IN), .A(n22316), .ZN(n22322) );
  INV_X1 U23920 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22311) );
  AOI211_X1 U23921 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(HOLD), .A(n22323), .B(
        n22311), .ZN(n22313) );
  AOI211_X1 U23922 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(n22317), .A(n22313), 
        .B(n22312), .ZN(n22314) );
  OAI21_X1 U23923 ( .B1(n22322), .B2(n22315), .A(n22314), .ZN(P2_U3210) );
  AOI22_X1 U23924 ( .A1(n22317), .A2(n22336), .B1(n22316), .B2(n22315), .ZN(
        n22321) );
  OAI33_X1 U23925 ( .A1(n22323), .A2(n22322), .A3(n22321), .B1(n22320), .B2(
        n22319), .B3(n22318), .ZN(P2_U3211) );
  NOR2_X1 U23926 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22342)
         );
  OAI21_X1 U23927 ( .B1(n22334), .B2(n22335), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n22326) );
  NOR2_X1 U23928 ( .A1(n22332), .A2(n22324), .ZN(n22337) );
  INV_X1 U23929 ( .A(n22337), .ZN(n22325) );
  OAI21_X1 U23930 ( .B1(n22342), .B2(n22326), .A(n22325), .ZN(n22329) );
  OAI211_X1 U23931 ( .C1(n22334), .C2(n22335), .A(P3_STATE_REG_0__SCAN_IN), 
        .B(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22327) );
  AOI21_X1 U23932 ( .B1(n22327), .B2(n22330), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n22328) );
  AOI21_X1 U23933 ( .B1(n22330), .B2(n22329), .A(n22328), .ZN(n22331) );
  OAI221_X1 U23934 ( .B1(n22333), .B2(P3_STATE_REG_2__SCAN_IN), .C1(n22333), 
        .C2(n22332), .A(n22331), .ZN(P3_U3030) );
  OAI22_X1 U23935 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n22335), .B2(n22334), .ZN(n22338)
         );
  OAI221_X1 U23936 ( .B1(n22338), .B2(n22337), .C1(n22338), .C2(n22336), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n22341) );
  OAI22_X1 U23937 ( .A1(n22342), .A2(n22341), .B1(n22340), .B2(n22339), .ZN(
        P3_U3031) );
  NOR2_X1 U23938 ( .A1(n22373), .A2(n22343), .ZN(n22345) );
  AOI21_X1 U23939 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n22377), .A(n22345), 
        .ZN(n22344) );
  OAI21_X1 U23940 ( .B1(n13442), .B2(n22379), .A(n22344), .ZN(P1_U2945) );
  AOI21_X1 U23941 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n22377), .A(n22345), 
        .ZN(n22346) );
  OAI21_X1 U23942 ( .B1(n16199), .B2(n22379), .A(n22346), .ZN(P1_U2960) );
  INV_X1 U23943 ( .A(n22347), .ZN(n22348) );
  NOR2_X1 U23944 ( .A1(n22373), .A2(n22348), .ZN(n22350) );
  AOI21_X1 U23945 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n22377), .A(n22350), 
        .ZN(n22349) );
  OAI21_X1 U23946 ( .B1(n13465), .B2(n22379), .A(n22349), .ZN(P1_U2946) );
  AOI21_X1 U23947 ( .B1(P1_LWORD_REG_9__SCAN_IN), .B2(n22377), .A(n22350), 
        .ZN(n22351) );
  OAI21_X1 U23948 ( .B1(n22352), .B2(n22379), .A(n22351), .ZN(P1_U2961) );
  NOR2_X1 U23949 ( .A1(n22373), .A2(n22353), .ZN(n22355) );
  AOI21_X1 U23950 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n22377), .A(n22355), 
        .ZN(n22354) );
  OAI21_X1 U23951 ( .B1(n13488), .B2(n22379), .A(n22354), .ZN(P1_U2947) );
  AOI21_X1 U23952 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n22377), .A(n22355), 
        .ZN(n22356) );
  OAI21_X1 U23953 ( .B1(n16271), .B2(n22379), .A(n22356), .ZN(P1_U2962) );
  NOR2_X1 U23954 ( .A1(n22373), .A2(n22357), .ZN(n22359) );
  AOI21_X1 U23955 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n22377), .A(n22359), 
        .ZN(n22358) );
  OAI21_X1 U23956 ( .B1(n13511), .B2(n22379), .A(n22358), .ZN(P1_U2948) );
  AOI21_X1 U23957 ( .B1(P1_LWORD_REG_11__SCAN_IN), .B2(n22377), .A(n22359), 
        .ZN(n22360) );
  OAI21_X1 U23958 ( .B1(n16279), .B2(n22379), .A(n22360), .ZN(P1_U2963) );
  INV_X1 U23959 ( .A(n22361), .ZN(n22362) );
  NOR2_X1 U23960 ( .A1(n22373), .A2(n22362), .ZN(n22364) );
  AOI21_X1 U23961 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n22377), .A(n22364), 
        .ZN(n22363) );
  OAI21_X1 U23962 ( .B1(n13533), .B2(n22379), .A(n22363), .ZN(P1_U2949) );
  AOI21_X1 U23963 ( .B1(P1_LWORD_REG_12__SCAN_IN), .B2(n22377), .A(n22364), 
        .ZN(n22365) );
  OAI21_X1 U23964 ( .B1(n22366), .B2(n22379), .A(n22365), .ZN(P1_U2964) );
  NOR2_X1 U23965 ( .A1(n22373), .A2(n22367), .ZN(n22370) );
  AOI21_X1 U23966 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n22377), .A(n22370), 
        .ZN(n22368) );
  OAI21_X1 U23967 ( .B1(n22369), .B2(n22379), .A(n22368), .ZN(P1_U2950) );
  AOI21_X1 U23968 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n22377), .A(n22370), 
        .ZN(n22371) );
  OAI21_X1 U23969 ( .B1(n16790), .B2(n22379), .A(n22371), .ZN(P1_U2965) );
  NOR2_X1 U23970 ( .A1(n22373), .A2(n22372), .ZN(n22376) );
  AOI21_X1 U23971 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n22377), .A(n22376), 
        .ZN(n22374) );
  OAI21_X1 U23972 ( .B1(n22375), .B2(n22379), .A(n22374), .ZN(P1_U2951) );
  AOI21_X1 U23973 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(n22377), .A(n22376), 
        .ZN(n22378) );
  OAI21_X1 U23974 ( .B1(n16786), .B2(n22379), .A(n22378), .ZN(P1_U2966) );
  NAND2_X1 U23975 ( .A1(n22700), .A2(n22497), .ZN(n22382) );
  NOR2_X1 U23976 ( .A1(n22506), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22471) );
  INV_X1 U23977 ( .A(n22471), .ZN(n22381) );
  OAI21_X1 U23978 ( .B1(n22708), .B2(n22382), .A(n22381), .ZN(n22391) );
  OR2_X1 U23979 ( .A1(n22384), .A2(n22383), .ZN(n22419) );
  NOR2_X1 U23980 ( .A1(n22419), .A2(n22501), .ZN(n22389) );
  NAND3_X1 U23981 ( .A1(n22409), .A2(n22408), .A3(n22476), .ZN(n22398) );
  OR2_X1 U23982 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22398), .ZN(
        n22698) );
  OAI22_X1 U23983 ( .A1(n22700), .A2(n22386), .B1(n22698), .B2(n22385), .ZN(
        n22387) );
  INV_X1 U23984 ( .A(n22387), .ZN(n22395) );
  INV_X1 U23985 ( .A(n22389), .ZN(n22390) );
  AOI22_X1 U23986 ( .A1(n22391), .A2(n22390), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22698), .ZN(n22392) );
  AOI22_X1 U23987 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22702), .B1(
        n22708), .B2(n22477), .ZN(n22394) );
  OAI211_X1 U23988 ( .C1(n22705), .C2(n22485), .A(n22395), .B(n22394), .ZN(
        P1_U3033) );
  INV_X1 U23989 ( .A(n22486), .ZN(n22396) );
  INV_X1 U23990 ( .A(n22419), .ZN(n22397) );
  NOR2_X1 U23991 ( .A1(n22487), .A2(n22398), .ZN(n22706) );
  AOI21_X1 U23992 ( .B1(n22397), .B2(n22488), .A(n22706), .ZN(n22399) );
  OAI22_X1 U23993 ( .A1(n22399), .A2(n22506), .B1(n22398), .B2(n22489), .ZN(
        n22707) );
  AOI22_X1 U23994 ( .A1(n22707), .A2(n22507), .B1(n22706), .B2(n22508), .ZN(
        n22404) );
  INV_X1 U23995 ( .A(n22398), .ZN(n22402) );
  INV_X1 U23996 ( .A(n22417), .ZN(n22400) );
  OAI211_X1 U23997 ( .C1(n22400), .C2(n22492), .A(n22497), .B(n22399), .ZN(
        n22401) );
  OAI211_X1 U23998 ( .C1(n22497), .C2(n22402), .A(n22401), .B(n22495), .ZN(
        n22709) );
  AOI22_X1 U23999 ( .A1(n22709), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n22708), .B2(n22515), .ZN(n22403) );
  OAI211_X1 U24000 ( .C1(n22518), .C2(n22712), .A(n22404), .B(n22403), .ZN(
        P1_U3041) );
  NOR3_X1 U24001 ( .A1(n22714), .A2(n22721), .A3(n22506), .ZN(n22406) );
  NOR2_X1 U24002 ( .A1(n22406), .A2(n22471), .ZN(n22413) );
  INV_X1 U24003 ( .A(n22413), .ZN(n22407) );
  NOR2_X1 U24004 ( .A1(n22419), .A2(n15965), .ZN(n22412) );
  NOR2_X1 U24005 ( .A1(n22445), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22433) );
  NAND3_X1 U24006 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n22409), .A3(
        n22408), .ZN(n22420) );
  NOR2_X1 U24007 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22420), .ZN(
        n22713) );
  AOI22_X1 U24008 ( .A1(n22721), .A2(n22477), .B1(n22508), .B2(n22713), .ZN(
        n22415) );
  INV_X1 U24009 ( .A(n22713), .ZN(n22410) );
  NOR2_X1 U24010 ( .A1(n22433), .A2(n22489), .ZN(n22436) );
  AOI21_X1 U24011 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22410), .A(n22436), 
        .ZN(n22411) );
  OAI211_X1 U24012 ( .C1(n22413), .C2(n22412), .A(n22465), .B(n22411), .ZN(
        n22715) );
  AOI22_X1 U24013 ( .A1(n22715), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n22714), .B2(n22515), .ZN(n22414) );
  OAI211_X1 U24014 ( .C1(n22718), .C2(n22485), .A(n22415), .B(n22414), .ZN(
        P1_U3049) );
  INV_X1 U24015 ( .A(n22420), .ZN(n22424) );
  AOI21_X1 U24016 ( .B1(n22417), .B2(n22416), .A(n22506), .ZN(n22427) );
  OR2_X1 U24017 ( .A1(n22419), .A2(n22418), .ZN(n22422) );
  NOR2_X1 U24018 ( .A1(n22487), .A2(n22420), .ZN(n22719) );
  INV_X1 U24019 ( .A(n22719), .ZN(n22421) );
  NAND2_X1 U24020 ( .A1(n22422), .A2(n22421), .ZN(n22423) );
  AOI22_X1 U24021 ( .A1(n22721), .A2(n22515), .B1(n22719), .B2(n22508), .ZN(
        n22430) );
  INV_X1 U24022 ( .A(n22423), .ZN(n22426) );
  OAI21_X1 U24023 ( .B1(n22497), .B2(n22424), .A(n22495), .ZN(n22425) );
  AOI21_X1 U24024 ( .B1(n22427), .B2(n22426), .A(n22425), .ZN(n22428) );
  AOI22_X1 U24025 ( .A1(n22722), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n22477), .B2(n22720), .ZN(n22429) );
  OAI211_X1 U24026 ( .C1(n22725), .C2(n22485), .A(n22430), .B(n22429), .ZN(
        P1_U3057) );
  NOR3_X1 U24027 ( .A1(n22728), .A2(n22727), .A3(n22506), .ZN(n22431) );
  NOR2_X1 U24028 ( .A1(n22431), .A2(n22471), .ZN(n22440) );
  INV_X1 U24029 ( .A(n22440), .ZN(n22434) );
  AND2_X1 U24030 ( .A1(n22432), .A2(n22501), .ZN(n22439) );
  NOR2_X1 U24031 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22435), .ZN(
        n22726) );
  AOI22_X1 U24032 ( .A1(n22727), .A2(n22515), .B1(n22726), .B2(n22508), .ZN(
        n22442) );
  INV_X1 U24033 ( .A(n22726), .ZN(n22437) );
  AOI21_X1 U24034 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22437), .A(n22436), 
        .ZN(n22438) );
  OAI211_X1 U24035 ( .C1(n22440), .C2(n22439), .A(n22512), .B(n22438), .ZN(
        n22729) );
  AOI22_X1 U24036 ( .A1(n22729), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n22477), .B2(n22728), .ZN(n22441) );
  OAI211_X1 U24037 ( .C1(n22732), .C2(n22485), .A(n22442), .B(n22441), .ZN(
        P1_U3081) );
  INV_X1 U24038 ( .A(n22456), .ZN(n22444) );
  NOR2_X1 U24039 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22443), .ZN(
        n22733) );
  AOI21_X1 U24040 ( .B1(n22444), .B2(n15965), .A(n22733), .ZN(n22449) );
  NAND2_X1 U24041 ( .A1(n22446), .A2(n22445), .ZN(n22479) );
  INV_X1 U24042 ( .A(n22459), .ZN(n22447) );
  OAI22_X1 U24043 ( .A1(n22449), .A2(n22506), .B1(n22479), .B2(n22447), .ZN(
        n22734) );
  AOI22_X1 U24044 ( .A1(n22734), .A2(n22507), .B1(n22733), .B2(n22508), .ZN(
        n22454) );
  INV_X1 U24045 ( .A(n22744), .ZN(n22448) );
  OAI21_X1 U24046 ( .B1(n22448), .B2(n22735), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n22450) );
  NAND2_X1 U24047 ( .A1(n22450), .A2(n22449), .ZN(n22451) );
  AOI22_X1 U24048 ( .A1(n22736), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n22735), .B2(n22515), .ZN(n22453) );
  OAI211_X1 U24049 ( .C1(n22518), .C2(n22744), .A(n22454), .B(n22453), .ZN(
        P1_U3097) );
  NOR3_X1 U24050 ( .A1(n22747), .A2(n22746), .A3(n22506), .ZN(n22455) );
  NOR2_X1 U24051 ( .A1(n22455), .A2(n22471), .ZN(n22467) );
  INV_X1 U24052 ( .A(n22467), .ZN(n22460) );
  NOR2_X1 U24053 ( .A1(n22456), .A2(n15965), .ZN(n22466) );
  NAND2_X1 U24054 ( .A1(n22457), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22504) );
  INV_X1 U24055 ( .A(n22504), .ZN(n22458) );
  NOR2_X1 U24056 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22461), .ZN(
        n22745) );
  AOI22_X1 U24057 ( .A1(n22746), .A2(n22477), .B1(n22508), .B2(n22745), .ZN(
        n22469) );
  INV_X1 U24058 ( .A(n22745), .ZN(n22463) );
  NAND2_X1 U24059 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22504), .ZN(n22513) );
  INV_X1 U24060 ( .A(n22513), .ZN(n22462) );
  AOI21_X1 U24061 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22463), .A(n22462), 
        .ZN(n22464) );
  OAI211_X1 U24062 ( .C1(n22467), .C2(n22466), .A(n22465), .B(n22464), .ZN(
        n22748) );
  AOI22_X1 U24063 ( .A1(n22748), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n22747), .B2(n22515), .ZN(n22468) );
  OAI211_X1 U24064 ( .C1(n22751), .C2(n22485), .A(n22469), .B(n22468), .ZN(
        P1_U3113) );
  NOR2_X1 U24065 ( .A1(n22762), .A2(n22506), .ZN(n22473) );
  AOI21_X1 U24066 ( .B1(n22473), .B2(n22472), .A(n22471), .ZN(n22482) );
  INV_X1 U24067 ( .A(n22482), .ZN(n22475) );
  AND2_X1 U24068 ( .A1(n22502), .A2(n15965), .ZN(n22481) );
  INV_X1 U24069 ( .A(n22479), .ZN(n22474) );
  NAND3_X1 U24070 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n22476), .ZN(n22490) );
  NOR2_X1 U24071 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22490), .ZN(
        n22752) );
  AOI22_X1 U24072 ( .A1(n22762), .A2(n22477), .B1(n22508), .B2(n22752), .ZN(
        n22484) );
  INV_X1 U24073 ( .A(n22752), .ZN(n22478) );
  AOI22_X1 U24074 ( .A1(n22479), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n22478), .ZN(n22480) );
  OAI211_X1 U24075 ( .C1(n22482), .C2(n22481), .A(n22512), .B(n22480), .ZN(
        n22755) );
  AOI22_X1 U24076 ( .A1(n22755), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n22754), .B2(n22515), .ZN(n22483) );
  OAI211_X1 U24077 ( .C1(n22759), .C2(n22485), .A(n22484), .B(n22483), .ZN(
        P1_U3129) );
  NOR2_X1 U24078 ( .A1(n22487), .A2(n22490), .ZN(n22760) );
  AOI21_X1 U24079 ( .B1(n22502), .B2(n22488), .A(n22760), .ZN(n22491) );
  OAI22_X1 U24080 ( .A1(n22491), .A2(n22506), .B1(n22490), .B2(n22489), .ZN(
        n22761) );
  AOI22_X1 U24081 ( .A1(n22507), .A2(n22761), .B1(n22508), .B2(n22760), .ZN(
        n22499) );
  INV_X1 U24082 ( .A(n22490), .ZN(n22496) );
  OAI211_X1 U24083 ( .C1(n22493), .C2(n22492), .A(n22497), .B(n22491), .ZN(
        n22494) );
  OAI211_X1 U24084 ( .C1(n22497), .C2(n22496), .A(n22495), .B(n22494), .ZN(
        n22763) );
  AOI22_X1 U24085 ( .A1(n22763), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n22762), .B2(n22515), .ZN(n22498) );
  OAI211_X1 U24086 ( .C1(n22518), .C2(n22766), .A(n22499), .B(n22498), .ZN(
        P1_U3137) );
  NOR2_X1 U24087 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22500), .ZN(
        n22769) );
  NAND2_X1 U24088 ( .A1(n22502), .A2(n22501), .ZN(n22510) );
  INV_X1 U24089 ( .A(n22503), .ZN(n22505) );
  OAI22_X1 U24090 ( .A1(n22510), .A2(n22506), .B1(n22505), .B2(n22504), .ZN(
        n22767) );
  AOI22_X1 U24091 ( .A1(n22508), .A2(n22769), .B1(n22507), .B2(n22767), .ZN(
        n22517) );
  INV_X1 U24092 ( .A(n22776), .ZN(n22509) );
  OAI21_X1 U24093 ( .B1(n22509), .B2(n22772), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n22511) );
  AOI21_X1 U24094 ( .B1(n22511), .B2(n22510), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n22514) );
  AOI22_X1 U24095 ( .A1(n22773), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n22772), .B2(n22515), .ZN(n22516) );
  OAI211_X1 U24096 ( .C1(n22518), .C2(n22776), .A(n22517), .B(n22516), .ZN(
        P1_U3145) );
  OAI22_X1 U24097 ( .A1(n22700), .A2(n11303), .B1(n22519), .B2(n22698), .ZN(
        n22520) );
  INV_X1 U24098 ( .A(n22520), .ZN(n22522) );
  AOI22_X1 U24099 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22702), .B1(
        n22708), .B2(n11302), .ZN(n22521) );
  OAI211_X1 U24100 ( .C1(n22705), .C2(n22541), .A(n22522), .B(n22521), .ZN(
        P1_U3034) );
  AOI22_X1 U24101 ( .A1(n22707), .A2(n22544), .B1(n22545), .B2(n22706), .ZN(
        n22524) );
  AOI22_X1 U24102 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n22709), .B1(
        n22708), .B2(n11304), .ZN(n22523) );
  OAI211_X1 U24103 ( .C1(n11301), .C2(n22712), .A(n22524), .B(n22523), .ZN(
        P1_U3042) );
  AOI22_X1 U24104 ( .A1(n22721), .A2(n11302), .B1(n22545), .B2(n22713), .ZN(
        n22526) );
  AOI22_X1 U24105 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n22715), .B1(
        n22714), .B2(n11304), .ZN(n22525) );
  OAI211_X1 U24106 ( .C1(n22718), .C2(n22541), .A(n22526), .B(n22525), .ZN(
        P1_U3050) );
  AOI22_X1 U24107 ( .A1(n22720), .A2(n11302), .B1(n22545), .B2(n22719), .ZN(
        n22528) );
  AOI22_X1 U24108 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n22722), .B1(
        n22721), .B2(n11304), .ZN(n22527) );
  OAI211_X1 U24109 ( .C1(n22725), .C2(n22541), .A(n22528), .B(n22527), .ZN(
        P1_U3058) );
  AOI22_X1 U24110 ( .A1(n22728), .A2(n11302), .B1(n22545), .B2(n22726), .ZN(
        n22530) );
  AOI22_X1 U24111 ( .A1(n22729), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11304), .B2(n22727), .ZN(n22529) );
  OAI211_X1 U24112 ( .C1(n22732), .C2(n22541), .A(n22530), .B(n22529), .ZN(
        P1_U3082) );
  AOI22_X1 U24113 ( .A1(n22734), .A2(n22544), .B1(n22545), .B2(n22733), .ZN(
        n22532) );
  AOI22_X1 U24114 ( .A1(n22736), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11304), .B2(n22735), .ZN(n22531) );
  OAI211_X1 U24115 ( .C1(n11301), .C2(n22744), .A(n22532), .B(n22531), .ZN(
        P1_U3098) );
  AOI22_X1 U24116 ( .A1(n22740), .A2(n22544), .B1(n22545), .B2(n22739), .ZN(
        n22535) );
  AOI22_X1 U24117 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n22741), .B1(
        n22747), .B2(n11302), .ZN(n22534) );
  OAI211_X1 U24118 ( .C1(n11303), .C2(n22744), .A(n22535), .B(n22534), .ZN(
        P1_U3106) );
  AOI22_X1 U24119 ( .A1(n22746), .A2(n11302), .B1(n22545), .B2(n22745), .ZN(
        n22537) );
  AOI22_X1 U24120 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22748), .B1(
        n22747), .B2(n11304), .ZN(n22536) );
  OAI211_X1 U24121 ( .C1(n22751), .C2(n22541), .A(n22537), .B(n22536), .ZN(
        P1_U3114) );
  AOI22_X1 U24122 ( .A1(n22762), .A2(n11302), .B1(n22545), .B2(n22752), .ZN(
        n22540) );
  AOI22_X1 U24123 ( .A1(n22755), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11304), .B2(n22754), .ZN(n22539) );
  OAI211_X1 U24124 ( .C1(n22759), .C2(n22541), .A(n22540), .B(n22539), .ZN(
        P1_U3130) );
  AOI22_X1 U24125 ( .A1(n22544), .A2(n22761), .B1(n22545), .B2(n22760), .ZN(
        n22543) );
  AOI22_X1 U24126 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n22763), .B1(
        n22762), .B2(n11304), .ZN(n22542) );
  OAI211_X1 U24127 ( .C1(n11301), .C2(n22766), .A(n22543), .B(n22542), .ZN(
        P1_U3138) );
  AOI22_X1 U24128 ( .A1(n22545), .A2(n22769), .B1(n22544), .B2(n22767), .ZN(
        n22548) );
  AOI22_X1 U24129 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n22773), .B1(
        n22772), .B2(n11304), .ZN(n22547) );
  OAI211_X1 U24130 ( .C1(n11301), .C2(n22776), .A(n22548), .B(n22547), .ZN(
        P1_U3146) );
  OAI22_X1 U24131 ( .A1(n22700), .A2(n22565), .B1(n22549), .B2(n22698), .ZN(
        n22550) );
  INV_X1 U24132 ( .A(n22550), .ZN(n22552) );
  AOI22_X1 U24133 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22702), .B1(
        n22708), .B2(n22568), .ZN(n22551) );
  OAI211_X1 U24134 ( .C1(n22705), .C2(n22571), .A(n22552), .B(n22551), .ZN(
        P1_U3035) );
  AOI22_X1 U24135 ( .A1(n22707), .A2(n22574), .B1(n22575), .B2(n22706), .ZN(
        n22554) );
  AOI22_X1 U24136 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n22709), .B1(
        n22708), .B2(n22576), .ZN(n22553) );
  OAI211_X1 U24137 ( .C1(n22579), .C2(n22712), .A(n22554), .B(n22553), .ZN(
        P1_U3043) );
  AOI22_X1 U24138 ( .A1(n22714), .A2(n22576), .B1(n22575), .B2(n22713), .ZN(
        n22556) );
  AOI22_X1 U24139 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22715), .B1(
        n22721), .B2(n22568), .ZN(n22555) );
  OAI211_X1 U24140 ( .C1(n22718), .C2(n22571), .A(n22556), .B(n22555), .ZN(
        P1_U3051) );
  AOI22_X1 U24141 ( .A1(n22720), .A2(n22568), .B1(n22575), .B2(n22719), .ZN(
        n22558) );
  AOI22_X1 U24142 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n22722), .B1(
        n22721), .B2(n22576), .ZN(n22557) );
  OAI211_X1 U24143 ( .C1(n22725), .C2(n22571), .A(n22558), .B(n22557), .ZN(
        P1_U3059) );
  AOI22_X1 U24144 ( .A1(n22727), .A2(n22576), .B1(n22575), .B2(n22726), .ZN(
        n22560) );
  AOI22_X1 U24145 ( .A1(n22729), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n22568), .B2(n22728), .ZN(n22559) );
  OAI211_X1 U24146 ( .C1(n22732), .C2(n22571), .A(n22560), .B(n22559), .ZN(
        P1_U3083) );
  AOI22_X1 U24147 ( .A1(n22734), .A2(n22574), .B1(n22575), .B2(n22733), .ZN(
        n22562) );
  AOI22_X1 U24148 ( .A1(n22736), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n22576), .B2(n22735), .ZN(n22561) );
  OAI211_X1 U24149 ( .C1(n22579), .C2(n22744), .A(n22562), .B(n22561), .ZN(
        P1_U3099) );
  AOI22_X1 U24150 ( .A1(n22740), .A2(n22574), .B1(n22575), .B2(n22739), .ZN(
        n22564) );
  AOI22_X1 U24151 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n22741), .B1(
        n22568), .B2(n22747), .ZN(n22563) );
  OAI211_X1 U24152 ( .C1(n22565), .C2(n22744), .A(n22564), .B(n22563), .ZN(
        P1_U3107) );
  AOI22_X1 U24153 ( .A1(n22747), .A2(n22576), .B1(n22575), .B2(n22745), .ZN(
        n22567) );
  AOI22_X1 U24154 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22748), .B1(
        n22746), .B2(n22568), .ZN(n22566) );
  OAI211_X1 U24155 ( .C1(n22751), .C2(n22571), .A(n22567), .B(n22566), .ZN(
        P1_U3115) );
  AOI22_X1 U24156 ( .A1(n22762), .A2(n22568), .B1(n22575), .B2(n22752), .ZN(
        n22570) );
  AOI22_X1 U24157 ( .A1(n22755), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n22576), .B2(n22754), .ZN(n22569) );
  OAI211_X1 U24158 ( .C1(n22759), .C2(n22571), .A(n22570), .B(n22569), .ZN(
        P1_U3131) );
  AOI22_X1 U24159 ( .A1(n22574), .A2(n22761), .B1(n22575), .B2(n22760), .ZN(
        n22573) );
  AOI22_X1 U24160 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n22763), .B1(
        n22762), .B2(n22576), .ZN(n22572) );
  OAI211_X1 U24161 ( .C1(n22579), .C2(n22766), .A(n22573), .B(n22572), .ZN(
        P1_U3139) );
  AOI22_X1 U24162 ( .A1(n22575), .A2(n22769), .B1(n22574), .B2(n22767), .ZN(
        n22578) );
  AOI22_X1 U24163 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n22773), .B1(
        n22772), .B2(n22576), .ZN(n22577) );
  OAI211_X1 U24164 ( .C1(n22579), .C2(n22776), .A(n22578), .B(n22577), .ZN(
        P1_U3147) );
  OAI22_X1 U24165 ( .A1(n22700), .A2(n22581), .B1(n22698), .B2(n22580), .ZN(
        n22582) );
  INV_X1 U24166 ( .A(n22582), .ZN(n22584) );
  AOI22_X1 U24167 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22702), .B1(
        n22597), .B2(n22708), .ZN(n22583) );
  OAI211_X1 U24168 ( .C1(n22705), .C2(n22600), .A(n22584), .B(n22583), .ZN(
        P1_U3036) );
  AOI22_X1 U24169 ( .A1(n22707), .A2(n22603), .B1(n22706), .B2(n22604), .ZN(
        n22586) );
  AOI22_X1 U24170 ( .A1(n22709), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n22708), .B2(n22605), .ZN(n22585) );
  OAI211_X1 U24171 ( .C1(n22608), .C2(n22712), .A(n22586), .B(n22585), .ZN(
        P1_U3044) );
  AOI22_X1 U24172 ( .A1(n22721), .A2(n22597), .B1(n22604), .B2(n22713), .ZN(
        n22588) );
  AOI22_X1 U24173 ( .A1(n22715), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n22714), .B2(n22605), .ZN(n22587) );
  OAI211_X1 U24174 ( .C1(n22718), .C2(n22600), .A(n22588), .B(n22587), .ZN(
        P1_U3052) );
  AOI22_X1 U24175 ( .A1(n22721), .A2(n22605), .B1(n22719), .B2(n22604), .ZN(
        n22590) );
  AOI22_X1 U24176 ( .A1(n22722), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n22597), .B2(n22720), .ZN(n22589) );
  OAI211_X1 U24177 ( .C1(n22725), .C2(n22600), .A(n22590), .B(n22589), .ZN(
        P1_U3060) );
  AOI22_X1 U24178 ( .A1(n22728), .A2(n22597), .B1(n22604), .B2(n22726), .ZN(
        n22592) );
  AOI22_X1 U24179 ( .A1(n22729), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n22727), .B2(n22605), .ZN(n22591) );
  OAI211_X1 U24180 ( .C1(n22732), .C2(n22600), .A(n22592), .B(n22591), .ZN(
        P1_U3084) );
  AOI22_X1 U24181 ( .A1(n22734), .A2(n22603), .B1(n22733), .B2(n22604), .ZN(
        n22594) );
  AOI22_X1 U24182 ( .A1(n22736), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n22735), .B2(n22605), .ZN(n22593) );
  OAI211_X1 U24183 ( .C1(n22608), .C2(n22744), .A(n22594), .B(n22593), .ZN(
        P1_U3100) );
  AOI22_X1 U24184 ( .A1(n22746), .A2(n22597), .B1(n22604), .B2(n22745), .ZN(
        n22596) );
  AOI22_X1 U24185 ( .A1(n22748), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n22747), .B2(n22605), .ZN(n22595) );
  OAI211_X1 U24186 ( .C1(n22751), .C2(n22600), .A(n22596), .B(n22595), .ZN(
        P1_U3116) );
  AOI22_X1 U24187 ( .A1(n22762), .A2(n22597), .B1(n22604), .B2(n22752), .ZN(
        n22599) );
  AOI22_X1 U24188 ( .A1(n22755), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n22754), .B2(n22605), .ZN(n22598) );
  OAI211_X1 U24189 ( .C1(n22759), .C2(n22600), .A(n22599), .B(n22598), .ZN(
        P1_U3132) );
  AOI22_X1 U24190 ( .A1(n22603), .A2(n22761), .B1(n22604), .B2(n22760), .ZN(
        n22602) );
  AOI22_X1 U24191 ( .A1(n22763), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n22762), .B2(n22605), .ZN(n22601) );
  OAI211_X1 U24192 ( .C1(n22608), .C2(n22766), .A(n22602), .B(n22601), .ZN(
        P1_U3140) );
  AOI22_X1 U24193 ( .A1(n22604), .A2(n22769), .B1(n22603), .B2(n22767), .ZN(
        n22607) );
  AOI22_X1 U24194 ( .A1(n22773), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n22772), .B2(n22605), .ZN(n22606) );
  OAI211_X1 U24195 ( .C1(n22608), .C2(n22776), .A(n22607), .B(n22606), .ZN(
        P1_U3148) );
  OAI22_X1 U24196 ( .A1(n22700), .A2(n11309), .B1(n22609), .B2(n22698), .ZN(
        n22610) );
  INV_X1 U24197 ( .A(n22610), .ZN(n22612) );
  AOI22_X1 U24198 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22702), .B1(
        n22708), .B2(n22627), .ZN(n22611) );
  OAI211_X1 U24199 ( .C1(n22705), .C2(n22630), .A(n22612), .B(n22611), .ZN(
        P1_U3037) );
  AOI22_X1 U24200 ( .A1(n22707), .A2(n22633), .B1(n22634), .B2(n22706), .ZN(
        n22614) );
  AOI22_X1 U24201 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22709), .B1(
        n22708), .B2(n11310), .ZN(n22613) );
  OAI211_X1 U24202 ( .C1(n22638), .C2(n22712), .A(n22614), .B(n22613), .ZN(
        P1_U3045) );
  AOI22_X1 U24203 ( .A1(n22721), .A2(n22627), .B1(n22634), .B2(n22713), .ZN(
        n22616) );
  AOI22_X1 U24204 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22715), .B1(
        n22714), .B2(n11310), .ZN(n22615) );
  OAI211_X1 U24205 ( .C1(n22718), .C2(n22630), .A(n22616), .B(n22615), .ZN(
        P1_U3053) );
  AOI22_X1 U24206 ( .A1(n22721), .A2(n11310), .B1(n22634), .B2(n22719), .ZN(
        n22618) );
  AOI22_X1 U24207 ( .A1(n22722), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n22720), .B2(n22627), .ZN(n22617) );
  OAI211_X1 U24208 ( .C1(n22725), .C2(n22630), .A(n22618), .B(n22617), .ZN(
        P1_U3061) );
  AOI22_X1 U24209 ( .A1(n22727), .A2(n11310), .B1(n22634), .B2(n22726), .ZN(
        n22620) );
  AOI22_X1 U24210 ( .A1(n22729), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n22627), .B2(n22728), .ZN(n22619) );
  OAI211_X1 U24211 ( .C1(n22732), .C2(n22630), .A(n22620), .B(n22619), .ZN(
        P1_U3085) );
  AOI22_X1 U24212 ( .A1(n22734), .A2(n22633), .B1(n22634), .B2(n22733), .ZN(
        n22622) );
  AOI22_X1 U24213 ( .A1(n22736), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11310), .B2(n22735), .ZN(n22621) );
  OAI211_X1 U24214 ( .C1(n22638), .C2(n22744), .A(n22622), .B(n22621), .ZN(
        P1_U3101) );
  AOI22_X1 U24215 ( .A1(n22740), .A2(n22633), .B1(n22634), .B2(n22739), .ZN(
        n22624) );
  AOI22_X1 U24216 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22741), .B1(
        n22627), .B2(n22747), .ZN(n22623) );
  OAI211_X1 U24217 ( .C1(n11309), .C2(n22744), .A(n22624), .B(n22623), .ZN(
        P1_U3109) );
  AOI22_X1 U24218 ( .A1(n22747), .A2(n11310), .B1(n22634), .B2(n22745), .ZN(
        n22626) );
  AOI22_X1 U24219 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22748), .B1(
        n22746), .B2(n22627), .ZN(n22625) );
  OAI211_X1 U24220 ( .C1(n22751), .C2(n22630), .A(n22626), .B(n22625), .ZN(
        P1_U3117) );
  AOI22_X1 U24221 ( .A1(n22762), .A2(n22627), .B1(n22634), .B2(n22752), .ZN(
        n22629) );
  AOI22_X1 U24222 ( .A1(n22755), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11310), .B2(n22754), .ZN(n22628) );
  OAI211_X1 U24223 ( .C1(n22759), .C2(n22630), .A(n22629), .B(n22628), .ZN(
        P1_U3133) );
  AOI22_X1 U24224 ( .A1(n22633), .A2(n22761), .B1(n22634), .B2(n22760), .ZN(
        n22632) );
  AOI22_X1 U24225 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22763), .B1(
        n22762), .B2(n11310), .ZN(n22631) );
  OAI211_X1 U24226 ( .C1(n22638), .C2(n22766), .A(n22632), .B(n22631), .ZN(
        P1_U3141) );
  AOI22_X1 U24227 ( .A1(n22634), .A2(n22769), .B1(n22633), .B2(n22767), .ZN(
        n22637) );
  AOI22_X1 U24228 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22773), .B1(
        n22772), .B2(n11310), .ZN(n22636) );
  OAI211_X1 U24229 ( .C1(n22638), .C2(n22776), .A(n22637), .B(n22636), .ZN(
        P1_U3149) );
  OAI22_X1 U24230 ( .A1(n22700), .A2(n11305), .B1(n22639), .B2(n22698), .ZN(
        n22640) );
  INV_X1 U24231 ( .A(n22640), .ZN(n22642) );
  AOI22_X1 U24232 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22702), .B1(
        n22708), .B2(n22657), .ZN(n22641) );
  OAI211_X1 U24233 ( .C1(n22705), .C2(n22660), .A(n22642), .B(n22641), .ZN(
        P1_U3038) );
  AOI22_X1 U24234 ( .A1(n22707), .A2(n22663), .B1(n22664), .B2(n22706), .ZN(
        n22644) );
  AOI22_X1 U24235 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n22709), .B1(
        n22708), .B2(n11306), .ZN(n22643) );
  OAI211_X1 U24236 ( .C1(n22668), .C2(n22712), .A(n22644), .B(n22643), .ZN(
        P1_U3046) );
  AOI22_X1 U24237 ( .A1(n22721), .A2(n22657), .B1(n22664), .B2(n22713), .ZN(
        n22646) );
  AOI22_X1 U24238 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22715), .B1(
        n22714), .B2(n11306), .ZN(n22645) );
  OAI211_X1 U24239 ( .C1(n22718), .C2(n22660), .A(n22646), .B(n22645), .ZN(
        P1_U3054) );
  AOI22_X1 U24240 ( .A1(n22720), .A2(n22657), .B1(n22664), .B2(n22719), .ZN(
        n22648) );
  AOI22_X1 U24241 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n22722), .B1(
        n22721), .B2(n11306), .ZN(n22647) );
  OAI211_X1 U24242 ( .C1(n22725), .C2(n22660), .A(n22648), .B(n22647), .ZN(
        P1_U3062) );
  AOI22_X1 U24243 ( .A1(n22728), .A2(n22657), .B1(n22664), .B2(n22726), .ZN(
        n22650) );
  AOI22_X1 U24244 ( .A1(n22729), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11306), .B2(n22727), .ZN(n22649) );
  OAI211_X1 U24245 ( .C1(n22732), .C2(n22660), .A(n22650), .B(n22649), .ZN(
        P1_U3086) );
  AOI22_X1 U24246 ( .A1(n22734), .A2(n22663), .B1(n22664), .B2(n22733), .ZN(
        n22652) );
  AOI22_X1 U24247 ( .A1(n22736), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11306), .B2(n22735), .ZN(n22651) );
  OAI211_X1 U24248 ( .C1(n22668), .C2(n22744), .A(n22652), .B(n22651), .ZN(
        P1_U3102) );
  AOI22_X1 U24249 ( .A1(n22740), .A2(n22663), .B1(n22664), .B2(n22739), .ZN(
        n22654) );
  AOI22_X1 U24250 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n22741), .B1(
        n22747), .B2(n22657), .ZN(n22653) );
  OAI211_X1 U24251 ( .C1(n11305), .C2(n22744), .A(n22654), .B(n22653), .ZN(
        P1_U3110) );
  AOI22_X1 U24252 ( .A1(n22747), .A2(n11306), .B1(n22664), .B2(n22745), .ZN(
        n22656) );
  AOI22_X1 U24253 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n22748), .B1(
        n22746), .B2(n22657), .ZN(n22655) );
  OAI211_X1 U24254 ( .C1(n22751), .C2(n22660), .A(n22656), .B(n22655), .ZN(
        P1_U3118) );
  AOI22_X1 U24255 ( .A1(n22762), .A2(n22657), .B1(n22664), .B2(n22752), .ZN(
        n22659) );
  AOI22_X1 U24256 ( .A1(n22755), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11306), .B2(n22754), .ZN(n22658) );
  OAI211_X1 U24257 ( .C1(n22759), .C2(n22660), .A(n22659), .B(n22658), .ZN(
        P1_U3134) );
  AOI22_X1 U24258 ( .A1(n22663), .A2(n22761), .B1(n22664), .B2(n22760), .ZN(
        n22662) );
  AOI22_X1 U24259 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n22763), .B1(
        n22762), .B2(n11306), .ZN(n22661) );
  OAI211_X1 U24260 ( .C1(n22668), .C2(n22766), .A(n22662), .B(n22661), .ZN(
        P1_U3142) );
  AOI22_X1 U24261 ( .A1(n22664), .A2(n22769), .B1(n22663), .B2(n22767), .ZN(
        n22667) );
  AOI22_X1 U24262 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n22773), .B1(
        n22772), .B2(n11306), .ZN(n22666) );
  OAI211_X1 U24263 ( .C1(n22668), .C2(n22776), .A(n22667), .B(n22666), .ZN(
        P1_U3150) );
  OAI22_X1 U24264 ( .A1(n22700), .A2(n22670), .B1(n22698), .B2(n22669), .ZN(
        n22671) );
  INV_X1 U24265 ( .A(n22671), .ZN(n22673) );
  AOI22_X1 U24266 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22702), .B1(
        n22708), .B2(n22686), .ZN(n22672) );
  OAI211_X1 U24267 ( .C1(n22705), .C2(n22689), .A(n22673), .B(n22672), .ZN(
        P1_U3039) );
  AOI22_X1 U24268 ( .A1(n22707), .A2(n22692), .B1(n22706), .B2(n22693), .ZN(
        n22675) );
  AOI22_X1 U24269 ( .A1(n22709), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n22708), .B2(n22694), .ZN(n22674) );
  OAI211_X1 U24270 ( .C1(n22697), .C2(n22712), .A(n22675), .B(n22674), .ZN(
        P1_U3047) );
  AOI22_X1 U24271 ( .A1(n22714), .A2(n22694), .B1(n22713), .B2(n22693), .ZN(
        n22677) );
  AOI22_X1 U24272 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n22715), .B1(
        n22721), .B2(n22686), .ZN(n22676) );
  OAI211_X1 U24273 ( .C1(n22718), .C2(n22689), .A(n22677), .B(n22676), .ZN(
        P1_U3055) );
  AOI22_X1 U24274 ( .A1(n22720), .A2(n22686), .B1(n22693), .B2(n22719), .ZN(
        n22679) );
  AOI22_X1 U24275 ( .A1(n22722), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n22721), .B2(n22694), .ZN(n22678) );
  OAI211_X1 U24276 ( .C1(n22725), .C2(n22689), .A(n22679), .B(n22678), .ZN(
        P1_U3063) );
  AOI22_X1 U24277 ( .A1(n22728), .A2(n22686), .B1(n22693), .B2(n22726), .ZN(
        n22681) );
  AOI22_X1 U24278 ( .A1(n22729), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n22727), .B2(n22694), .ZN(n22680) );
  OAI211_X1 U24279 ( .C1(n22732), .C2(n22689), .A(n22681), .B(n22680), .ZN(
        P1_U3087) );
  AOI22_X1 U24280 ( .A1(n22734), .A2(n22692), .B1(n22733), .B2(n22693), .ZN(
        n22683) );
  AOI22_X1 U24281 ( .A1(n22736), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n22735), .B2(n22694), .ZN(n22682) );
  OAI211_X1 U24282 ( .C1(n22697), .C2(n22744), .A(n22683), .B(n22682), .ZN(
        P1_U3103) );
  AOI22_X1 U24283 ( .A1(n22747), .A2(n22694), .B1(n22693), .B2(n22745), .ZN(
        n22685) );
  AOI22_X1 U24284 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22748), .B1(
        n22686), .B2(n22746), .ZN(n22684) );
  OAI211_X1 U24285 ( .C1(n22751), .C2(n22689), .A(n22685), .B(n22684), .ZN(
        P1_U3119) );
  AOI22_X1 U24286 ( .A1(n22762), .A2(n22686), .B1(n22693), .B2(n22752), .ZN(
        n22688) );
  AOI22_X1 U24287 ( .A1(n22755), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n22754), .B2(n22694), .ZN(n22687) );
  OAI211_X1 U24288 ( .C1(n22759), .C2(n22689), .A(n22688), .B(n22687), .ZN(
        P1_U3135) );
  AOI22_X1 U24289 ( .A1(n22692), .A2(n22761), .B1(n22693), .B2(n22760), .ZN(
        n22691) );
  AOI22_X1 U24290 ( .A1(n22763), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n22762), .B2(n22694), .ZN(n22690) );
  OAI211_X1 U24291 ( .C1(n22697), .C2(n22766), .A(n22691), .B(n22690), .ZN(
        P1_U3143) );
  AOI22_X1 U24292 ( .A1(n22693), .A2(n22769), .B1(n22692), .B2(n22767), .ZN(
        n22696) );
  AOI22_X1 U24293 ( .A1(n22773), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n22772), .B2(n22694), .ZN(n22695) );
  OAI211_X1 U24294 ( .C1(n22697), .C2(n22776), .A(n22696), .B(n22695), .ZN(
        P1_U3151) );
  OAI22_X1 U24295 ( .A1(n22700), .A2(n11307), .B1(n22699), .B2(n22698), .ZN(
        n22701) );
  INV_X1 U24296 ( .A(n22701), .ZN(n22704) );
  AOI22_X1 U24297 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22702), .B1(
        n22708), .B2(n22753), .ZN(n22703) );
  OAI211_X1 U24298 ( .C1(n22705), .C2(n22758), .A(n22704), .B(n22703), .ZN(
        P1_U3040) );
  AOI22_X1 U24299 ( .A1(n22707), .A2(n22768), .B1(n22770), .B2(n22706), .ZN(
        n22711) );
  AOI22_X1 U24300 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22709), .B1(
        n22708), .B2(n11308), .ZN(n22710) );
  OAI211_X1 U24301 ( .C1(n22777), .C2(n22712), .A(n22711), .B(n22710), .ZN(
        P1_U3048) );
  AOI22_X1 U24302 ( .A1(n22721), .A2(n22753), .B1(n22770), .B2(n22713), .ZN(
        n22717) );
  AOI22_X1 U24303 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22715), .B1(
        n22714), .B2(n11308), .ZN(n22716) );
  OAI211_X1 U24304 ( .C1(n22718), .C2(n22758), .A(n22717), .B(n22716), .ZN(
        P1_U3056) );
  AOI22_X1 U24305 ( .A1(n22720), .A2(n22753), .B1(n22770), .B2(n22719), .ZN(
        n22724) );
  AOI22_X1 U24306 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n22722), .B1(
        n22721), .B2(n11308), .ZN(n22723) );
  OAI211_X1 U24307 ( .C1(n22725), .C2(n22758), .A(n22724), .B(n22723), .ZN(
        P1_U3064) );
  AOI22_X1 U24308 ( .A1(n22727), .A2(n11308), .B1(n22770), .B2(n22726), .ZN(
        n22731) );
  AOI22_X1 U24309 ( .A1(n22729), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n22753), .B2(n22728), .ZN(n22730) );
  OAI211_X1 U24310 ( .C1(n22732), .C2(n22758), .A(n22731), .B(n22730), .ZN(
        P1_U3088) );
  AOI22_X1 U24311 ( .A1(n22734), .A2(n22768), .B1(n22770), .B2(n22733), .ZN(
        n22738) );
  AOI22_X1 U24312 ( .A1(n22736), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11308), .B2(n22735), .ZN(n22737) );
  OAI211_X1 U24313 ( .C1(n22777), .C2(n22744), .A(n22738), .B(n22737), .ZN(
        P1_U3104) );
  AOI22_X1 U24314 ( .A1(n22740), .A2(n22768), .B1(n22770), .B2(n22739), .ZN(
        n22743) );
  AOI22_X1 U24315 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22741), .B1(
        n22747), .B2(n22753), .ZN(n22742) );
  OAI211_X1 U24316 ( .C1(n11307), .C2(n22744), .A(n22743), .B(n22742), .ZN(
        P1_U3112) );
  AOI22_X1 U24317 ( .A1(n22746), .A2(n22753), .B1(n22770), .B2(n22745), .ZN(
        n22750) );
  AOI22_X1 U24318 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22748), .B1(
        n22747), .B2(n11308), .ZN(n22749) );
  OAI211_X1 U24319 ( .C1(n22751), .C2(n22758), .A(n22750), .B(n22749), .ZN(
        P1_U3120) );
  AOI22_X1 U24320 ( .A1(n22762), .A2(n22753), .B1(n22770), .B2(n22752), .ZN(
        n22757) );
  AOI22_X1 U24321 ( .A1(n22755), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11308), .B2(n22754), .ZN(n22756) );
  OAI211_X1 U24322 ( .C1(n22759), .C2(n22758), .A(n22757), .B(n22756), .ZN(
        P1_U3136) );
  AOI22_X1 U24323 ( .A1(n22768), .A2(n22761), .B1(n22770), .B2(n22760), .ZN(
        n22765) );
  AOI22_X1 U24324 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22763), .B1(
        n22762), .B2(n11308), .ZN(n22764) );
  OAI211_X1 U24325 ( .C1(n22777), .C2(n22766), .A(n22765), .B(n22764), .ZN(
        P1_U3144) );
  AOI22_X1 U24326 ( .A1(n22770), .A2(n22769), .B1(n22768), .B2(n22767), .ZN(
        n22775) );
  AOI22_X1 U24327 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22773), .B1(
        n22772), .B2(n11308), .ZN(n22774) );
  OAI211_X1 U24328 ( .C1(n22777), .C2(n22776), .A(n22775), .B(n22774), .ZN(
        P1_U3152) );
  INV_X1 U24329 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n22781) );
  AOI22_X1 U24330 ( .A1(n20780), .A2(n22781), .B1(n22779), .B2(n22778), .ZN(
        P1_U3486) );
  OAI21_X1 U24331 ( .B1(n22782), .B2(n22781), .A(n22780), .ZN(P1_U2801) );
  AND3_X1 U14652 ( .A1(n12780), .A2(n12779), .A3(n12778), .ZN(n12781) );
  AND2_X1 U13458 ( .A1(n14497), .A2(n11791), .ZN(n14487) );
  CLKBUF_X1 U11293 ( .A(n12829), .Z(n13578) );
  AND2_X1 U11307 ( .A1(n12025), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12063) );
  AND2_X1 U11328 ( .A1(n14497), .A2(n11792), .ZN(n14489) );
  CLKBUF_X1 U11591 ( .A(n19178), .Z(n11172) );
  CLKBUF_X1 U11825 ( .A(n16435), .Z(n11165) );
  CLKBUF_X1 U12554 ( .A(n13808), .Z(n13818) );
  CLKBUF_X1 U12556 ( .A(n18949), .Z(n18956) );
  CLKBUF_X1 U12985 ( .A(n20808), .Z(n20841) );
  CLKBUF_X2 U13461 ( .A(n21452), .Z(n11152) );
  INV_X2 U13716 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15673) );
endmodule

