

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987;

  INV_X4 U4767 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  CLKBUF_X2 U4769 ( .A(n5703), .Z(n8122) );
  CLKBUF_X2 U4770 ( .A(n5709), .Z(n4273) );
  CLKBUF_X2 U4771 ( .A(n5703), .Z(n7868) );
  INV_X1 U4772 ( .A(n8126), .ZN(n5703) );
  CLKBUF_X1 U4773 ( .A(n5708), .Z(n4272) );
  NAND4_X1 U4774 ( .A1(n5696), .A2(n5694), .A3(n5693), .A4(n5695), .ZN(n6578)
         );
  CLKBUF_X2 U4776 ( .A(n4989), .Z(n7899) );
  CLKBUF_X1 U4777 ( .A(n8223), .Z(n4262) );
  OAI21_X1 U4778 ( .B1(n5611), .B2(n5464), .A(n8587), .ZN(n8223) );
  OR2_X1 U4779 ( .A1(n5118), .A2(n5117), .ZN(n5133) );
  INV_X1 U4780 ( .A(n7899), .ZN(n5223) );
  AND2_X1 U4781 ( .A1(n4627), .A2(n9351), .ZN(n5709) );
  NOR2_X1 U4782 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5621) );
  INV_X2 U4783 ( .A(n7909), .ZN(n6567) );
  OR2_X1 U4784 ( .A1(n5238), .A2(n4803), .ZN(n5248) );
  NAND2_X1 U4786 ( .A1(n5549), .A2(n5548), .ZN(n8252) );
  BUF_X1 U4787 ( .A(n5697), .Z(n6173) );
  XNOR2_X1 U4788 ( .A(n4532), .B(n4972), .ZN(n6295) );
  INV_X1 U4789 ( .A(n5675), .ZN(n5676) );
  AND2_X2 U4790 ( .A1(n5676), .A2(n6170), .ZN(n8126) );
  NAND2_X1 U4791 ( .A1(n5675), .A2(n6583), .ZN(n5865) );
  OAI22_X1 U4792 ( .A1(n8727), .A2(n4613), .B1(n4301), .B2(n4615), .ZN(n8776)
         );
  AOI211_X2 U4793 ( .C1(P1_ADDR_REG_19__SCAN_IN), .C2(n9495), .A(n8943), .B(
        n8942), .ZN(n8944) );
  AOI211_X2 U4794 ( .C1(n9722), .C2(n8606), .A(n8605), .B(n8604), .ZN(n8607)
         );
  AND2_X2 U4795 ( .A1(n7280), .A2(n7452), .ZN(n7391) );
  AOI211_X2 U4796 ( .C1(n9722), .C2(n8616), .A(n8615), .B(n8614), .ZN(n8617)
         );
  INV_X4 U4797 ( .A(n5011), .ZN(n5354) );
  AOI211_X2 U4798 ( .C1(n8379), .C2(n9746), .A(n8384), .B(n8378), .ZN(n5454)
         );
  OR2_X2 U4799 ( .A1(n5701), .A2(n5702), .ZN(n4626) );
  XNOR2_X2 U4800 ( .A(n5364), .B(n5363), .ZN(n5430) );
  INV_X1 U4801 ( .A(n6888), .ZN(n9743) );
  OAI211_X2 U4802 ( .C1(n6283), .C2(n6307), .A(n5052), .B(n5051), .ZN(n6888)
         );
  CLKBUF_X1 U4803 ( .A(n5359), .Z(n4263) );
  BUF_X2 U4805 ( .A(n4997), .Z(n5359) );
  XNOR2_X2 U4806 ( .A(n6578), .B(n7773), .ZN(n6580) );
  BUF_X1 U4807 ( .A(n5692), .Z(n4265) );
  XNOR2_X2 U4808 ( .A(n5716), .B(n5715), .ZN(n6416) );
  NAND2_X2 U4809 ( .A1(n5714), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5716) );
  AOI22_X1 U4810 ( .A1(n9064), .A2(n9065), .B1(n8972), .B2(n9088), .ZN(n9050)
         );
  NAND2_X1 U4811 ( .A1(n8971), .A2(n8970), .ZN(n9064) );
  OAI21_X1 U4812 ( .B1(n9190), .B2(n9214), .A(n9204), .ZN(n8958) );
  NAND2_X1 U4813 ( .A1(n7926), .A2(n7928), .ZN(n5371) );
  NAND2_X1 U4814 ( .A1(n4856), .A2(n4855), .ZN(n5049) );
  INV_X2 U4815 ( .A(n6984), .ZN(n9639) );
  CLKBUF_X3 U4816 ( .A(n5724), .Z(n4266) );
  AND2_X1 U4817 ( .A1(n7771), .A2(n4434), .ZN(n7809) );
  BUF_X2 U4818 ( .A(n5343), .Z(n6261) );
  INV_X1 U4819 ( .A(n8575), .ZN(n9731) );
  CLKBUF_X1 U4820 ( .A(n6144), .Z(n4269) );
  INV_X4 U4821 ( .A(n6216), .ZN(n7538) );
  NAND2_X1 U4822 ( .A1(n6216), .A2(P1_U3084), .ZN(n9349) );
  INV_X2 U4823 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  OAI21_X1 U4824 ( .B1(n7890), .B2(n8060), .A(n8052), .ZN(n7896) );
  AOI211_X1 U4825 ( .C1(n9722), .C2(n8611), .A(n8610), .B(n8609), .ZN(n8612)
         );
  AND2_X1 U4826 ( .A1(n9245), .A2(n9246), .ZN(n4664) );
  NAND2_X1 U4827 ( .A1(n8826), .A2(n8827), .ZN(n6047) );
  AOI21_X1 U4828 ( .B1(n9050), .B2(n8974), .A(n4756), .ZN(n9034) );
  NAND2_X1 U4829 ( .A1(n8745), .A2(n5983), .ZN(n8803) );
  OAI21_X1 U4830 ( .B1(n9162), .B2(n4742), .A(n4739), .ZN(n4738) );
  AOI21_X2 U4831 ( .B1(n8960), .B2(n7567), .A(n9299), .ZN(n9162) );
  OAI21_X1 U4832 ( .B1(n9307), .B2(n8959), .A(n8958), .ZN(n9176) );
  INV_X1 U4833 ( .A(n4740), .ZN(n4739) );
  OAI21_X1 U4834 ( .B1(n7202), .B2(n4693), .A(n4690), .ZN(n4700) );
  NAND2_X1 U4835 ( .A1(n4744), .A2(n9131), .ZN(n4742) );
  NAND2_X1 U4836 ( .A1(n4763), .A2(n4761), .ZN(n8957) );
  NAND2_X1 U4837 ( .A1(n5872), .A2(n8762), .ZN(n8817) );
  NOR2_X1 U4838 ( .A1(n8911), .A2(n9565), .ZN(n8912) );
  NAND2_X1 U4839 ( .A1(n6831), .A2(n6832), .ZN(n6830) );
  NAND2_X1 U4840 ( .A1(n5160), .A2(n5159), .ZN(n7421) );
  AOI22_X1 U4841 ( .A1(n4598), .A2(n4600), .B1(n4596), .B2(n4277), .ZN(n4594)
         );
  OAI21_X1 U4842 ( .B1(n4600), .B2(n4275), .A(n7061), .ZN(n4599) );
  AND2_X1 U4843 ( .A1(n4293), .A2(n5740), .ZN(n4275) );
  OR2_X1 U4844 ( .A1(n4277), .A2(n7060), .ZN(n4600) );
  AND2_X1 U4845 ( .A1(n7947), .A2(n7948), .ZN(n8076) );
  NAND2_X1 U4846 ( .A1(n5104), .A2(n5103), .ZN(n7103) );
  NOR2_X1 U4847 ( .A1(n5375), .A2(n7915), .ZN(n4714) );
  NAND2_X1 U4848 ( .A1(n5084), .A2(n5083), .ZN(n6935) );
  NAND2_X1 U4849 ( .A1(n6858), .A2(n6862), .ZN(n6959) );
  INV_X1 U4850 ( .A(n6743), .ZN(n6797) );
  INV_X2 U4851 ( .A(n9424), .ZN(n9451) );
  AND2_X1 U4852 ( .A1(n4347), .A2(n4346), .ZN(n5701) );
  INV_X2 U4853 ( .A(n8567), .ZN(n8462) );
  NAND2_X1 U4854 ( .A1(n6979), .A2(n6785), .ZN(n6978) );
  NAND3_X1 U4855 ( .A1(n5036), .A2(n4449), .A3(n4302), .ZN(n6821) );
  AND2_X1 U4856 ( .A1(n6774), .A2(n6773), .ZN(n6979) );
  XNOR2_X1 U4857 ( .A(n5049), .B(n5048), .ZN(n6224) );
  CLKBUF_X1 U4858 ( .A(n6578), .Z(n8885) );
  AND4_X1 U4859 ( .A1(n5728), .A2(n5727), .A3(n5726), .A4(n5725), .ZN(n7839)
         );
  AND4_X1 U4860 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n6950)
         );
  AND4_X1 U4861 ( .A1(n5031), .A2(n5030), .A3(n5029), .A4(n5028), .ZN(n6726)
         );
  AND4_X1 U4862 ( .A1(n5060), .A2(n5059), .A3(n5058), .A4(n5057), .ZN(n6851)
         );
  AND4_X1 U4863 ( .A1(n5016), .A2(n5015), .A3(n5014), .A4(n5013), .ZN(n5023)
         );
  NAND3_X1 U4864 ( .A1(n4779), .A2(n5001), .A3(n5000), .ZN(n8314) );
  NAND2_X1 U4865 ( .A1(n4409), .A2(n4852), .ZN(n5035) );
  OAI211_X1 U4866 ( .C1(n6173), .C2(n6228), .A(n5674), .B(n5673), .ZN(n6984)
         );
  AND3_X1 U4867 ( .A1(n5009), .A2(n5008), .A3(n5007), .ZN(n5475) );
  BUF_X2 U4868 ( .A(n5708), .Z(n4270) );
  OR2_X2 U4869 ( .A1(n5606), .A2(n6701), .ZN(n7909) );
  CLKBUF_X1 U4870 ( .A(n5772), .Z(n5967) );
  BUF_X2 U4871 ( .A(n4982), .Z(n5343) );
  AND2_X1 U4872 ( .A1(n7520), .A2(n8114), .ZN(n4982) );
  AND2_X1 U4873 ( .A1(n4829), .A2(n4830), .ZN(n4997) );
  NAND2_X1 U4874 ( .A1(n5637), .A2(n9345), .ZN(n9351) );
  NAND2_X2 U4875 ( .A1(n5697), .A2(n6216), .ZN(n7562) );
  NAND2_X1 U4876 ( .A1(n5697), .A2(n7538), .ZN(n5771) );
  INV_X1 U4877 ( .A(n8114), .ZN(n4829) );
  NAND2_X1 U4878 ( .A1(n6144), .A2(n9488), .ZN(n5697) );
  XNOR2_X1 U4879 ( .A(n4828), .B(P2_IR_REG_30__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U4880 ( .A1(n5669), .A2(n5668), .ZN(n9488) );
  NAND2_X1 U4881 ( .A1(n4778), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U4882 ( .A1(n4826), .A2(n4827), .ZN(n8114) );
  MUX2_X1 U4883 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5666), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5669) );
  XNOR2_X1 U4884 ( .A(n5664), .B(n5663), .ZN(n6144) );
  NAND2_X1 U4885 ( .A1(n4827), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4828) );
  MUX2_X1 U4886 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4823), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n4826) );
  OR2_X1 U4887 ( .A1(n5667), .A2(n5801), .ZN(n5664) );
  INV_X2 U4888 ( .A(n8721), .ZN(n7519) );
  INV_X2 U4889 ( .A(n9344), .ZN(n8117) );
  XNOR2_X1 U4890 ( .A(n4850), .B(SI_4_), .ZN(n5019) );
  AND2_X1 U4891 ( .A1(n5631), .A2(n4632), .ZN(n5667) );
  INV_X2 U4892 ( .A(n6563), .ZN(n4267) );
  INV_X1 U4893 ( .A(n4716), .ZN(n4715) );
  AND2_X1 U4894 ( .A1(n4784), .A2(n4773), .ZN(n4772) );
  NOR3_X1 U4895 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(n4634), .A3(n4794), .ZN(
        n4633) );
  AND4_X1 U4896 ( .A1(n4586), .A2(n4585), .A3(n5624), .A4(n4584), .ZN(n4784)
         );
  INV_X1 U4897 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5643) );
  NOR2_X1 U4898 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4585) );
  NOR2_X1 U4899 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4586) );
  INV_X1 U4900 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8363) );
  NOR2_X1 U4901 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4987) );
  NOR2_X1 U4902 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4816) );
  INV_X1 U4903 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4960) );
  INV_X1 U4904 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5156) );
  INV_X1 U4905 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5363) );
  INV_X1 U4906 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5220) );
  INV_X1 U4907 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5153) );
  INV_X1 U4908 ( .A(n7524), .ZN(n4621) );
  AOI21_X2 U4909 ( .B1(n5389), .B2(n5388), .A(n5387), .ZN(n8466) );
  AND2_X2 U4910 ( .A1(n8275), .A2(n8427), .ZN(n8413) );
  NAND4_X2 U4911 ( .A1(n4976), .A2(n4975), .A3(n4974), .A4(n4973), .ZN(n5369)
         );
  NAND2_X1 U4912 ( .A1(n5677), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5678) );
  XNOR2_X2 U4913 ( .A(n5698), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6480) );
  XNOR2_X2 U4914 ( .A(n4579), .B(n4822), .ZN(n5394) );
  AND3_X2 U4915 ( .A1(n5670), .A2(n5621), .A3(n5622), .ZN(n5732) );
  AOI22_X2 U4916 ( .A1(n8957), .A2(n8956), .B1(n8955), .B2(n9312), .ZN(n9204)
         );
  NAND2_X2 U4917 ( .A1(n6049), .A2(n6048), .ZN(n8735) );
  OAI21_X4 U4918 ( .B1(n7346), .B2(n5817), .A(n5816), .ZN(n7299) );
  AND2_X1 U4919 ( .A1(n8115), .A2(n5638), .ZN(n5724) );
  BUF_X2 U4920 ( .A(n5708), .Z(n4271) );
  AND3_X1 U4921 ( .A1(n5637), .A2(n9345), .A3(n4627), .ZN(n5708) );
  NOR2_X2 U4922 ( .A1(n8485), .A2(n8471), .ZN(n8470) );
  OR2_X2 U4923 ( .A1(n8501), .A2(n8487), .ZN(n8485) );
  OR2_X1 U4924 ( .A1(n8590), .A2(n9715), .ZN(n8592) );
  OAI21_X2 U4925 ( .B1(n7299), .B2(n4604), .A(n4602), .ZN(n8763) );
  XNOR2_X2 U4926 ( .A(n5633), .B(n9346), .ZN(n8115) );
  INV_X4 U4927 ( .A(n6283), .ZN(n4560) );
  NAND2_X1 U4928 ( .A1(n4516), .A2(n4515), .ZN(n4514) );
  NAND2_X1 U4929 ( .A1(n7667), .A2(n7752), .ZN(n4515) );
  NAND2_X1 U4930 ( .A1(n7666), .A2(n7753), .ZN(n4516) );
  NAND2_X1 U4931 ( .A1(n4905), .A2(n4904), .ZN(n4908) );
  AOI21_X1 U4932 ( .B1(n5128), .B2(n4892), .A(n4408), .ZN(n4407) );
  INV_X1 U4933 ( .A(n4786), .ZN(n4408) );
  NAND2_X1 U4934 ( .A1(n5567), .A2(n5566), .ZN(n5571) );
  AOI21_X1 U4935 ( .B1(n4657), .B2(n4655), .A(n4320), .ZN(n4654) );
  NAND2_X1 U4936 ( .A1(n8966), .A2(n9109), .ZN(n8970) );
  INV_X1 U4937 ( .A(n4769), .ZN(n4767) );
  OR2_X1 U4938 ( .A1(n6339), .A2(n6338), .ZN(n4530) );
  INV_X1 U4939 ( .A(n4509), .ZN(n4508) );
  AOI21_X1 U4940 ( .B1(n7684), .B2(n4510), .A(n7683), .ZN(n4509) );
  INV_X1 U4941 ( .A(n7708), .ZN(n4500) );
  NOR2_X1 U4942 ( .A1(n4473), .A2(n8452), .ZN(n8016) );
  NOR2_X1 U4943 ( .A1(n8535), .A2(n8552), .ZN(n4446) );
  INV_X1 U4944 ( .A(n5217), .ZN(n4389) );
  NAND2_X1 U4945 ( .A1(n4411), .A2(n4414), .ZN(n4874) );
  INV_X1 U4946 ( .A(n4415), .ZN(n4414) );
  OAI21_X1 U4947 ( .B1(n4417), .B2(n4416), .A(n4785), .ZN(n4415) );
  NAND2_X1 U4948 ( .A1(n4717), .A2(n4719), .ZN(n7890) );
  AND2_X1 U4949 ( .A1(n4720), .A2(n8041), .ZN(n4719) );
  NAND2_X1 U4950 ( .A1(n4722), .A2(n4721), .ZN(n4720) );
  NOR2_X1 U4951 ( .A1(n7885), .A2(n6771), .ZN(n8060) );
  NAND2_X1 U4952 ( .A1(n4805), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5273) );
  INV_X1 U4953 ( .A(n5258), .ZN(n4805) );
  OR2_X1 U4954 ( .A1(n8471), .A2(n8156), .ZN(n8015) );
  OR2_X1 U4955 ( .A1(n7421), .A2(n7388), .ZN(n7976) );
  AND2_X1 U4956 ( .A1(n8084), .A2(n7967), .ZN(n4732) );
  NAND2_X1 U4957 ( .A1(n8417), .A2(n8109), .ZN(n8064) );
  INV_X1 U4958 ( .A(n8696), .ZN(n8487) );
  NAND2_X1 U4959 ( .A1(n4606), .A2(n4609), .ZN(n6044) );
  AND2_X1 U4960 ( .A1(n4610), .A2(n6021), .ZN(n4609) );
  OR2_X1 U4961 ( .A1(n9140), .A2(n9290), .ZN(n4557) );
  OAI21_X1 U4962 ( .B1(n4743), .B2(n4741), .A(n4336), .ZN(n4740) );
  INV_X1 U4963 ( .A(n9131), .ZN(n4741) );
  NAND2_X1 U4964 ( .A1(n5697), .A2(n4480), .ZN(n4481) );
  NOR2_X1 U4965 ( .A1(n6217), .A2(n6216), .ZN(n4480) );
  NAND2_X1 U4966 ( .A1(n4916), .A2(n4915), .ZN(n5186) );
  NAND2_X1 U4967 ( .A1(n4402), .A2(n4400), .ZN(n4916) );
  AOI21_X1 U4968 ( .B1(n4298), .B2(n4406), .A(n4401), .ZN(n4400) );
  NAND2_X1 U4969 ( .A1(n4908), .A2(n4907), .ZN(n5170) );
  XNOR2_X1 U4970 ( .A(n4900), .B(SI_14_), .ZN(n5151) );
  NAND2_X1 U4971 ( .A1(n4403), .A2(n4407), .ZN(n4899) );
  NAND2_X1 U4972 ( .A1(n5129), .A2(n4892), .ZN(n4403) );
  NAND2_X1 U4973 ( .A1(n4868), .A2(n4867), .ZN(n5078) );
  NOR2_X1 U4974 ( .A1(n7414), .A2(n4696), .ZN(n4695) );
  OR2_X1 U4975 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  OR2_X1 U4976 ( .A1(n8145), .A2(n5589), .ZN(n4701) );
  NOR2_X1 U4977 ( .A1(n8145), .A2(n8262), .ZN(n4703) );
  OAI21_X1 U4978 ( .B1(n8062), .B2(n4455), .A(n4452), .ZN(n8065) );
  NAND2_X1 U4979 ( .A1(n4456), .A2(n8058), .ZN(n4455) );
  INV_X1 U4980 ( .A(n4453), .ZN(n4452) );
  AND2_X1 U4981 ( .A1(n4835), .A2(n4834), .ZN(n8157) );
  AND3_X1 U4982 ( .A1(n5252), .A2(n5251), .A3(n5250), .ZN(n8244) );
  XNOR2_X1 U4983 ( .A(n8346), .B(n8342), .ZN(n8338) );
  OR2_X1 U4984 ( .A1(n8552), .A2(n8253), .ZN(n8527) );
  OR2_X1 U4985 ( .A1(n7210), .A2(n7218), .ZN(n7967) );
  OR2_X1 U4986 ( .A1(n7210), .A2(n8305), .ZN(n5139) );
  CLKBUF_X2 U4987 ( .A(n4450), .Z(n7898) );
  AND2_X1 U4988 ( .A1(n7056), .A2(n8099), .ZN(n9716) );
  NOR2_X1 U4989 ( .A1(n5834), .A2(n7296), .ZN(n4603) );
  NOR2_X1 U4990 ( .A1(n8115), .A2(n4629), .ZN(n4628) );
  NAND2_X1 U4991 ( .A1(n7549), .A2(n7548), .ZN(n9242) );
  OAI21_X1 U4992 ( .B1(n4758), .B2(n4760), .A(n4755), .ZN(n4751) );
  AOI21_X1 U4993 ( .B1(n4757), .B2(n9033), .A(n4321), .ZN(n4755) );
  AND2_X1 U4994 ( .A1(n9273), .A2(n9123), .ZN(n8964) );
  INV_X1 U4995 ( .A(n4766), .ZN(n4765) );
  OAI21_X1 U4996 ( .B1(n4280), .B2(n4770), .A(n7501), .ZN(n4766) );
  NAND2_X1 U4997 ( .A1(n8822), .A2(n8873), .ZN(n4769) );
  OR2_X1 U4998 ( .A1(n8822), .A2(n8873), .ZN(n4770) );
  INV_X1 U4999 ( .A(n9430), .ZN(n4363) );
  INV_X1 U5000 ( .A(n7562), .ZN(n5968) );
  NAND2_X1 U5001 ( .A1(n6861), .A2(n7780), .ZN(n6947) );
  OAI21_X1 U5002 ( .B1(n5129), .B2(n5128), .A(n4892), .ZN(n5140) );
  NAND2_X1 U5003 ( .A1(n4530), .A2(n4529), .ZN(n4528) );
  NAND2_X1 U5004 ( .A1(n6273), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4529) );
  NAND2_X1 U5005 ( .A1(n7936), .A2(n4476), .ZN(n4479) );
  NAND2_X1 U5006 ( .A1(n4479), .A2(n4477), .ZN(n7941) );
  NOR2_X1 U5007 ( .A1(n7663), .A2(n4521), .ZN(n4520) );
  INV_X1 U5008 ( .A(n7659), .ZN(n4521) );
  NAND2_X1 U5009 ( .A1(n4518), .A2(n4520), .ZN(n4517) );
  AOI21_X1 U5010 ( .B1(n7958), .B2(n4462), .A(n4460), .ZN(n4459) );
  OAI21_X1 U5011 ( .B1(n7966), .B2(n7959), .A(n4461), .ZN(n4460) );
  AND2_X1 U5012 ( .A1(n8083), .A2(n4463), .ZN(n4462) );
  AOI21_X1 U5013 ( .B1(n7964), .B2(n7963), .A(n4464), .ZN(n4469) );
  NOR2_X1 U5014 ( .A1(n4468), .A2(n4478), .ZN(n4467) );
  NOR2_X1 U5015 ( .A1(n7968), .A2(n7969), .ZN(n4468) );
  OAI21_X1 U5016 ( .B1(n4514), .B2(n7673), .A(n7672), .ZN(n4513) );
  NOR2_X1 U5017 ( .A1(n4500), .A2(n4495), .ZN(n4494) );
  NOR2_X1 U5018 ( .A1(n4497), .A2(n4496), .ZN(n4495) );
  INV_X1 U5019 ( .A(n9206), .ZN(n4496) );
  INV_X1 U5020 ( .A(n7707), .ZN(n4497) );
  NOR2_X1 U5021 ( .A1(n4500), .A2(n4499), .ZN(n4498) );
  NAND2_X1 U5022 ( .A1(n7704), .A2(n9177), .ZN(n4499) );
  OAI21_X1 U5023 ( .B1(n8016), .B2(n4471), .A(n8021), .ZN(n4470) );
  NAND2_X1 U5024 ( .A1(n4490), .A2(n9073), .ZN(n4487) );
  NOR2_X1 U5025 ( .A1(n7731), .A2(n7753), .ZN(n4490) );
  NAND2_X1 U5026 ( .A1(n9055), .A2(n9073), .ZN(n4488) );
  OR2_X1 U5027 ( .A1(n8679), .A2(n7905), .ZN(n8063) );
  NAND2_X1 U5028 ( .A1(n4446), .A2(n8703), .ZN(n4445) );
  NOR2_X1 U5029 ( .A1(n9315), .A2(n9312), .ZN(n4545) );
  INV_X1 U5030 ( .A(n4638), .ZN(n4401) );
  AOI21_X1 U5031 ( .B1(n4640), .B2(n4289), .A(n4639), .ZN(n4638) );
  INV_X1 U5032 ( .A(n4957), .ZN(n4639) );
  NAND2_X1 U5033 ( .A1(n4407), .A2(n4405), .ZN(n4404) );
  INV_X1 U5034 ( .A(n4892), .ZN(n4405) );
  INV_X1 U5035 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4423) );
  INV_X1 U5036 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4422) );
  NOR2_X1 U5037 ( .A1(n7216), .A2(n4699), .ZN(n4698) );
  INV_X1 U5038 ( .A(n5525), .ZN(n4699) );
  INV_X1 U5039 ( .A(n4698), .ZN(n4692) );
  AND2_X1 U5040 ( .A1(n7885), .A2(n6771), .ZN(n8047) );
  OR2_X1 U5041 ( .A1(n8503), .A2(n8173), .ZN(n8008) );
  OR2_X1 U5042 ( .A1(n8287), .A2(n7466), .ZN(n7980) );
  NAND2_X1 U5043 ( .A1(n4799), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5118) );
  INV_X1 U5044 ( .A(n5105), .ZN(n4799) );
  INV_X1 U5045 ( .A(n6226), .ZN(n4451) );
  NOR2_X1 U5046 ( .A1(n8436), .A2(n8616), .ZN(n8427) );
  INV_X1 U5047 ( .A(n5017), .ZN(n4811) );
  NOR2_X1 U5048 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4709) );
  NAND2_X1 U5049 ( .A1(n4599), .A2(n4597), .ZN(n4595) );
  OAI21_X1 U5050 ( .B1(n4619), .B2(n4617), .A(n5915), .ZN(n4616) );
  INV_X1 U5051 ( .A(n4618), .ZN(n4617) );
  OR2_X1 U5052 ( .A1(n6076), .A2(n6161), .ZN(n6077) );
  NOR2_X1 U5053 ( .A1(n8998), .A2(n4368), .ZN(n4364) );
  INV_X1 U5054 ( .A(n4662), .ZN(n4368) );
  OR2_X1 U5055 ( .A1(n9252), .A2(n9058), .ZN(n8999) );
  AND2_X1 U5056 ( .A1(n4660), .A2(n4370), .ZN(n4369) );
  INV_X1 U5057 ( .A(n9056), .ZN(n4370) );
  OR2_X1 U5058 ( .A1(n9278), .A2(n9108), .ZN(n8991) );
  OR2_X1 U5059 ( .A1(n9307), .A2(n9190), .ZN(n9182) );
  AND2_X1 U5060 ( .A1(n4765), .A2(n4297), .ZN(n4764) );
  NAND2_X1 U5061 ( .A1(n4379), .A2(n4380), .ZN(n4378) );
  INV_X1 U5062 ( .A(n7504), .ZN(n4379) );
  INV_X1 U5063 ( .A(n7590), .ZN(n4361) );
  AOI21_X1 U5064 ( .B1(n4360), .B2(n7574), .A(n4358), .ZN(n4357) );
  INV_X1 U5065 ( .A(n7687), .ZN(n4358) );
  OR2_X1 U5066 ( .A1(n8771), .A2(n9436), .ZN(n7688) );
  NAND2_X1 U5067 ( .A1(n8882), .A2(n6957), .ZN(n7583) );
  NAND2_X1 U5068 ( .A1(n8986), .A2(n4635), .ZN(n9130) );
  NOR2_X1 U5069 ( .A1(n4636), .A2(n8987), .ZN(n4635) );
  XNOR2_X1 U5070 ( .A(n7535), .B(n7534), .ZN(n7532) );
  OR2_X1 U5071 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4794) );
  NAND2_X1 U5072 ( .A1(n4425), .A2(n4424), .ZN(n7518) );
  AOI21_X1 U5073 ( .B1(n4426), .B2(n4428), .A(n4343), .ZN(n4424) );
  NAND2_X1 U5074 ( .A1(n5305), .A2(n5304), .ZN(n5316) );
  OAI21_X1 U5075 ( .B1(n5285), .B2(n5284), .A(n5283), .ZN(n5299) );
  NAND2_X1 U5076 ( .A1(n5269), .A2(n4946), .ZN(n5285) );
  OAI21_X1 U5077 ( .B1(n5245), .B2(n4429), .A(n4937), .ZN(n5255) );
  INV_X1 U5078 ( .A(n5244), .ZN(n4429) );
  NAND2_X1 U5079 ( .A1(n4934), .A2(n4933), .ZN(n5245) );
  NAND2_X1 U5080 ( .A1(n5234), .A2(n5233), .ZN(n4934) );
  AOI21_X1 U5081 ( .B1(n4394), .B2(n4393), .A(n4337), .ZN(n4392) );
  INV_X1 U5082 ( .A(n4920), .ZN(n4393) );
  INV_X1 U5083 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4773) );
  XNOR2_X1 U5084 ( .A(n4883), .B(SI_11_), .ZN(n5111) );
  NAND2_X1 U5085 ( .A1(n4878), .A2(n4877), .ZN(n4881) );
  NAND2_X1 U5086 ( .A1(n4874), .A2(n4873), .ZN(n5100) );
  NOR2_X1 U5087 ( .A1(n5078), .A2(n4418), .ZN(n4417) );
  INV_X1 U5088 ( .A(n4863), .ZN(n4418) );
  NAND2_X1 U5089 ( .A1(n4860), .A2(n4859), .ZN(n5066) );
  OAI21_X1 U5090 ( .B1(n7538), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4410), .ZN(
        n4850) );
  OR2_X1 U5091 ( .A1(n6216), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4410) );
  NOR2_X2 U5092 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5670) );
  NAND2_X1 U5093 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n4474) );
  NOR2_X1 U5094 ( .A1(n5529), .A2(n5528), .ZN(n4696) );
  NAND2_X1 U5095 ( .A1(n4806), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5291) );
  XNOR2_X1 U5096 ( .A(n5571), .B(n5569), .ZN(n8238) );
  INV_X1 U5097 ( .A(n5545), .ZN(n4687) );
  NAND2_X1 U5098 ( .A1(n5541), .A2(n5540), .ZN(n8195) );
  INV_X1 U5099 ( .A(n6629), .ZN(n4673) );
  AND2_X1 U5100 ( .A1(n6725), .A2(n4313), .ZN(n4671) );
  AND2_X1 U5101 ( .A1(n5265), .A2(n5264), .ZN(n8156) );
  AND4_X1 U5102 ( .A1(n5167), .A2(n5166), .A3(n5165), .A4(n5164), .ZN(n7388)
         );
  AND4_X1 U5103 ( .A1(n5138), .A2(n5137), .A3(n5136), .A4(n5135), .ZN(n7218)
         );
  AND2_X1 U5104 ( .A1(n4534), .A2(n4533), .ZN(n9954) );
  NAND2_X1 U5105 ( .A1(n6460), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4533) );
  NAND2_X1 U5106 ( .A1(n6891), .A2(n4526), .ZN(n6892) );
  OR2_X1 U5107 ( .A1(n6895), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4526) );
  NOR2_X1 U5108 ( .A1(n6892), .A2(n6893), .ZN(n6995) );
  OR2_X1 U5109 ( .A1(n7441), .A2(n7440), .ZN(n4525) );
  NOR2_X1 U5110 ( .A1(n8336), .A2(n4539), .ZN(n8346) );
  AND2_X1 U5111 ( .A1(n8337), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4539) );
  NAND2_X1 U5112 ( .A1(n8338), .A2(n9895), .ZN(n8347) );
  INV_X1 U5113 ( .A(n7890), .ZN(n7889) );
  NOR2_X1 U5114 ( .A1(n8060), .A2(n8047), .ZN(n8094) );
  NAND2_X1 U5115 ( .A1(n4708), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5221) );
  AND2_X1 U5116 ( .A1(n4295), .A2(n4815), .ZN(n4706) );
  OR2_X1 U5117 ( .A1(n8616), .A2(n8265), .ZN(n8408) );
  NAND2_X1 U5118 ( .A1(n4723), .A2(n4727), .ZN(n4730) );
  NAND2_X1 U5119 ( .A1(n8442), .A2(n5390), .ZN(n4723) );
  NOR2_X1 U5120 ( .A1(n8454), .A2(n8620), .ZN(n5402) );
  NOR2_X1 U5121 ( .A1(n8435), .A2(n4577), .ZN(n4576) );
  INV_X1 U5122 ( .A(n4780), .ZN(n4577) );
  NOR2_X1 U5123 ( .A1(n8696), .A2(n8244), .ZN(n5253) );
  NOR2_X1 U5124 ( .A1(n8535), .A2(n8300), .ZN(n5215) );
  NAND2_X1 U5125 ( .A1(n8715), .A2(n8302), .ZN(n4582) );
  AND2_X1 U5126 ( .A1(n5380), .A2(n7985), .ZN(n4737) );
  OR2_X1 U5127 ( .A1(n7469), .A2(n7983), .ZN(n4583) );
  NOR2_X1 U5128 ( .A1(n4798), .A2(n7250), .ZN(n7280) );
  NAND2_X1 U5129 ( .A1(n7072), .A2(n7968), .ZN(n4733) );
  NAND2_X1 U5130 ( .A1(n5127), .A2(n4571), .ZN(n4570) );
  NOR2_X1 U5131 ( .A1(n8083), .A2(n4572), .ZN(n4571) );
  INV_X1 U5132 ( .A(n5126), .ZN(n4572) );
  AND2_X1 U5133 ( .A1(n7967), .A2(n7911), .ZN(n8083) );
  NAND2_X1 U5134 ( .A1(n6920), .A2(n4306), .ZN(n7150) );
  NAND2_X1 U5135 ( .A1(n6920), .A2(n5087), .ZN(n7169) );
  OAI22_X1 U5136 ( .A1(n6923), .A2(n5085), .B1(n9751), .B2(n8309), .ZN(n7166)
         );
  INV_X1 U5137 ( .A(n4563), .ZN(n4562) );
  OAI21_X1 U5138 ( .B1(n8076), .B2(n4564), .A(n5069), .ZN(n4563) );
  NAND2_X1 U5139 ( .A1(n6881), .A2(n6883), .ZN(n6882) );
  NOR2_X1 U5140 ( .A1(n6822), .A2(n6821), .ZN(n6875) );
  NAND2_X1 U5141 ( .A1(n6641), .A2(n8070), .ZN(n6640) );
  NAND2_X1 U5142 ( .A1(n6283), .A2(n7538), .ZN(n4989) );
  INV_X1 U5143 ( .A(n9716), .ZN(n6701) );
  NAND2_X1 U5144 ( .A1(n5225), .A2(n5224), .ZN(n8517) );
  NAND2_X1 U5146 ( .A1(n7815), .A2(n7809), .ZN(n5682) );
  AND2_X1 U5147 ( .A1(n6130), .A2(n6129), .ZN(n7858) );
  AOI21_X1 U5148 ( .B1(n7764), .B2(n7765), .A(n4434), .ZN(n4433) );
  OR2_X1 U5149 ( .A1(n7762), .A2(n7763), .ZN(n4486) );
  NAND2_X1 U5150 ( .A1(n4485), .A2(n7808), .ZN(n4484) );
  NAND2_X1 U5151 ( .A1(n7766), .A2(n4434), .ZN(n4485) );
  AND4_X1 U5152 ( .A1(n5756), .A2(n5755), .A3(n5754), .A4(n5753), .ZN(n7840)
         );
  INV_X1 U5153 ( .A(n8896), .ZN(n4348) );
  NOR2_X1 U5154 ( .A1(n9242), .A2(n9020), .ZN(n9010) );
  OR2_X1 U5155 ( .A1(n9247), .A2(n9035), .ZN(n9020) );
  AND2_X1 U5156 ( .A1(n6148), .A2(n6089), .ZN(n9053) );
  NOR2_X1 U5157 ( .A1(n9069), .A2(n9090), .ZN(n9072) );
  NAND2_X1 U5158 ( .A1(n4556), .A2(n9103), .ZN(n4555) );
  NAND2_X1 U5159 ( .A1(n8963), .A2(n8962), .ZN(n9098) );
  NAND2_X1 U5160 ( .A1(n9130), .A2(n8988), .ZN(n9134) );
  AOI21_X1 U5161 ( .B1(n4744), .B2(n4749), .A(n4312), .ZN(n4743) );
  INV_X1 U5162 ( .A(n4299), .ZN(n4746) );
  NAND2_X1 U5163 ( .A1(n8961), .A2(n9166), .ZN(n4747) );
  NAND2_X1 U5164 ( .A1(n7721), .A2(n8989), .ZN(n9131) );
  OR2_X1 U5165 ( .A1(n9132), .A2(n8987), .ZN(n9150) );
  NAND2_X1 U5166 ( .A1(n4666), .A2(n8984), .ZN(n9163) );
  NAND2_X1 U5167 ( .A1(n4322), .A2(n4373), .ZN(n4372) );
  AND2_X1 U5168 ( .A1(n7709), .A2(n8985), .ZN(n9164) );
  OR2_X1 U5169 ( .A1(n7624), .A2(n7623), .ZN(n9218) );
  CLKBUF_X1 U5170 ( .A(n9403), .Z(n9404) );
  NOR2_X1 U5171 ( .A1(n4551), .A2(n8771), .ZN(n4550) );
  AND2_X1 U5172 ( .A1(n7688), .A2(n7687), .ZN(n7638) );
  OR2_X1 U5173 ( .A1(n5822), .A2(n6407), .ZN(n5842) );
  OAI21_X1 U5174 ( .B1(n7319), .B2(n7318), .A(n7575), .ZN(n9430) );
  NAND2_X1 U5175 ( .A1(n5784), .A2(n5783), .ZN(n7344) );
  AND2_X1 U5176 ( .A1(n7668), .A2(n7184), .ZN(n7631) );
  INV_X1 U5177 ( .A(n7226), .ZN(n7114) );
  OAI22_X1 U5178 ( .A1(n7822), .A2(n7830), .B1(n8880), .B2(n7824), .ZN(n6964)
         );
  OR2_X1 U5179 ( .A1(n6965), .A2(n7852), .ZN(n7836) );
  NAND2_X1 U5180 ( .A1(n4774), .A2(n6959), .ZN(n7851) );
  AND2_X1 U5181 ( .A1(n6961), .A2(n6958), .ZN(n4774) );
  NAND2_X1 U5182 ( .A1(n6786), .A2(n7777), .ZN(n7582) );
  INV_X1 U5183 ( .A(n8949), .ZN(n9237) );
  NAND2_X1 U5184 ( .A1(n5807), .A2(n5806), .ZN(n7287) );
  INV_X1 U5186 ( .A(n9635), .ZN(n7812) );
  AND2_X1 U5187 ( .A1(n6118), .A2(n5662), .ZN(n6168) );
  AND2_X1 U5188 ( .A1(n4776), .A2(n5632), .ZN(n4775) );
  XNOR2_X1 U5189 ( .A(n5285), .B(n5280), .ZN(n7198) );
  NAND2_X1 U5190 ( .A1(n4637), .A2(n4640), .ZN(n4958) );
  OR2_X1 U5191 ( .A1(n4899), .A2(n4289), .ZN(n4637) );
  NAND2_X1 U5192 ( .A1(n4643), .A2(n4902), .ZN(n5171) );
  NAND2_X1 U5193 ( .A1(n4899), .A2(n4644), .ZN(n4643) );
  CLKBUF_X1 U5194 ( .A(n5757), .Z(n5758) );
  XNOR2_X1 U5195 ( .A(n4853), .B(SI_5_), .ZN(n5034) );
  NAND2_X1 U5196 ( .A1(n4345), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5672) );
  INV_X1 U5197 ( .A(n5670), .ZN(n4345) );
  NAND2_X1 U5198 ( .A1(n4684), .A2(n4682), .ZN(n8163) );
  NAND2_X1 U5199 ( .A1(n8252), .A2(n8251), .ZN(n4684) );
  NOR2_X1 U5200 ( .A1(n8144), .A2(n5594), .ZN(n5603) );
  AOI21_X1 U5201 ( .B1(n4276), .B2(n4683), .A(n4317), .ZN(n4675) );
  NAND2_X1 U5202 ( .A1(n5132), .A2(n5131), .ZN(n7210) );
  NAND3_X1 U5203 ( .A1(n5580), .A2(n5579), .A3(n5578), .ZN(n8181) );
  NAND2_X1 U5204 ( .A1(n8216), .A2(n8215), .ZN(n5578) );
  NAND2_X1 U5205 ( .A1(n5193), .A2(n5192), .ZN(n8552) );
  NAND2_X1 U5206 ( .A1(n4677), .A2(n4679), .ZN(n8227) );
  NAND2_X1 U5207 ( .A1(n4678), .A2(n4682), .ZN(n4677) );
  INV_X1 U5208 ( .A(n8252), .ZN(n4678) );
  OAI21_X1 U5209 ( .B1(n7896), .B2(n8373), .A(n4793), .ZN(n7904) );
  OR2_X1 U5210 ( .A1(n8102), .A2(n8101), .ZN(n4783) );
  NAND2_X1 U5211 ( .A1(n5335), .A2(n5334), .ZN(n8293) );
  XNOR2_X1 U5212 ( .A(n6295), .B(n6271), .ZN(n6371) );
  NOR2_X1 U5213 ( .A1(n9354), .A2(n4296), .ZN(n6339) );
  AND2_X1 U5214 ( .A1(n4528), .A2(n4527), .ZN(n6350) );
  INV_X1 U5215 ( .A(n6351), .ZN(n4527) );
  OR2_X1 U5216 ( .A1(n6287), .A2(n6286), .ZN(n4536) );
  NAND2_X1 U5217 ( .A1(n7260), .A2(n7259), .ZN(n7437) );
  NAND2_X1 U5218 ( .A1(n5190), .A2(n4295), .ZN(n5219) );
  OR2_X1 U5219 ( .A1(n5610), .A2(n6280), .ZN(n8587) );
  OAI22_X1 U5220 ( .A1(n4560), .A2(n4558), .B1(n6283), .B2(n6295), .ZN(n8590)
         );
  INV_X1 U5221 ( .A(n4559), .ZN(n4558) );
  OAI22_X1 U5222 ( .A1(n6217), .A2(n7538), .B1(n6214), .B2(n6216), .ZN(n4559)
         );
  OR3_X1 U5223 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5004) );
  NAND2_X1 U5224 ( .A1(n5890), .A2(n5889), .ZN(n9322) );
  INV_X1 U5225 ( .A(n9103), .ZN(n9273) );
  NAND2_X1 U5226 ( .A1(n5970), .A2(n5969), .ZN(n9295) );
  AOI21_X1 U5227 ( .B1(n8838), .B2(n4603), .A(n4305), .ZN(n4602) );
  NAND2_X1 U5228 ( .A1(n8838), .A2(n4605), .ZN(n4604) );
  AND4_X1 U5229 ( .A1(n6040), .A2(n6039), .A3(n6038), .A4(n6037), .ZN(n9089)
         );
  NAND2_X1 U5230 ( .A1(n5875), .A2(n5874), .ZN(n8822) );
  AND4_X1 U5231 ( .A1(n6014), .A2(n6013), .A3(n6012), .A4(n6011), .ZN(n9154)
         );
  AND4_X1 U5232 ( .A1(n5770), .A2(n5769), .A3(n5768), .A4(n5767), .ZN(n7132)
         );
  INV_X1 U5233 ( .A(n9089), .ZN(n9123) );
  AND2_X1 U5234 ( .A1(n5639), .A2(n4631), .ZN(n4630) );
  INV_X1 U5235 ( .A(n4751), .ZN(n4750) );
  NAND2_X1 U5236 ( .A1(n9009), .A2(n9008), .ZN(n9241) );
  AND2_X1 U5237 ( .A1(n4543), .A2(n4542), .ZN(n9475) );
  AOI21_X1 U5238 ( .B1(n9454), .B2(n9455), .A(n9453), .ZN(n4542) );
  OR2_X1 U5239 ( .A1(n9452), .A2(n9679), .ZN(n4543) );
  NAND2_X1 U5240 ( .A1(n4475), .A2(n7940), .ZN(n7942) );
  INV_X1 U5241 ( .A(n7912), .ZN(n7916) );
  AND2_X1 U5242 ( .A1(n7662), .A2(n7661), .ZN(n4522) );
  NOR2_X1 U5243 ( .A1(n4465), .A2(n4464), .ZN(n4463) );
  INV_X1 U5244 ( .A(n7957), .ZN(n4465) );
  AND2_X1 U5245 ( .A1(n7967), .A2(n4478), .ZN(n4461) );
  OAI21_X1 U5246 ( .B1(n4514), .B2(n7678), .A(n7677), .ZN(n4510) );
  AOI21_X1 U5247 ( .B1(n4466), .B2(n4457), .A(n7974), .ZN(n7979) );
  OAI21_X1 U5248 ( .B1(n4469), .B2(n7970), .A(n4467), .ZN(n4466) );
  NOR2_X1 U5249 ( .A1(n4459), .A2(n4458), .ZN(n4457) );
  OAI211_X1 U5250 ( .C1(n4512), .C2(n7676), .A(n4511), .B(n4508), .ZN(n7702)
         );
  INV_X1 U5251 ( .A(n7701), .ZN(n4511) );
  AND2_X1 U5252 ( .A1(n4513), .A2(n7681), .ZN(n4512) );
  AND2_X1 U5253 ( .A1(n4493), .A2(n4491), .ZN(n7714) );
  INV_X1 U5254 ( .A(n4494), .ZN(n4491) );
  NAND2_X1 U5255 ( .A1(n4493), .A2(n4492), .ZN(n7712) );
  NOR2_X1 U5256 ( .A1(n4494), .A2(n4314), .ZN(n4492) );
  NAND2_X1 U5257 ( .A1(n8435), .A2(n4472), .ZN(n4471) );
  NAND2_X1 U5258 ( .A1(n8457), .A2(n8017), .ZN(n4472) );
  OAI21_X1 U5259 ( .B1(n4504), .B2(n4503), .A(n4502), .ZN(n4501) );
  AND2_X1 U5260 ( .A1(n8991), .A2(n7752), .ZN(n4502) );
  NOR2_X1 U5261 ( .A1(n7724), .A2(n7723), .ZN(n4504) );
  OAI21_X1 U5262 ( .B1(n4507), .B2(n7720), .A(n4506), .ZN(n4505) );
  NOR2_X1 U5263 ( .A1(n7752), .A2(n8990), .ZN(n4506) );
  AOI21_X1 U5264 ( .B1(n7724), .B2(n7719), .A(n4351), .ZN(n4507) );
  OAI21_X1 U5265 ( .B1(n7736), .B2(n4488), .A(n4315), .ZN(n4489) );
  AND2_X1 U5266 ( .A1(n8364), .A2(n8291), .ZN(n8057) );
  INV_X1 U5267 ( .A(n8040), .ZN(n4721) );
  NOR2_X1 U5268 ( .A1(n8092), .A2(n8388), .ZN(n4718) );
  NOR2_X1 U5269 ( .A1(n4612), .A2(n4608), .ZN(n4607) );
  INV_X1 U5270 ( .A(n8805), .ZN(n4608) );
  INV_X1 U5271 ( .A(n8755), .ZN(n4612) );
  NAND2_X1 U5272 ( .A1(n8755), .A2(n4611), .ZN(n4610) );
  AND2_X1 U5273 ( .A1(n7710), .A2(n9182), .ZN(n8982) );
  AND2_X1 U5274 ( .A1(n7662), .A2(n6948), .ZN(n7581) );
  INV_X1 U5275 ( .A(n4427), .ZN(n4426) );
  OAI21_X1 U5276 ( .B1(n5321), .B2(n4428), .A(n5347), .ZN(n4427) );
  INV_X1 U5277 ( .A(n5336), .ZN(n4428) );
  INV_X1 U5278 ( .A(n4407), .ZN(n4406) );
  NOR2_X1 U5279 ( .A1(n4656), .A2(n4653), .ZN(n4652) );
  INV_X1 U5280 ( .A(n4873), .ZN(n4653) );
  INV_X1 U5281 ( .A(n4657), .ZN(n4656) );
  NOR2_X1 U5282 ( .A1(n4885), .A2(n4658), .ZN(n4657) );
  INV_X1 U5283 ( .A(n4881), .ZN(n4658) );
  INV_X1 U5284 ( .A(n5111), .ZN(n4885) );
  INV_X1 U5285 ( .A(n4788), .ZN(n4655) );
  AND2_X1 U5286 ( .A1(n5506), .A2(n5500), .ZN(n4688) );
  INV_X1 U5287 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5025) );
  INV_X2 U5288 ( .A(n5590), .ZN(n5568) );
  OAI21_X1 U5289 ( .B1(n8061), .B2(n4454), .A(n5430), .ZN(n4453) );
  NAND2_X1 U5290 ( .A1(n4456), .A2(n8045), .ZN(n4454) );
  OR2_X1 U5291 ( .A1(n8063), .A2(n4478), .ZN(n4456) );
  AND2_X1 U5292 ( .A1(n4440), .A2(n4441), .ZN(n4439) );
  NOR2_X1 U5293 ( .A1(n8044), .A2(n8606), .ZN(n4441) );
  NOR2_X1 U5294 ( .A1(n8068), .A2(n8030), .ZN(n4729) );
  NOR2_X1 U5295 ( .A1(n8422), .A2(n4728), .ZN(n4727) );
  AND2_X1 U5296 ( .A1(n8443), .A2(n5390), .ZN(n4728) );
  OR2_X1 U5297 ( .A1(n5162), .A2(n5161), .ZN(n5177) );
  NAND2_X1 U5298 ( .A1(n4800), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5144) );
  AND2_X1 U5299 ( .A1(n4437), .A2(n6929), .ZN(n7091) );
  NOR2_X1 U5300 ( .A1(n7360), .A2(n7103), .ZN(n4437) );
  NAND2_X1 U5301 ( .A1(n4292), .A2(n5053), .ZN(n4564) );
  NOR2_X1 U5302 ( .A1(n8076), .A2(n4566), .ZN(n4565) );
  INV_X1 U5303 ( .A(n5053), .ZN(n4566) );
  AND2_X1 U5304 ( .A1(n4438), .A2(n6876), .ZN(n6929) );
  NOR2_X1 U5305 ( .A1(n6935), .A2(n6743), .ZN(n4438) );
  NAND2_X1 U5306 ( .A1(n8315), .A2(n9731), .ZN(n7926) );
  NOR2_X1 U5307 ( .A1(n8503), .A2(n4445), .ZN(n4443) );
  NOR2_X1 U5308 ( .A1(n8551), .A2(n4444), .ZN(n8533) );
  INV_X1 U5309 ( .A(n4446), .ZN(n4444) );
  NOR2_X1 U5310 ( .A1(n8551), .A2(n8552), .ZN(n8550) );
  OR2_X1 U5311 ( .A1(n6643), .A2(n6644), .ZN(n6822) );
  NOR2_X1 U5312 ( .A1(n4735), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4734) );
  NAND2_X1 U5313 ( .A1(n4822), .A2(n4736), .ZN(n4735) );
  INV_X1 U5314 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4948) );
  OR2_X1 U5315 ( .A1(n5089), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5101) );
  INV_X1 U5316 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4810) );
  OR2_X1 U5318 ( .A1(n9237), .A2(n8947), .ZN(n7747) );
  NAND2_X1 U5319 ( .A1(n4398), .A2(n4397), .ZN(n7802) );
  NOR2_X1 U5320 ( .A1(n9552), .A2(n4340), .ZN(n8910) );
  INV_X1 U5321 ( .A(n6168), .ZN(n6170) );
  INV_X1 U5322 ( .A(n9001), .ZN(n4649) );
  NAND2_X1 U5323 ( .A1(n7740), .A2(n9033), .ZN(n4647) );
  OR2_X1 U5324 ( .A1(n6670), .A2(n6669), .ZN(n7550) );
  AND2_X1 U5325 ( .A1(n7728), .A2(n8993), .ZN(n4662) );
  OAI22_X1 U5326 ( .A1(n9130), .A2(n4349), .B1(n4316), .B2(n8990), .ZN(n9104)
         );
  NAND2_X1 U5327 ( .A1(n4352), .A2(n8989), .ZN(n4349) );
  OR2_X1 U5328 ( .A1(n8988), .A2(n4351), .ZN(n4350) );
  OR2_X1 U5329 ( .A1(n6025), .A2(n6024), .ZN(n6035) );
  NOR2_X1 U5330 ( .A1(n9278), .A2(n4557), .ZN(n4556) );
  NAND2_X1 U5331 ( .A1(n4374), .A2(n8983), .ZN(n4373) );
  INV_X1 U5332 ( .A(n4375), .ZN(n4374) );
  AOI21_X1 U5333 ( .B1(n4376), .B2(n7640), .A(n7623), .ZN(n4375) );
  OR2_X1 U5334 ( .A1(n7567), .A2(n9208), .ZN(n7710) );
  NAND2_X1 U5335 ( .A1(n9368), .A2(n4552), .ZN(n4551) );
  INV_X1 U5336 ( .A(n7344), .ZN(n4552) );
  OR2_X1 U5337 ( .A1(n5796), .A2(n5785), .ZN(n5822) );
  INV_X1 U5338 ( .A(n7581), .ZN(n6949) );
  INV_X1 U5339 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5764) );
  AND2_X1 U5340 ( .A1(n9644), .A2(n6586), .ZN(n4546) );
  OR2_X1 U5341 ( .A1(n9099), .A2(n8967), .ZN(n9090) );
  NAND2_X1 U5342 ( .A1(n9195), .A2(n9173), .ZN(n9167) );
  NAND2_X1 U5343 ( .A1(n9226), .A2(n4545), .ZN(n9209) );
  OAI21_X1 U5344 ( .B1(n7518), .B2(n7517), .A(n7516), .ZN(n7535) );
  AND2_X1 U5345 ( .A1(n5663), .A2(n4777), .ZN(n4776) );
  INV_X1 U5346 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4777) );
  NAND2_X1 U5347 ( .A1(n5663), .A2(n5660), .ZN(n4634) );
  NOR3_X1 U5348 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .A3(
        n4794), .ZN(n4632) );
  NOR2_X1 U5349 ( .A1(n4794), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4540) );
  NAND2_X1 U5350 ( .A1(n5316), .A2(n5315), .ZN(n5322) );
  OAI21_X1 U5351 ( .B1(n5299), .B2(n5298), .A(n5297), .ZN(n5305) );
  NAND2_X1 U5352 ( .A1(n5647), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5649) );
  OAI21_X2 U5353 ( .B1(n5679), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U5354 ( .A1(n4386), .A2(n4387), .ZN(n5234) );
  AOI21_X1 U5355 ( .B1(n4278), .B2(n4395), .A(n4388), .ZN(n4387) );
  INV_X1 U5356 ( .A(n4928), .ZN(n4388) );
  AND2_X1 U5357 ( .A1(n4933), .A2(n4932), .ZN(n5233) );
  INV_X1 U5358 ( .A(n4902), .ZN(n4642) );
  INV_X1 U5359 ( .A(n4641), .ZN(n4640) );
  OAI21_X1 U5360 ( .B1(n4644), .B2(n4289), .A(n4908), .ZN(n4641) );
  NOR2_X1 U5361 ( .A1(n4903), .A2(n4645), .ZN(n4644) );
  INV_X1 U5362 ( .A(n4898), .ZN(n4645) );
  INV_X1 U5363 ( .A(n5151), .ZN(n4903) );
  NAND2_X1 U5364 ( .A1(n4889), .A2(n4888), .ZN(n4892) );
  XNOR2_X1 U5365 ( .A(n4862), .B(SI_7_), .ZN(n5065) );
  INV_X1 U5366 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4420) );
  NAND2_X1 U5367 ( .A1(n7202), .A2(n4698), .ZN(n4697) );
  INV_X1 U5368 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5070) );
  OR2_X1 U5369 ( .A1(n5071), .A2(n5070), .ZN(n5094) );
  INV_X1 U5370 ( .A(n8226), .ZN(n4676) );
  NAND2_X1 U5371 ( .A1(n4804), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5258) );
  OAI21_X1 U5372 ( .B1(n8216), .B2(n8295), .A(n4331), .ZN(n5573) );
  OR2_X1 U5373 ( .A1(n5179), .A2(n7430), .ZN(n5195) );
  NAND2_X1 U5374 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5026) );
  INV_X1 U5375 ( .A(n6623), .ZN(n5482) );
  NAND2_X1 U5376 ( .A1(n6850), .A2(n6849), .ZN(n4689) );
  AOI21_X1 U5377 ( .B1(n4682), .B2(n4681), .A(n4680), .ZN(n4679) );
  INV_X1 U5378 ( .A(n5558), .ZN(n4680) );
  INV_X1 U5379 ( .A(n8251), .ZN(n4681) );
  INV_X1 U5380 ( .A(n8316), .ZN(n4978) );
  NOR2_X1 U5381 ( .A1(n5026), .A2(n5025), .ZN(n5039) );
  INV_X1 U5382 ( .A(n8228), .ZN(n8264) );
  AOI21_X1 U5383 ( .B1(n4695), .B2(n4692), .A(n4691), .ZN(n4690) );
  INV_X1 U5384 ( .A(n4695), .ZN(n4693) );
  INV_X1 U5385 ( .A(n5535), .ZN(n4691) );
  INV_X1 U5386 ( .A(n8065), .ZN(n8102) );
  AND3_X1 U5387 ( .A1(n5242), .A2(n5241), .A3(n5240), .ZN(n8173) );
  AND4_X1 U5388 ( .A1(n4956), .A2(n4955), .A3(n4954), .A4(n4953), .ZN(n8206)
         );
  AND4_X1 U5389 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n5146), .ZN(n7277)
         );
  AND4_X1 U5390 ( .A1(n5123), .A2(n5122), .A3(n5121), .A4(n5120), .ZN(n7075)
         );
  AND4_X1 U5391 ( .A1(n5110), .A2(n5109), .A3(n5108), .A4(n5107), .ZN(n7033)
         );
  AND4_X1 U5392 ( .A1(n5099), .A2(n5098), .A3(n5097), .A4(n5096), .ZN(n7015)
         );
  OR2_X1 U5393 ( .A1(n6325), .A2(n6324), .ZN(n4534) );
  NOR2_X1 U5394 ( .A1(n6605), .A2(n4537), .ZN(n6608) );
  AND2_X1 U5395 ( .A1(n6606), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4537) );
  NOR2_X1 U5396 ( .A1(n6608), .A2(n6607), .ZN(n6660) );
  NOR2_X1 U5397 ( .A1(n6995), .A2(n4341), .ZN(n6999) );
  NAND2_X1 U5398 ( .A1(n6999), .A2(n6998), .ZN(n7045) );
  INV_X1 U5399 ( .A(n4308), .ZN(n8374) );
  NAND2_X1 U5400 ( .A1(n8413), .A2(n8403), .ZN(n8396) );
  AND2_X1 U5401 ( .A1(n7881), .A2(n5342), .ZN(n8380) );
  NAND2_X1 U5402 ( .A1(n4726), .A2(n4724), .ZN(n8410) );
  NAND2_X1 U5403 ( .A1(n4725), .A2(n4729), .ZN(n4724) );
  NAND2_X1 U5404 ( .A1(n8442), .A2(n4304), .ZN(n4726) );
  INV_X1 U5405 ( .A(n4727), .ZN(n4725) );
  AOI21_X1 U5406 ( .B1(n4576), .B2(n4574), .A(n4318), .ZN(n4573) );
  INV_X1 U5407 ( .A(n4576), .ZN(n4575) );
  NOR2_X1 U5408 ( .A1(n8442), .A2(n8443), .ZN(n8441) );
  INV_X1 U5409 ( .A(n8480), .ZN(n5388) );
  NAND2_X1 U5410 ( .A1(n8495), .A2(n8008), .ZN(n8481) );
  OR2_X1 U5411 ( .A1(n8517), .A2(n8299), .ZN(n5231) );
  AOI21_X1 U5412 ( .B1(n4279), .B2(n7983), .A(n4311), .ZN(n4581) );
  NAND2_X1 U5413 ( .A1(n7465), .A2(n7985), .ZN(n8545) );
  OAI21_X1 U5414 ( .B1(n7270), .B2(n7272), .A(n5169), .ZN(n7384) );
  NAND2_X1 U5415 ( .A1(n7384), .A2(n8086), .ZN(n7383) );
  OR2_X1 U5416 ( .A1(n7152), .A2(n7210), .ZN(n4798) );
  CLKBUF_X1 U5417 ( .A(n7072), .Z(n7073) );
  OR2_X1 U5418 ( .A1(n5124), .A2(n7088), .ZN(n7149) );
  NAND2_X1 U5419 ( .A1(n6929), .A2(n7179), .ZN(n7174) );
  AND2_X1 U5420 ( .A1(n7963), .A2(n7960), .ZN(n8077) );
  NAND2_X1 U5421 ( .A1(n5086), .A2(n5085), .ZN(n6920) );
  INV_X1 U5422 ( .A(n8075), .ZN(n5085) );
  INV_X1 U5423 ( .A(n4714), .ZN(n4713) );
  INV_X1 U5424 ( .A(n7948), .ZN(n4711) );
  NAND2_X1 U5425 ( .A1(n6876), .A2(n6797), .ZN(n6930) );
  AND2_X1 U5426 ( .A1(n6875), .A2(n9743), .ZN(n6876) );
  NAND2_X1 U5427 ( .A1(n4451), .A2(n4450), .ZN(n4449) );
  AND2_X1 U5428 ( .A1(n7914), .A2(n7913), .ZN(n4731) );
  NAND2_X1 U5429 ( .A1(n6545), .A2(n5010), .ZN(n6641) );
  OR2_X1 U5430 ( .A1(n6277), .A2(P2_U3152), .ZN(n6280) );
  NAND2_X1 U5431 ( .A1(n7894), .A2(n7893), .ZN(n8373) );
  NAND2_X1 U5432 ( .A1(n5257), .A2(n5256), .ZN(n8471) );
  AND2_X1 U5433 ( .A1(n4820), .A2(n4821), .ZN(n4435) );
  NAND2_X1 U5434 ( .A1(n5190), .A2(n5189), .ZN(n5204) );
  AND2_X1 U5435 ( .A1(n4959), .A2(n4960), .ZN(n5190) );
  NOR2_X1 U5436 ( .A1(n4716), .A2(n5017), .ZN(n4959) );
  OR2_X1 U5437 ( .A1(n5101), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5113) );
  INV_X1 U5438 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5061) );
  INV_X1 U5439 ( .A(n4599), .ZN(n4598) );
  AND2_X1 U5440 ( .A1(n8794), .A2(n6077), .ZN(n7863) );
  OR2_X1 U5441 ( .A1(n7859), .A2(n7858), .ZN(n7861) );
  AND2_X1 U5442 ( .A1(n8825), .A2(n6042), .ZN(n6046) );
  INV_X1 U5443 ( .A(n8128), .ZN(n6096) );
  INV_X1 U5444 ( .A(n8747), .ZN(n5981) );
  INV_X1 U5445 ( .A(n5835), .ZN(n4605) );
  INV_X1 U5446 ( .A(n6160), .ZN(n4592) );
  OR2_X1 U5447 ( .A1(n4617), .A2(n4301), .ZN(n4613) );
  INV_X1 U5448 ( .A(n4616), .ZN(n4615) );
  OR2_X1 U5449 ( .A1(n6035), .A2(n6034), .ZN(n6052) );
  OR2_X1 U5450 ( .A1(n6052), .A2(n8797), .ZN(n6063) );
  NAND2_X1 U5451 ( .A1(n8803), .A2(n8805), .ZN(n8802) );
  INV_X1 U5452 ( .A(n4626), .ZN(n7522) );
  INV_X1 U5453 ( .A(n6614), .ZN(n4623) );
  NAND2_X1 U5454 ( .A1(n7522), .A2(n4621), .ZN(n4624) );
  OR2_X1 U5455 ( .A1(n6084), .A2(n6083), .ZN(n6129) );
  AND2_X1 U5456 ( .A1(n6145), .A2(n9490), .ZN(n8848) );
  NAND2_X1 U5457 ( .A1(n4620), .A2(n8724), .ZN(n4619) );
  INV_X1 U5458 ( .A(n8725), .ZN(n4620) );
  NAND2_X1 U5459 ( .A1(n8725), .A2(n5899), .ZN(n4618) );
  AND2_X1 U5460 ( .A1(n6405), .A2(n6404), .ZN(n6503) );
  AOI21_X1 U5461 ( .B1(n9545), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9540), .ZN(
        n9554) );
  XNOR2_X1 U5462 ( .A(n8910), .B(n8924), .ZN(n9567) );
  NOR2_X1 U5463 ( .A1(n8913), .A2(n9577), .ZN(n9590) );
  XNOR2_X1 U5464 ( .A(n9242), .B(n9027), .ZN(n9002) );
  NOR2_X1 U5465 ( .A1(n4758), .A2(n4754), .ZN(n4753) );
  INV_X1 U5466 ( .A(n8974), .ZN(n4754) );
  OR2_X1 U5467 ( .A1(n9041), .A2(n9000), .ZN(n4650) );
  INV_X1 U5468 ( .A(n4650), .ZN(n9026) );
  NAND2_X1 U5469 ( .A1(n4367), .A2(n4365), .ZN(n9043) );
  NAND2_X1 U5470 ( .A1(n8997), .A2(n4366), .ZN(n4365) );
  INV_X1 U5471 ( .A(n4369), .ZN(n4366) );
  NAND2_X1 U5472 ( .A1(n9040), .A2(n9051), .ZN(n9035) );
  NAND2_X1 U5473 ( .A1(n4661), .A2(n7728), .ZN(n4660) );
  INV_X1 U5474 ( .A(n4663), .ZN(n4661) );
  NAND2_X1 U5475 ( .A1(n8994), .A2(n4662), .ZN(n4371) );
  AND2_X1 U5476 ( .A1(n9055), .A2(n9072), .ZN(n9051) );
  NAND2_X1 U5477 ( .A1(n8997), .A2(n7621), .ZN(n9056) );
  NAND2_X1 U5478 ( .A1(n7728), .A2(n7731), .ZN(n9065) );
  NAND2_X1 U5479 ( .A1(n9083), .A2(n8995), .ZN(n9066) );
  NOR2_X1 U5480 ( .A1(n9065), .A2(n7653), .ZN(n4663) );
  NAND2_X1 U5481 ( .A1(n8994), .A2(n8993), .ZN(n9083) );
  NAND2_X1 U5482 ( .A1(n9104), .A2(n9105), .ZN(n9111) );
  AND2_X1 U5483 ( .A1(n8992), .A2(n7622), .ZN(n9105) );
  NOR2_X1 U5484 ( .A1(n9167), .A2(n4554), .ZN(n9117) );
  INV_X1 U5485 ( .A(n4556), .ZN(n4554) );
  AND2_X1 U5486 ( .A1(n7710), .A2(n8984), .ZN(n9184) );
  AND2_X1 U5487 ( .A1(n9226), .A2(n4544), .ZN(n9195) );
  AND2_X1 U5488 ( .A1(n4283), .A2(n9193), .ZN(n4544) );
  AND2_X1 U5489 ( .A1(n8977), .A2(n9182), .ZN(n9206) );
  OR2_X1 U5490 ( .A1(n5905), .A2(n5904), .ZN(n5920) );
  NAND2_X1 U5491 ( .A1(n4378), .A2(n4376), .ZN(n8981) );
  AND4_X1 U5492 ( .A1(n5940), .A2(n5939), .A3(n5938), .A4(n5937), .ZN(n9190)
         );
  AOI21_X1 U5493 ( .B1(n4765), .B2(n4307), .A(n4762), .ZN(n4761) );
  NOR2_X1 U5494 ( .A1(n9232), .A2(n8780), .ZN(n4762) );
  NAND2_X1 U5495 ( .A1(n9226), .A2(n9232), .ZN(n9227) );
  NAND2_X1 U5496 ( .A1(n4378), .A2(n7700), .ZN(n9219) );
  NOR2_X1 U5497 ( .A1(n9406), .A2(n9322), .ZN(n9226) );
  OR2_X1 U5498 ( .A1(n9405), .A2(n8822), .ZN(n9406) );
  INV_X1 U5499 ( .A(n4357), .ZN(n4356) );
  AOI21_X1 U5500 ( .B1(n4357), .B2(n4359), .A(n4355), .ZN(n4354) );
  NAND2_X1 U5501 ( .A1(n4353), .A2(n4357), .ZN(n9410) );
  NAND2_X1 U5502 ( .A1(n9430), .A2(n4360), .ZN(n4353) );
  AND2_X1 U5503 ( .A1(n5857), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5876) );
  NOR2_X1 U5504 ( .A1(n5842), .A2(n5841), .ZN(n5857) );
  OR2_X1 U5505 ( .A1(n7330), .A2(n7329), .ZN(n9427) );
  NOR2_X1 U5506 ( .A1(n7140), .A2(n4551), .ZN(n9444) );
  NAND2_X1 U5507 ( .A1(n7119), .A2(n4382), .ZN(n7185) );
  NOR2_X1 U5508 ( .A1(n7678), .A2(n4383), .ZN(n4382) );
  INV_X1 U5509 ( .A(n7661), .ZN(n4383) );
  NOR2_X1 U5510 ( .A1(n7140), .A2(n7344), .ZN(n7192) );
  NAND2_X1 U5511 ( .A1(n7119), .A2(n7661), .ZN(n7131) );
  NAND2_X1 U5512 ( .A1(n6949), .A2(n4518), .ZN(n6954) );
  NAND2_X1 U5513 ( .A1(n7842), .A2(n7659), .ZN(n7831) );
  NOR2_X1 U5514 ( .A1(n7836), .A2(n7824), .ZN(n7823) );
  AND3_X1 U5515 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U5516 ( .A1(n4546), .A2(n4547), .ZN(n6866) );
  NAND2_X1 U5517 ( .A1(n7780), .A2(n7579), .ZN(n6859) );
  OR2_X1 U5518 ( .A1(n7562), .A2(n6229), .ZN(n5674) );
  NAND2_X1 U5519 ( .A1(n7625), .A2(n6782), .ZN(n4381) );
  INV_X1 U5520 ( .A(n6785), .ZN(n7626) );
  NAND2_X1 U5521 ( .A1(n7778), .A2(n7777), .ZN(n6785) );
  NAND2_X1 U5522 ( .A1(n6586), .A2(n7773), .ZN(n6980) );
  AND2_X1 U5523 ( .A1(n6715), .A2(n6615), .ZN(n6782) );
  NAND2_X1 U5524 ( .A1(n7891), .A2(n5779), .ZN(n4399) );
  NAND2_X1 U5525 ( .A1(n7564), .A2(n7563), .ZN(n9252) );
  NAND2_X1 U5526 ( .A1(n6593), .A2(n5779), .ZN(n4667) );
  NAND2_X1 U5527 ( .A1(n5919), .A2(n5918), .ZN(n9312) );
  INV_X1 U5528 ( .A(n9681), .ZN(n9324) );
  NAND2_X1 U5529 ( .A1(n7658), .A2(n7657), .ZN(n7838) );
  INV_X1 U5530 ( .A(n9679), .ZN(n9661) );
  INV_X1 U5531 ( .A(n6715), .ZN(n6586) );
  XNOR2_X1 U5532 ( .A(n7518), .B(n5351), .ZN(n8113) );
  XNOR2_X1 U5533 ( .A(n5654), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U5534 ( .A1(n5657), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U5535 ( .A1(n5631), .A2(n5660), .ZN(n5652) );
  OAI21_X1 U5536 ( .B1(n5255), .B2(n5254), .A(n4942), .ZN(n5267) );
  AND2_X1 U5537 ( .A1(n4946), .A2(n4945), .ZN(n5266) );
  NAND2_X1 U5538 ( .A1(n4390), .A2(n4392), .ZN(n5218) );
  NAND2_X1 U5539 ( .A1(n4391), .A2(n4394), .ZN(n4390) );
  INV_X1 U5540 ( .A(n5186), .ZN(n4391) );
  XNOR2_X1 U5541 ( .A(n5186), .B(n5185), .ZN(n6593) );
  NAND2_X1 U5542 ( .A1(n5886), .A2(n5644), .ZN(n5916) );
  NAND2_X1 U5543 ( .A1(n4899), .A2(n4898), .ZN(n5152) );
  INV_X1 U5544 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4584) );
  NAND2_X1 U5545 ( .A1(n4659), .A2(n4881), .ZN(n5112) );
  NAND2_X1 U5546 ( .A1(n5100), .A2(n4788), .ZN(n4659) );
  OR2_X1 U5547 ( .A1(n5818), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5836) );
  XNOR2_X1 U5548 ( .A(n5100), .B(n4788), .ZN(n6251) );
  INV_X1 U5549 ( .A(n4413), .ZN(n5088) );
  AOI21_X1 U5550 ( .B1(n4412), .B2(n4417), .A(n4416), .ZN(n4413) );
  NAND2_X1 U5551 ( .A1(n4412), .A2(n4863), .ZN(n5079) );
  XNOR2_X1 U5552 ( .A(n4857), .B(SI_6_), .ZN(n5048) );
  AND2_X1 U5553 ( .A1(n5670), .A2(n5621), .ZN(n5729) );
  INV_X1 U5554 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5622) );
  OAI21_X1 U5555 ( .B1(n4673), .B2(n4670), .A(n4668), .ZN(n6758) );
  AOI21_X1 U5556 ( .B1(n4671), .B2(n6628), .A(n4669), .ZN(n4668) );
  INV_X1 U5557 ( .A(n4671), .ZN(n4670) );
  INV_X1 U5558 ( .A(n5494), .ZN(n4669) );
  AND2_X1 U5559 ( .A1(n4705), .A2(n5589), .ZN(n8146) );
  NAND2_X1 U5560 ( .A1(n4697), .A2(n4694), .ZN(n7413) );
  INV_X1 U5561 ( .A(n4696), .ZN(n4694) );
  NAND2_X1 U5562 ( .A1(n5271), .A2(n5270), .ZN(n8626) );
  OAI22_X1 U5563 ( .A1(n6441), .A2(n6442), .B1(n5474), .B2(n5473), .ZN(n6451)
         );
  OR2_X1 U5564 ( .A1(n5598), .A2(n5597), .ZN(n5599) );
  AND2_X1 U5565 ( .A1(n5472), .A2(n5470), .ZN(n6430) );
  NAND2_X1 U5566 ( .A1(n6430), .A2(n6429), .ZN(n6428) );
  NAND2_X1 U5567 ( .A1(n8195), .A2(n5545), .ZN(n8205) );
  NAND2_X1 U5568 ( .A1(n4951), .A2(n4950), .ZN(n8620) );
  NAND2_X1 U5569 ( .A1(n6451), .A2(n6450), .ZN(n4685) );
  NAND2_X1 U5570 ( .A1(n7202), .A2(n5525), .ZN(n7217) );
  NAND2_X1 U5571 ( .A1(n5142), .A2(n5141), .ZN(n7250) );
  AND2_X1 U5572 ( .A1(n5607), .A2(n8107), .ZN(n8281) );
  NOR2_X1 U5573 ( .A1(n8204), .A2(n4687), .ZN(n4686) );
  AND2_X1 U5574 ( .A1(n4672), .A2(n4313), .ZN(n6724) );
  NAND2_X1 U5575 ( .A1(n4673), .A2(n5488), .ZN(n4672) );
  NAND2_X1 U5576 ( .A1(n5586), .A2(n5585), .ZN(n8261) );
  AND2_X1 U5577 ( .A1(n5327), .A2(n5310), .ZN(n8415) );
  NAND2_X1 U5578 ( .A1(n5175), .A2(n5174), .ZN(n8287) );
  INV_X1 U5579 ( .A(n6280), .ZN(n9706) );
  NOR2_X1 U5580 ( .A1(n6371), .A2(n4531), .ZN(n6370) );
  NAND2_X1 U5581 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n4531) );
  AND2_X1 U5582 ( .A1(n4536), .A2(n4535), .ZN(n6325) );
  NAND2_X1 U5583 ( .A1(n6326), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4535) );
  INV_X1 U5584 ( .A(n4534), .ZN(n6455) );
  NOR2_X1 U5585 ( .A1(n9952), .A2(n4538), .ZN(n6458) );
  AND2_X1 U5586 ( .A1(n6459), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4538) );
  NOR2_X1 U5587 ( .A1(n6458), .A2(n6457), .ZN(n6605) );
  NAND2_X1 U5588 ( .A1(n7437), .A2(n7438), .ZN(n7441) );
  INV_X1 U5589 ( .A(n4525), .ZN(n8318) );
  AND2_X1 U5590 ( .A1(n4525), .A2(n4524), .ZN(n8321) );
  NAND2_X1 U5591 ( .A1(n8322), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4524) );
  NAND2_X1 U5592 ( .A1(n8347), .A2(n8348), .ZN(n8349) );
  AND2_X1 U5593 ( .A1(n6289), .A2(n6285), .ZN(n9697) );
  OR2_X1 U5594 ( .A1(n5341), .A2(n5340), .ZN(n7881) );
  INV_X1 U5595 ( .A(n5399), .ZN(n5400) );
  AOI22_X1 U5596 ( .A1(n8292), .A2(n8228), .B1(n8366), .B2(n8291), .ZN(n5399)
         );
  AOI21_X1 U5597 ( .B1(n8390), .B2(n8040), .A(n8092), .ZN(n5450) );
  AND2_X1 U5598 ( .A1(n5222), .A2(n5362), .ZN(n8417) );
  NAND2_X1 U5599 ( .A1(n5308), .A2(n5307), .ZN(n8611) );
  NAND2_X1 U5600 ( .A1(n5290), .A2(n5289), .ZN(n8616) );
  NAND2_X1 U5601 ( .A1(n8624), .A2(n4780), .ZN(n8434) );
  NAND2_X1 U5602 ( .A1(n8453), .A2(n8452), .ZN(n8624) );
  NAND2_X1 U5603 ( .A1(n4583), .A2(n4279), .ZN(n8542) );
  AND2_X1 U5604 ( .A1(n4583), .A2(n4582), .ZN(n8543) );
  NAND2_X1 U5605 ( .A1(n4733), .A2(n7967), .ZN(n7243) );
  NAND2_X1 U5606 ( .A1(n4570), .A2(n5139), .ZN(n7249) );
  NAND2_X1 U5607 ( .A1(n5127), .A2(n5126), .ZN(n7078) );
  NAND2_X1 U5608 ( .A1(n6882), .A2(n7946), .ZN(n6734) );
  NAND2_X1 U5609 ( .A1(n6640), .A2(n5024), .ZN(n6812) );
  INV_X1 U5610 ( .A(n8370), .ZN(n8572) );
  AND2_X1 U5611 ( .A1(n8567), .A2(n6700), .ZN(n8582) );
  AND2_X1 U5612 ( .A1(n8567), .A2(n6702), .ZN(n8581) );
  NAND2_X1 U5613 ( .A1(n7901), .A2(n7900), .ZN(n8679) );
  NAND2_X1 U5614 ( .A1(n7897), .A2(n7898), .ZN(n7901) );
  AND2_X1 U5615 ( .A1(n5247), .A2(n5246), .ZN(n8696) );
  INV_X1 U5616 ( .A(n8517), .ZN(n8703) );
  NAND2_X1 U5617 ( .A1(n4965), .A2(n4964), .ZN(n8715) );
  INV_X1 U5618 ( .A(n8287), .ZN(n7495) );
  INV_X1 U5619 ( .A(n8417), .ZN(n8357) );
  INV_X1 U5620 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6238) );
  INV_X1 U5621 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9822) );
  NAND2_X1 U5622 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4532) );
  AND4_X1 U5623 ( .A1(n5800), .A2(n5799), .A3(n5798), .A4(n5797), .ZN(n7231)
         );
  AND2_X1 U5624 ( .A1(n6670), .A2(n6149), .ZN(n9038) );
  AND4_X1 U5625 ( .A1(n6030), .A2(n6029), .A3(n6028), .A4(n6027), .ZN(n9108)
         );
  OR2_X1 U5626 ( .A1(n8133), .A2(n8132), .ZN(n8120) );
  NAND2_X1 U5627 ( .A1(n7558), .A2(n7557), .ZN(n9247) );
  NAND2_X1 U5628 ( .A1(n4626), .A2(n4625), .ZN(n6613) );
  NOR2_X1 U5629 ( .A1(n6161), .A2(n4589), .ZN(n4588) );
  INV_X1 U5630 ( .A(n8794), .ZN(n4589) );
  OAI22_X1 U5631 ( .A1(n6161), .A2(n4592), .B1(n6162), .B2(n4591), .ZN(n4590)
         );
  NOR2_X1 U5632 ( .A1(n8794), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U5633 ( .A1(n6830), .A2(n5740), .ZN(n6911) );
  AND4_X1 U5634 ( .A1(n5924), .A2(n5923), .A3(n5922), .A4(n5921), .ZN(n9220)
         );
  AND2_X1 U5635 ( .A1(n6051), .A2(n6050), .ZN(n8966) );
  AND4_X1 U5636 ( .A1(n5827), .A2(n5826), .A3(n5825), .A4(n5824), .ZN(n9434)
         );
  INV_X1 U5637 ( .A(n8850), .ZN(n8860) );
  INV_X1 U5638 ( .A(n4346), .ZN(n6538) );
  NAND2_X1 U5639 ( .A1(n8763), .A2(n8761), .ZN(n5872) );
  OAI21_X1 U5640 ( .B1(n7299), .B2(n5835), .A(n4601), .ZN(n8839) );
  INV_X1 U5641 ( .A(n4603), .ZN(n4601) );
  AND4_X1 U5642 ( .A1(n5862), .A2(n5861), .A3(n5860), .A4(n5859), .ZN(n9436)
         );
  NAND2_X1 U5643 ( .A1(n4622), .A2(n4624), .ZN(n7523) );
  AOI21_X1 U5644 ( .B1(n6830), .B2(n4275), .A(n4277), .ZN(n7059) );
  INV_X1 U5645 ( .A(n8848), .ZN(n8864) );
  NAND2_X1 U5646 ( .A1(n4614), .A2(n4618), .ZN(n8859) );
  NAND2_X1 U5647 ( .A1(n8727), .A2(n4619), .ZN(n4614) );
  AOI21_X1 U5648 ( .B1(n4486), .B2(n7770), .A(n4484), .ZN(n4483) );
  AND4_X1 U5649 ( .A1(n6675), .A2(n6674), .A3(n6673), .A4(n6672), .ZN(n9044)
         );
  AND4_X1 U5650 ( .A1(n6068), .A2(n6067), .A3(n6066), .A4(n6065), .ZN(n9088)
         );
  INV_X1 U5651 ( .A(n7840), .ZN(n8880) );
  INV_X1 U5652 ( .A(n7839), .ZN(n8882) );
  INV_X1 U5653 ( .A(n6777), .ZN(n8883) );
  AOI21_X1 U5654 ( .B1(n9521), .B2(n6385), .A(n6386), .ZN(n6388) );
  NOR2_X1 U5655 ( .A1(n6488), .A2(n6489), .ZN(n6487) );
  AND2_X1 U5656 ( .A1(n6490), .A2(n6204), .ZN(n8901) );
  AND2_X1 U5657 ( .A1(n6500), .A2(n6499), .ZN(n6502) );
  AOI21_X1 U5658 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6504), .A(n6503), .ZN(
        n6507) );
  AOI21_X1 U5659 ( .B1(n7897), .B2(n5779), .A(n7542), .ZN(n8949) );
  XNOR2_X1 U5660 ( .A(n9010), .B(n4398), .ZN(n9452) );
  AOI21_X1 U5661 ( .B1(n4385), .B2(n4384), .A(n9029), .ZN(n9250) );
  NAND2_X1 U5662 ( .A1(n4787), .A2(n9028), .ZN(n9029) );
  NAND2_X1 U5663 ( .A1(n9026), .A2(n9025), .ZN(n4385) );
  AOI21_X1 U5664 ( .B1(n4650), .B2(n7740), .A(n9433), .ZN(n4384) );
  OAI21_X1 U5665 ( .B1(n9019), .B2(n9025), .A(n9018), .ZN(n9251) );
  AND2_X1 U5666 ( .A1(n4759), .A2(n4294), .ZN(n9019) );
  NAND2_X1 U5667 ( .A1(n4759), .A2(n4757), .ZN(n9018) );
  NAND2_X1 U5668 ( .A1(n9034), .A2(n9042), .ZN(n4759) );
  NAND2_X1 U5669 ( .A1(n6060), .A2(n6059), .ZN(n9069) );
  INV_X1 U5670 ( .A(n8966), .ZN(n8967) );
  AND2_X1 U5671 ( .A1(n6033), .A2(n6032), .ZN(n9103) );
  NAND2_X1 U5672 ( .A1(n9134), .A2(n8989), .ZN(n9122) );
  OAI21_X1 U5673 ( .B1(n9162), .B2(n4745), .A(n4743), .ZN(n9129) );
  NAND2_X1 U5674 ( .A1(n6006), .A2(n6005), .ZN(n9140) );
  NAND2_X1 U5675 ( .A1(n8986), .A2(n8985), .ZN(n9151) );
  OAI21_X1 U5676 ( .B1(n9404), .B2(n4280), .A(n4765), .ZN(n9222) );
  NAND2_X1 U5677 ( .A1(n9404), .A2(n4770), .ZN(n4768) );
  NAND2_X1 U5678 ( .A1(n4362), .A2(n7590), .ZN(n7456) );
  NAND2_X1 U5679 ( .A1(n4363), .A2(n7686), .ZN(n4362) );
  NAND2_X1 U5680 ( .A1(n5856), .A2(n5855), .ZN(n8771) );
  NAND2_X1 U5681 ( .A1(n7116), .A2(n7115), .ZN(n7135) );
  OR2_X1 U5682 ( .A1(n9456), .A2(n6678), .ZN(n9419) );
  INV_X1 U5683 ( .A(n9419), .ZN(n9439) );
  OAI211_X1 U5684 ( .C1(n6173), .C2(n6225), .A(n5748), .B(n5747), .ZN(n7852)
         );
  NAND2_X1 U5685 ( .A1(n6959), .A2(n6958), .ZN(n7849) );
  INV_X1 U5686 ( .A(n9418), .ZN(n9441) );
  INV_X2 U5687 ( .A(n9693), .ZN(n9696) );
  INV_X1 U5688 ( .A(n9241), .ZN(n4665) );
  INV_X2 U5689 ( .A(n9683), .ZN(n9685) );
  XNOR2_X1 U5690 ( .A(n5348), .B(n5347), .ZN(n7555) );
  NAND2_X1 U5691 ( .A1(n5337), .A2(n5336), .ZN(n5348) );
  INV_X1 U5692 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6241) );
  OR2_X1 U5693 ( .A1(n5805), .A2(n5804), .ZN(n6239) );
  INV_X1 U5694 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9837) );
  INV_X1 U5695 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5759) );
  NOR2_X1 U5696 ( .A1(n9397), .A2(n9980), .ZN(n9798) );
  INV_X1 U5697 ( .A(n4530), .ZN(n6337) );
  INV_X1 U5698 ( .A(n4528), .ZN(n6352) );
  INV_X1 U5699 ( .A(n4536), .ZN(n6322) );
  NOR2_X1 U5700 ( .A1(n5437), .A2(n4334), .ZN(n5438) );
  NOR2_X1 U5701 ( .A1(n9770), .A2(n5436), .ZN(n5437) );
  OAI21_X1 U5702 ( .B1(n9055), .B2(n8813), .A(n6156), .ZN(n6157) );
  MUX2_X1 U5703 ( .A(n8941), .B(n8940), .S(n9157), .Z(n8942) );
  AOI21_X1 U5704 ( .B1(n9475), .B2(n9685), .A(n4342), .ZN(P1_U3521) );
  AND2_X1 U5705 ( .A1(n4679), .A2(n4676), .ZN(n4276) );
  NAND2_X1 U5706 ( .A1(n4396), .A2(n4922), .ZN(n4395) );
  NAND2_X1 U5707 ( .A1(n9001), .A2(n7742), .ZN(n9025) );
  AND2_X1 U5708 ( .A1(n6909), .A2(n6908), .ZN(n4277) );
  INV_X1 U5709 ( .A(n4268), .ZN(n5719) );
  AND2_X1 U5710 ( .A1(n4392), .A2(n4389), .ZN(n4278) );
  AND2_X1 U5711 ( .A1(n8544), .A2(n4582), .ZN(n4279) );
  XNOR2_X1 U5712 ( .A(n8626), .B(n8243), .ZN(n8452) );
  INV_X1 U5713 ( .A(n8452), .ZN(n4574) );
  OR2_X1 U5714 ( .A1(n7502), .A2(n4767), .ZN(n4280) );
  NAND2_X1 U5715 ( .A1(n4811), .A2(n4810), .ZN(n5032) );
  AND2_X1 U5716 ( .A1(n4482), .A2(n4481), .ZN(n4281) );
  INV_X1 U5717 ( .A(n4758), .ZN(n4757) );
  NAND2_X1 U5718 ( .A1(n9025), .A2(n4294), .ZN(n4758) );
  INV_X1 U5719 ( .A(n8092), .ZN(n4722) );
  NAND2_X1 U5720 ( .A1(n8041), .A2(n8037), .ZN(n8092) );
  OR2_X1 U5721 ( .A1(n9257), .A2(n9073), .ZN(n8997) );
  NAND2_X1 U5722 ( .A1(n8999), .A2(n7738), .ZN(n9042) );
  NAND2_X1 U5723 ( .A1(n7914), .A2(n6814), .ZN(n8070) );
  NAND2_X1 U5724 ( .A1(n4399), .A2(n7543), .ZN(n9454) );
  INV_X1 U5725 ( .A(n9454), .ZN(n4398) );
  OR2_X1 U5726 ( .A1(n4791), .A2(n7808), .ZN(n4282) );
  AND2_X1 U5727 ( .A1(n4545), .A2(n9214), .ZN(n4283) );
  AND2_X1 U5728 ( .A1(n6216), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4284) );
  AND2_X1 U5729 ( .A1(n9469), .A2(n4550), .ZN(n4285) );
  AND2_X1 U5730 ( .A1(n5386), .A2(n7998), .ZN(n4286) );
  INV_X1 U5731 ( .A(n4749), .ZN(n4748) );
  NOR2_X1 U5732 ( .A1(n9173), .A2(n9153), .ZN(n4749) );
  AND2_X1 U5733 ( .A1(n7117), .A2(n7115), .ZN(n4287) );
  NOR2_X1 U5734 ( .A1(n7624), .A2(n4377), .ZN(n4376) );
  NAND2_X1 U5735 ( .A1(n8417), .A2(n7910), .ZN(n8045) );
  OR2_X1 U5736 ( .A1(n9167), .A2(n4557), .ZN(n4288) );
  INV_X1 U5737 ( .A(n7640), .ZN(n4380) );
  INV_X1 U5738 ( .A(n4395), .ZN(n4394) );
  INV_X1 U5739 ( .A(n8985), .ZN(n4636) );
  NAND2_X1 U5740 ( .A1(n4771), .A2(n4784), .ZN(n5853) );
  AND2_X1 U5741 ( .A1(n9278), .A2(n9108), .ZN(n8990) );
  NAND2_X1 U5742 ( .A1(n4381), .A2(n6784), .ZN(n6974) );
  AND4_X1 U5743 ( .A1(n6093), .A2(n6092), .A3(n6091), .A4(n6090), .ZN(n9073)
         );
  INV_X1 U5744 ( .A(n9073), .ZN(n8973) );
  OR2_X1 U5745 ( .A1(n8620), .A2(n8157), .ZN(n5390) );
  OR2_X1 U5746 ( .A1(n5170), .A2(n4642), .ZN(n4289) );
  INV_X1 U5747 ( .A(n8590), .ZN(n4979) );
  XNOR2_X1 U5748 ( .A(n5035), .B(n5034), .ZN(n6226) );
  XNOR2_X1 U5749 ( .A(n7541), .B(n7540), .ZN(n7897) );
  NAND2_X1 U5750 ( .A1(n5552), .A2(n5551), .ZN(n4290) );
  AND2_X1 U5751 ( .A1(n8413), .A2(n4441), .ZN(n4291) );
  INV_X1 U5752 ( .A(n4981), .ZN(n5398) );
  AND4_X1 U5753 ( .A1(n5713), .A2(n5712), .A3(n5711), .A4(n5710), .ZN(n6777)
         );
  NAND2_X1 U5754 ( .A1(n5839), .A2(n5838), .ZN(n9442) );
  INV_X1 U5755 ( .A(n4683), .ZN(n4682) );
  NAND2_X1 U5756 ( .A1(n8164), .A2(n4290), .ZN(n4683) );
  AND2_X1 U5757 ( .A1(n6023), .A2(n6022), .ZN(n9120) );
  INV_X1 U5758 ( .A(n9120), .ZN(n9278) );
  OAI21_X1 U5759 ( .B1(n4749), .B2(n4746), .A(n4747), .ZN(n4745) );
  NOR2_X1 U5760 ( .A1(n8311), .A2(n6888), .ZN(n4292) );
  OR2_X1 U5761 ( .A1(n6909), .A2(n6908), .ZN(n4293) );
  XNOR2_X1 U5762 ( .A(n8606), .B(n8293), .ZN(n8391) );
  NAND2_X1 U5763 ( .A1(n8802), .A2(n8804), .ZN(n8754) );
  OR2_X1 U5764 ( .A1(n9252), .A2(n8975), .ZN(n4294) );
  AND2_X1 U5765 ( .A1(n5189), .A2(n4707), .ZN(n4295) );
  OR2_X1 U5766 ( .A1(n9069), .A2(n9088), .ZN(n7728) );
  AND2_X1 U5767 ( .A1(n9358), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4296) );
  OR2_X1 U5768 ( .A1(n9315), .A2(n8871), .ZN(n4297) );
  AND2_X1 U5769 ( .A1(n4404), .A2(n4640), .ZN(n4298) );
  NOR2_X1 U5770 ( .A1(n9295), .A2(n9187), .ZN(n4299) );
  INV_X1 U5771 ( .A(n7962), .ZN(n4464) );
  NAND4_X1 U5772 ( .A1(n5686), .A2(n5685), .A3(n5684), .A4(n5683), .ZN(n6579)
         );
  NAND2_X1 U5773 ( .A1(n5903), .A2(n5902), .ZN(n9315) );
  NAND2_X1 U5774 ( .A1(n5985), .A2(n5984), .ZN(n9290) );
  NAND2_X1 U5775 ( .A1(n5932), .A2(n5645), .ZN(n5679) );
  NAND3_X1 U5776 ( .A1(n4715), .A2(n4811), .A3(n4819), .ZN(n4300) );
  NAND2_X1 U5777 ( .A1(n6283), .A2(n6216), .ZN(n5050) );
  INV_X1 U5778 ( .A(n5050), .ZN(n4450) );
  NOR2_X1 U5779 ( .A1(n8856), .A2(n8857), .ZN(n4301) );
  NAND2_X1 U5780 ( .A1(n5207), .A2(n5206), .ZN(n8535) );
  OR2_X1 U5781 ( .A1(n6283), .A2(n6319), .ZN(n4302) );
  AND2_X1 U5782 ( .A1(n4523), .A2(n7657), .ZN(n4303) );
  NAND2_X1 U5783 ( .A1(n5385), .A2(n7998), .ZN(n8496) );
  NAND2_X1 U5784 ( .A1(n6947), .A2(n7583), .ZN(n7658) );
  INV_X1 U5785 ( .A(n5631), .ZN(n5659) );
  AND2_X1 U5786 ( .A1(n4729), .A2(n5390), .ZN(n4304) );
  AND2_X1 U5787 ( .A1(n5850), .A2(n5852), .ZN(n4305) );
  AND2_X1 U5788 ( .A1(n4782), .A2(n5087), .ZN(n4306) );
  INV_X1 U5789 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5415) );
  INV_X1 U5790 ( .A(n8262), .ZN(n4704) );
  INV_X1 U5791 ( .A(n8606), .ZN(n8403) );
  NAND2_X1 U5792 ( .A1(n5325), .A2(n5324), .ZN(n8606) );
  AND2_X1 U5793 ( .A1(n4297), .A2(n4280), .ZN(n4307) );
  AND2_X1 U5794 ( .A1(n8413), .A2(n4439), .ZN(n4308) );
  AND2_X1 U5795 ( .A1(n8624), .A2(n4576), .ZN(n4309) );
  INV_X1 U5796 ( .A(n4597), .ZN(n4596) );
  OAI21_X1 U5797 ( .B1(n4275), .B2(n4277), .A(n7060), .ZN(n4597) );
  AND2_X1 U5798 ( .A1(n4371), .A2(n4369), .ZN(n4310) );
  INV_X1 U5799 ( .A(n4868), .ZN(n4416) );
  NAND2_X1 U5800 ( .A1(n4865), .A2(n4864), .ZN(n4868) );
  INV_X1 U5801 ( .A(n8084), .ZN(n4458) );
  AND2_X1 U5802 ( .A1(n5201), .A2(n8253), .ZN(n4311) );
  NOR2_X1 U5803 ( .A1(n8961), .A2(n9166), .ZN(n4312) );
  INV_X1 U5804 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U5805 ( .A1(n5487), .A2(n5486), .ZN(n4313) );
  AND2_X1 U5806 ( .A1(n7976), .A2(n7975), .ZN(n7272) );
  INV_X1 U5807 ( .A(n9411), .ZN(n4355) );
  NAND2_X1 U5808 ( .A1(n4702), .A2(n4701), .ZN(n8144) );
  INV_X1 U5809 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4707) );
  NAND2_X1 U5810 ( .A1(n7709), .A2(n7710), .ZN(n4314) );
  AND2_X1 U5811 ( .A1(n7730), .A2(n4487), .ZN(n4315) );
  AND2_X1 U5812 ( .A1(n4350), .A2(n8991), .ZN(n4316) );
  AND2_X1 U5813 ( .A1(n5562), .A2(n5561), .ZN(n4317) );
  AND2_X1 U5814 ( .A1(n8440), .A2(n8157), .ZN(n4318) );
  OR2_X1 U5815 ( .A1(n8441), .A2(n8023), .ZN(n4319) );
  INV_X1 U5816 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6215) );
  AND2_X1 U5817 ( .A1(n4884), .A2(SI_11_), .ZN(n4320) );
  INV_X1 U5818 ( .A(n8435), .ZN(n8443) );
  AND2_X1 U5819 ( .A1(n5390), .A2(n8021), .ZN(n8435) );
  NOR2_X1 U5820 ( .A1(n9024), .A2(n9044), .ZN(n4321) );
  INV_X1 U5821 ( .A(n9055), .ZN(n9257) );
  AND2_X1 U5822 ( .A1(n6086), .A2(n6085), .ZN(n9055) );
  OR2_X1 U5823 ( .A1(n9247), .A2(n9044), .ZN(n9001) );
  INV_X1 U5824 ( .A(n9442), .ZN(n9469) );
  INV_X1 U5825 ( .A(n4745), .ZN(n4744) );
  INV_X1 U5826 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4822) );
  OR2_X1 U5827 ( .A1(n8979), .A2(n8978), .ZN(n4322) );
  AND2_X1 U5828 ( .A1(n8983), .A2(n4376), .ZN(n4323) );
  AND2_X1 U5829 ( .A1(n9083), .A2(n4663), .ZN(n4324) );
  AND2_X1 U5830 ( .A1(n7986), .A2(n7985), .ZN(n7983) );
  AND2_X1 U5831 ( .A1(n4547), .A2(n6957), .ZN(n4325) );
  AND2_X1 U5832 ( .A1(n7971), .A2(n7273), .ZN(n8084) );
  AOI21_X1 U5833 ( .B1(n7740), .B2(n9000), .A(n4649), .ZN(n4648) );
  AND2_X1 U5834 ( .A1(n4861), .A2(n4868), .ZN(n4326) );
  AND2_X1 U5835 ( .A1(n5482), .A2(n5479), .ZN(n4327) );
  OR2_X1 U5836 ( .A1(n6239), .A2(n6187), .ZN(n4328) );
  AND2_X1 U5837 ( .A1(n4458), .A2(n5139), .ZN(n4329) );
  NAND2_X1 U5838 ( .A1(n9737), .A2(n8312), .ZN(n7936) );
  INV_X1 U5839 ( .A(n7567), .ZN(n9193) );
  NAND2_X1 U5840 ( .A1(n5952), .A2(n5951), .ZN(n7567) );
  INV_X1 U5841 ( .A(n8424), .ZN(n8422) );
  AND2_X1 U5842 ( .A1(n8408), .A2(n8028), .ZN(n8424) );
  OR2_X1 U5843 ( .A1(n8044), .A2(n8149), .ZN(n8041) );
  NAND2_X1 U5844 ( .A1(n5707), .A2(n5706), .ZN(n4330) );
  NOR2_X1 U5845 ( .A1(n8243), .A2(n6567), .ZN(n4331) );
  AND2_X1 U5846 ( .A1(n9226), .A2(n4283), .ZN(n4332) );
  INV_X1 U5847 ( .A(n4700), .ZN(n8190) );
  NAND2_X1 U5848 ( .A1(n5339), .A2(n5338), .ZN(n8044) );
  NOR2_X1 U5849 ( .A1(n9167), .A2(n9290), .ZN(n4333) );
  INV_X1 U5850 ( .A(n4996), .ZN(n5011) );
  NOR2_X1 U5851 ( .A1(n4440), .A2(n8667), .ZN(n4334) );
  INV_X1 U5852 ( .A(n7722), .ZN(n4503) );
  NAND2_X1 U5853 ( .A1(n5353), .A2(n5352), .ZN(n7885) );
  INV_X1 U5854 ( .A(n7885), .ZN(n4440) );
  NAND2_X1 U5855 ( .A1(n4768), .A2(n4769), .ZN(n7503) );
  INV_X1 U5856 ( .A(n7700), .ZN(n4377) );
  NAND2_X1 U5857 ( .A1(n4667), .A2(n5934), .ZN(n9307) );
  INV_X1 U5858 ( .A(n9307), .ZN(n9214) );
  INV_X1 U5859 ( .A(n8989), .ZN(n4351) );
  AND2_X1 U5860 ( .A1(n4697), .A2(n4695), .ZN(n4335) );
  INV_X1 U5861 ( .A(n4448), .ZN(n8515) );
  NOR2_X1 U5862 ( .A1(n8551), .A2(n4445), .ZN(n4448) );
  NOR2_X1 U5863 ( .A1(n9167), .A2(n4555), .ZN(n4553) );
  NAND2_X1 U5864 ( .A1(n9140), .A2(n9124), .ZN(n4336) );
  AND2_X1 U5865 ( .A1(n4923), .A2(SI_18_), .ZN(n4337) );
  INV_X1 U5866 ( .A(n4760), .ZN(n4756) );
  NAND2_X1 U5867 ( .A1(n9257), .A2(n8973), .ZN(n4760) );
  OR2_X1 U5868 ( .A1(n6162), .A2(n4592), .ZN(n4338) );
  AND2_X1 U5869 ( .A1(n4684), .A2(n4290), .ZN(n4339) );
  NAND2_X1 U5870 ( .A1(n5236), .A2(n5235), .ZN(n8503) );
  INV_X1 U5871 ( .A(n8503), .ZN(n4447) );
  NAND2_X1 U5872 ( .A1(n6126), .A2(n6143), .ZN(n8868) );
  INV_X1 U5873 ( .A(n8868), .ZN(n8806) );
  AND2_X1 U5874 ( .A1(n9557), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4340) );
  INV_X1 U5875 ( .A(n7815), .ZN(n7768) );
  AND2_X1 U5876 ( .A1(n6996), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4341) );
  OAI21_X1 U5877 ( .B1(n6874), .B2(n4292), .A(n5053), .ZN(n6737) );
  NAND2_X1 U5878 ( .A1(n6549), .A2(n7913), .ZN(n6645) );
  INV_X1 U5879 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4736) );
  AND2_X1 U5880 ( .A1(n9683), .A2(n9890), .ZN(n4342) );
  INV_X1 U5881 ( .A(n8804), .ZN(n4611) );
  NAND2_X1 U5882 ( .A1(n4672), .A2(n4671), .ZN(n6723) );
  NAND2_X1 U5883 ( .A1(n4689), .A2(n5500), .ZN(n7020) );
  OR2_X1 U5884 ( .A1(n7141), .A2(n7287), .ZN(n7140) );
  NAND2_X1 U5885 ( .A1(n6953), .A2(n7629), .ZN(n7119) );
  INV_X1 U5886 ( .A(n4360), .ZN(n4359) );
  NOR2_X1 U5887 ( .A1(n4361), .A2(n7455), .ZN(n4360) );
  INV_X1 U5888 ( .A(n4549), .ZN(n9443) );
  NOR3_X1 U5889 ( .A1(n7140), .A2(n9442), .A3(n4551), .ZN(n4549) );
  AND2_X1 U5890 ( .A1(n5350), .A2(n9800), .ZN(n4343) );
  NOR2_X1 U5891 ( .A1(n6984), .A2(n6783), .ZN(n4547) );
  INV_X1 U5892 ( .A(n9767), .ZN(n9770) );
  INV_X1 U5893 ( .A(n9005), .ZN(n4397) );
  NAND2_X1 U5894 ( .A1(n4685), .A2(n5479), .ZN(n6620) );
  NAND2_X1 U5895 ( .A1(n7659), .A2(n6960), .ZN(n6961) );
  INV_X1 U5896 ( .A(n7808), .ZN(n7771) );
  INV_X1 U5897 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n4629) );
  AOI21_X1 U5898 ( .B1(n5401), .B2(n8585), .A(n5400), .ZN(n7888) );
  AOI21_X1 U5899 ( .B1(n8018), .B2(n8045), .A(n4470), .ZN(n8019) );
  AOI21_X1 U5900 ( .B1(n8007), .B2(n8011), .A(n8045), .ZN(n4473) );
  AND2_X1 U5901 ( .A1(n6814), .A2(n8045), .ZN(n4476) );
  NAND2_X1 U5902 ( .A1(n7134), .A2(n7118), .ZN(n7325) );
  NAND2_X1 U5903 ( .A1(n5631), .A2(n4540), .ZN(n4541) );
  INV_X1 U5904 ( .A(n8115), .ZN(n4627) );
  NAND2_X1 U5905 ( .A1(n4665), .A2(n4664), .ZN(n9327) );
  NAND2_X1 U5906 ( .A1(n4752), .A2(n4750), .ZN(n8976) );
  INV_X1 U5907 ( .A(n4738), .ZN(n9116) );
  NAND2_X1 U5908 ( .A1(n7116), .A2(n4287), .ZN(n7134) );
  NAND3_X1 U5909 ( .A1(n4344), .A2(n6132), .A3(n8806), .ZN(n6159) );
  NAND2_X1 U5910 ( .A1(n6127), .A2(n6128), .ZN(n4344) );
  AOI21_X2 U5911 ( .B1(n6750), .B2(n6746), .A(n6747), .ZN(n6831) );
  AND3_X2 U5912 ( .A1(n4624), .A2(n4622), .A3(n4330), .ZN(n6750) );
  AND2_X2 U5913 ( .A1(n4771), .A2(n4772), .ZN(n5642) );
  NAND2_X1 U5914 ( .A1(n5885), .A2(n5884), .ZN(n8727) );
  NAND2_X1 U5915 ( .A1(n9516), .A2(n9517), .ZN(n9521) );
  AOI21_X1 U5916 ( .B1(n8892), .B2(n4328), .A(n4348), .ZN(n8893) );
  NOR2_X1 U5917 ( .A1(n9541), .A2(n9542), .ZN(n9540) );
  NOR2_X1 U5918 ( .A1(n6183), .A2(n6388), .ZN(n6522) );
  NOR2_X1 U5919 ( .A1(n9616), .A2(n9615), .ZN(n9614) );
  AOI21_X1 U5920 ( .B1(n9593), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9588), .ZN(
        n9602) );
  AND3_X4 U5921 ( .A1(n4771), .A2(n4772), .A3(n5630), .ZN(n5631) );
  NOR2_X2 U5922 ( .A1(n8965), .A2(n8964), .ZN(n9082) );
  NAND2_X1 U5923 ( .A1(n6046), .A2(n6047), .ZN(n8736) );
  NAND2_X1 U5924 ( .A1(n5379), .A2(n7983), .ZN(n7465) );
  NAND2_X1 U5925 ( .A1(n8511), .A2(n8512), .ZN(n5385) );
  NAND2_X1 U5926 ( .A1(n5020), .A2(n5019), .ZN(n4409) );
  NOR2_X2 U5927 ( .A1(n8410), .A2(n5391), .ZN(n8392) );
  OR2_X1 U5928 ( .A1(n6539), .A2(n4265), .ZN(n4346) );
  NAND2_X1 U5929 ( .A1(n4265), .A2(n5865), .ZN(n4347) );
  NAND2_X1 U5930 ( .A1(n8776), .A2(n8775), .ZN(n8774) );
  NOR2_X2 U5931 ( .A1(n5916), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5932) );
  INV_X1 U5932 ( .A(n8990), .ZN(n4352) );
  OAI21_X1 U5933 ( .B1(n9430), .B2(n4356), .A(n4354), .ZN(n9409) );
  NAND2_X1 U5934 ( .A1(n8994), .A2(n4364), .ZN(n4367) );
  NAND2_X1 U5935 ( .A1(n4371), .A2(n4660), .ZN(n9057) );
  AOI21_X1 U5936 ( .B1(n7504), .B2(n4323), .A(n4372), .ZN(n4666) );
  INV_X2 U5937 ( .A(n5757), .ZN(n4771) );
  NAND2_X1 U5938 ( .A1(n5186), .A2(n4278), .ZN(n4386) );
  OAI21_X1 U5939 ( .B1(n5186), .B2(n4921), .A(n4920), .ZN(n5203) );
  NAND2_X1 U5940 ( .A1(n4921), .A2(n4920), .ZN(n4396) );
  XNOR2_X1 U5941 ( .A(n7532), .B(SI_30_), .ZN(n7891) );
  NAND2_X1 U5942 ( .A1(n5129), .A2(n4298), .ZN(n4402) );
  NAND2_X1 U5943 ( .A1(n5066), .A2(n4326), .ZN(n4411) );
  NAND2_X1 U5944 ( .A1(n5066), .A2(n4861), .ZN(n4412) );
  NAND2_X2 U5945 ( .A1(n4421), .A2(n4419), .ZN(n4849) );
  NAND3_X1 U5946 ( .A1(n4420), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4419) );
  NAND3_X1 U5947 ( .A1(n8363), .A2(n4423), .A3(n4422), .ZN(n4421) );
  NAND2_X1 U5948 ( .A1(n5322), .A2(n4426), .ZN(n4425) );
  NAND2_X1 U5949 ( .A1(n5322), .A2(n5321), .ZN(n5337) );
  NAND2_X1 U5950 ( .A1(n4486), .A2(n7764), .ZN(n4432) );
  NAND2_X1 U5951 ( .A1(n4430), .A2(n4282), .ZN(n7821) );
  NAND2_X1 U5952 ( .A1(n4483), .A2(n4431), .ZN(n4430) );
  NAND2_X1 U5953 ( .A1(n4432), .A2(n4433), .ZN(n4431) );
  AND4_X1 U5954 ( .A1(n4715), .A2(n4436), .A3(n4819), .A4(n4820), .ZN(n5413)
         );
  NAND4_X1 U5955 ( .A1(n4435), .A2(n4436), .A3(n4819), .A4(n4715), .ZN(n5411)
         );
  NAND3_X1 U5956 ( .A1(n4715), .A2(n4819), .A3(n4436), .ZN(n5366) );
  NOR2_X2 U5957 ( .A1(n5017), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n4436) );
  NOR2_X2 U5958 ( .A1(n4817), .A2(n4818), .ZN(n4819) );
  NAND2_X1 U5959 ( .A1(n4308), .A2(n8364), .ZN(n8371) );
  INV_X1 U5960 ( .A(n8551), .ZN(n4442) );
  NAND2_X1 U5961 ( .A1(n4442), .A2(n4443), .ZN(n8501) );
  INV_X2 U5962 ( .A(n4849), .ZN(n6216) );
  XNOR2_X1 U5963 ( .A(n4838), .B(n4837), .ZN(n4971) );
  OAI21_X1 U5964 ( .B1(n4849), .B2(n4474), .A(n5689), .ZN(n4838) );
  NAND3_X1 U5965 ( .A1(n4479), .A2(n4477), .A3(n7936), .ZN(n4475) );
  AND2_X1 U5966 ( .A1(n7936), .A2(n6814), .ZN(n7937) );
  NAND3_X1 U5967 ( .A1(n7914), .A2(n7912), .A3(n4478), .ZN(n4477) );
  INV_X1 U5968 ( .A(n8045), .ZN(n4478) );
  NAND2_X1 U5969 ( .A1(n5697), .A2(n4284), .ZN(n4482) );
  NAND2_X1 U5970 ( .A1(n7737), .A2(n4489), .ZN(n7741) );
  NAND2_X1 U5971 ( .A1(n7705), .A2(n4498), .ZN(n4493) );
  NAND4_X1 U5972 ( .A1(n4505), .A2(n7725), .A3(n4501), .A4(n9105), .ZN(n7726)
         );
  INV_X1 U5973 ( .A(n7658), .ZN(n4518) );
  NAND2_X1 U5974 ( .A1(n4303), .A2(n7658), .ZN(n7842) );
  OAI211_X1 U5975 ( .C1(n4303), .C2(n4519), .A(n4517), .B(n4522), .ZN(n7665)
         );
  INV_X1 U5976 ( .A(n4520), .ZN(n4519) );
  INV_X1 U5977 ( .A(n6961), .ZN(n4523) );
  NAND2_X1 U5978 ( .A1(n4541), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5666) );
  INV_X1 U5979 ( .A(n4541), .ZN(n5665) );
  NAND2_X1 U5980 ( .A1(n4325), .A2(n4546), .ZN(n6965) );
  AND2_X1 U5981 ( .A1(n4547), .A2(n6586), .ZN(n6982) );
  INV_X1 U5982 ( .A(n7140), .ZN(n4548) );
  NAND2_X1 U5983 ( .A1(n4548), .A2(n4285), .ZN(n9405) );
  INV_X1 U5984 ( .A(n4553), .ZN(n9099) );
  NAND2_X1 U5985 ( .A1(n6874), .A2(n4565), .ZN(n4561) );
  NAND2_X1 U5986 ( .A1(n4561), .A2(n4562), .ZN(n6918) );
  INV_X1 U5987 ( .A(n8070), .ZN(n4567) );
  NAND2_X1 U5988 ( .A1(n4567), .A2(n5024), .ZN(n4568) );
  NAND3_X1 U5989 ( .A1(n4569), .A2(n8073), .A3(n4568), .ZN(n5038) );
  NAND3_X1 U5990 ( .A1(n6545), .A2(n5024), .A3(n5010), .ZN(n4569) );
  NAND2_X1 U5991 ( .A1(n4570), .A2(n4329), .ZN(n7247) );
  OAI21_X1 U5992 ( .B1(n8453), .B2(n4575), .A(n4573), .ZN(n4578) );
  INV_X1 U5993 ( .A(n4578), .ZN(n8423) );
  OAI21_X2 U5994 ( .B1(n5411), .B2(P2_IR_REG_26__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4579) );
  NAND2_X1 U5995 ( .A1(n7469), .A2(n4279), .ZN(n4580) );
  NAND2_X1 U5996 ( .A1(n4580), .A2(n4581), .ZN(n8525) );
  INV_X1 U5997 ( .A(n4583), .ZN(n7471) );
  OAI211_X1 U5998 ( .C1(n8795), .C2(n4338), .A(n4590), .B(n4587), .ZN(n6167)
         );
  NAND2_X1 U5999 ( .A1(n8795), .A2(n4588), .ZN(n4587) );
  NAND2_X2 U6000 ( .A1(n7860), .A2(n8735), .ZN(n8795) );
  NAND2_X1 U6001 ( .A1(n6830), .A2(n4595), .ZN(n4593) );
  NAND2_X1 U6002 ( .A1(n4593), .A2(n4594), .ZN(n7233) );
  NAND2_X1 U6003 ( .A1(n8803), .A2(n4607), .ZN(n4606) );
  NAND4_X1 U6004 ( .A1(n4621), .A2(n4626), .A3(n4623), .A4(n4625), .ZN(n4622)
         );
  XNOR2_X1 U6005 ( .A(n5704), .B(n5705), .ZN(n7524) );
  NAND2_X1 U6006 ( .A1(n5701), .A2(n5702), .ZN(n4625) );
  NAND3_X1 U6007 ( .A1(n4628), .A2(n9345), .A3(n5637), .ZN(n4631) );
  NAND3_X1 U6008 ( .A1(n5640), .A2(n4630), .A3(n5641), .ZN(n8884) );
  NAND2_X1 U6009 ( .A1(n5631), .A2(n4633), .ZN(n5634) );
  NOR2_X1 U6010 ( .A1(n9043), .A2(n9042), .ZN(n9041) );
  INV_X1 U6011 ( .A(n4646), .ZN(n9003) );
  OAI21_X1 U6012 ( .B1(n9043), .B2(n4647), .A(n4648), .ZN(n4646) );
  NAND2_X1 U6013 ( .A1(n4874), .A2(n4652), .ZN(n4651) );
  NAND2_X1 U6014 ( .A1(n4651), .A2(n4654), .ZN(n5129) );
  NAND2_X1 U6015 ( .A1(n8252), .A2(n4276), .ZN(n4674) );
  NAND2_X1 U6016 ( .A1(n4674), .A2(n4675), .ZN(n8172) );
  NAND2_X1 U6017 ( .A1(n4685), .A2(n4327), .ZN(n6621) );
  NAND2_X1 U6018 ( .A1(n8195), .A2(n4686), .ZN(n5549) );
  NAND3_X1 U6019 ( .A1(n6701), .A2(n8099), .A3(n8064), .ZN(n5458) );
  NAND2_X1 U6020 ( .A1(n4689), .A2(n4688), .ZN(n7010) );
  NAND3_X1 U6021 ( .A1(n5586), .A2(n5585), .A3(n4703), .ZN(n4702) );
  NAND3_X1 U6022 ( .A1(n5586), .A2(n4704), .A3(n5585), .ZN(n4705) );
  INV_X1 U6023 ( .A(n4705), .ZN(n8260) );
  NAND2_X1 U6024 ( .A1(n5190), .A2(n4706), .ZN(n4708) );
  NAND4_X1 U6025 ( .A1(n4709), .A2(n4812), .A3(n4814), .A4(n4813), .ZN(n4716)
         );
  INV_X1 U6026 ( .A(n6883), .ZN(n4712) );
  OAI21_X2 U6027 ( .B1(n6881), .B2(n4713), .A(n4710), .ZN(n6923) );
  AOI21_X1 U6028 ( .B1(n4712), .B2(n4714), .A(n4711), .ZN(n4710) );
  NAND2_X1 U6029 ( .A1(n8392), .A2(n8391), .ZN(n8390) );
  NAND2_X1 U6030 ( .A1(n8392), .A2(n4718), .ZN(n4717) );
  NAND2_X1 U6031 ( .A1(n5385), .A2(n4286), .ZN(n8495) );
  NAND2_X1 U6032 ( .A1(n4731), .A2(n6549), .ZN(n6813) );
  NAND2_X1 U6033 ( .A1(n6813), .A2(n7937), .ZN(n5374) );
  NAND2_X1 U6034 ( .A1(n4732), .A2(n4733), .ZN(n7242) );
  OR2_X2 U6035 ( .A1(n4947), .A2(n5415), .ZN(n4949) );
  AND2_X2 U6036 ( .A1(n5413), .A2(n4734), .ZN(n4947) );
  NAND2_X1 U6037 ( .A1(n7465), .A2(n4737), .ZN(n8526) );
  NAND2_X1 U6038 ( .A1(n8526), .A2(n5382), .ZN(n5383) );
  OAI21_X1 U6039 ( .B1(n9162), .B2(n4299), .A(n4748), .ZN(n9149) );
  NAND2_X1 U6040 ( .A1(n9050), .A2(n4753), .ZN(n4752) );
  NAND2_X1 U6041 ( .A1(n9403), .A2(n4764), .ZN(n4763) );
  NAND2_X1 U6042 ( .A1(n6964), .A2(n6963), .ZN(n7116) );
  NAND2_X1 U6043 ( .A1(n5665), .A2(n4775), .ZN(n4778) );
  INV_X1 U6044 ( .A(n4778), .ZN(n5636) );
  NOR2_X1 U6045 ( .A1(n9250), .A2(n9451), .ZN(n9030) );
  NAND2_X1 U6046 ( .A1(n7867), .A2(n7866), .ZN(n8121) );
  OR2_X1 U6047 ( .A1(n7765), .A2(n7809), .ZN(n6683) );
  NAND2_X1 U6048 ( .A1(n8795), .A2(n7863), .ZN(n6131) );
  NAND2_X1 U6049 ( .A1(n5649), .A2(n5648), .ZN(n5677) );
  NAND2_X1 U6050 ( .A1(n7815), .A2(n9157), .ZN(n7752) );
  OAI21_X1 U6051 ( .B1(n6615), .B2(n8128), .A(n5691), .ZN(n6539) );
  NAND2_X1 U6052 ( .A1(n6099), .A2(n7771), .ZN(n5675) );
  NAND2_X1 U6053 ( .A1(n5267), .A2(n5266), .ZN(n5269) );
  XNOR2_X1 U6054 ( .A(n5203), .B(n5202), .ZN(n6766) );
  NAND2_X1 U6055 ( .A1(n8236), .A2(n5572), .ZN(n5577) );
  OR2_X1 U6056 ( .A1(n4825), .A2(n5415), .ZN(n4823) );
  INV_X1 U6057 ( .A(n8884), .ZN(n6775) );
  XNOR2_X1 U6058 ( .A(n5651), .B(P1_IR_REG_20__SCAN_IN), .ZN(n7808) );
  NOR2_X1 U6059 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4809) );
  INV_X1 U6060 ( .A(n8181), .ZN(n5584) );
  CLKBUF_X1 U6061 ( .A(n7242), .Z(n7274) );
  NAND2_X1 U6062 ( .A1(n8238), .A2(n8237), .ZN(n8236) );
  AOI22_X1 U6063 ( .A1(n5445), .A2(n8092), .B1(n8382), .B2(n8149), .ZN(n5361)
         );
  NOR2_X1 U6064 ( .A1(n5577), .A2(n5576), .ZN(n8214) );
  AND4_X2 U6065 ( .A1(n4986), .A2(n4985), .A3(n4984), .A4(n4983), .ZN(n4994)
         );
  NOR2_X1 U6066 ( .A1(n8592), .A2(n8575), .ZN(n6553) );
  NAND4_X2 U6067 ( .A1(n4969), .A2(n4968), .A3(n4967), .A4(n4966), .ZN(n8316)
         );
  AND2_X2 U6068 ( .A1(n4830), .A2(n8114), .ZN(n4996) );
  XNOR2_X1 U6069 ( .A(n5299), .B(n5298), .ZN(n7399) );
  NAND2_X1 U6070 ( .A1(n4270), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5694) );
  NAND2_X2 U6071 ( .A1(n7232), .A2(n7236), .ZN(n7346) );
  NOR2_X1 U6072 ( .A1(n9176), .A2(n9184), .ZN(n9299) );
  NAND2_X4 U6073 ( .A1(n5392), .A2(n5394), .ZN(n6283) );
  INV_X1 U6074 ( .A(n7631), .ZN(n7117) );
  AND2_X1 U6075 ( .A1(n4999), .A2(n4998), .ZN(n4779) );
  AND2_X1 U6076 ( .A1(n6589), .A2(n6588), .ZN(n9433) );
  INV_X1 U6077 ( .A(n8667), .ZN(n5451) );
  OR2_X1 U6078 ( .A1(n8457), .A2(n8243), .ZN(n4780) );
  OR2_X1 U6079 ( .A1(n8703), .A2(n5384), .ZN(n4781) );
  NOR2_X1 U6080 ( .A1(n8077), .A2(n5124), .ZN(n4782) );
  AND2_X1 U6081 ( .A1(n4873), .A2(n4872), .ZN(n4785) );
  AND2_X1 U6082 ( .A1(n4898), .A2(n4897), .ZN(n4786) );
  OR2_X1 U6083 ( .A1(n9058), .A2(n9435), .ZN(n4787) );
  AND2_X1 U6084 ( .A1(n4881), .A2(n4880), .ZN(n4788) );
  OR3_X1 U6085 ( .A1(n8065), .A2(n8098), .A3(n9716), .ZN(n4789) );
  AND2_X1 U6086 ( .A1(n7747), .A2(n7620), .ZN(n4790) );
  OR2_X1 U6087 ( .A1(n7810), .A2(n4434), .ZN(n4791) );
  OR2_X1 U6088 ( .A1(n9120), .A2(n9108), .ZN(n4792) );
  AND2_X1 U6089 ( .A1(n7905), .A2(n7925), .ZN(n4793) );
  AND4_X1 U6090 ( .A1(n9002), .A2(n7740), .A3(n9033), .A4(n7646), .ZN(n4795)
         );
  AND2_X1 U6091 ( .A1(n5443), .A2(n5442), .ZN(n4796) );
  NAND2_X1 U6092 ( .A1(n8503), .A2(n8298), .ZN(n4797) );
  INV_X1 U6093 ( .A(n5402), .ZN(n8436) );
  INV_X1 U6094 ( .A(n8552), .ZN(n5201) );
  INV_X1 U6095 ( .A(n8544), .ZN(n5380) );
  INV_X1 U6096 ( .A(n8044), .ZN(n8382) );
  NAND2_X1 U6097 ( .A1(n8023), .A2(n8045), .ZN(n8024) );
  NAND2_X1 U6098 ( .A1(n8424), .A2(n8024), .ZN(n8025) );
  NAND2_X1 U6099 ( .A1(n8022), .A2(n8045), .ZN(n8026) );
  AOI21_X1 U6100 ( .B1(n8027), .B2(n8026), .A(n8025), .ZN(n8033) );
  OAI21_X1 U6101 ( .B1(n8052), .B2(n4478), .A(n8051), .ZN(n8053) );
  NOR2_X1 U6102 ( .A1(n8057), .A2(n8053), .ZN(n8054) );
  AND2_X1 U6103 ( .A1(n8055), .A2(n8054), .ZN(n8056) );
  INV_X1 U6104 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5624) );
  INV_X1 U6105 ( .A(n8497), .ZN(n5386) );
  INV_X1 U6106 ( .A(n8057), .ZN(n7895) );
  INV_X1 U6107 ( .A(n5133), .ZN(n4800) );
  NOR2_X1 U6108 ( .A1(n5629), .A2(n5628), .ZN(n5630) );
  INV_X1 U6109 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5623) );
  INV_X1 U6110 ( .A(n5195), .ZN(n4802) );
  AND2_X1 U6111 ( .A1(n8316), .A2(n7909), .ZN(n5469) );
  INV_X1 U6112 ( .A(n5275), .ZN(n4806) );
  INV_X1 U6113 ( .A(n5177), .ZN(n4801) );
  OR2_X1 U6114 ( .A1(n5273), .A2(n5272), .ZN(n5275) );
  INV_X1 U6115 ( .A(n5851), .ZN(n5852) );
  OR2_X1 U6116 ( .A1(n9278), .A2(n9138), .ZN(n8962) );
  NOR2_X1 U6117 ( .A1(n5765), .A2(n5764), .ZN(n5794) );
  INV_X1 U6118 ( .A(n7728), .ZN(n8996) );
  AND2_X1 U6119 ( .A1(n7680), .A2(n7693), .ZN(n9411) );
  NAND2_X1 U6120 ( .A1(n5651), .A2(n5646), .ZN(n5647) );
  INV_X1 U6121 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5947) );
  INV_X1 U6122 ( .A(n5065), .ZN(n4861) );
  INV_X1 U6123 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U6124 ( .A1(n4802), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5209) );
  INV_X1 U6125 ( .A(n5248), .ZN(n4804) );
  INV_X1 U6126 ( .A(n5573), .ZN(n5574) );
  INV_X1 U6127 ( .A(n7204), .ZN(n5523) );
  NAND2_X1 U6128 ( .A1(n4801), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5179) );
  INV_X1 U6129 ( .A(n8373), .ZN(n8364) );
  NAND2_X1 U6130 ( .A1(n4994), .A2(n8575), .ZN(n7928) );
  OR2_X1 U6131 ( .A1(n6088), .A2(n6087), .ZN(n6148) );
  INV_X1 U6132 ( .A(n5697), .ZN(n5772) );
  NAND2_X1 U6133 ( .A1(n8787), .A2(n5946), .ZN(n5962) );
  OAI22_X1 U6134 ( .A1(n9044), .A2(n9435), .B1(n9006), .B2(n9005), .ZN(n9007)
         );
  AND2_X1 U6135 ( .A1(n5876), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5891) );
  AND2_X1 U6136 ( .A1(n9242), .A2(n9455), .ZN(n9243) );
  OR2_X1 U6137 ( .A1(n9322), .A2(n8872), .ZN(n7501) );
  OR2_X1 U6138 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  INV_X1 U6139 ( .A(n5932), .ZN(n5933) );
  NAND2_X1 U6140 ( .A1(n4895), .A2(n4894), .ZN(n4898) );
  NAND2_X1 U6141 ( .A1(n4870), .A2(n4869), .ZN(n4873) );
  OR2_X1 U6142 ( .A1(n5055), .A2(n5054), .ZN(n5071) );
  OR2_X1 U6143 ( .A1(n5209), .A2(n5208), .ZN(n5238) );
  OR2_X1 U6144 ( .A1(n5291), .A2(n8185), .ZN(n5309) );
  XNOR2_X1 U6145 ( .A(n8620), .B(n5590), .ZN(n8216) );
  AND2_X1 U6146 ( .A1(n5393), .A2(n6279), .ZN(n8228) );
  OR2_X1 U6147 ( .A1(n5309), .A2(n8268), .ZN(n5327) );
  INV_X1 U6148 ( .A(n8478), .ZN(n8479) );
  AND2_X1 U6149 ( .A1(n8001), .A2(n7998), .ZN(n8512) );
  INV_X1 U6150 ( .A(n8267), .ZN(n8242) );
  AND2_X1 U6151 ( .A1(n5433), .A2(n9709), .ZN(n6696) );
  INV_X1 U6152 ( .A(n8626), .ZN(n8457) );
  INV_X1 U6153 ( .A(n9752), .ZN(n8670) );
  OR2_X1 U6154 ( .A1(n9752), .A2(n8357), .ZN(n5610) );
  NAND2_X1 U6155 ( .A1(n8817), .A2(n5883), .ZN(n5885) );
  OR2_X1 U6156 ( .A1(n7865), .A2(n7864), .ZN(n7866) );
  NOR2_X1 U6157 ( .A1(n5920), .A2(n8778), .ZN(n5935) );
  OR2_X1 U6158 ( .A1(n5739), .A2(n5738), .ZN(n5740) );
  AOI22_X1 U6159 ( .A1(n8126), .A2(n6715), .B1(n6168), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U6160 ( .A1(n5953), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5990) );
  OR2_X1 U6161 ( .A1(n9455), .A2(n6530), .ZN(n6138) );
  AND2_X1 U6162 ( .A1(n7550), .A2(n6671), .ZN(n9022) );
  INV_X1 U6163 ( .A(n9252), .ZN(n9040) );
  INV_X1 U6164 ( .A(n9315), .ZN(n9232) );
  INV_X1 U6165 ( .A(n8872), .ZN(n9412) );
  AND2_X1 U6166 ( .A1(n7681), .A2(n7674), .ZN(n7637) );
  NOR2_X1 U6167 ( .A1(n9244), .A2(n9243), .ZN(n9245) );
  INV_X1 U6168 ( .A(n6780), .ZN(n9644) );
  INV_X1 U6169 ( .A(n9188), .ZN(n9437) );
  AND2_X1 U6170 ( .A1(n4915), .A2(n4914), .ZN(n4957) );
  NAND2_X1 U6171 ( .A1(n4892), .A2(n4891), .ZN(n5128) );
  NOR2_X1 U6172 ( .A1(n5616), .A2(n8285), .ZN(n5617) );
  INV_X1 U6173 ( .A(n8285), .ZN(n8271) );
  NAND2_X1 U6174 ( .A1(n4789), .A2(n4783), .ZN(n8103) );
  OR2_X1 U6175 ( .A1(n8399), .A2(n5329), .ZN(n5335) );
  AND4_X1 U6176 ( .A1(n5200), .A2(n5199), .A3(n5198), .A4(n5197), .ZN(n8253)
         );
  INV_X1 U6177 ( .A(n9697), .ZN(n9951) );
  NAND2_X1 U6178 ( .A1(n6739), .A2(n8587), .ZN(n8567) );
  AND2_X1 U6179 ( .A1(n5606), .A2(n9716), .ZN(n9722) );
  AND2_X1 U6180 ( .A1(n9759), .A2(n9722), .ZN(n8714) );
  OR2_X1 U6181 ( .A1(n5462), .A2(n5432), .ZN(n6694) );
  AND4_X1 U6182 ( .A1(n6153), .A2(n6152), .A3(n6151), .A4(n6150), .ZN(n9058)
         );
  AND4_X1 U6183 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n9109)
         );
  AND4_X1 U6184 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n9208)
         );
  AND2_X1 U6185 ( .A1(n4352), .A2(n8991), .ZN(n9121) );
  INV_X1 U6186 ( .A(n9433), .ZN(n9414) );
  AND2_X1 U6187 ( .A1(n7662), .A2(n7660), .ZN(n7830) );
  AND2_X1 U6188 ( .A1(n9424), .A2(n6714), .ZN(n9446) );
  OR2_X1 U6189 ( .A1(n6713), .A2(n7808), .ZN(n9679) );
  OR2_X1 U6190 ( .A1(n7752), .A2(n7808), .ZN(n9456) );
  INV_X1 U6191 ( .A(n6113), .ZN(n9630) );
  INV_X1 U6192 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5887) );
  INV_X1 U6193 ( .A(n8362), .ZN(n9960) );
  AND4_X1 U6194 ( .A1(n5183), .A2(n5182), .A3(n5181), .A4(n5180), .ZN(n7466)
         );
  INV_X1 U6195 ( .A(n6726), .ZN(n8312) );
  INV_X1 U6196 ( .A(n8581), .ZN(n8556) );
  INV_X1 U6197 ( .A(n8582), .ZN(n8559) );
  INV_X1 U6198 ( .A(n9767), .ZN(n8676) );
  OR2_X1 U6199 ( .A1(n6694), .A2(n5435), .ZN(n9767) );
  INV_X1 U6200 ( .A(n8535), .ZN(n8707) );
  INV_X1 U6201 ( .A(n8714), .ZN(n8711) );
  OR2_X1 U6202 ( .A1(n6694), .A2(n5440), .ZN(n9758) );
  INV_X1 U6203 ( .A(n7925), .ZN(n8099) );
  INV_X1 U6204 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6250) );
  INV_X1 U6205 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9820) );
  NAND2_X1 U6206 ( .A1(n8121), .A2(n8120), .ZN(n8143) );
  INV_X1 U6207 ( .A(n6157), .ZN(n6158) );
  INV_X1 U6208 ( .A(n7231), .ZN(n8878) );
  OR2_X1 U6209 ( .A1(P1_U3083), .A2(n9504), .ZN(n9628) );
  OR2_X1 U6210 ( .A1(n6535), .A2(n6679), .ZN(n9693) );
  OR2_X1 U6211 ( .A1(n6535), .A2(n9343), .ZN(n9683) );
  INV_X1 U6212 ( .A(n9631), .ZN(n9632) );
  OR3_X1 U6213 ( .A1(n6168), .A2(n7100), .A3(P1_U3084), .ZN(n9635) );
  INV_X1 U6214 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6247) );
  INV_X1 U6215 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6220) );
  NOR2_X1 U6216 ( .A1(n9798), .A2(n9797), .ZN(n9796) );
  NAND2_X1 U6217 ( .A1(n5039), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5055) );
  INV_X1 U6218 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5093) );
  OR2_X2 U6219 ( .A1(n5094), .A2(n5093), .ZN(n5105) );
  INV_X1 U6220 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5117) );
  INV_X1 U6221 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5143) );
  OR2_X2 U6222 ( .A1(n5144), .A2(n5143), .ZN(n5162) );
  INV_X1 U6223 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5161) );
  INV_X1 U6224 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7430) );
  INV_X1 U6225 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U6226 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n4803) );
  INV_X1 U6227 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5272) );
  INV_X1 U6228 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n4807) );
  NAND2_X1 U6229 ( .A1(n5275), .A2(n4807), .ZN(n4808) );
  NAND2_X1 U6230 ( .A1(n5291), .A2(n4808), .ZN(n8437) );
  NAND2_X1 U6231 ( .A1(n4987), .A2(n4809), .ZN(n5017) );
  NOR2_X1 U6232 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4814) );
  NOR2_X1 U6233 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4813) );
  NOR2_X1 U6234 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4812) );
  INV_X1 U6235 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4815) );
  NAND4_X1 U6236 ( .A1(n4816), .A2(n4815), .A3(n4960), .A4(n5153), .ZN(n4818)
         );
  NAND4_X1 U6237 ( .A1(n5220), .A2(n4707), .A3(n5156), .A4(n5363), .ZN(n4817)
         );
  NOR3_X1 U6238 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n4820) );
  INV_X1 U6239 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4821) );
  AND2_X2 U6240 ( .A1(n4947), .A2(n4948), .ZN(n4825) );
  INV_X1 U6241 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4824) );
  NAND2_X1 U6242 ( .A1(n4825), .A2(n4824), .ZN(n4827) );
  INV_X1 U6243 ( .A(n4264), .ZN(n5329) );
  OR2_X1 U6244 ( .A1(n8437), .A2(n5329), .ZN(n4835) );
  INV_X1 U6245 ( .A(n4830), .ZN(n7520) );
  INV_X1 U6246 ( .A(n6261), .ZN(n5357) );
  INV_X1 U6247 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9846) );
  AND2_X2 U6248 ( .A1(n7520), .A2(n4829), .ZN(n4981) );
  INV_X2 U6249 ( .A(n5398), .ZN(n6260) );
  NAND2_X1 U6250 ( .A1(n6260), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n4832) );
  NAND2_X1 U6251 ( .A1(n5354), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n4831) );
  OAI211_X1 U6252 ( .C1(n5357), .C2(n9846), .A(n4832), .B(n4831), .ZN(n4833)
         );
  INV_X1 U6253 ( .A(n4833), .ZN(n4834) );
  AND2_X1 U6254 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4836) );
  NAND2_X1 U6255 ( .A1(n4849), .A2(n4836), .ZN(n5689) );
  INV_X1 U6256 ( .A(SI_1_), .ZN(n4837) );
  MUX2_X1 U6257 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4849), .Z(n4970) );
  NAND2_X1 U6258 ( .A1(n4971), .A2(n4970), .ZN(n4840) );
  NAND2_X1 U6259 ( .A1(n4838), .A2(SI_1_), .ZN(n4839) );
  NAND2_X1 U6260 ( .A1(n4840), .A2(n4839), .ZN(n4991) );
  INV_X1 U6261 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6232) );
  INV_X1 U6262 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6229) );
  MUX2_X1 U6263 ( .A(n6232), .B(n6229), .S(n4849), .Z(n4841) );
  XNOR2_X1 U6264 ( .A(n4841), .B(SI_2_), .ZN(n4990) );
  NAND2_X1 U6265 ( .A1(n4991), .A2(n4990), .ZN(n4844) );
  INV_X1 U6266 ( .A(n4841), .ZN(n4842) );
  NAND2_X1 U6267 ( .A1(n4842), .A2(SI_2_), .ZN(n4843) );
  NAND2_X1 U6268 ( .A1(n4844), .A2(n4843), .ZN(n5003) );
  INV_X1 U6269 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6222) );
  MUX2_X1 U6270 ( .A(n9822), .B(n6222), .S(n4849), .Z(n4845) );
  XNOR2_X1 U6271 ( .A(n4845), .B(SI_3_), .ZN(n5002) );
  NAND2_X1 U6272 ( .A1(n5003), .A2(n5002), .ZN(n4848) );
  INV_X1 U6273 ( .A(n4845), .ZN(n4846) );
  NAND2_X1 U6274 ( .A1(n4846), .A2(SI_3_), .ZN(n4847) );
  NAND2_X1 U6275 ( .A1(n4848), .A2(n4847), .ZN(n5020) );
  INV_X1 U6276 ( .A(n4850), .ZN(n4851) );
  NAND2_X1 U6277 ( .A1(n4851), .A2(SI_4_), .ZN(n4852) );
  INV_X1 U6278 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6223) );
  INV_X1 U6279 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6227) );
  MUX2_X1 U6280 ( .A(n6223), .B(n6227), .S(n7538), .Z(n4853) );
  NAND2_X1 U6281 ( .A1(n5035), .A2(n5034), .ZN(n4856) );
  INV_X1 U6282 ( .A(n4853), .ZN(n4854) );
  NAND2_X1 U6283 ( .A1(n4854), .A2(SI_5_), .ZN(n4855) );
  MUX2_X1 U6284 ( .A(n9820), .B(n9837), .S(n7538), .Z(n4857) );
  NAND2_X1 U6285 ( .A1(n5049), .A2(n5048), .ZN(n4860) );
  INV_X1 U6286 ( .A(n4857), .ZN(n4858) );
  NAND2_X1 U6287 ( .A1(n4858), .A2(SI_6_), .ZN(n4859) );
  MUX2_X1 U6288 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7538), .Z(n4862) );
  NAND2_X1 U6289 ( .A1(n4862), .A2(SI_7_), .ZN(n4863) );
  MUX2_X1 U6290 ( .A(n6238), .B(n6241), .S(n7538), .Z(n4865) );
  INV_X1 U6291 ( .A(SI_8_), .ZN(n4864) );
  INV_X1 U6292 ( .A(n4865), .ZN(n4866) );
  NAND2_X1 U6293 ( .A1(n4866), .A2(SI_8_), .ZN(n4867) );
  MUX2_X1 U6294 ( .A(n6250), .B(n6247), .S(n7538), .Z(n4870) );
  INV_X1 U6295 ( .A(SI_9_), .ZN(n4869) );
  INV_X1 U6296 ( .A(n4870), .ZN(n4871) );
  NAND2_X1 U6297 ( .A1(n4871), .A2(SI_9_), .ZN(n4872) );
  INV_X1 U6298 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n4876) );
  INV_X1 U6299 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n4875) );
  MUX2_X1 U6300 ( .A(n4876), .B(n4875), .S(n7538), .Z(n4878) );
  INV_X1 U6301 ( .A(SI_10_), .ZN(n4877) );
  INV_X1 U6302 ( .A(n4878), .ZN(n4879) );
  NAND2_X1 U6303 ( .A1(n4879), .A2(SI_10_), .ZN(n4880) );
  INV_X1 U6304 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n4882) );
  INV_X1 U6305 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6258) );
  MUX2_X1 U6306 ( .A(n4882), .B(n6258), .S(n7538), .Z(n4883) );
  INV_X1 U6307 ( .A(n4883), .ZN(n4884) );
  INV_X1 U6308 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n4887) );
  INV_X1 U6309 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n4886) );
  MUX2_X1 U6310 ( .A(n4887), .B(n4886), .S(n7538), .Z(n4889) );
  INV_X1 U6311 ( .A(SI_12_), .ZN(n4888) );
  INV_X1 U6312 ( .A(n4889), .ZN(n4890) );
  NAND2_X1 U6313 ( .A1(n4890), .A2(SI_12_), .ZN(n4891) );
  INV_X1 U6314 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6393) );
  INV_X1 U6315 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4893) );
  MUX2_X1 U6316 ( .A(n6393), .B(n4893), .S(n7538), .Z(n4895) );
  INV_X1 U6317 ( .A(SI_13_), .ZN(n4894) );
  INV_X1 U6318 ( .A(n4895), .ZN(n4896) );
  NAND2_X1 U6319 ( .A1(n4896), .A2(SI_13_), .ZN(n4897) );
  INV_X1 U6320 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6449) );
  INV_X1 U6321 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6415) );
  MUX2_X1 U6322 ( .A(n6449), .B(n6415), .S(n7538), .Z(n4900) );
  INV_X1 U6323 ( .A(n4900), .ZN(n4901) );
  NAND2_X1 U6324 ( .A1(n4901), .A2(SI_14_), .ZN(n4902) );
  INV_X1 U6325 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6577) );
  INV_X1 U6326 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6575) );
  MUX2_X1 U6327 ( .A(n6577), .B(n6575), .S(n7538), .Z(n4905) );
  INV_X1 U6328 ( .A(SI_15_), .ZN(n4904) );
  INV_X1 U6329 ( .A(n4905), .ZN(n4906) );
  NAND2_X1 U6330 ( .A1(n4906), .A2(SI_15_), .ZN(n4907) );
  INV_X1 U6331 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n4910) );
  INV_X1 U6332 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n4909) );
  MUX2_X1 U6333 ( .A(n4910), .B(n4909), .S(n7538), .Z(n4912) );
  INV_X1 U6334 ( .A(SI_16_), .ZN(n4911) );
  NAND2_X1 U6335 ( .A1(n4912), .A2(n4911), .ZN(n4915) );
  INV_X1 U6336 ( .A(n4912), .ZN(n4913) );
  NAND2_X1 U6337 ( .A1(n4913), .A2(SI_16_), .ZN(n4914) );
  INV_X1 U6338 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6639) );
  INV_X1 U6339 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n4917) );
  MUX2_X1 U6340 ( .A(n6639), .B(n4917), .S(n7538), .Z(n4918) );
  XNOR2_X1 U6341 ( .A(n4918), .B(SI_17_), .ZN(n5185) );
  INV_X1 U6342 ( .A(n5185), .ZN(n4921) );
  INV_X1 U6343 ( .A(n4918), .ZN(n4919) );
  NAND2_X1 U6344 ( .A1(n4919), .A2(SI_17_), .ZN(n4920) );
  MUX2_X1 U6345 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7538), .Z(n4923) );
  XNOR2_X1 U6346 ( .A(n4923), .B(SI_18_), .ZN(n5202) );
  INV_X1 U6347 ( .A(n5202), .ZN(n4922) );
  INV_X1 U6348 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6809) );
  INV_X1 U6349 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6811) );
  MUX2_X1 U6350 ( .A(n6809), .B(n6811), .S(n7538), .Z(n4925) );
  INV_X1 U6351 ( .A(SI_19_), .ZN(n4924) );
  NAND2_X1 U6352 ( .A1(n4925), .A2(n4924), .ZN(n4928) );
  INV_X1 U6353 ( .A(n4925), .ZN(n4926) );
  NAND2_X1 U6354 ( .A1(n4926), .A2(SI_19_), .ZN(n4927) );
  NAND2_X1 U6355 ( .A1(n4928), .A2(n4927), .ZN(n5217) );
  INV_X1 U6356 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7512) );
  INV_X1 U6357 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6973) );
  MUX2_X1 U6358 ( .A(n7512), .B(n6973), .S(n7538), .Z(n4930) );
  INV_X1 U6359 ( .A(SI_20_), .ZN(n4929) );
  NAND2_X1 U6360 ( .A1(n4930), .A2(n4929), .ZN(n4933) );
  INV_X1 U6361 ( .A(n4930), .ZN(n4931) );
  NAND2_X1 U6362 ( .A1(n4931), .A2(SI_20_), .ZN(n4932) );
  INV_X1 U6363 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7009) );
  INV_X1 U6364 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7006) );
  MUX2_X1 U6365 ( .A(n7009), .B(n7006), .S(n7538), .Z(n4935) );
  XNOR2_X1 U6366 ( .A(n4935), .B(SI_21_), .ZN(n5244) );
  INV_X1 U6367 ( .A(n4935), .ZN(n4936) );
  NAND2_X1 U6368 ( .A1(n4936), .A2(SI_21_), .ZN(n4937) );
  INV_X1 U6369 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7058) );
  INV_X1 U6370 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9862) );
  MUX2_X1 U6371 ( .A(n7058), .B(n9862), .S(n7538), .Z(n4939) );
  INV_X1 U6372 ( .A(SI_22_), .ZN(n4938) );
  NAND2_X1 U6373 ( .A1(n4939), .A2(n4938), .ZN(n4942) );
  INV_X1 U6374 ( .A(n4939), .ZN(n4940) );
  NAND2_X1 U6375 ( .A1(n4940), .A2(SI_22_), .ZN(n4941) );
  NAND2_X1 U6376 ( .A1(n4942), .A2(n4941), .ZN(n5254) );
  INV_X1 U6377 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7148) );
  INV_X1 U6378 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n6031) );
  MUX2_X1 U6379 ( .A(n7148), .B(n6031), .S(n7538), .Z(n4943) );
  INV_X1 U6380 ( .A(SI_23_), .ZN(n9881) );
  NAND2_X1 U6381 ( .A1(n4943), .A2(n9881), .ZN(n4946) );
  INV_X1 U6382 ( .A(n4943), .ZN(n4944) );
  NAND2_X1 U6383 ( .A1(n4944), .A2(SI_23_), .ZN(n4945) );
  INV_X1 U6384 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7213) );
  INV_X1 U6385 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7199) );
  MUX2_X1 U6386 ( .A(n7213), .B(n7199), .S(n7538), .Z(n5281) );
  XNOR2_X1 U6387 ( .A(n5281), .B(SI_24_), .ZN(n5280) );
  XNOR2_X2 U6388 ( .A(n4949), .B(n4948), .ZN(n5392) );
  NAND2_X1 U6389 ( .A1(n7198), .A2(n7898), .ZN(n4951) );
  OR2_X1 U6390 ( .A1(n7899), .A2(n7213), .ZN(n4950) );
  INV_X1 U6391 ( .A(n8620), .ZN(n8440) );
  NAND2_X1 U6392 ( .A1(n5354), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4956) );
  NAND2_X1 U6393 ( .A1(n6260), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4955) );
  NAND2_X1 U6394 ( .A1(n5179), .A2(n7430), .ZN(n4952) );
  AND2_X1 U6395 ( .A1(n5195), .A2(n4952), .ZN(n8199) );
  NAND2_X1 U6396 ( .A1(n4264), .A2(n8199), .ZN(n4954) );
  NAND2_X1 U6397 ( .A1(n5343), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n4953) );
  INV_X1 U6398 ( .A(n8206), .ZN(n8302) );
  XNOR2_X1 U6399 ( .A(n4958), .B(n4957), .ZN(n6562) );
  NAND2_X1 U6400 ( .A1(n6562), .A2(n7898), .ZN(n4965) );
  INV_X1 U6401 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4961) );
  AND3_X1 U6402 ( .A1(n5153), .A2(n5156), .A3(n4961), .ZN(n5188) );
  NAND2_X1 U6403 ( .A1(n5190), .A2(n5188), .ZN(n4962) );
  NAND2_X1 U6404 ( .A1(n4962), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4963) );
  XNOR2_X1 U6405 ( .A(n4963), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8322) );
  AOI22_X1 U6406 ( .A1(n5223), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4560), .B2(
        n8322), .ZN(n4964) );
  NAND2_X1 U6407 ( .A1(n4997), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4969) );
  NAND2_X1 U6408 ( .A1(n4981), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4968) );
  NAND2_X1 U6409 ( .A1(n4982), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4967) );
  NAND2_X1 U6410 ( .A1(n4996), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4966) );
  INV_X1 U6411 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6214) );
  XNOR2_X1 U6412 ( .A(n4971), .B(n4970), .ZN(n6217) );
  INV_X1 U6413 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4972) );
  NAND2_X1 U6414 ( .A1(n4978), .A2(n8590), .ZN(n7919) );
  NAND2_X1 U6415 ( .A1(n8316), .A2(n4979), .ZN(n7927) );
  NAND2_X1 U6416 ( .A1(n7919), .A2(n7927), .ZN(n8069) );
  NAND2_X1 U6417 ( .A1(n4996), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U6418 ( .A1(n4981), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4975) );
  NAND2_X1 U6419 ( .A1(n4982), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U6420 ( .A1(n4997), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U6421 ( .A1(n6216), .A2(SI_0_), .ZN(n4977) );
  XNOR2_X1 U6422 ( .A(n4977), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8723) );
  MUX2_X1 U6423 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8723), .S(n6283), .Z(n9715) );
  NAND2_X1 U6424 ( .A1(n5369), .A2(n9715), .ZN(n8580) );
  NAND2_X1 U6425 ( .A1(n8069), .A2(n8580), .ZN(n8579) );
  NAND2_X1 U6426 ( .A1(n4978), .A2(n4979), .ZN(n4980) );
  NAND2_X1 U6427 ( .A1(n8579), .A2(n4980), .ZN(n8574) );
  NAND2_X1 U6428 ( .A1(n4996), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U6429 ( .A1(n4981), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U6430 ( .A1(n4982), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6431 ( .A1(n4997), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n4983) );
  INV_X1 U6432 ( .A(n4994), .ZN(n8315) );
  OR2_X1 U6433 ( .A1(n4987), .A2(n5415), .ZN(n4988) );
  XNOR2_X1 U6434 ( .A(n4988), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9358) );
  INV_X1 U6435 ( .A(n9358), .ZN(n6230) );
  OR2_X1 U6436 ( .A1(n4989), .A2(n6232), .ZN(n4993) );
  XNOR2_X1 U6437 ( .A(n4991), .B(n4990), .ZN(n6231) );
  OR2_X1 U6438 ( .A1(n5050), .A2(n6231), .ZN(n4992) );
  OAI211_X2 U6439 ( .C1(n6283), .C2(n6230), .A(n4993), .B(n4992), .ZN(n8575)
         );
  NAND2_X1 U6440 ( .A1(n8574), .A2(n5371), .ZN(n8573) );
  NAND2_X1 U6441 ( .A1(n4994), .A2(n9731), .ZN(n4995) );
  NAND2_X1 U6442 ( .A1(n8573), .A2(n4995), .ZN(n6547) );
  NAND2_X1 U6443 ( .A1(n4996), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4999) );
  INV_X1 U6444 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U6445 ( .A1(n4997), .A2(n6343), .ZN(n4998) );
  NAND2_X1 U6446 ( .A1(n4981), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U6447 ( .A1(n5343), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5000) );
  XNOR2_X1 U6448 ( .A(n5003), .B(n5002), .ZN(n6221) );
  OR2_X1 U6449 ( .A1(n5050), .A2(n6221), .ZN(n5009) );
  OR2_X1 U6450 ( .A1(n7899), .A2(n9822), .ZN(n5008) );
  INV_X1 U6451 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U6452 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5004), .ZN(n5005) );
  XNOR2_X1 U6453 ( .A(n5006), .B(n5005), .ZN(n6347) );
  OR2_X1 U6454 ( .A1(n6283), .A2(n6347), .ZN(n5007) );
  XNOR2_X1 U6455 ( .A(n8314), .B(n5475), .ZN(n6546) );
  NAND2_X1 U6456 ( .A1(n6547), .A2(n6546), .ZN(n6545) );
  INV_X1 U6457 ( .A(n8314), .ZN(n7939) );
  NAND2_X1 U6458 ( .A1(n7939), .A2(n5475), .ZN(n5010) );
  NAND2_X1 U6459 ( .A1(n5354), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5016) );
  NAND2_X1 U6460 ( .A1(n4981), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5015) );
  INV_X1 U6461 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U6462 ( .A1(n6343), .A2(n6356), .ZN(n5012) );
  AND2_X1 U6463 ( .A1(n5012), .A2(n5026), .ZN(n6841) );
  NAND2_X1 U6464 ( .A1(n4264), .A2(n6841), .ZN(n5014) );
  NAND2_X1 U6465 ( .A1(n5343), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U6466 ( .A1(n5017), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5018) );
  XNOR2_X1 U6467 ( .A(n5018), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6292) );
  INV_X1 U6468 ( .A(n6292), .ZN(n6360) );
  XNOR2_X1 U6469 ( .A(n5020), .B(n5019), .ZN(n6219) );
  OR2_X1 U6470 ( .A1(n5050), .A2(n6219), .ZN(n5022) );
  OR2_X1 U6471 ( .A1(n7899), .A2(n6215), .ZN(n5021) );
  OAI211_X1 U6472 ( .C1(n6283), .C2(n6360), .A(n5022), .B(n5021), .ZN(n6644)
         );
  NAND2_X1 U6473 ( .A1(n5023), .A2(n6644), .ZN(n7914) );
  INV_X1 U6474 ( .A(n5023), .ZN(n8313) );
  INV_X1 U6475 ( .A(n6644), .ZN(n6844) );
  NAND2_X1 U6476 ( .A1(n8313), .A2(n6844), .ZN(n6814) );
  NAND2_X1 U6477 ( .A1(n5023), .A2(n6844), .ZN(n5024) );
  NAND2_X1 U6478 ( .A1(n4996), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U6479 ( .A1(n6260), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5030) );
  AND2_X1 U6480 ( .A1(n5026), .A2(n5025), .ZN(n5027) );
  NOR2_X1 U6481 ( .A1(n5039), .A2(n5027), .ZN(n6630) );
  NAND2_X1 U6482 ( .A1(n4264), .A2(n6630), .ZN(n5029) );
  NAND2_X1 U6483 ( .A1(n6261), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U6484 ( .A1(n5032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5033) );
  XNOR2_X1 U6485 ( .A(n5033), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6290) );
  INV_X1 U6486 ( .A(n6290), .ZN(n6319) );
  OR2_X1 U6487 ( .A1(n7899), .A2(n6223), .ZN(n5036) );
  NAND2_X1 U6488 ( .A1(n6726), .A2(n6821), .ZN(n7912) );
  INV_X1 U6489 ( .A(n6821), .ZN(n9737) );
  NAND2_X1 U6490 ( .A1(n7912), .A2(n7936), .ZN(n8073) );
  NAND2_X1 U6491 ( .A1(n6726), .A2(n9737), .ZN(n5037) );
  NAND2_X1 U6492 ( .A1(n5038), .A2(n5037), .ZN(n6874) );
  NAND2_X1 U6493 ( .A1(n4981), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5047) );
  INV_X1 U6494 ( .A(n5039), .ZN(n5041) );
  INV_X1 U6495 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U6496 ( .A1(n5041), .A2(n5040), .ZN(n5042) );
  NAND2_X1 U6497 ( .A1(n5055), .A2(n5042), .ZN(n6878) );
  INV_X1 U6498 ( .A(n6878), .ZN(n5043) );
  NAND2_X1 U6499 ( .A1(n4263), .A2(n5043), .ZN(n5046) );
  NAND2_X1 U6500 ( .A1(n4996), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U6501 ( .A1(n5343), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5044) );
  NAND4_X1 U6502 ( .A1(n5047), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n8311)
         );
  NOR2_X1 U6503 ( .A1(n5032), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5081) );
  OR2_X1 U6504 ( .A1(n5081), .A2(n5415), .ZN(n5062) );
  XNOR2_X1 U6505 ( .A(n5062), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6326) );
  INV_X1 U6506 ( .A(n6326), .ZN(n6307) );
  OR2_X1 U6507 ( .A1(n5050), .A2(n6224), .ZN(n5052) );
  OR2_X1 U6508 ( .A1(n7899), .A2(n9820), .ZN(n5051) );
  NAND2_X1 U6509 ( .A1(n8311), .A2(n6888), .ZN(n5053) );
  NAND2_X1 U6510 ( .A1(n5354), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6511 ( .A1(n6260), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6512 ( .A1(n5055), .A2(n5054), .ZN(n5056) );
  AND2_X1 U6513 ( .A1(n5071), .A2(n5056), .ZN(n6762) );
  NAND2_X1 U6514 ( .A1(n4264), .A2(n6762), .ZN(n5058) );
  NAND2_X1 U6515 ( .A1(n6261), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U6516 ( .A1(n5062), .A2(n5061), .ZN(n5063) );
  NAND2_X1 U6517 ( .A1(n5063), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5064) );
  XNOR2_X1 U6518 ( .A(n5064), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6460) );
  AOI22_X1 U6519 ( .A1(n5223), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n4560), .B2(
        n6460), .ZN(n5068) );
  XNOR2_X1 U6520 ( .A(n5066), .B(n5065), .ZN(n6233) );
  NAND2_X1 U6521 ( .A1(n6233), .A2(n4450), .ZN(n5067) );
  NAND2_X1 U6522 ( .A1(n5068), .A2(n5067), .ZN(n6743) );
  NAND2_X1 U6523 ( .A1(n6851), .A2(n6743), .ZN(n7947) );
  INV_X1 U6524 ( .A(n6851), .ZN(n8310) );
  NAND2_X1 U6525 ( .A1(n8310), .A2(n6797), .ZN(n7948) );
  NAND2_X1 U6526 ( .A1(n6851), .A2(n6797), .ZN(n5069) );
  INV_X1 U6527 ( .A(n6918), .ZN(n5086) );
  NAND2_X1 U6528 ( .A1(n6260), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U6529 ( .A1(n5071), .A2(n5070), .ZN(n5072) );
  NAND2_X1 U6530 ( .A1(n5094), .A2(n5072), .ZN(n6927) );
  INV_X1 U6531 ( .A(n6927), .ZN(n5073) );
  NAND2_X1 U6532 ( .A1(n4264), .A2(n5073), .ZN(n5076) );
  NAND2_X1 U6533 ( .A1(n5354), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6534 ( .A1(n5343), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5074) );
  NAND4_X1 U6535 ( .A1(n5077), .A2(n5076), .A3(n5075), .A4(n5074), .ZN(n8309)
         );
  XNOR2_X1 U6536 ( .A(n5079), .B(n5078), .ZN(n6237) );
  NAND2_X1 U6537 ( .A1(n6237), .A2(n4450), .ZN(n5084) );
  NOR2_X1 U6538 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5080) );
  NAND2_X1 U6539 ( .A1(n5081), .A2(n5080), .ZN(n5089) );
  NAND2_X1 U6540 ( .A1(n5089), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5082) );
  XNOR2_X1 U6541 ( .A(n5082), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6459) );
  AOI22_X1 U6542 ( .A1(n5223), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4560), .B2(
        n6459), .ZN(n5083) );
  XNOR2_X1 U6543 ( .A(n8309), .B(n6935), .ZN(n8075) );
  NAND2_X1 U6544 ( .A1(n6935), .A2(n8309), .ZN(n5087) );
  XNOR2_X1 U6545 ( .A(n5088), .B(n4785), .ZN(n6246) );
  NAND2_X1 U6546 ( .A1(n6246), .A2(n7898), .ZN(n5092) );
  NAND2_X1 U6547 ( .A1(n5101), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5090) );
  XNOR2_X1 U6548 ( .A(n5090), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6606) );
  AOI22_X1 U6549 ( .A1(n5223), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4560), .B2(
        n6606), .ZN(n5091) );
  NAND2_X1 U6550 ( .A1(n5092), .A2(n5091), .ZN(n7360) );
  NAND2_X1 U6551 ( .A1(n6260), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6552 ( .A1(n6261), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U6553 ( .A1(n5094), .A2(n5093), .ZN(n5095) );
  AND2_X1 U6554 ( .A1(n5105), .A2(n5095), .ZN(n7177) );
  NAND2_X1 U6555 ( .A1(n4264), .A2(n7177), .ZN(n5097) );
  NAND2_X1 U6556 ( .A1(n5354), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5096) );
  OR2_X1 U6557 ( .A1(n7360), .A2(n7015), .ZN(n7963) );
  NAND2_X1 U6558 ( .A1(n7360), .A2(n7015), .ZN(n7960) );
  NAND2_X1 U6559 ( .A1(n6251), .A2(n7898), .ZN(n5104) );
  NAND2_X1 U6560 ( .A1(n5113), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5102) );
  XNOR2_X1 U6561 ( .A(n5102), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6661) );
  AOI22_X1 U6562 ( .A1(n5223), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4560), .B2(
        n6661), .ZN(n5103) );
  NAND2_X1 U6563 ( .A1(n6260), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6564 ( .A1(n5354), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5109) );
  INV_X1 U6565 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U6566 ( .A1(n5105), .A2(n6595), .ZN(n5106) );
  AND2_X1 U6567 ( .A1(n5118), .A2(n5106), .ZN(n7014) );
  NAND2_X1 U6568 ( .A1(n4264), .A2(n7014), .ZN(n5108) );
  NAND2_X1 U6569 ( .A1(n6261), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5107) );
  INV_X1 U6570 ( .A(n7033), .ZN(n8307) );
  AND2_X1 U6571 ( .A1(n7103), .A2(n8307), .ZN(n5124) );
  XNOR2_X1 U6572 ( .A(n5112), .B(n5111), .ZN(n6255) );
  NAND2_X1 U6573 ( .A1(n6255), .A2(n7898), .ZN(n5116) );
  OAI21_X1 U6574 ( .B1(n5113), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5114) );
  XNOR2_X1 U6575 ( .A(n5114), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6895) );
  AOI22_X1 U6576 ( .A1(n5223), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4560), .B2(
        n6895), .ZN(n5115) );
  NAND2_X1 U6577 ( .A1(n5116), .A2(n5115), .ZN(n8669) );
  NAND2_X1 U6578 ( .A1(n6260), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6579 ( .A1(n6261), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6580 ( .A1(n5118), .A2(n5117), .ZN(n5119) );
  AND2_X1 U6581 ( .A1(n5133), .A2(n5119), .ZN(n7155) );
  NAND2_X1 U6582 ( .A1(n4264), .A2(n7155), .ZN(n5121) );
  NAND2_X1 U6583 ( .A1(n5354), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5120) );
  OR2_X1 U6584 ( .A1(n8669), .A2(n7075), .ZN(n7966) );
  NAND2_X1 U6585 ( .A1(n8669), .A2(n7075), .ZN(n7957) );
  NAND2_X1 U6586 ( .A1(n7966), .A2(n7957), .ZN(n7159) );
  OR2_X1 U6587 ( .A1(n7103), .A2(n7033), .ZN(n7965) );
  NAND2_X1 U6588 ( .A1(n7103), .A2(n7033), .ZN(n7962) );
  NAND2_X1 U6589 ( .A1(n7965), .A2(n7962), .ZN(n8079) );
  INV_X1 U6590 ( .A(n7015), .ZN(n8308) );
  OR2_X1 U6591 ( .A1(n7360), .A2(n8308), .ZN(n7087) );
  AND2_X1 U6592 ( .A1(n8079), .A2(n7087), .ZN(n7088) );
  AND2_X1 U6593 ( .A1(n7159), .A2(n7149), .ZN(n5125) );
  NAND2_X1 U6594 ( .A1(n7150), .A2(n5125), .ZN(n5127) );
  INV_X1 U6595 ( .A(n7075), .ZN(n8306) );
  NAND2_X1 U6596 ( .A1(n8669), .A2(n8306), .ZN(n5126) );
  XNOR2_X1 U6597 ( .A(n5129), .B(n5128), .ZN(n6267) );
  NAND2_X1 U6598 ( .A1(n6267), .A2(n7898), .ZN(n5132) );
  OR2_X1 U6599 ( .A1(n4959), .A2(n5415), .ZN(n5130) );
  XNOR2_X1 U6600 ( .A(n5130), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6996) );
  AOI22_X1 U6601 ( .A1(n5223), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n4560), .B2(
        n6996), .ZN(n5131) );
  NAND2_X1 U6602 ( .A1(n6260), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6603 ( .A1(n5354), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5137) );
  INV_X1 U6604 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6900) );
  NAND2_X1 U6605 ( .A1(n5133), .A2(n6900), .ZN(n5134) );
  AND2_X1 U6606 ( .A1(n5144), .A2(n5134), .ZN(n7205) );
  NAND2_X1 U6607 ( .A1(n4264), .A2(n7205), .ZN(n5136) );
  NAND2_X1 U6608 ( .A1(n5343), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5135) );
  NAND2_X1 U6609 ( .A1(n7210), .A2(n7218), .ZN(n7911) );
  INV_X1 U6610 ( .A(n7218), .ZN(n8305) );
  XNOR2_X1 U6611 ( .A(n5140), .B(n4786), .ZN(n6377) );
  NAND2_X1 U6612 ( .A1(n6377), .A2(n7898), .ZN(n5142) );
  OR2_X1 U6613 ( .A1(n5190), .A2(n5415), .ZN(n5154) );
  XNOR2_X1 U6614 ( .A(n5154), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7046) );
  AOI22_X1 U6615 ( .A1(n5223), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n4560), .B2(
        n7046), .ZN(n5141) );
  NAND2_X1 U6616 ( .A1(n6260), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6617 ( .A1(n5354), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6618 ( .A1(n5144), .A2(n5143), .ZN(n5145) );
  AND2_X1 U6619 ( .A1(n5162), .A2(n5145), .ZN(n7251) );
  NAND2_X1 U6620 ( .A1(n4264), .A2(n7251), .ZN(n5147) );
  NAND2_X1 U6621 ( .A1(n6261), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5146) );
  OR2_X1 U6622 ( .A1(n7250), .A2(n7277), .ZN(n7971) );
  NAND2_X1 U6623 ( .A1(n7250), .A2(n7277), .ZN(n7273) );
  INV_X1 U6624 ( .A(n7277), .ZN(n8304) );
  NAND2_X1 U6625 ( .A1(n7250), .A2(n8304), .ZN(n5150) );
  NAND2_X1 U6626 ( .A1(n7247), .A2(n5150), .ZN(n7270) );
  XNOR2_X1 U6627 ( .A(n5152), .B(n5151), .ZN(n6414) );
  NAND2_X1 U6628 ( .A1(n6414), .A2(n7898), .ZN(n5160) );
  NAND2_X1 U6629 ( .A1(n5154), .A2(n5153), .ZN(n5155) );
  NAND2_X1 U6630 ( .A1(n5155), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5157) );
  OR2_X1 U6631 ( .A1(n5157), .A2(n5156), .ZN(n5158) );
  NAND2_X1 U6632 ( .A1(n5157), .A2(n5156), .ZN(n5172) );
  AND2_X1 U6633 ( .A1(n5158), .A2(n5172), .ZN(n7258) );
  AOI22_X1 U6634 ( .A1(n5223), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n4560), .B2(
        n7258), .ZN(n5159) );
  NAND2_X1 U6635 ( .A1(n6260), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6636 ( .A1(n5354), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6637 ( .A1(n5162), .A2(n5161), .ZN(n5163) );
  AND2_X1 U6638 ( .A1(n5177), .A2(n5163), .ZN(n7415) );
  NAND2_X1 U6639 ( .A1(n4264), .A2(n7415), .ZN(n5165) );
  NAND2_X1 U6640 ( .A1(n5343), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5164) );
  NAND2_X1 U6641 ( .A1(n7421), .A2(n7388), .ZN(n7975) );
  INV_X1 U6642 ( .A(n7272), .ZN(n5168) );
  INV_X1 U6643 ( .A(n7388), .ZN(n8303) );
  OR2_X1 U6644 ( .A1(n7421), .A2(n8303), .ZN(n5169) );
  XNOR2_X1 U6645 ( .A(n5171), .B(n5170), .ZN(n6574) );
  NAND2_X1 U6646 ( .A1(n6574), .A2(n7898), .ZN(n5175) );
  NAND2_X1 U6647 ( .A1(n5172), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5173) );
  XNOR2_X1 U6648 ( .A(n5173), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7425) );
  AOI22_X1 U6649 ( .A1(n5223), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n4560), .B2(
        n7425), .ZN(n5174) );
  NAND2_X1 U6650 ( .A1(n6260), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6651 ( .A1(n6261), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5182) );
  INV_X1 U6652 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6653 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  AND2_X1 U6654 ( .A1(n5179), .A2(n5178), .ZN(n8279) );
  NAND2_X1 U6655 ( .A1(n4264), .A2(n8279), .ZN(n5181) );
  NAND2_X1 U6656 ( .A1(n5354), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6657 ( .A1(n8287), .A2(n7466), .ZN(n7981) );
  NAND2_X1 U6658 ( .A1(n7980), .A2(n7981), .ZN(n8086) );
  NAND2_X1 U6659 ( .A1(n7495), .A2(n7466), .ZN(n5184) );
  NAND2_X1 U6660 ( .A1(n7383), .A2(n5184), .ZN(n7469) );
  OR2_X1 U6661 ( .A1(n8715), .A2(n8206), .ZN(n7986) );
  NAND2_X1 U6662 ( .A1(n8715), .A2(n8206), .ZN(n7985) );
  NAND2_X1 U6663 ( .A1(n6593), .A2(n7898), .ZN(n5193) );
  INV_X1 U6664 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5187) );
  AND2_X1 U6665 ( .A1(n5188), .A2(n5187), .ZN(n5189) );
  NAND2_X1 U6666 ( .A1(n5204), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5191) );
  XNOR2_X1 U6667 ( .A(n5191), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8337) );
  AOI22_X1 U6668 ( .A1(n5223), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4560), .B2(
        n8337), .ZN(n5192) );
  NAND2_X1 U6669 ( .A1(n6260), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6670 ( .A1(n5343), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5199) );
  INV_X1 U6671 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6672 ( .A1(n5195), .A2(n5194), .ZN(n5196) );
  AND2_X1 U6673 ( .A1(n5209), .A2(n5196), .ZN(n8553) );
  NAND2_X1 U6674 ( .A1(n4264), .A2(n8553), .ZN(n5198) );
  NAND2_X1 U6675 ( .A1(n5354), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6676 ( .A1(n8552), .A2(n8253), .ZN(n7989) );
  NAND2_X1 U6677 ( .A1(n8527), .A2(n7989), .ZN(n8544) );
  INV_X1 U6678 ( .A(n8253), .ZN(n8301) );
  NAND2_X1 U6679 ( .A1(n6766), .A2(n7898), .ZN(n5207) );
  NAND2_X1 U6680 ( .A1(n5219), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5205) );
  XNOR2_X1 U6681 ( .A(n5205), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8342) );
  AOI22_X1 U6682 ( .A1(n5223), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4560), .B2(
        n8342), .ZN(n5206) );
  NAND2_X1 U6683 ( .A1(n5209), .A2(n5208), .ZN(n5210) );
  AND2_X1 U6684 ( .A1(n5238), .A2(n5210), .ZN(n8536) );
  NAND2_X1 U6685 ( .A1(n8536), .A2(n4264), .ZN(n5214) );
  NAND2_X1 U6686 ( .A1(n5354), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6687 ( .A1(n6260), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U6688 ( .A1(n6261), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5211) );
  NAND4_X1 U6689 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n8300)
         );
  NAND2_X1 U6690 ( .A1(n8535), .A2(n8300), .ZN(n5216) );
  INV_X1 U6691 ( .A(n8300), .ZN(n8166) );
  AOI21_X1 U6692 ( .B1(n8525), .B2(n5216), .A(n5215), .ZN(n8510) );
  XNOR2_X1 U6693 ( .A(n5218), .B(n5217), .ZN(n6808) );
  NAND2_X1 U6694 ( .A1(n6808), .A2(n7898), .ZN(n5225) );
  NAND2_X1 U6695 ( .A1(n5221), .A2(n5220), .ZN(n5362) );
  OR2_X1 U6696 ( .A1(n5221), .A2(n5220), .ZN(n5222) );
  AOI22_X1 U6697 ( .A1(n5223), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8417), .B2(
        n4560), .ZN(n5224) );
  INV_X1 U6698 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5230) );
  XNOR2_X1 U6699 ( .A(n5238), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U6700 ( .A1(n8518), .A2(n4264), .ZN(n5229) );
  NAND2_X1 U6701 ( .A1(n6260), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6702 ( .A1(n6261), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5226) );
  AND2_X1 U6703 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  OAI211_X1 U6704 ( .C1(n5011), .C2(n5230), .A(n5229), .B(n5228), .ZN(n8299)
         );
  NAND2_X1 U6705 ( .A1(n8510), .A2(n5231), .ZN(n5232) );
  INV_X1 U6706 ( .A(n8299), .ZN(n5384) );
  NAND2_X1 U6707 ( .A1(n5232), .A2(n4781), .ZN(n8494) );
  INV_X1 U6708 ( .A(n8494), .ZN(n5243) );
  XNOR2_X1 U6709 ( .A(n5234), .B(n5233), .ZN(n6972) );
  NAND2_X1 U6710 ( .A1(n6972), .A2(n7898), .ZN(n5236) );
  OR2_X1 U6711 ( .A1(n7899), .A2(n7512), .ZN(n5235) );
  INV_X1 U6712 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5237) );
  INV_X1 U6713 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8231) );
  OAI21_X1 U6714 ( .B1(n5238), .B2(n5237), .A(n8231), .ZN(n5239) );
  AND2_X1 U6715 ( .A1(n5248), .A2(n5239), .ZN(n8504) );
  NAND2_X1 U6716 ( .A1(n8504), .A2(n4264), .ZN(n5242) );
  AOI22_X1 U6717 ( .A1(n5354), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n6260), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6718 ( .A1(n6261), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6719 ( .A1(n8503), .A2(n8173), .ZN(n8005) );
  NAND2_X1 U6720 ( .A1(n8008), .A2(n8005), .ZN(n8497) );
  INV_X1 U6721 ( .A(n8173), .ZN(n8298) );
  OAI21_X1 U6722 ( .B1(n5243), .B2(n5386), .A(n4797), .ZN(n8478) );
  XNOR2_X1 U6723 ( .A(n5245), .B(n5244), .ZN(n7005) );
  NAND2_X1 U6724 ( .A1(n7005), .A2(n7898), .ZN(n5247) );
  OR2_X1 U6725 ( .A1(n7899), .A2(n7009), .ZN(n5246) );
  INV_X1 U6726 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9845) );
  NAND2_X1 U6727 ( .A1(n5248), .A2(n9845), .ZN(n5249) );
  AND2_X1 U6728 ( .A1(n5258), .A2(n5249), .ZN(n8488) );
  NAND2_X1 U6729 ( .A1(n8488), .A2(n4264), .ZN(n5252) );
  AOI22_X1 U6730 ( .A1(n5354), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n6260), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6731 ( .A1(n6261), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5250) );
  INV_X1 U6732 ( .A(n8244), .ZN(n8297) );
  OAI22_X1 U6733 ( .A1(n8478), .A2(n5253), .B1(n8297), .B2(n8487), .ZN(n8464)
         );
  XNOR2_X1 U6734 ( .A(n5255), .B(n5254), .ZN(n7055) );
  NAND2_X1 U6735 ( .A1(n7055), .A2(n7898), .ZN(n5257) );
  OR2_X1 U6736 ( .A1(n7899), .A2(n7058), .ZN(n5256) );
  INV_X1 U6737 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8247) );
  NAND2_X1 U6738 ( .A1(n5258), .A2(n8247), .ZN(n5259) );
  NAND2_X1 U6739 ( .A1(n5273), .A2(n5259), .ZN(n8241) );
  OR2_X1 U6740 ( .A1(n8241), .A2(n5329), .ZN(n5265) );
  INV_X1 U6741 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6742 ( .A1(n6260), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U6743 ( .A1(n5343), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5260) );
  OAI211_X1 U6744 ( .C1(n5262), .C2(n5011), .A(n5261), .B(n5260), .ZN(n5263)
         );
  INV_X1 U6745 ( .A(n5263), .ZN(n5264) );
  NAND2_X1 U6746 ( .A1(n8471), .A2(n8156), .ZN(n8011) );
  NAND2_X1 U6747 ( .A1(n8015), .A2(n8011), .ZN(n8463) );
  INV_X1 U6748 ( .A(n8471), .ZN(n8692) );
  AOI22_X1 U6749 ( .A1(n8464), .A2(n8463), .B1(n8156), .B2(n8692), .ZN(n8453)
         );
  OR2_X1 U6750 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  NAND2_X1 U6751 ( .A1(n5269), .A2(n5268), .ZN(n7146) );
  NAND2_X1 U6752 ( .A1(n7146), .A2(n7898), .ZN(n5271) );
  OR2_X1 U6753 ( .A1(n7899), .A2(n7148), .ZN(n5270) );
  NAND2_X1 U6754 ( .A1(n5273), .A2(n5272), .ZN(n5274) );
  AND2_X1 U6755 ( .A1(n5275), .A2(n5274), .ZN(n8455) );
  INV_X1 U6756 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6757 ( .A1(n6260), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6758 ( .A1(n5354), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5276) );
  OAI211_X1 U6759 ( .C1(n5357), .C2(n5278), .A(n5277), .B(n5276), .ZN(n5279)
         );
  AOI21_X1 U6760 ( .B1(n8455), .B2(n4264), .A(n5279), .ZN(n8243) );
  NAND2_X1 U6761 ( .A1(n8620), .A2(n8157), .ZN(n8021) );
  INV_X1 U6762 ( .A(n5280), .ZN(n5284) );
  INV_X1 U6763 ( .A(n5281), .ZN(n5282) );
  NAND2_X1 U6764 ( .A1(n5282), .A2(SI_24_), .ZN(n5283) );
  INV_X1 U6765 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7401) );
  INV_X1 U6766 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7404) );
  MUX2_X1 U6767 ( .A(n7401), .B(n7404), .S(n7538), .Z(n5286) );
  INV_X1 U6768 ( .A(SI_25_), .ZN(n9836) );
  NAND2_X1 U6769 ( .A1(n5286), .A2(n9836), .ZN(n5297) );
  INV_X1 U6770 ( .A(n5286), .ZN(n5287) );
  NAND2_X1 U6771 ( .A1(n5287), .A2(SI_25_), .ZN(n5288) );
  NAND2_X1 U6772 ( .A1(n5297), .A2(n5288), .ZN(n5298) );
  NAND2_X1 U6773 ( .A1(n7399), .A2(n7898), .ZN(n5290) );
  OR2_X1 U6774 ( .A1(n7899), .A2(n7401), .ZN(n5289) );
  INV_X1 U6775 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8185) );
  NAND2_X1 U6776 ( .A1(n5291), .A2(n8185), .ZN(n5292) );
  AND2_X1 U6777 ( .A1(n5309), .A2(n5292), .ZN(n8428) );
  INV_X1 U6778 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6779 ( .A1(n5343), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6780 ( .A1(n4981), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5293) );
  OAI211_X1 U6781 ( .C1(n5011), .C2(n5295), .A(n5294), .B(n5293), .ZN(n5296)
         );
  AOI21_X1 U6782 ( .B1(n8428), .B2(n4264), .A(n5296), .ZN(n8265) );
  NAND2_X1 U6783 ( .A1(n8616), .A2(n8265), .ZN(n8028) );
  INV_X1 U6784 ( .A(n8265), .ZN(n8294) );
  OAI22_X1 U6785 ( .A1(n8423), .A2(n8424), .B1(n8294), .B2(n8616), .ZN(n8406)
         );
  INV_X1 U6786 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9806) );
  INV_X1 U6787 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7483) );
  MUX2_X1 U6788 ( .A(n9806), .B(n7483), .S(n7538), .Z(n5301) );
  INV_X1 U6789 ( .A(SI_26_), .ZN(n5300) );
  NAND2_X1 U6790 ( .A1(n5301), .A2(n5300), .ZN(n5315) );
  INV_X1 U6791 ( .A(n5301), .ZN(n5302) );
  NAND2_X1 U6792 ( .A1(n5302), .A2(SI_26_), .ZN(n5303) );
  AND2_X1 U6793 ( .A1(n5315), .A2(n5303), .ZN(n5304) );
  OR2_X1 U6794 ( .A1(n5305), .A2(n5304), .ZN(n5306) );
  NAND2_X1 U6795 ( .A1(n5316), .A2(n5306), .ZN(n7479) );
  NAND2_X1 U6796 ( .A1(n7479), .A2(n7898), .ZN(n5308) );
  OR2_X1 U6797 ( .A1(n7899), .A2(n9806), .ZN(n5307) );
  INV_X1 U6798 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8268) );
  NAND2_X1 U6799 ( .A1(n5309), .A2(n8268), .ZN(n5310) );
  INV_X1 U6800 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6801 ( .A1(n5354), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U6802 ( .A1(n4981), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5311) );
  OAI211_X1 U6803 ( .C1(n5313), .C2(n5357), .A(n5312), .B(n5311), .ZN(n5314)
         );
  AOI21_X1 U6804 ( .B1(n8415), .B2(n4264), .A(n5314), .ZN(n8182) );
  OR2_X1 U6805 ( .A1(n8611), .A2(n8182), .ZN(n8034) );
  NAND2_X1 U6806 ( .A1(n8611), .A2(n8182), .ZN(n8035) );
  NAND2_X1 U6807 ( .A1(n8034), .A2(n8035), .ZN(n8068) );
  INV_X1 U6808 ( .A(n8611), .ZN(n8275) );
  AOI22_X1 U6809 ( .A1(n8406), .A2(n8068), .B1(n8275), .B2(n8182), .ZN(n8389)
         );
  INV_X1 U6810 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9869) );
  INV_X1 U6811 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7561) );
  MUX2_X1 U6812 ( .A(n9869), .B(n7561), .S(n7538), .Z(n5318) );
  INV_X1 U6813 ( .A(SI_27_), .ZN(n5317) );
  NAND2_X1 U6814 ( .A1(n5318), .A2(n5317), .ZN(n5336) );
  INV_X1 U6815 ( .A(n5318), .ZN(n5319) );
  NAND2_X1 U6816 ( .A1(n5319), .A2(SI_27_), .ZN(n5320) );
  AND2_X1 U6817 ( .A1(n5336), .A2(n5320), .ZN(n5321) );
  OR2_X1 U6818 ( .A1(n5322), .A2(n5321), .ZN(n5323) );
  NAND2_X1 U6819 ( .A1(n5337), .A2(n5323), .ZN(n7560) );
  NAND2_X1 U6820 ( .A1(n7560), .A2(n7898), .ZN(n5325) );
  OR2_X1 U6821 ( .A1(n7899), .A2(n9869), .ZN(n5324) );
  INV_X1 U6822 ( .A(n5327), .ZN(n5326) );
  NAND2_X1 U6823 ( .A1(n5326), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5341) );
  INV_X1 U6824 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9934) );
  NAND2_X1 U6825 ( .A1(n5327), .A2(n9934), .ZN(n5328) );
  NAND2_X1 U6826 ( .A1(n5341), .A2(n5328), .ZN(n8399) );
  INV_X1 U6827 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6828 ( .A1(n5354), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6829 ( .A1(n6260), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5330) );
  OAI211_X1 U6830 ( .C1(n5332), .C2(n5357), .A(n5331), .B(n5330), .ZN(n5333)
         );
  INV_X1 U6831 ( .A(n5333), .ZN(n5334) );
  OAI22_X1 U6832 ( .A1(n8389), .A2(n8391), .B1(n8606), .B2(n8293), .ZN(n5445)
         );
  MUX2_X1 U6833 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7538), .Z(n5349) );
  INV_X1 U6834 ( .A(SI_28_), .ZN(n9800) );
  XNOR2_X1 U6835 ( .A(n5349), .B(n9800), .ZN(n5347) );
  NAND2_X1 U6836 ( .A1(n7555), .A2(n7898), .ZN(n5339) );
  INV_X1 U6837 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7499) );
  OR2_X1 U6838 ( .A1(n7899), .A2(n7499), .ZN(n5338) );
  INV_X1 U6839 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6840 ( .A1(n5341), .A2(n5340), .ZN(n5342) );
  INV_X1 U6841 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U6842 ( .A1(n5354), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U6843 ( .A1(n5343), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5344) );
  OAI211_X1 U6844 ( .C1(n5398), .C2(n9834), .A(n5345), .B(n5344), .ZN(n5346)
         );
  AOI21_X1 U6845 ( .B1(n8380), .B2(n4264), .A(n5346), .ZN(n8149) );
  NAND2_X1 U6846 ( .A1(n8044), .A2(n8149), .ZN(n8037) );
  INV_X1 U6847 ( .A(n5349), .ZN(n5350) );
  INV_X1 U6848 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9866) );
  INV_X1 U6849 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9350) );
  MUX2_X1 U6850 ( .A(n9866), .B(n9350), .S(n7538), .Z(n7514) );
  XNOR2_X1 U6851 ( .A(n7514), .B(SI_29_), .ZN(n5351) );
  NAND2_X1 U6852 ( .A1(n8113), .A2(n7898), .ZN(n5353) );
  OR2_X1 U6853 ( .A1(n7899), .A2(n9866), .ZN(n5352) );
  INV_X1 U6854 ( .A(n7881), .ZN(n5360) );
  INV_X1 U6855 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6856 ( .A1(n5354), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6857 ( .A1(n6260), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5355) );
  OAI211_X1 U6858 ( .C1(n5441), .C2(n5357), .A(n5356), .B(n5355), .ZN(n5358)
         );
  AOI21_X1 U6859 ( .B1(n5360), .B2(n4264), .A(n5358), .ZN(n6771) );
  XNOR2_X1 U6860 ( .A(n5361), .B(n8094), .ZN(n7879) );
  NAND2_X1 U6861 ( .A1(n5362), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6862 ( .A1(n4300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5365) );
  XNOR2_X1 U6863 ( .A(n5365), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U6864 ( .A1(n5430), .A2(n7925), .ZN(n6699) );
  NAND2_X1 U6865 ( .A1(n5366), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5419) );
  XNOR2_X1 U6866 ( .A(n5419), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8109) );
  XNOR2_X1 U6867 ( .A(n6699), .B(n8109), .ZN(n5367) );
  NAND2_X1 U6868 ( .A1(n5367), .A2(n8357), .ZN(n7170) );
  NOR2_X1 U6869 ( .A1(n8357), .A2(n8109), .ZN(n5368) );
  NAND2_X1 U6870 ( .A1(n5430), .A2(n5368), .ZN(n9748) );
  NAND2_X1 U6871 ( .A1(n7170), .A2(n9748), .ZN(n9746) );
  INV_X1 U6872 ( .A(n5369), .ZN(n5370) );
  NAND2_X1 U6873 ( .A1(n5370), .A2(n9715), .ZN(n8583) );
  NAND2_X1 U6874 ( .A1(n7919), .A2(n8583), .ZN(n7923) );
  NAND2_X1 U6875 ( .A1(n7923), .A2(n7927), .ZN(n8562) );
  INV_X1 U6876 ( .A(n8562), .ZN(n5373) );
  INV_X1 U6877 ( .A(n5371), .ZN(n5372) );
  NAND2_X1 U6878 ( .A1(n5373), .A2(n5372), .ZN(n8561) );
  NAND2_X1 U6879 ( .A1(n8561), .A2(n7928), .ZN(n6550) );
  INV_X1 U6880 ( .A(n6546), .ZN(n6548) );
  NAND2_X1 U6881 ( .A1(n6550), .A2(n6548), .ZN(n6549) );
  INV_X1 U6882 ( .A(n5475), .ZN(n7938) );
  NAND2_X1 U6883 ( .A1(n7939), .A2(n7938), .ZN(n7913) );
  NAND2_X1 U6884 ( .A1(n5374), .A2(n7912), .ZN(n6881) );
  INV_X1 U6885 ( .A(n8311), .ZN(n6735) );
  NAND2_X1 U6886 ( .A1(n6735), .A2(n6888), .ZN(n7946) );
  NAND2_X1 U6887 ( .A1(n8311), .A2(n9743), .ZN(n7944) );
  AND2_X1 U6888 ( .A1(n7946), .A2(n7944), .ZN(n6883) );
  INV_X1 U6889 ( .A(n7947), .ZN(n5375) );
  INV_X1 U6890 ( .A(n6935), .ZN(n9751) );
  NAND2_X1 U6891 ( .A1(n7166), .A2(n7963), .ZN(n5376) );
  NAND2_X1 U6892 ( .A1(n5376), .A2(n7960), .ZN(n7084) );
  NAND2_X1 U6893 ( .A1(n7084), .A2(n7965), .ZN(n7158) );
  NAND2_X1 U6894 ( .A1(n7158), .A2(n7962), .ZN(n5377) );
  INV_X1 U6895 ( .A(n7159), .ZN(n8082) );
  NAND2_X1 U6896 ( .A1(n5377), .A2(n8082), .ZN(n7072) );
  AND2_X1 U6897 ( .A1(n7911), .A2(n7957), .ZN(n7968) );
  INV_X1 U6898 ( .A(n7273), .ZN(n7972) );
  NOR2_X1 U6899 ( .A1(n5168), .A2(n7972), .ZN(n5378) );
  NAND2_X1 U6900 ( .A1(n7242), .A2(n5378), .ZN(n7271) );
  NAND2_X1 U6901 ( .A1(n7271), .A2(n7976), .ZN(n7386) );
  INV_X1 U6902 ( .A(n8086), .ZN(n7978) );
  NAND2_X1 U6903 ( .A1(n7386), .A2(n7978), .ZN(n7385) );
  NAND2_X1 U6904 ( .A1(n7385), .A2(n7980), .ZN(n7463) );
  INV_X1 U6905 ( .A(n7463), .ZN(n5379) );
  INV_X1 U6906 ( .A(n7983), .ZN(n8087) );
  OR2_X1 U6907 ( .A1(n8535), .A2(n8166), .ZN(n7993) );
  NAND2_X1 U6908 ( .A1(n8535), .A2(n8166), .ZN(n7997) );
  NAND2_X1 U6909 ( .A1(n7993), .A2(n7997), .ZN(n8524) );
  INV_X1 U6910 ( .A(n8527), .ZN(n5381) );
  NOR2_X1 U6911 ( .A1(n8524), .A2(n5381), .ZN(n5382) );
  NAND2_X1 U6912 ( .A1(n5383), .A2(n7997), .ZN(n8511) );
  OR2_X1 U6913 ( .A1(n8517), .A2(n5384), .ZN(n8001) );
  NAND2_X1 U6914 ( .A1(n8517), .A2(n5384), .ZN(n7998) );
  INV_X1 U6915 ( .A(n8481), .ZN(n5389) );
  XNOR2_X1 U6916 ( .A(n8487), .B(n8244), .ZN(n8480) );
  NAND2_X1 U6917 ( .A1(n8487), .A2(n8244), .ZN(n8010) );
  INV_X1 U6918 ( .A(n8010), .ZN(n5387) );
  INV_X1 U6919 ( .A(n8463), .ZN(n8467) );
  NAND2_X1 U6920 ( .A1(n8466), .A2(n8467), .ZN(n8465) );
  NAND2_X1 U6921 ( .A1(n8465), .A2(n8015), .ZN(n8449) );
  NAND2_X1 U6922 ( .A1(n8626), .A2(n8243), .ZN(n8020) );
  OAI21_X2 U6923 ( .B1(n8449), .B2(n8452), .A(n8020), .ZN(n8442) );
  INV_X1 U6924 ( .A(n5390), .ZN(n8023) );
  INV_X1 U6925 ( .A(n8408), .ZN(n8030) );
  INV_X1 U6926 ( .A(n8035), .ZN(n5391) );
  NAND2_X1 U6927 ( .A1(n8403), .A2(n8293), .ZN(n8040) );
  XNOR2_X1 U6928 ( .A(n7889), .B(n8094), .ZN(n5401) );
  INV_X1 U6929 ( .A(n5430), .ZN(n5463) );
  NAND2_X1 U6930 ( .A1(n5463), .A2(n7925), .ZN(n7908) );
  NAND2_X1 U6931 ( .A1(n7908), .A2(n8064), .ZN(n8585) );
  INV_X1 U6932 ( .A(n8149), .ZN(n8292) );
  INV_X1 U6933 ( .A(n6288), .ZN(n5393) );
  AND2_X1 U6934 ( .A1(n8109), .A2(n7925), .ZN(n6279) );
  AND2_X1 U6935 ( .A1(n6288), .A2(n6279), .ZN(n8267) );
  INV_X1 U6936 ( .A(n5394), .ZN(n8106) );
  NAND2_X1 U6937 ( .A1(n8106), .A2(P2_B_REG_SCAN_IN), .ZN(n5395) );
  AND2_X1 U6938 ( .A1(n8267), .A2(n5395), .ZN(n8366) );
  INV_X1 U6939 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U6940 ( .A1(n4996), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6941 ( .A1(n6261), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5396) );
  OAI211_X1 U6942 ( .C1(n5398), .C2(n9830), .A(n5397), .B(n5396), .ZN(n8291)
         );
  NAND2_X1 U6943 ( .A1(n6553), .A2(n5475), .ZN(n6643) );
  INV_X1 U6944 ( .A(n8669), .ZN(n7157) );
  NAND2_X1 U6945 ( .A1(n7091), .A2(n7157), .ZN(n7152) );
  INV_X1 U6946 ( .A(n7421), .ZN(n7452) );
  NAND2_X1 U6947 ( .A1(n7391), .A2(n7495), .ZN(n7472) );
  OR2_X2 U6948 ( .A1(n7472), .A2(n8715), .ZN(n8551) );
  NAND2_X1 U6949 ( .A1(n8470), .A2(n8457), .ZN(n8454) );
  INV_X1 U6950 ( .A(n8109), .ZN(n7056) );
  NAND2_X1 U6951 ( .A1(n5430), .A2(n9716), .ZN(n9752) );
  OAI211_X1 U6952 ( .C1(n4440), .C2(n4291), .A(n8374), .B(n8670), .ZN(n7882)
         );
  NAND2_X1 U6953 ( .A1(n7888), .A2(n7882), .ZN(n5403) );
  AOI21_X1 U6954 ( .B1(n7879), .B2(n9746), .A(n5403), .ZN(n5444) );
  NOR4_X1 U6955 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5407) );
  NOR4_X1 U6956 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5406) );
  NOR4_X1 U6957 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n5405) );
  NOR4_X1 U6958 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5404) );
  AND4_X1 U6959 ( .A1(n5407), .A2(n5406), .A3(n5405), .A4(n5404), .ZN(n5429)
         );
  NOR2_X1 U6960 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .ZN(
        n9923) );
  NOR4_X1 U6961 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5410) );
  NOR4_X1 U6962 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5409) );
  NOR4_X1 U6963 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n5408) );
  AND4_X1 U6964 ( .A1(n9923), .A2(n5410), .A3(n5409), .A4(n5408), .ZN(n5428)
         );
  NAND2_X1 U6965 ( .A1(n5411), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5412) );
  XNOR2_X1 U6966 ( .A(n5412), .B(n4736), .ZN(n7480) );
  INV_X1 U6967 ( .A(n7480), .ZN(n5427) );
  NOR2_X1 U6968 ( .A1(n5413), .A2(n5415), .ZN(n5414) );
  MUX2_X1 U6969 ( .A(n5415), .B(n5414), .S(P2_IR_REG_25__SCAN_IN), .Z(n5416)
         );
  INV_X1 U6970 ( .A(n5416), .ZN(n5417) );
  NAND2_X1 U6971 ( .A1(n5417), .A2(n5411), .ZN(n7400) );
  INV_X1 U6972 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U6973 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  NAND2_X1 U6974 ( .A1(n5420), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5431) );
  INV_X1 U6975 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6976 ( .A1(n5431), .A2(n5421), .ZN(n5422) );
  NAND2_X1 U6977 ( .A1(n5422), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5424) );
  INV_X1 U6978 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5423) );
  XNOR2_X1 U6979 ( .A(n5424), .B(n5423), .ZN(n7215) );
  XNOR2_X1 U6980 ( .A(n7215), .B(P2_B_REG_SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6981 ( .A1(n7400), .A2(n5425), .ZN(n5426) );
  NAND2_X1 U6982 ( .A1(n5427), .A2(n5426), .ZN(n9705) );
  AOI21_X1 U6983 ( .B1(n5429), .B2(n5428), .A(n9705), .ZN(n5462) );
  NAND2_X1 U6984 ( .A1(n5430), .A2(n8357), .ZN(n5606) );
  NAND2_X1 U6985 ( .A1(n5606), .A2(n6279), .ZN(n5613) );
  XNOR2_X1 U6986 ( .A(n5431), .B(P2_IR_REG_23__SCAN_IN), .ZN(n6242) );
  NOR3_X1 U6987 ( .A1(n7215), .A2(n7400), .A3(n7480), .ZN(n6169) );
  OR2_X1 U6988 ( .A1(n6242), .A2(n6169), .ZN(n6277) );
  NAND2_X1 U6989 ( .A1(n5613), .A2(n9706), .ZN(n5432) );
  OR2_X1 U6990 ( .A1(n9705), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U6991 ( .A1(n7215), .A2(n7480), .ZN(n9709) );
  OR2_X1 U6992 ( .A1(n9705), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6993 ( .A1(n7400), .A2(n7480), .ZN(n9713) );
  NAND2_X1 U6994 ( .A1(n5434), .A2(n9713), .ZN(n6695) );
  NAND3_X1 U6995 ( .A1(n6696), .A2(n5610), .A3(n6695), .ZN(n5435) );
  INV_X1 U6996 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6997 ( .A1(n8676), .A2(n9722), .ZN(n8667) );
  OAI21_X1 U6998 ( .B1(n5444), .B2(n9767), .A(n5438), .ZN(P2_U3549) );
  INV_X1 U6999 ( .A(n6696), .ZN(n5439) );
  NAND3_X1 U7000 ( .A1(n5439), .A2(n5610), .A3(n6695), .ZN(n5440) );
  INV_X2 U7001 ( .A(n9758), .ZN(n9759) );
  NAND2_X1 U7002 ( .A1(n7885), .A2(n8714), .ZN(n5443) );
  NAND2_X1 U7003 ( .A1(n9758), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5442) );
  OAI21_X1 U7004 ( .B1(n5444), .B2(n9758), .A(n4796), .ZN(P2_U3517) );
  XNOR2_X1 U7005 ( .A(n5445), .B(n8092), .ZN(n8379) );
  AOI211_X1 U7006 ( .C1(n8044), .C2(n8396), .A(n9752), .B(n4291), .ZN(n8384)
         );
  NAND3_X1 U7007 ( .A1(n8390), .A2(n8092), .A3(n8040), .ZN(n5446) );
  NAND2_X1 U7008 ( .A1(n5446), .A2(n8585), .ZN(n5449) );
  OR2_X1 U7009 ( .A1(n6771), .A2(n8242), .ZN(n5448) );
  NAND2_X1 U7010 ( .A1(n8293), .A2(n8228), .ZN(n5447) );
  AND2_X1 U7011 ( .A1(n5448), .A2(n5447), .ZN(n5605) );
  OAI21_X1 U7012 ( .B1(n5450), .B2(n5449), .A(n5605), .ZN(n8378) );
  MUX2_X1 U7013 ( .A(n9834), .B(n5454), .S(n9770), .Z(n5453) );
  NAND2_X1 U7014 ( .A1(n8044), .A2(n5451), .ZN(n5452) );
  NAND2_X1 U7015 ( .A1(n5453), .A2(n5452), .ZN(P2_U3548) );
  INV_X1 U7016 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5455) );
  MUX2_X1 U7017 ( .A(n5455), .B(n5454), .S(n9759), .Z(n5457) );
  NAND2_X1 U7018 ( .A1(n8044), .A2(n8714), .ZN(n5456) );
  NAND2_X1 U7019 ( .A1(n5457), .A2(n5456), .ZN(P2_U3516) );
  OR2_X1 U7020 ( .A1(n8149), .A2(n6567), .ZN(n5459) );
  NAND2_X4 U7021 ( .A1(n5458), .A2(n6699), .ZN(n5590) );
  XNOR2_X1 U7022 ( .A(n5459), .B(n5590), .ZN(n5595) );
  INV_X1 U7023 ( .A(n5595), .ZN(n5596) );
  INV_X1 U7024 ( .A(n6695), .ZN(n5460) );
  NAND2_X1 U7025 ( .A1(n5460), .A2(n6696), .ZN(n5461) );
  OR2_X1 U7026 ( .A1(n5462), .A2(n5461), .ZN(n5611) );
  NAND3_X1 U7027 ( .A1(n5463), .A2(n9716), .A3(n9706), .ZN(n5464) );
  NOR3_X1 U7028 ( .A1(n8382), .A2(n5596), .A3(n4262), .ZN(n5465) );
  AOI21_X1 U7029 ( .B1(n5596), .B2(n8382), .A(n5465), .ZN(n5604) );
  INV_X1 U7030 ( .A(n5469), .ZN(n5467) );
  XNOR2_X1 U7031 ( .A(n8590), .B(n5590), .ZN(n5468) );
  INV_X1 U7032 ( .A(n5468), .ZN(n5466) );
  NAND2_X1 U7033 ( .A1(n5467), .A2(n5466), .ZN(n5472) );
  NAND2_X1 U7034 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  NAND2_X1 U7035 ( .A1(n5369), .A2(n7909), .ZN(n5471) );
  INV_X1 U7036 ( .A(n9715), .ZN(n6569) );
  MUX2_X1 U7037 ( .A(n5471), .B(n5590), .S(n6569), .Z(n6429) );
  NAND2_X1 U7038 ( .A1(n6428), .A2(n5472), .ZN(n6441) );
  OR2_X1 U7039 ( .A1(n4994), .A2(n6567), .ZN(n5473) );
  XNOR2_X1 U7040 ( .A(n8575), .B(n5568), .ZN(n5474) );
  XNOR2_X1 U7041 ( .A(n5473), .B(n5474), .ZN(n6442) );
  NAND2_X1 U7042 ( .A1(n8314), .A2(n7909), .ZN(n5476) );
  XNOR2_X1 U7043 ( .A(n5475), .B(n5568), .ZN(n5477) );
  XNOR2_X1 U7044 ( .A(n5476), .B(n5477), .ZN(n6450) );
  INV_X1 U7045 ( .A(n5476), .ZN(n5478) );
  NAND2_X1 U7046 ( .A1(n5478), .A2(n5477), .ZN(n5479) );
  OR2_X1 U7047 ( .A1(n5023), .A2(n6567), .ZN(n5481) );
  XNOR2_X1 U7048 ( .A(n6644), .B(n5568), .ZN(n5480) );
  NAND2_X1 U7049 ( .A1(n5481), .A2(n5480), .ZN(n5483) );
  OAI21_X1 U7050 ( .B1(n5481), .B2(n5480), .A(n5483), .ZN(n6623) );
  NAND2_X1 U7051 ( .A1(n6621), .A2(n5483), .ZN(n6629) );
  OR2_X1 U7052 ( .A1(n6726), .A2(n6567), .ZN(n5484) );
  XNOR2_X1 U7053 ( .A(n6821), .B(n5568), .ZN(n5485) );
  XNOR2_X1 U7054 ( .A(n5484), .B(n5485), .ZN(n6628) );
  INV_X1 U7055 ( .A(n6628), .ZN(n5488) );
  INV_X1 U7056 ( .A(n5484), .ZN(n5487) );
  INV_X1 U7057 ( .A(n5485), .ZN(n5486) );
  AND2_X1 U7058 ( .A1(n8311), .A2(n7909), .ZN(n5489) );
  XNOR2_X1 U7059 ( .A(n6888), .B(n5590), .ZN(n5490) );
  NAND2_X1 U7060 ( .A1(n5489), .A2(n5490), .ZN(n5493) );
  INV_X1 U7061 ( .A(n5489), .ZN(n5492) );
  INV_X1 U7062 ( .A(n5490), .ZN(n5491) );
  NAND2_X1 U7063 ( .A1(n5492), .A2(n5491), .ZN(n5494) );
  AND2_X1 U7064 ( .A1(n5493), .A2(n5494), .ZN(n6725) );
  OR2_X1 U7065 ( .A1(n6851), .A2(n6567), .ZN(n5495) );
  XNOR2_X1 U7066 ( .A(n6743), .B(n5568), .ZN(n5496) );
  XNOR2_X1 U7067 ( .A(n5495), .B(n5496), .ZN(n6757) );
  OAI22_X2 U7068 ( .A1(n6758), .A2(n6757), .B1(n5496), .B2(n5495), .ZN(n6850)
         );
  XNOR2_X1 U7069 ( .A(n6935), .B(n5590), .ZN(n5499) );
  NAND2_X1 U7070 ( .A1(n8309), .A2(n7909), .ZN(n5497) );
  XNOR2_X1 U7071 ( .A(n5499), .B(n5497), .ZN(n6849) );
  INV_X1 U7072 ( .A(n5497), .ZN(n5498) );
  NAND2_X1 U7073 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  XNOR2_X1 U7074 ( .A(n7360), .B(n5568), .ZN(n5501) );
  OR2_X1 U7075 ( .A1(n7015), .A2(n6567), .ZN(n5502) );
  NAND2_X1 U7076 ( .A1(n5501), .A2(n5502), .ZN(n7011) );
  INV_X1 U7077 ( .A(n5501), .ZN(n5504) );
  INV_X1 U7078 ( .A(n5502), .ZN(n5503) );
  NAND2_X1 U7079 ( .A1(n5504), .A2(n5503), .ZN(n5505) );
  NAND2_X1 U7080 ( .A1(n7011), .A2(n5505), .ZN(n7022) );
  INV_X1 U7081 ( .A(n7022), .ZN(n5506) );
  XNOR2_X1 U7082 ( .A(n7103), .B(n5590), .ZN(n5510) );
  NOR2_X1 U7083 ( .A1(n7033), .A2(n6567), .ZN(n5509) );
  XNOR2_X1 U7084 ( .A(n5510), .B(n5509), .ZN(n7012) );
  INV_X1 U7085 ( .A(n7012), .ZN(n5507) );
  AND2_X1 U7086 ( .A1(n5507), .A2(n7011), .ZN(n5508) );
  NAND2_X1 U7087 ( .A1(n7010), .A2(n5508), .ZN(n5512) );
  NAND2_X1 U7088 ( .A1(n5510), .A2(n5509), .ZN(n5511) );
  NAND2_X1 U7089 ( .A1(n5512), .A2(n5511), .ZN(n7031) );
  XNOR2_X1 U7090 ( .A(n8669), .B(n5568), .ZN(n5513) );
  NOR2_X1 U7091 ( .A1(n7075), .A2(n6567), .ZN(n5514) );
  XNOR2_X1 U7092 ( .A(n5513), .B(n5514), .ZN(n7032) );
  NAND2_X1 U7093 ( .A1(n7031), .A2(n7032), .ZN(n5517) );
  INV_X1 U7094 ( .A(n5513), .ZN(n5515) );
  NAND2_X1 U7095 ( .A1(n5515), .A2(n5514), .ZN(n5516) );
  NAND2_X1 U7096 ( .A1(n5517), .A2(n5516), .ZN(n7201) );
  INV_X1 U7097 ( .A(n7201), .ZN(n5524) );
  XNOR2_X1 U7098 ( .A(n7210), .B(n5568), .ZN(n5518) );
  OR2_X1 U7099 ( .A1(n7218), .A2(n6567), .ZN(n5519) );
  NAND2_X1 U7100 ( .A1(n5518), .A2(n5519), .ZN(n5525) );
  INV_X1 U7101 ( .A(n5518), .ZN(n5521) );
  INV_X1 U7102 ( .A(n5519), .ZN(n5520) );
  NAND2_X1 U7103 ( .A1(n5521), .A2(n5520), .ZN(n5522) );
  NAND2_X1 U7104 ( .A1(n5525), .A2(n5522), .ZN(n7204) );
  NAND2_X1 U7105 ( .A1(n5524), .A2(n5523), .ZN(n7202) );
  XNOR2_X1 U7106 ( .A(n7250), .B(n5590), .ZN(n5526) );
  NOR2_X1 U7107 ( .A1(n7277), .A2(n6567), .ZN(n5527) );
  XNOR2_X1 U7108 ( .A(n5526), .B(n5527), .ZN(n7216) );
  INV_X1 U7109 ( .A(n5526), .ZN(n5529) );
  INV_X1 U7110 ( .A(n5527), .ZN(n5528) );
  XNOR2_X1 U7111 ( .A(n7421), .B(n5568), .ZN(n5530) );
  OR2_X1 U7112 ( .A1(n7388), .A2(n6567), .ZN(n5531) );
  NAND2_X1 U7113 ( .A1(n5530), .A2(n5531), .ZN(n5535) );
  INV_X1 U7114 ( .A(n5530), .ZN(n5533) );
  INV_X1 U7115 ( .A(n5531), .ZN(n5532) );
  NAND2_X1 U7116 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  NAND2_X1 U7117 ( .A1(n5535), .A2(n5534), .ZN(n7414) );
  XNOR2_X1 U7118 ( .A(n8287), .B(n5568), .ZN(n8191) );
  OR2_X1 U7119 ( .A1(n7466), .A2(n6567), .ZN(n5537) );
  NAND2_X1 U7120 ( .A1(n8191), .A2(n5537), .ZN(n5536) );
  NAND2_X1 U7121 ( .A1(n8190), .A2(n5536), .ZN(n5541) );
  XNOR2_X1 U7122 ( .A(n8715), .B(n5568), .ZN(n5544) );
  NOR2_X1 U7123 ( .A1(n8206), .A2(n6567), .ZN(n5542) );
  XNOR2_X1 U7124 ( .A(n5544), .B(n5542), .ZN(n8193) );
  INV_X1 U7125 ( .A(n8191), .ZN(n5538) );
  INV_X1 U7126 ( .A(n5537), .ZN(n8278) );
  NAND2_X1 U7127 ( .A1(n5538), .A2(n8278), .ZN(n5539) );
  AND2_X1 U7128 ( .A1(n8193), .A2(n5539), .ZN(n5540) );
  INV_X1 U7129 ( .A(n5542), .ZN(n5543) );
  NAND2_X1 U7130 ( .A1(n5544), .A2(n5543), .ZN(n5545) );
  XNOR2_X1 U7131 ( .A(n8552), .B(n5590), .ZN(n5547) );
  NOR2_X1 U7132 ( .A1(n8253), .A2(n6567), .ZN(n5546) );
  XNOR2_X1 U7133 ( .A(n5547), .B(n5546), .ZN(n8204) );
  NAND2_X1 U7134 ( .A1(n5547), .A2(n5546), .ZN(n5548) );
  XNOR2_X1 U7135 ( .A(n8535), .B(n5590), .ZN(n5552) );
  NAND2_X1 U7136 ( .A1(n8300), .A2(n7909), .ZN(n5550) );
  XNOR2_X1 U7137 ( .A(n5552), .B(n5550), .ZN(n8251) );
  INV_X1 U7138 ( .A(n5550), .ZN(n5551) );
  XNOR2_X1 U7139 ( .A(n8517), .B(n5568), .ZN(n5553) );
  NAND2_X1 U7140 ( .A1(n8299), .A2(n7909), .ZN(n5554) );
  NAND2_X1 U7141 ( .A1(n5553), .A2(n5554), .ZN(n5558) );
  INV_X1 U7142 ( .A(n5553), .ZN(n5556) );
  INV_X1 U7143 ( .A(n5554), .ZN(n5555) );
  NAND2_X1 U7144 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  AND2_X1 U7145 ( .A1(n5558), .A2(n5557), .ZN(n8164) );
  XNOR2_X1 U7146 ( .A(n8503), .B(n5568), .ZN(n5559) );
  NAND2_X1 U7147 ( .A1(n8298), .A2(n7909), .ZN(n5560) );
  XNOR2_X1 U7148 ( .A(n5559), .B(n5560), .ZN(n8226) );
  INV_X1 U7149 ( .A(n5559), .ZN(n5562) );
  INV_X1 U7150 ( .A(n5560), .ZN(n5561) );
  XNOR2_X1 U7151 ( .A(n8696), .B(n5590), .ZN(n5563) );
  NOR2_X1 U7152 ( .A1(n8244), .A2(n6567), .ZN(n5564) );
  XNOR2_X1 U7153 ( .A(n5563), .B(n5564), .ZN(n8171) );
  NAND2_X1 U7154 ( .A1(n8172), .A2(n8171), .ZN(n5567) );
  INV_X1 U7155 ( .A(n5563), .ZN(n5565) );
  NAND2_X1 U7156 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  XNOR2_X1 U7157 ( .A(n8471), .B(n5568), .ZN(n5569) );
  INV_X1 U7158 ( .A(n8156), .ZN(n8296) );
  NAND2_X1 U7159 ( .A1(n8296), .A2(n7909), .ZN(n8237) );
  INV_X1 U7160 ( .A(n5569), .ZN(n5570) );
  XNOR2_X1 U7161 ( .A(n8626), .B(n5590), .ZN(n5575) );
  XNOR2_X1 U7162 ( .A(n5577), .B(n5575), .ZN(n8155) );
  INV_X1 U7163 ( .A(n8157), .ZN(n8295) );
  NAND2_X1 U7164 ( .A1(n8155), .A2(n5574), .ZN(n5580) );
  NOR2_X1 U7165 ( .A1(n8157), .A2(n6567), .ZN(n8215) );
  INV_X1 U7166 ( .A(n5575), .ZN(n5576) );
  OAI21_X1 U7167 ( .B1(n8215), .B2(n8216), .A(n8214), .ZN(n5579) );
  XOR2_X1 U7168 ( .A(n5590), .B(n8616), .Z(n5583) );
  INV_X1 U7169 ( .A(n5583), .ZN(n5581) );
  NAND2_X1 U7170 ( .A1(n8181), .A2(n5581), .ZN(n5582) );
  NAND2_X1 U7171 ( .A1(n8294), .A2(n7909), .ZN(n8179) );
  NAND2_X1 U7172 ( .A1(n5582), .A2(n8179), .ZN(n5586) );
  NAND2_X1 U7173 ( .A1(n5584), .A2(n5583), .ZN(n5585) );
  XNOR2_X1 U7174 ( .A(n8611), .B(n5590), .ZN(n5588) );
  NOR2_X1 U7175 ( .A1(n8182), .A2(n6567), .ZN(n5587) );
  NAND2_X1 U7176 ( .A1(n5588), .A2(n5587), .ZN(n5589) );
  OAI21_X1 U7177 ( .B1(n5588), .B2(n5587), .A(n5589), .ZN(n8262) );
  XNOR2_X1 U7178 ( .A(n8606), .B(n5590), .ZN(n5592) );
  AND2_X1 U7179 ( .A1(n8293), .A2(n7909), .ZN(n5591) );
  NAND2_X1 U7180 ( .A1(n5592), .A2(n5591), .ZN(n5593) );
  OAI21_X1 U7181 ( .B1(n5592), .B2(n5591), .A(n5593), .ZN(n8145) );
  INV_X1 U7182 ( .A(n5593), .ZN(n5594) );
  NOR3_X1 U7183 ( .A1(n8382), .A2(n4262), .A3(n5595), .ZN(n5598) );
  NOR2_X1 U7184 ( .A1(n8044), .A2(n5596), .ZN(n5597) );
  NAND2_X1 U7185 ( .A1(n5603), .A2(n5599), .ZN(n5602) );
  INV_X1 U7186 ( .A(n4262), .ZN(n8274) );
  NOR2_X1 U7187 ( .A1(n5611), .A2(n6280), .ZN(n5607) );
  NOR2_X1 U7188 ( .A1(n9722), .A2(n6279), .ZN(n5600) );
  NAND2_X1 U7189 ( .A1(n5607), .A2(n5600), .ZN(n8289) );
  OAI21_X1 U7190 ( .B1(n8382), .B2(n8274), .A(n8289), .ZN(n5601) );
  OAI211_X1 U7191 ( .C1(n5604), .C2(n5603), .A(n5602), .B(n5601), .ZN(n5620)
         );
  INV_X1 U7192 ( .A(n5605), .ZN(n5608) );
  INV_X1 U7193 ( .A(n5606), .ZN(n8107) );
  AOI22_X1 U7194 ( .A1(n5608), .A2(n8281), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5609) );
  INV_X1 U7195 ( .A(n5609), .ZN(n5618) );
  INV_X1 U7196 ( .A(n8380), .ZN(n5616) );
  NAND2_X1 U7197 ( .A1(n5611), .A2(n5610), .ZN(n5615) );
  INV_X1 U7198 ( .A(n6277), .ZN(n5612) );
  AND2_X1 U7199 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  NAND2_X1 U7200 ( .A1(n5615), .A2(n5614), .ZN(n6431) );
  NAND2_X1 U7201 ( .A1(n6431), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8285) );
  NOR2_X1 U7202 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  NAND2_X1 U7203 ( .A1(n5620), .A2(n5619), .ZN(P2_U3222) );
  NAND2_X1 U7204 ( .A1(n5732), .A2(n5623), .ZN(n5757) );
  NOR2_X1 U7205 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n6123) );
  NAND3_X1 U7206 ( .A1(n6123), .A2(n5887), .A3(n5947), .ZN(n5629) );
  NOR2_X1 U7207 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5627) );
  NOR2_X1 U7208 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5626) );
  NOR2_X1 U7209 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5625) );
  NAND4_X1 U7210 ( .A1(n5627), .A2(n5626), .A3(n5625), .A4(n5643), .ZN(n5628)
         );
  INV_X1 U7211 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5632) );
  INV_X1 U7212 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5663) );
  INV_X1 U7213 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U7214 ( .A1(n5634), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5635) );
  MUX2_X1 U7215 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5635), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5637) );
  INV_X1 U7216 ( .A(n5636), .ZN(n9345) );
  AND2_X4 U7217 ( .A1(n8115), .A2(n9351), .ZN(n5840) );
  NAND2_X1 U7218 ( .A1(n5840), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5641) );
  INV_X1 U7219 ( .A(n9351), .ZN(n5638) );
  NAND2_X1 U7220 ( .A1(n5724), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U7221 ( .A1(n5709), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5639) );
  AND2_X2 U7222 ( .A1(n5642), .A2(n5643), .ZN(n5886) );
  NOR2_X1 U7223 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5644) );
  NOR2_X1 U7224 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5645) );
  INV_X1 U7225 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5646) );
  INV_X1 U7226 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5648) );
  AND2_X2 U7227 ( .A1(n5650), .A2(n5677), .ZN(n6099) );
  NAND2_X1 U7228 ( .A1(n5652), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5655) );
  INV_X1 U7229 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7230 ( .A1(n5655), .A2(n5653), .ZN(n5657) );
  INV_X1 U7231 ( .A(n5655), .ZN(n5656) );
  NAND2_X1 U7232 ( .A1(n5656), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U7233 ( .A1(n5658), .A2(n5657), .ZN(n7402) );
  NAND2_X1 U7234 ( .A1(n5659), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5661) );
  XNOR2_X1 U7235 ( .A(n5661), .B(n5660), .ZN(n7200) );
  NOR2_X1 U7236 ( .A1(n7402), .A2(n7200), .ZN(n5662) );
  INV_X1 U7237 ( .A(n5667), .ZN(n5668) );
  INV_X1 U7238 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7239 ( .A1(n5672), .A2(n5671), .ZN(n5714) );
  OAI21_X1 U7240 ( .B1(n5672), .B2(n5671), .A(n5714), .ZN(n6228) );
  OR2_X1 U7241 ( .A1(n5771), .A2(n6231), .ZN(n5673) );
  AND2_X2 U7242 ( .A1(n5675), .A2(n6170), .ZN(n5897) );
  INV_X2 U7243 ( .A(n5897), .ZN(n6094) );
  OAI22_X1 U7244 ( .A1(n6775), .A2(n5703), .B1(n9639), .B2(n6094), .ZN(n5681)
         );
  INV_X1 U7245 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6121) );
  XNOR2_X2 U7246 ( .A(n5678), .B(n6121), .ZN(n7815) );
  NAND2_X1 U7247 ( .A1(n5679), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5680) );
  XNOR2_X2 U7248 ( .A(n5680), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U7249 ( .A1(n7768), .A2(n4434), .ZN(n6583) );
  XNOR2_X1 U7250 ( .A(n5681), .B(n5865), .ZN(n5704) );
  INV_X1 U7251 ( .A(n5704), .ZN(n5707) );
  NAND2_X4 U7252 ( .A1(n5682), .A2(n5897), .ZN(n8128) );
  OAI22_X1 U7253 ( .A1(n6775), .A2(n8128), .B1(n9639), .B2(n5703), .ZN(n5705)
         );
  INV_X1 U7254 ( .A(n5705), .ZN(n5706) );
  NAND2_X1 U7255 ( .A1(n4271), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7256 ( .A1(n5840), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7257 ( .A1(n5709), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7258 ( .A1(n5724), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7259 ( .A1(n7538), .A2(SI_0_), .ZN(n5688) );
  INV_X1 U7260 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U7261 ( .A1(n5688), .A2(n5687), .ZN(n5690) );
  AND2_X1 U7262 ( .A1(n5690), .A2(n5689), .ZN(n9353) );
  MUX2_X1 U7263 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9353), .S(n6173), .Z(n6715) );
  AOI222_X1 U7264 ( .A1(n6579), .A2(n8126), .B1(n6715), .B2(n5897), .C1(n6168), 
        .C2(P1_REG1_REG_0__SCAN_IN), .ZN(n5692) );
  INV_X1 U7265 ( .A(n6579), .ZN(n6615) );
  NAND2_X1 U7266 ( .A1(n5840), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U7267 ( .A1(n5709), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7268 ( .A1(n5724), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5693) );
  INV_X1 U7269 ( .A(n8885), .ZN(n7526) );
  INV_X1 U7270 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7271 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5698) );
  NAND2_X1 U7272 ( .A1(n5772), .A2(n6480), .ZN(n5699) );
  OAI22_X1 U7273 ( .A1(n7526), .A2(n7868), .B1(n7773), .B2(n6094), .ZN(n5700)
         );
  XNOR2_X1 U7274 ( .A(n5700), .B(n5865), .ZN(n5702) );
  OAI22_X1 U7275 ( .A1(n7526), .A2(n8128), .B1(n7773), .B2(n8122), .ZN(n6614)
         );
  INV_X1 U7276 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U7277 ( .A1(n4272), .A2(n6779), .ZN(n5713) );
  NAND2_X1 U7278 ( .A1(n5840), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7279 ( .A1(n5709), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U7280 ( .A1(n5724), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5710) );
  INV_X1 U7281 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5715) );
  OR2_X1 U7282 ( .A1(n7562), .A2(n6222), .ZN(n5718) );
  OR2_X1 U7283 ( .A1(n5771), .A2(n6221), .ZN(n5717) );
  OAI211_X1 U7284 ( .C1(n6173), .C2(n6416), .A(n5718), .B(n5717), .ZN(n6780)
         );
  OAI22_X1 U7285 ( .A1(n6777), .A2(n7868), .B1(n9644), .B2(n6094), .ZN(n5720)
         );
  XNOR2_X1 U7286 ( .A(n5720), .B(n4268), .ZN(n5722) );
  OAI22_X1 U7287 ( .A1(n6777), .A2(n8128), .B1(n9644), .B2(n8122), .ZN(n5721)
         );
  OR2_X1 U7288 ( .A1(n5722), .A2(n5721), .ZN(n6746) );
  AND2_X1 U7289 ( .A1(n5722), .A2(n5721), .ZN(n6747) );
  NAND2_X1 U7290 ( .A1(n5840), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7291 ( .A1(n4273), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5727) );
  INV_X1 U7292 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5723) );
  XNOR2_X1 U7293 ( .A(n5723), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6940) );
  NAND2_X1 U7294 ( .A1(n4271), .A2(n6940), .ZN(n5726) );
  NAND2_X1 U7295 ( .A1(n4266), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5725) );
  INV_X1 U7296 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5801) );
  NOR2_X1 U7297 ( .A1(n5729), .A2(n5801), .ZN(n5730) );
  MUX2_X1 U7298 ( .A(n5801), .B(n5730), .S(P1_IR_REG_4__SCAN_IN), .Z(n5731) );
  INV_X1 U7299 ( .A(n5731), .ZN(n5734) );
  INV_X1 U7300 ( .A(n5732), .ZN(n5733) );
  NAND2_X1 U7301 ( .A1(n5734), .A2(n5733), .ZN(n9522) );
  OR2_X1 U7302 ( .A1(n7562), .A2(n6220), .ZN(n5736) );
  OR2_X1 U7303 ( .A1(n5771), .A2(n6219), .ZN(n5735) );
  OAI211_X1 U7304 ( .C1(n6173), .C2(n9522), .A(n5736), .B(n5735), .ZN(n6867)
         );
  INV_X1 U7305 ( .A(n6867), .ZN(n6957) );
  OAI22_X1 U7306 ( .A1(n7839), .A2(n8128), .B1(n6957), .B2(n8122), .ZN(n5739)
         );
  OAI22_X1 U7307 ( .A1(n7839), .A2(n7868), .B1(n6957), .B2(n6094), .ZN(n5737)
         );
  XNOR2_X1 U7308 ( .A(n5737), .B(n5865), .ZN(n5738) );
  XOR2_X1 U7309 ( .A(n5739), .B(n5738), .Z(n6832) );
  NAND2_X1 U7310 ( .A1(n5840), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U7311 ( .A1(n4266), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5744) );
  AOI21_X1 U7312 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5741) );
  NOR2_X1 U7313 ( .A1(n5741), .A2(n5752), .ZN(n7846) );
  NAND2_X1 U7314 ( .A1(n4270), .A2(n7846), .ZN(n5743) );
  NAND2_X1 U7315 ( .A1(n4273), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5742) );
  OR2_X1 U7316 ( .A1(n5732), .A2(n5801), .ZN(n5746) );
  XNOR2_X1 U7317 ( .A(n5746), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6384) );
  INV_X1 U7318 ( .A(n6384), .ZN(n6225) );
  OR2_X1 U7319 ( .A1(n5771), .A2(n6226), .ZN(n5748) );
  OR2_X1 U7320 ( .A1(n7562), .A2(n6227), .ZN(n5747) );
  INV_X1 U7321 ( .A(n7852), .ZN(n9653) );
  OAI22_X1 U7322 ( .A1(n6950), .A2(n7868), .B1(n9653), .B2(n6094), .ZN(n5749)
         );
  XNOR2_X1 U7323 ( .A(n5749), .B(n5865), .ZN(n6909) );
  OR2_X1 U7324 ( .A1(n8128), .A2(n6950), .ZN(n5751) );
  OR2_X1 U7325 ( .A1(n9653), .A2(n8122), .ZN(n5750) );
  NAND2_X1 U7326 ( .A1(n5751), .A2(n5750), .ZN(n6908) );
  NAND2_X1 U7327 ( .A1(n5840), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U7328 ( .A1(n4273), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U7329 ( .A1(n5752), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5765) );
  OAI21_X1 U7330 ( .B1(n5752), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5765), .ZN(
        n7826) );
  INV_X1 U7331 ( .A(n7826), .ZN(n7066) );
  NAND2_X1 U7332 ( .A1(n4272), .A2(n7066), .ZN(n5754) );
  NAND2_X1 U7333 ( .A1(n4266), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U7334 ( .A1(n5758), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5760) );
  XNOR2_X1 U7335 ( .A(n5760), .B(n5759), .ZN(n6517) );
  OR2_X1 U7336 ( .A1(n6224), .A2(n5771), .ZN(n5762) );
  OR2_X1 U7337 ( .A1(n7562), .A2(n9837), .ZN(n5761) );
  OAI211_X1 U7338 ( .C1(n6173), .C2(n6517), .A(n5762), .B(n5761), .ZN(n7824)
         );
  INV_X1 U7339 ( .A(n7824), .ZN(n7825) );
  OAI22_X1 U7340 ( .A1(n7840), .A2(n8128), .B1(n7825), .B2(n8122), .ZN(n7060)
         );
  OAI22_X1 U7341 ( .A1(n7840), .A2(n7868), .B1(n7825), .B2(n6094), .ZN(n5763)
         );
  XNOR2_X1 U7342 ( .A(n5763), .B(n4268), .ZN(n7061) );
  NAND2_X1 U7343 ( .A1(n4266), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U7344 ( .A1(n5840), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5769) );
  AND2_X1 U7345 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  NOR2_X1 U7346 ( .A1(n5794), .A2(n5766), .ZN(n7228) );
  NAND2_X1 U7347 ( .A1(n4272), .A2(n7228), .ZN(n5768) );
  NAND2_X1 U7348 ( .A1(n4273), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5767) );
  INV_X2 U7349 ( .A(n5771), .ZN(n5779) );
  NAND2_X1 U7350 ( .A1(n6233), .A2(n5779), .ZN(n5775) );
  OR2_X1 U7351 ( .A1(n5758), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7352 ( .A1(n5780), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5773) );
  XNOR2_X1 U7353 ( .A(n5773), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6234) );
  AOI22_X1 U7354 ( .A1(n5968), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5967), .B2(
        n6234), .ZN(n5774) );
  NAND2_X1 U7355 ( .A1(n5775), .A2(n5774), .ZN(n7226) );
  OAI22_X1 U7356 ( .A1(n7132), .A2(n7868), .B1(n7114), .B2(n6094), .ZN(n5776)
         );
  XNOR2_X1 U7357 ( .A(n5776), .B(n4268), .ZN(n5778) );
  OAI22_X1 U7358 ( .A1(n7132), .A2(n8128), .B1(n7114), .B2(n8122), .ZN(n5777)
         );
  OR2_X1 U7359 ( .A1(n5778), .A2(n5777), .ZN(n7234) );
  NAND2_X1 U7360 ( .A1(n7233), .A2(n7234), .ZN(n7232) );
  NAND2_X1 U7361 ( .A1(n5778), .A2(n5777), .ZN(n7236) );
  NAND2_X1 U7362 ( .A1(n6246), .A2(n5779), .ZN(n5784) );
  NOR2_X1 U7363 ( .A1(n5780), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5802) );
  INV_X1 U7364 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U7365 ( .A1(n5802), .A2(n5781), .ZN(n5818) );
  NAND2_X1 U7366 ( .A1(n5818), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5782) );
  XNOR2_X1 U7367 ( .A(n5782), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6394) );
  AOI22_X1 U7368 ( .A1(n5968), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5967), .B2(
        n6394), .ZN(n5783) );
  NAND2_X1 U7369 ( .A1(n4266), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7370 ( .A1(n5840), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7371 ( .A1(n5794), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5796) );
  INV_X1 U7372 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7373 ( .A1(n5796), .A2(n5785), .ZN(n5786) );
  AND2_X1 U7374 ( .A1(n5822), .A2(n5786), .ZN(n7354) );
  NAND2_X1 U7375 ( .A1(n4271), .A2(n7354), .ZN(n5788) );
  NAND2_X1 U7376 ( .A1(n4273), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5787) );
  NAND4_X1 U7377 ( .A1(n5790), .A2(n5789), .A3(n5788), .A4(n5787), .ZN(n8877)
         );
  AOI22_X1 U7378 ( .A1(n7344), .A2(n5986), .B1(n4274), .B2(n8877), .ZN(n5791)
         );
  XNOR2_X1 U7379 ( .A(n5791), .B(n4268), .ZN(n7349) );
  NAND2_X1 U7380 ( .A1(n7344), .A2(n4274), .ZN(n5793) );
  NAND2_X1 U7381 ( .A1(n6096), .A2(n8877), .ZN(n5792) );
  NAND2_X1 U7382 ( .A1(n5793), .A2(n5792), .ZN(n5813) );
  INV_X1 U7383 ( .A(n5813), .ZN(n7348) );
  NAND2_X1 U7384 ( .A1(n4266), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7385 ( .A1(n5840), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5799) );
  OR2_X1 U7386 ( .A1(n5794), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5795) );
  AND2_X1 U7387 ( .A1(n5796), .A2(n5795), .ZN(n7375) );
  NAND2_X1 U7388 ( .A1(n4271), .A2(n7375), .ZN(n5798) );
  NAND2_X1 U7389 ( .A1(n4273), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5797) );
  OR2_X1 U7390 ( .A1(n8128), .A2(n7231), .ZN(n5809) );
  NAND2_X1 U7391 ( .A1(n6237), .A2(n5779), .ZN(n5807) );
  NOR2_X1 U7392 ( .A1(n5802), .A2(n5801), .ZN(n5803) );
  MUX2_X1 U7393 ( .A(n5801), .B(n5803), .S(P1_IR_REG_8__SCAN_IN), .Z(n5805) );
  INV_X1 U7394 ( .A(n5818), .ZN(n5804) );
  INV_X1 U7395 ( .A(n6239), .ZN(n8889) );
  AOI22_X1 U7396 ( .A1(n5968), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5967), .B2(
        n8889), .ZN(n5806) );
  NAND2_X1 U7397 ( .A1(n7287), .A2(n4274), .ZN(n5808) );
  NAND2_X1 U7398 ( .A1(n5809), .A2(n5808), .ZN(n7345) );
  INV_X1 U7399 ( .A(n7345), .ZN(n5812) );
  NAND2_X1 U7400 ( .A1(n7287), .A2(n5986), .ZN(n5810) );
  OAI21_X1 U7401 ( .B1(n7231), .B2(n8122), .A(n5810), .ZN(n5811) );
  XNOR2_X1 U7402 ( .A(n5811), .B(n4268), .ZN(n7371) );
  INV_X1 U7403 ( .A(n7371), .ZN(n7347) );
  OAI22_X1 U7404 ( .A1(n7349), .A2(n7348), .B1(n5812), .B2(n7347), .ZN(n5817)
         );
  OAI21_X1 U7405 ( .B1(n7371), .B2(n7345), .A(n5813), .ZN(n5815) );
  NOR3_X1 U7406 ( .A1(n7371), .A2(n7345), .A3(n5813), .ZN(n5814) );
  AOI21_X1 U7407 ( .B1(n7349), .B2(n5815), .A(n5814), .ZN(n5816) );
  NAND2_X1 U7408 ( .A1(n6251), .A2(n5779), .ZN(n5821) );
  NAND2_X1 U7409 ( .A1(n5836), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5819) );
  XNOR2_X1 U7410 ( .A(n5819), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6504) );
  AOI22_X1 U7411 ( .A1(n5968), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5967), .B2(
        n6504), .ZN(n5820) );
  NAND2_X1 U7412 ( .A1(n5821), .A2(n5820), .ZN(n7322) );
  NAND2_X1 U7413 ( .A1(n7322), .A2(n5986), .ZN(n5829) );
  INV_X1 U7414 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U7415 ( .A1(n5822), .A2(n6407), .ZN(n5823) );
  AND2_X1 U7416 ( .A1(n5842), .A2(n5823), .ZN(n7301) );
  NAND2_X1 U7417 ( .A1(n4270), .A2(n7301), .ZN(n5827) );
  NAND2_X1 U7418 ( .A1(n5840), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U7419 ( .A1(n4273), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U7420 ( .A1(n4266), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5824) );
  OR2_X1 U7421 ( .A1(n9434), .A2(n8122), .ZN(n5828) );
  NAND2_X1 U7422 ( .A1(n5829), .A2(n5828), .ZN(n5830) );
  XNOR2_X1 U7423 ( .A(n5830), .B(n4268), .ZN(n7297) );
  NAND2_X1 U7424 ( .A1(n7322), .A2(n4274), .ZN(n5832) );
  INV_X1 U7425 ( .A(n9434), .ZN(n8876) );
  NAND2_X1 U7426 ( .A1(n8876), .A2(n6096), .ZN(n5831) );
  NAND2_X1 U7427 ( .A1(n5832), .A2(n5831), .ZN(n5833) );
  NOR2_X1 U7428 ( .A1(n7297), .A2(n5833), .ZN(n5835) );
  INV_X1 U7429 ( .A(n7297), .ZN(n5834) );
  INV_X1 U7430 ( .A(n5833), .ZN(n7296) );
  NAND2_X1 U7431 ( .A1(n6255), .A2(n5779), .ZN(n5839) );
  OAI21_X1 U7432 ( .B1(n5836), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5837) );
  XNOR2_X1 U7433 ( .A(n5837), .B(P1_IR_REG_11__SCAN_IN), .ZN(n8908) );
  AOI22_X1 U7434 ( .A1(n5968), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5967), .B2(
        n8908), .ZN(n5838) );
  NAND2_X1 U7435 ( .A1(n5840), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U7436 ( .A1(n4273), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5846) );
  INV_X1 U7437 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5841) );
  AND2_X1 U7438 ( .A1(n5842), .A2(n5841), .ZN(n5843) );
  NOR2_X1 U7439 ( .A1(n5857), .A2(n5843), .ZN(n9440) );
  NAND2_X1 U7440 ( .A1(n4272), .A2(n9440), .ZN(n5845) );
  NAND2_X1 U7441 ( .A1(n4266), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5844) );
  NAND4_X1 U7442 ( .A1(n5847), .A2(n5846), .A3(n5845), .A4(n5844), .ZN(n8875)
         );
  INV_X1 U7443 ( .A(n8875), .ZN(n7320) );
  OAI22_X1 U7444 ( .A1(n9469), .A2(n6094), .B1(n7320), .B2(n8122), .ZN(n5848)
         );
  XNOR2_X1 U7445 ( .A(n5848), .B(n4268), .ZN(n5850) );
  AND2_X1 U7446 ( .A1(n6096), .A2(n8875), .ZN(n5849) );
  AOI21_X1 U7447 ( .B1(n9442), .B2(n4274), .A(n5849), .ZN(n5851) );
  XNOR2_X1 U7448 ( .A(n5850), .B(n5851), .ZN(n8838) );
  NAND2_X1 U7449 ( .A1(n6267), .A2(n5779), .ZN(n5856) );
  NAND2_X1 U7450 ( .A1(n5853), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5854) );
  XNOR2_X1 U7451 ( .A(n5854), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9545) );
  AOI22_X1 U7452 ( .A1(n5968), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5967), .B2(
        n9545), .ZN(n5855) );
  NAND2_X1 U7453 ( .A1(n8771), .A2(n5986), .ZN(n5864) );
  NAND2_X1 U7454 ( .A1(n5840), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7455 ( .A1(n4273), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5861) );
  NOR2_X1 U7456 ( .A1(n5857), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5858) );
  OR2_X1 U7457 ( .A1(n5876), .A2(n5858), .ZN(n7337) );
  INV_X1 U7458 ( .A(n7337), .ZN(n8766) );
  NAND2_X1 U7459 ( .A1(n4270), .A2(n8766), .ZN(n5860) );
  NAND2_X1 U7460 ( .A1(n4266), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5859) );
  OR2_X1 U7461 ( .A1(n9436), .A2(n8122), .ZN(n5863) );
  NAND2_X1 U7462 ( .A1(n5864), .A2(n5863), .ZN(n5866) );
  XNOR2_X1 U7463 ( .A(n5866), .B(n5719), .ZN(n5868) );
  NOR2_X1 U7464 ( .A1(n9436), .A2(n8128), .ZN(n5867) );
  AOI21_X1 U7465 ( .B1(n8771), .B2(n4274), .A(n5867), .ZN(n5869) );
  NAND2_X1 U7466 ( .A1(n5868), .A2(n5869), .ZN(n8761) );
  INV_X1 U7467 ( .A(n5868), .ZN(n5871) );
  INV_X1 U7468 ( .A(n5869), .ZN(n5870) );
  NAND2_X1 U7469 ( .A1(n5871), .A2(n5870), .ZN(n8762) );
  NAND2_X1 U7470 ( .A1(n6377), .A2(n5779), .ZN(n5875) );
  OR2_X1 U7471 ( .A1(n5642), .A2(n5801), .ZN(n5873) );
  XNOR2_X1 U7472 ( .A(n5873), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9557) );
  AOI22_X1 U7473 ( .A1(n5968), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5967), .B2(
        n9557), .ZN(n5874) );
  NAND2_X1 U7474 ( .A1(n5840), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7475 ( .A1(n4266), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5880) );
  NOR2_X1 U7476 ( .A1(n5876), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5877) );
  OR2_X1 U7477 ( .A1(n5891), .A2(n5877), .ZN(n9420) );
  INV_X1 U7478 ( .A(n9420), .ZN(n8818) );
  NAND2_X1 U7479 ( .A1(n4270), .A2(n8818), .ZN(n5879) );
  NAND2_X1 U7480 ( .A1(n4273), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5878) );
  NAND4_X1 U7481 ( .A1(n5881), .A2(n5880), .A3(n5879), .A4(n5878), .ZN(n8873)
         );
  AOI22_X1 U7482 ( .A1(n8822), .A2(n5986), .B1(n4274), .B2(n8873), .ZN(n5882)
         );
  XOR2_X1 U7483 ( .A(n4268), .B(n5882), .Z(n5883) );
  INV_X1 U7484 ( .A(n5883), .ZN(n8815) );
  INV_X1 U7485 ( .A(n8822), .ZN(n9457) );
  INV_X1 U7486 ( .A(n8873), .ZN(n8769) );
  OAI22_X1 U7487 ( .A1(n9457), .A2(n7868), .B1(n8769), .B2(n8128), .ZN(n8814)
         );
  OAI21_X1 U7488 ( .B1(n8817), .B2(n5883), .A(n8814), .ZN(n5884) );
  NAND2_X1 U7489 ( .A1(n6414), .A2(n5779), .ZN(n5890) );
  OR2_X1 U7490 ( .A1(n5886), .A2(n5801), .ZN(n5888) );
  NAND2_X1 U7491 ( .A1(n5888), .A2(n5887), .ZN(n5900) );
  OAI21_X1 U7492 ( .B1(n5888), .B2(n5887), .A(n5900), .ZN(n8924) );
  INV_X1 U7493 ( .A(n8924), .ZN(n9570) );
  AOI22_X1 U7494 ( .A1(n5968), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5967), .B2(
        n9570), .ZN(n5889) );
  INV_X1 U7495 ( .A(n9322), .ZN(n7460) );
  NAND2_X1 U7496 ( .A1(n4266), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7497 ( .A1(n5840), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5895) );
  OR2_X1 U7498 ( .A1(n5891), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7499 ( .A1(n5891), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5905) );
  AND2_X1 U7500 ( .A1(n5892), .A2(n5905), .ZN(n8729) );
  NAND2_X1 U7501 ( .A1(n4271), .A2(n8729), .ZN(n5894) );
  NAND2_X1 U7502 ( .A1(n4273), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5893) );
  NAND4_X1 U7503 ( .A1(n5896), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n8872)
         );
  OAI22_X1 U7504 ( .A1(n7460), .A2(n8122), .B1(n9412), .B2(n8128), .ZN(n5899)
         );
  INV_X1 U7505 ( .A(n5899), .ZN(n8724) );
  AOI22_X1 U7506 ( .A1(n9322), .A2(n5986), .B1(n4274), .B2(n8872), .ZN(n5898)
         );
  XOR2_X1 U7507 ( .A(n4268), .B(n5898), .Z(n8725) );
  NAND2_X1 U7508 ( .A1(n6574), .A2(n5779), .ZN(n5903) );
  NAND2_X1 U7509 ( .A1(n5900), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5901) );
  XNOR2_X1 U7510 ( .A(n5901), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9582) );
  AOI22_X1 U7511 ( .A1(n5968), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5967), .B2(
        n9582), .ZN(n5902) );
  NAND2_X1 U7512 ( .A1(n9315), .A2(n5986), .ZN(n5912) );
  NAND2_X1 U7513 ( .A1(n4266), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7514 ( .A1(n5840), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5909) );
  INV_X1 U7515 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7516 ( .A1(n5905), .A2(n5904), .ZN(n5906) );
  AND2_X1 U7517 ( .A1(n5920), .A2(n5906), .ZN(n9230) );
  NAND2_X1 U7518 ( .A1(n4272), .A2(n9230), .ZN(n5908) );
  NAND2_X1 U7519 ( .A1(n4273), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5907) );
  NAND4_X1 U7520 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(n8871)
         );
  NAND2_X1 U7521 ( .A1(n8871), .A2(n4274), .ZN(n5911) );
  NAND2_X1 U7522 ( .A1(n5912), .A2(n5911), .ZN(n5913) );
  XNOR2_X1 U7523 ( .A(n5913), .B(n5719), .ZN(n8856) );
  AND2_X1 U7524 ( .A1(n6096), .A2(n8871), .ZN(n5914) );
  AOI21_X1 U7525 ( .B1(n9315), .B2(n4274), .A(n5914), .ZN(n8857) );
  NAND2_X1 U7526 ( .A1(n8856), .A2(n8857), .ZN(n5915) );
  NAND2_X1 U7527 ( .A1(n6562), .A2(n5779), .ZN(n5919) );
  NAND2_X1 U7528 ( .A1(n5916), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5917) );
  XNOR2_X1 U7529 ( .A(n5917), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9593) );
  AOI22_X1 U7530 ( .A1(n5968), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5967), .B2(
        n9593), .ZN(n5918) );
  NAND2_X1 U7531 ( .A1(n5840), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7532 ( .A1(n4266), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5923) );
  INV_X1 U7533 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8778) );
  AOI21_X1 U7534 ( .B1(n5920), .B2(n8778), .A(n5935), .ZN(n8782) );
  NAND2_X1 U7535 ( .A1(n4272), .A2(n8782), .ZN(n5922) );
  NAND2_X1 U7536 ( .A1(n4273), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5921) );
  NOR2_X1 U7537 ( .A1(n9220), .A2(n8122), .ZN(n5925) );
  AOI21_X1 U7538 ( .B1(n9312), .B2(n5986), .A(n5925), .ZN(n5926) );
  XNOR2_X1 U7539 ( .A(n5926), .B(n4268), .ZN(n5929) );
  NOR2_X1 U7540 ( .A1(n9220), .A2(n8128), .ZN(n5927) );
  AOI21_X1 U7541 ( .B1(n9312), .B2(n4274), .A(n5927), .ZN(n5928) );
  NAND2_X1 U7542 ( .A1(n5929), .A2(n5928), .ZN(n5931) );
  OAI21_X1 U7543 ( .B1(n5929), .B2(n5928), .A(n5931), .ZN(n5930) );
  INV_X1 U7544 ( .A(n5930), .ZN(n8775) );
  NAND2_X1 U7545 ( .A1(n8774), .A2(n5931), .ZN(n8786) );
  NAND2_X1 U7546 ( .A1(n5933), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5948) );
  XNOR2_X1 U7547 ( .A(n5948), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9605) );
  AOI22_X1 U7548 ( .A1(n5968), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5967), .B2(
        n9605), .ZN(n5934) );
  NAND2_X1 U7549 ( .A1(n4266), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7550 ( .A1(n5840), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7551 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(n5935), .ZN(n5955) );
  OAI21_X1 U7552 ( .B1(P1_REG3_REG_17__SCAN_IN), .B2(n5935), .A(n5955), .ZN(
        n5936) );
  INV_X1 U7553 ( .A(n5936), .ZN(n9211) );
  NAND2_X1 U7554 ( .A1(n4270), .A2(n9211), .ZN(n5938) );
  NAND2_X1 U7555 ( .A1(n4273), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5937) );
  OAI22_X1 U7556 ( .A1(n9214), .A2(n7868), .B1(n9190), .B2(n8128), .ZN(n5943)
         );
  OAI22_X1 U7557 ( .A1(n9214), .A2(n6094), .B1(n9190), .B2(n8122), .ZN(n5941)
         );
  XNOR2_X1 U7558 ( .A(n5941), .B(n4268), .ZN(n5942) );
  XOR2_X1 U7559 ( .A(n5943), .B(n5942), .Z(n8788) );
  NAND2_X1 U7560 ( .A1(n8786), .A2(n8788), .ZN(n8787) );
  INV_X1 U7561 ( .A(n5942), .ZN(n5945) );
  INV_X1 U7562 ( .A(n5943), .ZN(n5944) );
  NAND2_X1 U7563 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  NAND2_X1 U7564 ( .A1(n6766), .A2(n5779), .ZN(n5952) );
  NAND2_X1 U7565 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  NAND2_X1 U7566 ( .A1(n5949), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U7567 ( .A(n5950), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9620) );
  AOI22_X1 U7568 ( .A1(n5968), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5967), .B2(
        n9620), .ZN(n5951) );
  NAND2_X1 U7569 ( .A1(n4266), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7570 ( .A1(n5840), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5959) );
  INV_X1 U7571 ( .A(n5955), .ZN(n5953) );
  INV_X1 U7572 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7573 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  AND2_X1 U7574 ( .A1(n5990), .A2(n5956), .ZN(n9196) );
  NAND2_X1 U7575 ( .A1(n4271), .A2(n9196), .ZN(n5958) );
  NAND2_X1 U7576 ( .A1(n4273), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5957) );
  OAI22_X1 U7577 ( .A1(n9193), .A2(n6094), .B1(n9208), .B2(n8122), .ZN(n5961)
         );
  XOR2_X1 U7578 ( .A(n4268), .B(n5961), .Z(n5963) );
  NAND2_X1 U7579 ( .A1(n5962), .A2(n5963), .ZN(n8844) );
  OAI22_X1 U7580 ( .A1(n9193), .A2(n7868), .B1(n9208), .B2(n8128), .ZN(n8847)
         );
  NAND2_X1 U7581 ( .A1(n8844), .A2(n8847), .ZN(n5966) );
  INV_X1 U7582 ( .A(n5962), .ZN(n5965) );
  INV_X1 U7583 ( .A(n5963), .ZN(n5964) );
  NAND2_X1 U7584 ( .A1(n5965), .A2(n5964), .ZN(n8845) );
  NAND2_X1 U7585 ( .A1(n5966), .A2(n8845), .ZN(n8744) );
  INV_X1 U7586 ( .A(n8744), .ZN(n5982) );
  NAND2_X1 U7587 ( .A1(n6808), .A2(n5779), .ZN(n5970) );
  AOI22_X1 U7588 ( .A1(n5968), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9157), .B2(
        n5967), .ZN(n5969) );
  NAND2_X1 U7589 ( .A1(n9295), .A2(n5986), .ZN(n5976) );
  NAND2_X1 U7590 ( .A1(n5840), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7591 ( .A1(n4273), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5973) );
  XNOR2_X1 U7592 ( .A(n5990), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n9170) );
  NAND2_X1 U7593 ( .A1(n4270), .A2(n9170), .ZN(n5972) );
  NAND2_X1 U7594 ( .A1(n4266), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5971) );
  NAND4_X1 U7595 ( .A1(n5974), .A2(n5973), .A3(n5972), .A4(n5971), .ZN(n9187)
         );
  NAND2_X1 U7596 ( .A1(n9187), .A2(n4274), .ZN(n5975) );
  NAND2_X1 U7597 ( .A1(n5976), .A2(n5975), .ZN(n5977) );
  XNOR2_X1 U7598 ( .A(n5977), .B(n5719), .ZN(n5980) );
  AND2_X1 U7599 ( .A1(n6096), .A2(n9187), .ZN(n5978) );
  AOI21_X1 U7600 ( .B1(n9295), .B2(n4274), .A(n5978), .ZN(n5979) );
  NAND2_X1 U7601 ( .A1(n5980), .A2(n5979), .ZN(n5983) );
  OAI21_X1 U7602 ( .B1(n5980), .B2(n5979), .A(n5983), .ZN(n8747) );
  NAND2_X1 U7603 ( .A1(n5982), .A2(n5981), .ZN(n8745) );
  NAND2_X1 U7604 ( .A1(n6972), .A2(n5779), .ZN(n5985) );
  OR2_X1 U7605 ( .A1(n7562), .A2(n6973), .ZN(n5984) );
  NAND2_X1 U7606 ( .A1(n9290), .A2(n5986), .ZN(n5997) );
  NAND2_X1 U7607 ( .A1(n5840), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7608 ( .A1(n4266), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5994) );
  INV_X1 U7609 ( .A(n5990), .ZN(n5988) );
  AND2_X1 U7610 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5987) );
  NAND2_X1 U7611 ( .A1(n5988), .A2(n5987), .ZN(n6009) );
  INV_X1 U7612 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8748) );
  INV_X1 U7613 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5989) );
  OAI21_X1 U7614 ( .B1(n5990), .B2(n8748), .A(n5989), .ZN(n5991) );
  AND2_X1 U7615 ( .A1(n6009), .A2(n5991), .ZN(n9155) );
  NAND2_X1 U7616 ( .A1(n4271), .A2(n9155), .ZN(n5993) );
  NAND2_X1 U7617 ( .A1(n4273), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5992) );
  NAND4_X1 U7618 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .ZN(n9137)
         );
  NAND2_X1 U7619 ( .A1(n9137), .A2(n4274), .ZN(n5996) );
  NAND2_X1 U7620 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  XNOR2_X1 U7621 ( .A(n5998), .B(n4268), .ZN(n6001) );
  NAND2_X1 U7622 ( .A1(n9290), .A2(n4274), .ZN(n6000) );
  NAND2_X1 U7623 ( .A1(n6096), .A2(n9137), .ZN(n5999) );
  NAND2_X1 U7624 ( .A1(n6000), .A2(n5999), .ZN(n6002) );
  NAND2_X1 U7625 ( .A1(n6001), .A2(n6002), .ZN(n8805) );
  INV_X1 U7626 ( .A(n6001), .ZN(n6004) );
  INV_X1 U7627 ( .A(n6002), .ZN(n6003) );
  NAND2_X1 U7628 ( .A1(n6004), .A2(n6003), .ZN(n8804) );
  NAND2_X1 U7629 ( .A1(n7005), .A2(n5779), .ZN(n6006) );
  OR2_X1 U7630 ( .A1(n7562), .A2(n7006), .ZN(n6005) );
  NAND2_X1 U7631 ( .A1(n9140), .A2(n5986), .ZN(n6016) );
  NAND2_X1 U7632 ( .A1(n4266), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7633 ( .A1(n5840), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6013) );
  INV_X1 U7634 ( .A(n6009), .ZN(n6007) );
  NAND2_X1 U7635 ( .A1(n6007), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6025) );
  INV_X1 U7636 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7637 ( .A1(n6009), .A2(n6008), .ZN(n6010) );
  AND2_X1 U7638 ( .A1(n6025), .A2(n6010), .ZN(n9142) );
  NAND2_X1 U7639 ( .A1(n4272), .A2(n9142), .ZN(n6012) );
  NAND2_X1 U7640 ( .A1(n4273), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6011) );
  OR2_X1 U7641 ( .A1(n9154), .A2(n8122), .ZN(n6015) );
  NAND2_X1 U7642 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  XNOR2_X1 U7643 ( .A(n6017), .B(n4268), .ZN(n6018) );
  INV_X1 U7644 ( .A(n9154), .ZN(n9124) );
  AOI22_X1 U7645 ( .A1(n9140), .A2(n4274), .B1(n6096), .B2(n9124), .ZN(n6019)
         );
  XNOR2_X1 U7646 ( .A(n6018), .B(n6019), .ZN(n8755) );
  INV_X1 U7647 ( .A(n6018), .ZN(n6020) );
  NAND2_X1 U7648 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  NAND2_X1 U7649 ( .A1(n7055), .A2(n5779), .ZN(n6023) );
  OR2_X1 U7650 ( .A1(n7562), .A2(n9862), .ZN(n6022) );
  NAND2_X1 U7651 ( .A1(n4266), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7652 ( .A1(n5840), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6029) );
  INV_X1 U7653 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7654 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  AND2_X1 U7655 ( .A1(n6035), .A2(n6026), .ZN(n9118) );
  NAND2_X1 U7656 ( .A1(n4270), .A2(n9118), .ZN(n6028) );
  NAND2_X1 U7657 ( .A1(n4273), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6027) );
  INV_X1 U7658 ( .A(n9108), .ZN(n9138) );
  AOI22_X1 U7659 ( .A1(n9278), .A2(n4274), .B1(n6096), .B2(n9138), .ZN(n6043)
         );
  NAND2_X1 U7660 ( .A1(n6044), .A2(n6043), .ZN(n8825) );
  NAND2_X1 U7661 ( .A1(n7146), .A2(n5779), .ZN(n6033) );
  OR2_X1 U7662 ( .A1(n7562), .A2(n6031), .ZN(n6032) );
  NAND2_X1 U7663 ( .A1(n5840), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7664 ( .A1(n4273), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6039) );
  INV_X1 U7665 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7666 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  AND2_X1 U7667 ( .A1(n6052), .A2(n6036), .ZN(n9101) );
  NAND2_X1 U7668 ( .A1(n4272), .A2(n9101), .ZN(n6038) );
  NAND2_X1 U7669 ( .A1(n4266), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6037) );
  OAI22_X1 U7670 ( .A1(n9103), .A2(n6094), .B1(n9089), .B2(n8122), .ZN(n6041)
         );
  XOR2_X1 U7671 ( .A(n6041), .B(n4268), .Z(n6048) );
  INV_X1 U7672 ( .A(n6048), .ZN(n6042) );
  OR2_X2 U7673 ( .A1(n6044), .A2(n6043), .ZN(n8826) );
  OAI22_X1 U7674 ( .A1(n9120), .A2(n6094), .B1(n9108), .B2(n8122), .ZN(n6045)
         );
  XOR2_X1 U7675 ( .A(n4268), .B(n6045), .Z(n8827) );
  AOI22_X1 U7676 ( .A1(n9273), .A2(n4274), .B1(n6096), .B2(n9123), .ZN(n8737)
         );
  NAND2_X1 U7677 ( .A1(n8736), .A2(n8737), .ZN(n7860) );
  NAND2_X1 U7678 ( .A1(n6047), .A2(n8825), .ZN(n6049) );
  NAND2_X1 U7679 ( .A1(n7198), .A2(n5779), .ZN(n6051) );
  OR2_X1 U7680 ( .A1(n7562), .A2(n7199), .ZN(n6050) );
  NAND2_X1 U7681 ( .A1(n4266), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7682 ( .A1(n5840), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6056) );
  INV_X1 U7683 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U7684 ( .A1(n6052), .A2(n8797), .ZN(n6053) );
  AND2_X1 U7685 ( .A1(n6063), .A2(n6053), .ZN(n9092) );
  NAND2_X1 U7686 ( .A1(n4270), .A2(n9092), .ZN(n6055) );
  NAND2_X1 U7687 ( .A1(n4273), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6054) );
  OAI22_X1 U7688 ( .A1(n8966), .A2(n7868), .B1(n9109), .B2(n8128), .ZN(n6079)
         );
  OAI22_X1 U7689 ( .A1(n8966), .A2(n6094), .B1(n9109), .B2(n8122), .ZN(n6058)
         );
  XNOR2_X1 U7690 ( .A(n6058), .B(n4268), .ZN(n6078) );
  XOR2_X1 U7691 ( .A(n6079), .B(n6078), .Z(n8794) );
  NAND2_X1 U7692 ( .A1(n7399), .A2(n5779), .ZN(n6060) );
  OR2_X1 U7693 ( .A1(n7562), .A2(n7404), .ZN(n6059) );
  NAND2_X1 U7694 ( .A1(n9069), .A2(n5986), .ZN(n6070) );
  NAND2_X1 U7695 ( .A1(n5840), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7696 ( .A1(n4273), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6067) );
  INV_X1 U7697 ( .A(n6063), .ZN(n6061) );
  NAND2_X1 U7698 ( .A1(n6061), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6088) );
  INV_X1 U7699 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7700 ( .A1(n6063), .A2(n6062), .ZN(n6064) );
  AND2_X1 U7701 ( .A1(n6088), .A2(n6064), .ZN(n9076) );
  NAND2_X1 U7702 ( .A1(n4271), .A2(n9076), .ZN(n6066) );
  NAND2_X1 U7703 ( .A1(n4266), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6065) );
  OR2_X1 U7704 ( .A1(n9088), .A2(n8122), .ZN(n6069) );
  NAND2_X1 U7705 ( .A1(n6070), .A2(n6069), .ZN(n6071) );
  XNOR2_X1 U7706 ( .A(n6071), .B(n4268), .ZN(n6074) );
  INV_X1 U7707 ( .A(n6074), .ZN(n6073) );
  INV_X1 U7708 ( .A(n9069), .ZN(n8972) );
  OAI22_X1 U7709 ( .A1(n8972), .A2(n7868), .B1(n9088), .B2(n8128), .ZN(n6075)
         );
  INV_X1 U7710 ( .A(n6075), .ZN(n6072) );
  NAND2_X1 U7711 ( .A1(n6073), .A2(n6072), .ZN(n6082) );
  INV_X1 U7712 ( .A(n6082), .ZN(n6076) );
  XOR2_X1 U7713 ( .A(n6075), .B(n6074), .Z(n6161) );
  INV_X1 U7714 ( .A(n6077), .ZN(n6084) );
  INV_X1 U7715 ( .A(n6078), .ZN(n6081) );
  INV_X1 U7716 ( .A(n6079), .ZN(n6080) );
  NAND2_X1 U7717 ( .A1(n6081), .A2(n6080), .ZN(n6160) );
  AND2_X1 U7718 ( .A1(n6160), .A2(n6082), .ZN(n6083) );
  NAND2_X1 U7719 ( .A1(n6131), .A2(n6129), .ZN(n6127) );
  NAND2_X1 U7720 ( .A1(n7479), .A2(n5779), .ZN(n6086) );
  OR2_X1 U7721 ( .A1(n7562), .A2(n7483), .ZN(n6085) );
  NAND2_X1 U7722 ( .A1(n4266), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7723 ( .A1(n5840), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6092) );
  INV_X1 U7724 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7725 ( .A1(n6088), .A2(n6087), .ZN(n6089) );
  NAND2_X1 U7726 ( .A1(n4271), .A2(n9053), .ZN(n6091) );
  NAND2_X1 U7727 ( .A1(n4273), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6090) );
  OAI22_X1 U7728 ( .A1(n9055), .A2(n6094), .B1(n9073), .B2(n8122), .ZN(n6095)
         );
  XNOR2_X1 U7729 ( .A(n6095), .B(n4268), .ZN(n7857) );
  OR2_X1 U7730 ( .A1(n9055), .A2(n8122), .ZN(n6098) );
  NAND2_X1 U7731 ( .A1(n8973), .A2(n6096), .ZN(n6097) );
  NAND2_X1 U7732 ( .A1(n6098), .A2(n6097), .ZN(n7856) );
  XNOR2_X1 U7733 ( .A(n7857), .B(n7856), .ZN(n6128) );
  INV_X1 U7734 ( .A(n6099), .ZN(n7647) );
  NAND2_X1 U7735 ( .A1(n7815), .A2(n7647), .ZN(n6713) );
  INV_X1 U7736 ( .A(n6713), .ZN(n6100) );
  INV_X1 U7737 ( .A(n7809), .ZN(n6712) );
  AND2_X2 U7738 ( .A1(n6100), .A2(n6712), .ZN(n9455) );
  NAND2_X1 U7739 ( .A1(n7768), .A2(n6099), .ZN(n7765) );
  INV_X1 U7740 ( .A(n7765), .ZN(n6530) );
  INV_X1 U7741 ( .A(n6138), .ZN(n6126) );
  NAND2_X1 U7742 ( .A1(n7402), .A2(P1_B_REG_SCAN_IN), .ZN(n6102) );
  INV_X1 U7743 ( .A(n7200), .ZN(n6101) );
  MUX2_X1 U7744 ( .A(n6102), .B(P1_B_REG_SCAN_IN), .S(n6101), .Z(n6103) );
  NAND2_X1 U7745 ( .A1(n6103), .A2(n6118), .ZN(n6113) );
  INV_X1 U7746 ( .A(n7402), .ZN(n6104) );
  OAI22_X1 U7747 ( .A1(n6113), .A2(P1_D_REG_1__SCAN_IN), .B1(n6118), .B2(n6104), .ZN(n6526) );
  INV_X1 U7748 ( .A(n6526), .ZN(n6116) );
  NOR4_X1 U7749 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6108) );
  NOR4_X1 U7750 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6107) );
  NOR4_X1 U7751 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6106) );
  NOR4_X1 U7752 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6105) );
  NAND4_X1 U7753 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n6115)
         );
  NOR2_X1 U7754 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .ZN(
        n6112) );
  NOR4_X1 U7755 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6111) );
  NOR4_X1 U7756 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6110) );
  NOR4_X1 U7757 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6109) );
  NAND4_X1 U7758 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n6114)
         );
  OAI21_X1 U7759 ( .B1(n6115), .B2(n6114), .A(n9630), .ZN(n6527) );
  NAND2_X1 U7760 ( .A1(n6116), .A2(n6527), .ZN(n6681) );
  INV_X1 U7761 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7762 ( .A1(n9630), .A2(n6117), .ZN(n6120) );
  INV_X1 U7763 ( .A(n6118), .ZN(n7481) );
  NAND2_X1 U7764 ( .A1(n7481), .A2(n7200), .ZN(n6119) );
  NAND2_X1 U7765 ( .A1(n6120), .A2(n6119), .ZN(n6679) );
  OR2_X1 U7766 ( .A1(n6681), .A2(n6679), .ZN(n6136) );
  INV_X1 U7767 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6122) );
  NAND3_X1 U7768 ( .A1(n6123), .A2(n6122), .A3(n6121), .ZN(n6124) );
  OAI21_X1 U7769 ( .B1(n5679), .B2(n6124), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6125) );
  XNOR2_X1 U7770 ( .A(n6125), .B(P1_IR_REG_23__SCAN_IN), .ZN(n7100) );
  NOR2_X1 U7771 ( .A1(n6136), .A2(n9635), .ZN(n6143) );
  INV_X1 U7772 ( .A(n6128), .ZN(n6130) );
  NAND2_X1 U7773 ( .A1(n6131), .A2(n7858), .ZN(n6132) );
  AND2_X1 U7774 ( .A1(n6136), .A2(n7812), .ZN(n6134) );
  OR2_X1 U7775 ( .A1(n5675), .A2(n6583), .ZN(n7818) );
  OR2_X1 U7776 ( .A1(n6713), .A2(n7771), .ZN(n6690) );
  NAND2_X1 U7777 ( .A1(n7818), .A2(n6690), .ZN(n6133) );
  NAND2_X1 U7778 ( .A1(n6134), .A2(n6133), .ZN(n6140) );
  AND2_X1 U7779 ( .A1(n6683), .A2(n7812), .ZN(n6135) );
  AND2_X1 U7780 ( .A1(n6140), .A2(n6135), .ZN(n7240) );
  NAND2_X1 U7781 ( .A1(n7240), .A2(n9455), .ZN(n8813) );
  INV_X1 U7782 ( .A(n6136), .ZN(n6540) );
  NOR2_X1 U7783 ( .A1(n7100), .A2(n6168), .ZN(n6137) );
  OAI211_X1 U7784 ( .C1(n6138), .C2(n6540), .A(n6137), .B(n6683), .ZN(n6139)
         );
  NAND2_X1 U7785 ( .A1(n6139), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6141) );
  NAND2_X2 U7786 ( .A1(n6141), .A2(n6140), .ZN(n8861) );
  INV_X1 U7787 ( .A(n7818), .ZN(n6142) );
  AND2_X1 U7788 ( .A1(n6143), .A2(n6142), .ZN(n6145) );
  INV_X1 U7789 ( .A(n4269), .ZN(n9490) );
  NAND2_X1 U7790 ( .A1(n6145), .A2(n4269), .ZN(n8850) );
  NAND2_X1 U7791 ( .A1(n5840), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7792 ( .A1(n4266), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6152) );
  INV_X1 U7793 ( .A(n6148), .ZN(n6146) );
  NAND2_X1 U7794 ( .A1(n6146), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6670) );
  INV_X1 U7795 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7796 ( .A1(n6148), .A2(n6147), .ZN(n6149) );
  NAND2_X1 U7797 ( .A1(n4272), .A2(n9038), .ZN(n6151) );
  NAND2_X1 U7798 ( .A1(n4273), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6150) );
  INV_X1 U7799 ( .A(n9058), .ZN(n8975) );
  AOI22_X1 U7800 ( .A1(n8860), .A2(n8975), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n6154) );
  OAI21_X1 U7801 ( .B1(n9088), .B2(n8864), .A(n6154), .ZN(n6155) );
  AOI21_X1 U7802 ( .B1(n9053), .B2(n8861), .A(n6155), .ZN(n6156) );
  NAND2_X1 U7803 ( .A1(n6159), .A2(n6158), .ZN(P1_U3238) );
  INV_X1 U7804 ( .A(n6161), .ZN(n6162) );
  AOI22_X1 U7805 ( .A1(n8860), .A2(n8973), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n6163) );
  OAI21_X1 U7806 ( .B1(n9109), .B2(n8864), .A(n6163), .ZN(n6165) );
  NAND2_X1 U7807 ( .A1(n9069), .A2(n9455), .ZN(n9262) );
  INV_X1 U7808 ( .A(n7240), .ZN(n8851) );
  NOR2_X1 U7809 ( .A1(n9262), .A2(n8851), .ZN(n6164) );
  AOI211_X1 U7810 ( .C1(n9076), .C2(n8861), .A(n6165), .B(n6164), .ZN(n6166)
         );
  OAI21_X1 U7811 ( .B1(n6167), .B2(n8868), .A(n6166), .ZN(P1_U3223) );
  INV_X1 U7812 ( .A(n7100), .ZN(n6171) );
  AND2_X1 U7813 ( .A1(n6171), .A2(n6168), .ZN(n9504) );
  AND2_X2 U7814 ( .A1(n9504), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NOR2_X1 U7815 ( .A1(n6242), .A2(P2_U3152), .ZN(n9708) );
  AND2_X1 U7816 ( .A1(n6169), .A2(n9708), .ZN(P2_U3966) );
  NAND2_X1 U7817 ( .A1(n7765), .A2(n6170), .ZN(n6172) );
  NAND2_X1 U7818 ( .A1(n6172), .A2(n6171), .ZN(n6191) );
  NAND2_X1 U7819 ( .A1(n6191), .A2(n6173), .ZN(n9486) );
  NAND2_X1 U7820 ( .A1(n9486), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U7821 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7353) );
  OR2_X1 U7822 ( .A1(n6394), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7823 ( .A1(n6394), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6401) );
  AND2_X1 U7824 ( .A1(n6174), .A2(n6401), .ZN(n6188) );
  INV_X1 U7825 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6187) );
  INV_X1 U7826 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6175) );
  OR2_X1 U7827 ( .A1(n6234), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6186) );
  MUX2_X1 U7828 ( .A(n6175), .B(P1_REG2_REG_7__SCAN_IN), .S(n6234), .Z(n6488)
         );
  INV_X1 U7829 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6184) );
  NOR2_X1 U7830 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6384), .ZN(n6183) );
  INV_X1 U7831 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6176) );
  MUX2_X1 U7832 ( .A(n6176), .B(P1_REG2_REG_3__SCAN_IN), .S(n6416), .Z(n6424)
         );
  XNOR2_X1 U7833 ( .A(n6228), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9499) );
  AND2_X1 U7834 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6177) );
  NAND2_X1 U7835 ( .A1(n6480), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6178) );
  OAI211_X1 U7836 ( .C1(n6480), .C2(P1_REG2_REG_1__SCAN_IN), .A(n6177), .B(
        n6178), .ZN(n6482) );
  NAND2_X1 U7837 ( .A1(n6482), .A2(n6178), .ZN(n9498) );
  NAND2_X1 U7838 ( .A1(n9499), .A2(n9498), .ZN(n6180) );
  INV_X1 U7839 ( .A(n6228), .ZN(n9511) );
  NAND2_X1 U7840 ( .A1(n9511), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7841 ( .A1(n6180), .A2(n6179), .ZN(n6423) );
  NAND2_X1 U7842 ( .A1(n6424), .A2(n6423), .ZN(n6422) );
  OR2_X1 U7843 ( .A1(n6416), .A2(n6176), .ZN(n6181) );
  AND2_X1 U7844 ( .A1(n6422), .A2(n6181), .ZN(n9516) );
  INV_X1 U7845 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6182) );
  MUX2_X1 U7846 ( .A(n6182), .B(P1_REG2_REG_4__SCAN_IN), .S(n9522), .Z(n9517)
         );
  NAND2_X1 U7847 ( .A1(n9522), .A2(n6182), .ZN(n6385) );
  INV_X1 U7848 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7848) );
  MUX2_X1 U7849 ( .A(n7848), .B(P1_REG2_REG_5__SCAN_IN), .S(n6384), .Z(n6386)
         );
  MUX2_X1 U7850 ( .A(n6184), .B(P1_REG2_REG_6__SCAN_IN), .S(n6517), .Z(n6521)
         );
  NAND2_X1 U7851 ( .A1(n6522), .A2(n6521), .ZN(n6520) );
  OAI21_X1 U7852 ( .B1(n6517), .B2(n6184), .A(n6520), .ZN(n6489) );
  INV_X1 U7853 ( .A(n6487), .ZN(n6185) );
  NAND2_X1 U7854 ( .A1(n6186), .A2(n6185), .ZN(n8892) );
  NAND2_X1 U7855 ( .A1(n6239), .A2(n6187), .ZN(n8896) );
  NOR2_X1 U7856 ( .A1(n9488), .A2(P1_U3084), .ZN(n7484) );
  NAND2_X1 U7857 ( .A1(n6191), .A2(n7484), .ZN(n8938) );
  OR2_X1 U7858 ( .A1(n8938), .A2(n4269), .ZN(n9613) );
  INV_X1 U7859 ( .A(n9613), .ZN(n8895) );
  NAND2_X1 U7860 ( .A1(n8893), .A2(n6188), .ZN(n6402) );
  OAI211_X1 U7861 ( .C1(n6188), .C2(n8893), .A(n8895), .B(n6402), .ZN(n6189)
         );
  INV_X1 U7862 ( .A(n6189), .ZN(n6213) );
  OR2_X1 U7863 ( .A1(n4269), .A2(P1_U3084), .ZN(n9484) );
  INV_X1 U7864 ( .A(n9488), .ZN(n9491) );
  NOR2_X1 U7865 ( .A1(n9484), .A2(n9491), .ZN(n6190) );
  NAND2_X1 U7866 ( .A1(n6191), .A2(n6190), .ZN(n9625) );
  XNOR2_X1 U7867 ( .A(n9522), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9526) );
  INV_X1 U7868 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6192) );
  OR2_X1 U7869 ( .A1(n6416), .A2(n6192), .ZN(n9524) );
  AND2_X1 U7870 ( .A1(n9526), .A2(n9524), .ZN(n6197) );
  MUX2_X1 U7871 ( .A(n6192), .B(P1_REG1_REG_3__SCAN_IN), .S(n6416), .Z(n6418)
         );
  XNOR2_X1 U7872 ( .A(n6228), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9508) );
  INV_X1 U7873 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6193) );
  XNOR2_X1 U7874 ( .A(n6480), .B(n6193), .ZN(n6472) );
  NAND2_X1 U7875 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6476) );
  INV_X1 U7876 ( .A(n6476), .ZN(n6194) );
  NAND2_X1 U7877 ( .A1(n6472), .A2(n6194), .ZN(n6473) );
  NAND2_X1 U7878 ( .A1(n6480), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7879 ( .A1(n6473), .A2(n6195), .ZN(n9507) );
  NAND2_X1 U7880 ( .A1(n9508), .A2(n9507), .ZN(n9506) );
  NAND2_X1 U7881 ( .A1(n9511), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7882 ( .A1(n9506), .A2(n6196), .ZN(n6417) );
  NAND2_X1 U7883 ( .A1(n6418), .A2(n6417), .ZN(n9525) );
  NAND2_X1 U7884 ( .A1(n6197), .A2(n9525), .ZN(n9529) );
  INV_X1 U7885 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7886 ( .A1(n9522), .A2(n6198), .ZN(n6199) );
  NAND2_X1 U7887 ( .A1(n9529), .A2(n6199), .ZN(n6382) );
  NAND2_X1 U7888 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6384), .ZN(n6200) );
  OAI21_X1 U7889 ( .B1(n6384), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6200), .ZN(
        n6381) );
  OR2_X1 U7890 ( .A1(n6382), .A2(n6381), .ZN(n6379) );
  AND2_X1 U7891 ( .A1(n6379), .A2(n6200), .ZN(n6514) );
  XNOR2_X1 U7892 ( .A(n6517), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n6515) );
  NAND2_X1 U7893 ( .A1(n6514), .A2(n6515), .ZN(n6513) );
  INV_X1 U7894 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7895 ( .A1(n6517), .A2(n6201), .ZN(n6202) );
  NAND2_X1 U7896 ( .A1(n6513), .A2(n6202), .ZN(n6491) );
  INV_X1 U7897 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6203) );
  MUX2_X1 U7898 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6203), .S(n6234), .Z(n6492)
         );
  NAND2_X1 U7899 ( .A1(n6491), .A2(n6492), .ZN(n6490) );
  OR2_X1 U7900 ( .A1(n6234), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6204) );
  INV_X1 U7901 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7902 ( .A1(n6239), .A2(n6205), .ZN(n8900) );
  NAND2_X1 U7903 ( .A1(n8901), .A2(n8900), .ZN(n6207) );
  NAND2_X1 U7904 ( .A1(n8889), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7905 ( .A1(n6207), .A2(n6206), .ZN(n8898) );
  INV_X1 U7906 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9694) );
  INV_X1 U7907 ( .A(n6394), .ZN(n6248) );
  AOI22_X1 U7908 ( .A1(n6394), .A2(n9694), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6248), .ZN(n6208) );
  NOR2_X1 U7909 ( .A1(n8898), .A2(n6208), .ZN(n6395) );
  AOI21_X1 U7910 ( .B1(n8898), .B2(n6208), .A(n6395), .ZN(n6209) );
  NOR2_X1 U7911 ( .A1(n9625), .A2(n6209), .ZN(n6212) );
  INV_X1 U7912 ( .A(n8938), .ZN(n6210) );
  AND2_X1 U7913 ( .A1(n6210), .A2(n4269), .ZN(n9619) );
  INV_X1 U7914 ( .A(n9619), .ZN(n8888) );
  INV_X1 U7915 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9982) );
  OAI22_X1 U7916 ( .A1(n8888), .A2(n6248), .B1(n9628), .B2(n9982), .ZN(n6211)
         );
  OR4_X1 U7917 ( .A1(n7353), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(P1_U3250)
         );
  AND2_X1 U7918 ( .A1(n7538), .A2(P2_U3152), .ZN(n6563) );
  NOR2_X1 U7919 ( .A1(n7538), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8721) );
  OAI222_X1 U7920 ( .A1(n4267), .A2(n9822), .B1(n7519), .B2(n6221), .C1(
        P2_U3152), .C2(n6347), .ZN(P2_U3355) );
  OAI222_X1 U7921 ( .A1(n4267), .A2(n6214), .B1(n7519), .B2(n6217), .C1(
        P2_U3152), .C2(n6295), .ZN(P2_U3357) );
  OAI222_X1 U7922 ( .A1(n4267), .A2(n6215), .B1(n7519), .B2(n6219), .C1(
        P2_U3152), .C2(n6360), .ZN(P2_U3354) );
  AND2_X1 U7923 ( .A1(n7538), .A2(P1_U3084), .ZN(n9344) );
  INV_X1 U7924 ( .A(n6480), .ZN(n6477) );
  OAI222_X1 U7925 ( .A1(n9349), .A2(n6218), .B1(n8117), .B2(n6217), .C1(
        P1_U3084), .C2(n6477), .ZN(P1_U3352) );
  OAI222_X1 U7926 ( .A1(n9349), .A2(n6220), .B1(n8117), .B2(n6219), .C1(
        P1_U3084), .C2(n9522), .ZN(P1_U3349) );
  OAI222_X1 U7927 ( .A1(n9349), .A2(n6222), .B1(n8117), .B2(n6221), .C1(
        P1_U3084), .C2(n6416), .ZN(P1_U3350) );
  OAI222_X1 U7928 ( .A1(n4267), .A2(n6223), .B1(n7519), .B2(n6226), .C1(
        P2_U3152), .C2(n6319), .ZN(P2_U3353) );
  OAI222_X1 U7929 ( .A1(n9349), .A2(n9837), .B1(n8117), .B2(n6224), .C1(
        P1_U3084), .C2(n6517), .ZN(P1_U3347) );
  OAI222_X1 U7930 ( .A1(n4267), .A2(n9820), .B1(n7519), .B2(n6224), .C1(
        P2_U3152), .C2(n6307), .ZN(P2_U3352) );
  OAI222_X1 U7931 ( .A1(n9349), .A2(n6227), .B1(n8117), .B2(n6226), .C1(
        P1_U3084), .C2(n6225), .ZN(P1_U3348) );
  OAI222_X1 U7932 ( .A1(n9349), .A2(n6229), .B1(n8117), .B2(n6231), .C1(
        P1_U3084), .C2(n6228), .ZN(P1_U3351) );
  OAI222_X1 U7933 ( .A1(n4267), .A2(n6232), .B1(n7519), .B2(n6231), .C1(
        P2_U3152), .C2(n6230), .ZN(P2_U3356) );
  INV_X1 U7934 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9821) );
  INV_X1 U7935 ( .A(n6233), .ZN(n6235) );
  INV_X1 U7936 ( .A(n6234), .ZN(n6493) );
  OAI222_X1 U7937 ( .A1(n9349), .A2(n9821), .B1(n8117), .B2(n6235), .C1(
        P1_U3084), .C2(n6493), .ZN(P1_U3346) );
  INV_X1 U7938 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6236) );
  INV_X1 U7939 ( .A(n6460), .ZN(n6334) );
  OAI222_X1 U7940 ( .A1(n4267), .A2(n6236), .B1(n7519), .B2(n6235), .C1(
        P2_U3152), .C2(n6334), .ZN(P2_U3351) );
  INV_X1 U7941 ( .A(n6237), .ZN(n6240) );
  INV_X1 U7942 ( .A(n6459), .ZN(n9963) );
  OAI222_X1 U7943 ( .A1(n4267), .A2(n6238), .B1(n7519), .B2(n6240), .C1(
        P2_U3152), .C2(n9963), .ZN(P2_U3350) );
  OAI222_X1 U7944 ( .A1(n9349), .A2(n6241), .B1(n8117), .B2(n6240), .C1(
        P1_U3084), .C2(n6239), .ZN(P1_U3345) );
  NAND2_X1 U7945 ( .A1(n6242), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8111) );
  OAI21_X1 U7946 ( .B1(n6283), .B2(n8111), .A(n6280), .ZN(n6245) );
  INV_X1 U7947 ( .A(n6279), .ZN(n6243) );
  NAND2_X1 U7948 ( .A1(n6283), .A2(n6243), .ZN(n6244) );
  NAND2_X1 U7949 ( .A1(n6245), .A2(n6244), .ZN(n8362) );
  NOR2_X1 U7950 ( .A1(P2_U3966), .A2(n9960), .ZN(P2_U3151) );
  INV_X1 U7951 ( .A(n6246), .ZN(n6249) );
  OAI222_X1 U7952 ( .A1(n8117), .A2(n6249), .B1(n6248), .B2(P1_U3084), .C1(
        n6247), .C2(n9349), .ZN(P1_U3344) );
  INV_X1 U7953 ( .A(n6606), .ZN(n6469) );
  OAI222_X1 U7954 ( .A1(n4267), .A2(n6250), .B1(n7519), .B2(n6249), .C1(n6469), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U7955 ( .A(n6251), .ZN(n6254) );
  INV_X1 U7956 ( .A(n9349), .ZN(n7485) );
  AOI22_X1 U7957 ( .A1(n6504), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7485), .ZN(n6252) );
  OAI21_X1 U7958 ( .B1(n6254), .B2(n8117), .A(n6252), .ZN(P1_U3343) );
  AOI22_X1 U7959 ( .A1(n6661), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n6563), .ZN(n6253) );
  OAI21_X1 U7960 ( .B1(n6254), .B2(n7519), .A(n6253), .ZN(P2_U3348) );
  INV_X1 U7961 ( .A(n6255), .ZN(n6259) );
  AOI22_X1 U7962 ( .A1(n6895), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n6563), .ZN(n6256) );
  OAI21_X1 U7963 ( .B1(n6259), .B2(n7519), .A(n6256), .ZN(P2_U3347) );
  INV_X2 U7964 ( .A(P2_U3966), .ZN(n8317) );
  NAND2_X1 U7965 ( .A1(n8317), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n6257) );
  OAI21_X1 U7966 ( .B1(n7466), .B2(n8317), .A(n6257), .ZN(P2_U3567) );
  INV_X1 U7967 ( .A(n8908), .ZN(n8920) );
  OAI222_X1 U7968 ( .A1(n8117), .A2(n6259), .B1(n8920), .B2(P1_U3084), .C1(
        n6258), .C2(n9349), .ZN(P1_U3342) );
  INV_X1 U7969 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7970 ( .A1(n6260), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6264) );
  NAND2_X1 U7971 ( .A1(n5354), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U7972 ( .A1(n6261), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6262) );
  AND3_X1 U7973 ( .A1(n6264), .A2(n6263), .A3(n6262), .ZN(n7905) );
  INV_X1 U7974 ( .A(n7905), .ZN(n8367) );
  NAND2_X1 U7975 ( .A1(n8367), .A2(P2_U3966), .ZN(n6265) );
  OAI21_X1 U7976 ( .B1(n6266), .B2(P2_U3966), .A(n6265), .ZN(P2_U3583) );
  INV_X1 U7977 ( .A(n6267), .ZN(n6270) );
  AOI22_X1 U7978 ( .A1(n6996), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n6563), .ZN(n6268) );
  OAI21_X1 U7979 ( .B1(n6270), .B2(n7519), .A(n6268), .ZN(P2_U3346) );
  AOI22_X1 U7980 ( .A1(n9545), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n7485), .ZN(n6269) );
  OAI21_X1 U7981 ( .B1(n6270), .B2(n8117), .A(n6269), .ZN(P1_U3341) );
  INV_X1 U7982 ( .A(n6347), .ZN(n6273) );
  INV_X1 U7983 ( .A(n6295), .ZN(n6375) );
  INV_X1 U7984 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6271) );
  INV_X1 U7985 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9878) );
  INV_X1 U7986 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9933) );
  AOI21_X1 U7987 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n6375), .A(n6370), .ZN(
        n9356) );
  XNOR2_X1 U7988 ( .A(n9358), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9355) );
  NOR2_X1 U7989 ( .A1(n9356), .A2(n9355), .ZN(n9354) );
  INV_X1 U7990 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6272) );
  MUX2_X1 U7991 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6272), .S(n6347), .Z(n6338)
         );
  NAND2_X1 U7992 ( .A1(n6292), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6274) );
  OAI21_X1 U7993 ( .B1(n6292), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6274), .ZN(
        n6351) );
  AOI21_X1 U7994 ( .B1(n6292), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6350), .ZN(
        n6312) );
  NAND2_X1 U7995 ( .A1(n6290), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6275) );
  OAI21_X1 U7996 ( .B1(n6290), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6275), .ZN(
        n6311) );
  NOR2_X1 U7997 ( .A1(n6312), .A2(n6311), .ZN(n6310) );
  AOI21_X1 U7998 ( .B1(n6290), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6310), .ZN(
        n6287) );
  NAND2_X1 U7999 ( .A1(n6326), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6276) );
  OAI21_X1 U8000 ( .B1(n6326), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6276), .ZN(
        n6286) );
  OR2_X1 U8001 ( .A1(n6288), .A2(P2_U3152), .ZN(n7497) );
  NAND2_X1 U8002 ( .A1(n7497), .A2(n8111), .ZN(n6278) );
  NAND2_X1 U8003 ( .A1(n6278), .A2(n6277), .ZN(n6282) );
  OR2_X1 U8004 ( .A1(n6280), .A2(n6279), .ZN(n6281) );
  NAND2_X1 U8005 ( .A1(n6282), .A2(n6281), .ZN(n6284) );
  NAND2_X1 U8006 ( .A1(n6284), .A2(n6283), .ZN(n6301) );
  NAND2_X1 U8007 ( .A1(n8317), .A2(n6301), .ZN(n6289) );
  NOR2_X1 U8008 ( .A1(n6288), .A2(n5394), .ZN(n6285) );
  AOI211_X1 U8009 ( .C1(n6287), .C2(n6286), .A(n6322), .B(n9951), .ZN(n6309)
         );
  NAND2_X1 U8010 ( .A1(n6289), .A2(n6288), .ZN(n9964) );
  NAND2_X1 U8011 ( .A1(n6290), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6299) );
  INV_X1 U8012 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6291) );
  MUX2_X1 U8013 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6291), .S(n6290), .Z(n6314)
         );
  NAND2_X1 U8014 ( .A1(n6292), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6298) );
  INV_X1 U8015 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6293) );
  MUX2_X1 U8016 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6293), .S(n6292), .Z(n6354)
         );
  INV_X1 U8017 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6558) );
  MUX2_X1 U8018 ( .A(n6558), .B(P2_REG1_REG_3__SCAN_IN), .S(n6347), .Z(n6341)
         );
  INV_X1 U8019 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6294) );
  MUX2_X1 U8020 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6294), .S(n9358), .Z(n9361)
         );
  XNOR2_X1 U8021 ( .A(n6295), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6367) );
  AND2_X1 U8022 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n6366) );
  NAND2_X1 U8023 ( .A1(n6367), .A2(n6366), .ZN(n6365) );
  NAND2_X1 U8024 ( .A1(n6375), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U8025 ( .A1(n6365), .A2(n6296), .ZN(n9362) );
  NAND2_X1 U8026 ( .A1(n9361), .A2(n9362), .ZN(n9360) );
  NAND2_X1 U8027 ( .A1(n9358), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U8028 ( .A1(n9360), .A2(n6297), .ZN(n6342) );
  NAND2_X1 U8029 ( .A1(n6341), .A2(n6342), .ZN(n6340) );
  OAI21_X1 U8030 ( .B1(n6347), .B2(n6558), .A(n6340), .ZN(n6355) );
  NAND2_X1 U8031 ( .A1(n6354), .A2(n6355), .ZN(n6353) );
  NAND2_X1 U8032 ( .A1(n6298), .A2(n6353), .ZN(n6315) );
  NAND2_X1 U8033 ( .A1(n6314), .A2(n6315), .ZN(n6313) );
  NAND2_X1 U8034 ( .A1(n6299), .A2(n6313), .ZN(n6303) );
  INV_X1 U8035 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6300) );
  MUX2_X1 U8036 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6300), .S(n6326), .Z(n6302)
         );
  OR2_X1 U8037 ( .A1(n6301), .A2(n8106), .ZN(n9699) );
  INV_X1 U8038 ( .A(n9699), .ZN(n9956) );
  NAND2_X1 U8039 ( .A1(n6302), .A2(n6303), .ZN(n6327) );
  OAI211_X1 U8040 ( .C1(n6303), .C2(n6302), .A(n9956), .B(n6327), .ZN(n6306)
         );
  NAND2_X1 U8041 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6728) );
  INV_X1 U8042 ( .A(n6728), .ZN(n6304) );
  AOI21_X1 U8043 ( .B1(n9960), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6304), .ZN(
        n6305) );
  OAI211_X1 U8044 ( .C1(n9964), .C2(n6307), .A(n6306), .B(n6305), .ZN(n6308)
         );
  OR2_X1 U8045 ( .A1(n6309), .A2(n6308), .ZN(P2_U3251) );
  AOI211_X1 U8046 ( .C1(n6312), .C2(n6311), .A(n6310), .B(n9951), .ZN(n6321)
         );
  OAI211_X1 U8047 ( .C1(n6315), .C2(n6314), .A(n9956), .B(n6313), .ZN(n6318)
         );
  AND2_X1 U8048 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6316) );
  AOI21_X1 U8049 ( .B1(n9960), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6316), .ZN(
        n6317) );
  OAI211_X1 U8050 ( .C1(n9964), .C2(n6319), .A(n6318), .B(n6317), .ZN(n6320)
         );
  OR2_X1 U8051 ( .A1(n6321), .A2(n6320), .ZN(P2_U3250) );
  INV_X1 U8052 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6323) );
  MUX2_X1 U8053 ( .A(n6323), .B(P2_REG2_REG_7__SCAN_IN), .S(n6460), .Z(n6324)
         );
  AOI211_X1 U8054 ( .C1(n6325), .C2(n6324), .A(n6455), .B(n9951), .ZN(n6336)
         );
  NAND2_X1 U8055 ( .A1(n6326), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U8056 ( .A1(n6328), .A2(n6327), .ZN(n6331) );
  INV_X1 U8057 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6329) );
  MUX2_X1 U8058 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6329), .S(n6460), .Z(n6330)
         );
  NAND2_X1 U8059 ( .A1(n6330), .A2(n6331), .ZN(n6461) );
  OAI211_X1 U8060 ( .C1(n6331), .C2(n6330), .A(n9956), .B(n6461), .ZN(n6333)
         );
  AND2_X1 U8061 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6760) );
  AOI21_X1 U8062 ( .B1(n9960), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6760), .ZN(
        n6332) );
  OAI211_X1 U8063 ( .C1(n9964), .C2(n6334), .A(n6333), .B(n6332), .ZN(n6335)
         );
  OR2_X1 U8064 ( .A1(n6336), .A2(n6335), .ZN(P2_U3252) );
  AOI211_X1 U8065 ( .C1(n6339), .C2(n6338), .A(n6337), .B(n9951), .ZN(n6349)
         );
  OAI211_X1 U8066 ( .C1(n6342), .C2(n6341), .A(n9956), .B(n6340), .ZN(n6346)
         );
  NOR2_X1 U8067 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6343), .ZN(n6344) );
  AOI21_X1 U8068 ( .B1(n9960), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6344), .ZN(
        n6345) );
  OAI211_X1 U8069 ( .C1(n9964), .C2(n6347), .A(n6346), .B(n6345), .ZN(n6348)
         );
  OR2_X1 U8070 ( .A1(n6349), .A2(n6348), .ZN(P2_U3248) );
  AOI211_X1 U8071 ( .C1(n6352), .C2(n6351), .A(n6350), .B(n9951), .ZN(n6362)
         );
  OAI211_X1 U8072 ( .C1(n6355), .C2(n6354), .A(n9956), .B(n6353), .ZN(n6359)
         );
  NOR2_X1 U8073 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6356), .ZN(n6357) );
  AOI21_X1 U8074 ( .B1(n9960), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6357), .ZN(
        n6358) );
  OAI211_X1 U8075 ( .C1(n9964), .C2(n6360), .A(n6359), .B(n6358), .ZN(n6361)
         );
  OR2_X1 U8076 ( .A1(n6362), .A2(n6361), .ZN(P2_U3249) );
  INV_X1 U8077 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U8078 ( .A1(n6579), .A2(P1_U4006), .ZN(n6363) );
  OAI21_X1 U8079 ( .B1(P1_U4006), .B2(n6364), .A(n6363), .ZN(P1_U3555) );
  INV_X1 U8080 ( .A(n9964), .ZN(n9359) );
  INV_X1 U8081 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8588) );
  OAI211_X1 U8082 ( .C1(n6367), .C2(n6366), .A(n9956), .B(n6365), .ZN(n6369)
         );
  INV_X1 U8083 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9378) );
  OR2_X1 U8084 ( .A1(n8362), .A2(n9378), .ZN(n6368) );
  OAI211_X1 U8085 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n8588), .A(n6369), .B(n6368), .ZN(n6374) );
  NAND2_X1 U8086 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n6372) );
  AOI211_X1 U8087 ( .C1(n6372), .C2(n6371), .A(n6370), .B(n9951), .ZN(n6373)
         );
  AOI211_X1 U8088 ( .C1(n9359), .C2(n6375), .A(n6374), .B(n6373), .ZN(n6376)
         );
  INV_X1 U8089 ( .A(n6376), .ZN(P2_U3246) );
  INV_X1 U8090 ( .A(n6377), .ZN(n6392) );
  AOI22_X1 U8091 ( .A1(n9557), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7485), .ZN(n6378) );
  OAI21_X1 U8092 ( .B1(n6392), .B2(n8117), .A(n6378), .ZN(P1_U3340) );
  INV_X1 U8093 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6391) );
  AND2_X1 U8094 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6912) );
  INV_X1 U8095 ( .A(n6379), .ZN(n6380) );
  AOI211_X1 U8096 ( .C1(n6382), .C2(n6381), .A(n6380), .B(n9625), .ZN(n6383)
         );
  AOI211_X1 U8097 ( .C1(n9619), .C2(n6384), .A(n6912), .B(n6383), .ZN(n6390)
         );
  AND3_X1 U8098 ( .A1(n9521), .A2(n6386), .A3(n6385), .ZN(n6387) );
  OAI21_X1 U8099 ( .B1(n6388), .B2(n6387), .A(n8895), .ZN(n6389) );
  OAI211_X1 U8100 ( .C1(n6391), .C2(n9628), .A(n6390), .B(n6389), .ZN(P1_U3246) );
  INV_X1 U8101 ( .A(n7046), .ZN(n7041) );
  OAI222_X1 U8102 ( .A1(n4267), .A2(n6393), .B1(n7519), .B2(n6392), .C1(n7041), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  NOR2_X1 U8103 ( .A1(n6394), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6396) );
  NOR2_X1 U8104 ( .A1(n6396), .A2(n6395), .ZN(n6400) );
  INV_X1 U8105 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6397) );
  MUX2_X1 U8106 ( .A(n6397), .B(P1_REG1_REG_10__SCAN_IN), .S(n6504), .Z(n6399)
         );
  OR2_X1 U8107 ( .A1(n6400), .A2(n6399), .ZN(n6500) );
  INV_X1 U8108 ( .A(n6500), .ZN(n6398) );
  AOI21_X1 U8109 ( .B1(n6400), .B2(n6399), .A(n6398), .ZN(n6413) );
  INV_X1 U8110 ( .A(n9628), .ZN(n9495) );
  NAND2_X1 U8111 ( .A1(n6402), .A2(n6401), .ZN(n6405) );
  INV_X1 U8112 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6403) );
  XNOR2_X1 U8113 ( .A(n6504), .B(n6403), .ZN(n6404) );
  NOR2_X1 U8114 ( .A1(n6405), .A2(n6404), .ZN(n6406) );
  OR2_X1 U8115 ( .A1(n6503), .A2(n6406), .ZN(n6410) );
  NAND2_X1 U8116 ( .A1(n9619), .A2(n6504), .ZN(n6409) );
  NOR2_X1 U8117 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6407), .ZN(n7300) );
  INV_X1 U8118 ( .A(n7300), .ZN(n6408) );
  OAI211_X1 U8119 ( .C1(n6410), .C2(n9613), .A(n6409), .B(n6408), .ZN(n6411)
         );
  AOI21_X1 U8120 ( .B1(n9495), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6411), .ZN(
        n6412) );
  OAI21_X1 U8121 ( .B1(n6413), .B2(n9625), .A(n6412), .ZN(P1_U3251) );
  INV_X1 U8122 ( .A(n6414), .ZN(n6448) );
  OAI222_X1 U8123 ( .A1(n8117), .A2(n6448), .B1(n8924), .B2(P1_U3084), .C1(
        n6415), .C2(n9349), .ZN(P1_U3339) );
  INV_X1 U8124 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6427) );
  INV_X1 U8125 ( .A(n6416), .ZN(n6421) );
  AND2_X1 U8126 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6751) );
  INV_X1 U8127 ( .A(n9625), .ZN(n9607) );
  OAI211_X1 U8128 ( .C1(n6418), .C2(n6417), .A(n9607), .B(n9525), .ZN(n6419)
         );
  INV_X1 U8129 ( .A(n6419), .ZN(n6420) );
  AOI211_X1 U8130 ( .C1(n9619), .C2(n6421), .A(n6751), .B(n6420), .ZN(n6426)
         );
  OAI211_X1 U8131 ( .C1(n6424), .C2(n6423), .A(n8895), .B(n6422), .ZN(n6425)
         );
  OAI211_X1 U8132 ( .C1(n6427), .C2(n9628), .A(n6426), .B(n6425), .ZN(P1_U3244) );
  INV_X1 U8133 ( .A(n8289), .ZN(n8239) );
  OAI21_X1 U8134 ( .B1(n6430), .B2(n6429), .A(n6428), .ZN(n6432) );
  OR2_X1 U8135 ( .A1(n6431), .A2(P2_U3152), .ZN(n6572) );
  AOI22_X1 U8136 ( .A1(n8239), .A2(n6432), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n6572), .ZN(n6435) );
  NAND2_X1 U8137 ( .A1(n5369), .A2(n8228), .ZN(n6433) );
  OAI21_X1 U8138 ( .B1(n4994), .B2(n8242), .A(n6433), .ZN(n8584) );
  AOI22_X1 U8139 ( .A1(n8281), .A2(n8584), .B1(n8590), .B2(n4262), .ZN(n6434)
         );
  NAND2_X1 U8140 ( .A1(n6435), .A2(n6434), .ZN(P2_U3224) );
  INV_X1 U8141 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U8142 ( .A1(n4266), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U8143 ( .A1(n4273), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U8144 ( .A1(n5840), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6436) );
  AND3_X1 U8145 ( .A1(n6438), .A2(n6437), .A3(n6436), .ZN(n8947) );
  INV_X1 U8146 ( .A(n8947), .ZN(n7609) );
  NAND2_X1 U8147 ( .A1(n7609), .A2(P1_U4006), .ZN(n6439) );
  OAI21_X1 U8148 ( .B1(P1_U4006), .B2(n6440), .A(n6439), .ZN(P1_U3586) );
  XNOR2_X1 U8149 ( .A(n6441), .B(n6442), .ZN(n6447) );
  OR2_X1 U8150 ( .A1(n4978), .A2(n8264), .ZN(n6444) );
  NAND2_X1 U8151 ( .A1(n8314), .A2(n8267), .ZN(n6443) );
  NAND2_X1 U8152 ( .A1(n6444), .A2(n6443), .ZN(n8564) );
  AOI22_X1 U8153 ( .A1(n8281), .A2(n8564), .B1(n8575), .B2(n4262), .ZN(n6446)
         );
  NAND2_X1 U8154 ( .A1(n6572), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6445) );
  OAI211_X1 U8155 ( .C1(n6447), .C2(n8289), .A(n6446), .B(n6445), .ZN(P2_U3239) );
  INV_X1 U8156 ( .A(n7258), .ZN(n7262) );
  OAI222_X1 U8157 ( .A1(n4267), .A2(n6449), .B1(n7519), .B2(n6448), .C1(n7262), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  XNOR2_X1 U8158 ( .A(n6451), .B(n6450), .ZN(n6454) );
  OAI22_X1 U8159 ( .A1(n4994), .A2(n8264), .B1(n5023), .B2(n8242), .ZN(n6551)
         );
  AOI22_X1 U8160 ( .A1(n8281), .A2(n6551), .B1(n7938), .B2(n4262), .ZN(n6453)
         );
  MUX2_X1 U8161 ( .A(n8285), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6452) );
  OAI211_X1 U8162 ( .C1(n6454), .C2(n8289), .A(n6453), .B(n6452), .ZN(P2_U3220) );
  INV_X1 U8163 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6928) );
  MUX2_X1 U8164 ( .A(n6928), .B(P2_REG2_REG_8__SCAN_IN), .S(n6459), .Z(n9953)
         );
  NOR2_X1 U8165 ( .A1(n9954), .A2(n9953), .ZN(n9952) );
  NAND2_X1 U8166 ( .A1(n6606), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6456) );
  OAI21_X1 U8167 ( .B1(n6606), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6456), .ZN(
        n6457) );
  AOI211_X1 U8168 ( .C1(n6458), .C2(n6457), .A(n6605), .B(n9951), .ZN(n6471)
         );
  INV_X1 U8169 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9768) );
  MUX2_X1 U8170 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9768), .S(n6459), .Z(n9957)
         );
  NAND2_X1 U8171 ( .A1(n6460), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U8172 ( .A1(n6462), .A2(n6461), .ZN(n9958) );
  NAND2_X1 U8173 ( .A1(n9957), .A2(n9958), .ZN(n9955) );
  OAI21_X1 U8174 ( .B1(n9963), .B2(n9768), .A(n9955), .ZN(n6465) );
  INV_X1 U8175 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6463) );
  MUX2_X1 U8176 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6463), .S(n6606), .Z(n6464)
         );
  NAND2_X1 U8177 ( .A1(n6464), .A2(n6465), .ZN(n6596) );
  OAI211_X1 U8178 ( .C1(n6465), .C2(n6464), .A(n9956), .B(n6596), .ZN(n6468)
         );
  NAND2_X1 U8179 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7025) );
  INV_X1 U8180 ( .A(n7025), .ZN(n6466) );
  AOI21_X1 U8181 ( .B1(n9960), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n6466), .ZN(
        n6467) );
  OAI211_X1 U8182 ( .C1(n9964), .C2(n6469), .A(n6468), .B(n6467), .ZN(n6470)
         );
  OR2_X1 U8183 ( .A1(n6471), .A2(n6470), .ZN(P2_U3254) );
  INV_X1 U8184 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6486) );
  INV_X1 U8185 ( .A(n6472), .ZN(n6475) );
  INV_X1 U8186 ( .A(n6473), .ZN(n6474) );
  AOI211_X1 U8187 ( .C1(n6476), .C2(n6475), .A(n6474), .B(n9625), .ZN(n6479)
         );
  NOR2_X1 U8188 ( .A1(n8888), .A2(n6477), .ZN(n6478) );
  AOI211_X1 U8189 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n6479), .B(
        n6478), .ZN(n6485) );
  NAND2_X1 U8190 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9487) );
  INV_X1 U8191 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6481) );
  MUX2_X1 U8192 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6481), .S(n6480), .Z(n6483)
         );
  OAI211_X1 U8193 ( .C1(n6177), .C2(n6483), .A(n8895), .B(n6482), .ZN(n6484)
         );
  OAI211_X1 U8194 ( .C1(n6486), .C2(n9628), .A(n6485), .B(n6484), .ZN(P1_U3242) );
  AOI21_X1 U8195 ( .B1(n6489), .B2(n6488), .A(n6487), .ZN(n6498) );
  OAI21_X1 U8196 ( .B1(n6492), .B2(n6491), .A(n6490), .ZN(n6495) );
  AND2_X1 U8197 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7227) );
  NOR2_X1 U8198 ( .A1(n8888), .A2(n6493), .ZN(n6494) );
  AOI211_X1 U8199 ( .C1(n9607), .C2(n6495), .A(n7227), .B(n6494), .ZN(n6497)
         );
  NAND2_X1 U8200 ( .A1(n9495), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6496) );
  OAI211_X1 U8201 ( .C1(n6498), .C2(n9613), .A(n6497), .B(n6496), .ZN(P1_U3248) );
  OR2_X1 U8202 ( .A1(n6504), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6499) );
  INV_X1 U8203 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9474) );
  AOI22_X1 U8204 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n8920), .B1(n8908), .B2(
        n9474), .ZN(n6501) );
  NOR2_X1 U8205 ( .A1(n6502), .A2(n6501), .ZN(n8919) );
  AOI21_X1 U8206 ( .B1(n6502), .B2(n6501), .A(n8919), .ZN(n6512) );
  NOR2_X1 U8207 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n8908), .ZN(n6505) );
  AOI21_X1 U8208 ( .B1(n8908), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6505), .ZN(
        n6506) );
  NAND2_X1 U8209 ( .A1(n6506), .A2(n6507), .ZN(n8907) );
  OAI21_X1 U8210 ( .B1(n6507), .B2(n6506), .A(n8907), .ZN(n6510) );
  INV_X1 U8211 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9817) );
  NOR2_X1 U8212 ( .A1(n9628), .A2(n9817), .ZN(n6509) );
  NAND2_X1 U8213 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8834) );
  OAI21_X1 U8214 ( .B1(n8888), .B2(n8920), .A(n8834), .ZN(n6508) );
  AOI211_X1 U8215 ( .C1(n8895), .C2(n6510), .A(n6509), .B(n6508), .ZN(n6511)
         );
  OAI21_X1 U8216 ( .B1(n6512), .B2(n9625), .A(n6511), .ZN(P1_U3252) );
  INV_X1 U8217 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6525) );
  OAI21_X1 U8218 ( .B1(n6515), .B2(n6514), .A(n6513), .ZN(n6519) );
  INV_X1 U8219 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6516) );
  NOR2_X1 U8220 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6516), .ZN(n7065) );
  NOR2_X1 U8221 ( .A1(n8888), .A2(n6517), .ZN(n6518) );
  AOI211_X1 U8222 ( .C1(n9607), .C2(n6519), .A(n7065), .B(n6518), .ZN(n6524)
         );
  OAI211_X1 U8223 ( .C1(n6522), .C2(n6521), .A(n8895), .B(n6520), .ZN(n6523)
         );
  OAI211_X1 U8224 ( .C1(n6525), .C2(n9628), .A(n6524), .B(n6523), .ZN(P1_U3247) );
  AND2_X1 U8225 ( .A1(n7812), .A2(n6526), .ZN(n9633) );
  AND2_X1 U8226 ( .A1(n9633), .A2(n6527), .ZN(n6528) );
  OAI211_X1 U8227 ( .C1(n9456), .C2(n6099), .A(n6528), .B(n6683), .ZN(n6535)
         );
  INV_X1 U8228 ( .A(n6679), .ZN(n9343) );
  INV_X1 U8229 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6534) );
  AND2_X1 U8230 ( .A1(n6579), .A2(n6586), .ZN(n7772) );
  NOR2_X1 U8231 ( .A1(n6782), .A2(n7772), .ZN(n7627) );
  NAND2_X1 U8232 ( .A1(n7818), .A2(n6713), .ZN(n6529) );
  OR2_X1 U8233 ( .A1(n7627), .A2(n6529), .ZN(n6532) );
  AND2_X1 U8234 ( .A1(n6530), .A2(n4269), .ZN(n9188) );
  NAND2_X1 U8235 ( .A1(n9188), .A2(n8885), .ZN(n6531) );
  AND2_X1 U8236 ( .A1(n6532), .A2(n6531), .ZN(n6709) );
  OAI21_X1 U8237 ( .B1(n6586), .B2(n6713), .A(n6709), .ZN(n6536) );
  NAND2_X1 U8238 ( .A1(n6536), .A2(n9685), .ZN(n6533) );
  OAI21_X1 U8239 ( .B1(n9685), .B2(n6534), .A(n6533), .ZN(P1_U3454) );
  INV_X1 U8240 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U8241 ( .A1(n6536), .A2(n9696), .ZN(n6537) );
  OAI21_X1 U8242 ( .B1(n9696), .B2(n9922), .A(n6537), .ZN(P1_U3523) );
  AOI21_X1 U8243 ( .B1(n4265), .B2(n6539), .A(n6538), .ZN(n9501) );
  INV_X1 U8244 ( .A(n8813), .ZN(n8866) );
  OAI21_X1 U8245 ( .B1(n9455), .B2(n6540), .A(n7240), .ZN(n7529) );
  AOI22_X1 U8246 ( .A1(n8866), .A2(n6715), .B1(n7529), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U8247 ( .A1(n8860), .A2(n8885), .ZN(n6541) );
  OAI211_X1 U8248 ( .C1(n9501), .C2(n8868), .A(n6542), .B(n6541), .ZN(P1_U3230) );
  INV_X1 U8249 ( .A(P1_U4006), .ZN(n8870) );
  NAND2_X1 U8250 ( .A1(n8870), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6543) );
  OAI21_X1 U8251 ( .B1(n9088), .B2(n8870), .A(n6543), .ZN(P1_U3580) );
  INV_X1 U8252 ( .A(n8243), .ZN(n8017) );
  NAND2_X1 U8253 ( .A1(n8017), .A2(P2_U3966), .ZN(n6544) );
  OAI21_X1 U8254 ( .B1(n6031), .B2(P2_U3966), .A(n6544), .ZN(P2_U3575) );
  OAI21_X1 U8255 ( .B1(n6547), .B2(n6546), .A(n6545), .ZN(n6703) );
  INV_X1 U8256 ( .A(n6703), .ZN(n6556) );
  INV_X1 U8257 ( .A(n9746), .ZN(n8674) );
  OAI21_X1 U8258 ( .B1(n6550), .B2(n6548), .A(n6549), .ZN(n6552) );
  AOI21_X1 U8259 ( .B1(n6552), .B2(n8585), .A(n6551), .ZN(n6708) );
  INV_X1 U8260 ( .A(n6553), .ZN(n8569) );
  INV_X1 U8261 ( .A(n6643), .ZN(n6554) );
  AOI21_X1 U8262 ( .B1(n7938), .B2(n8569), .A(n6554), .ZN(n6705) );
  AOI22_X1 U8263 ( .A1(n6705), .A2(n8670), .B1(n9722), .B2(n7938), .ZN(n6555)
         );
  OAI211_X1 U8264 ( .C1(n6556), .C2(n8674), .A(n6708), .B(n6555), .ZN(n6559)
         );
  NAND2_X1 U8265 ( .A1(n6559), .A2(n8676), .ZN(n6557) );
  OAI21_X1 U8266 ( .B1(n8676), .B2(n6558), .A(n6557), .ZN(P2_U3523) );
  INV_X1 U8267 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U8268 ( .A1(n6559), .A2(n9759), .ZN(n6560) );
  OAI21_X1 U8269 ( .B1(n9759), .B2(n6561), .A(n6560), .ZN(P2_U3460) );
  INV_X1 U8270 ( .A(n6562), .ZN(n6566) );
  AOI22_X1 U8271 ( .A1(n8322), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n6563), .ZN(n6564) );
  OAI21_X1 U8272 ( .B1(n6566), .B2(n7519), .A(n6564), .ZN(P2_U3342) );
  AOI22_X1 U8273 ( .A1(n9593), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7485), .ZN(n6565) );
  OAI21_X1 U8274 ( .B1(n6566), .B2(n8117), .A(n6565), .ZN(P1_U3337) );
  NAND2_X1 U8275 ( .A1(n5369), .A2(n6569), .ZN(n7924) );
  MUX2_X1 U8276 ( .A(n7924), .B(n6569), .S(n6567), .Z(n6568) );
  AOI21_X1 U8277 ( .B1(n8583), .B2(n6568), .A(n8289), .ZN(n6571) );
  INV_X1 U8278 ( .A(n8281), .ZN(n8269) );
  OR2_X1 U8279 ( .A1(n4978), .A2(n8242), .ZN(n6801) );
  OAI22_X1 U8280 ( .A1(n8269), .A2(n6801), .B1(n8274), .B2(n6569), .ZN(n6570)
         );
  AOI211_X1 U8281 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n6572), .A(n6571), .B(
        n6570), .ZN(n6573) );
  INV_X1 U8282 ( .A(n6573), .ZN(P2_U3234) );
  INV_X1 U8283 ( .A(n6574), .ZN(n6576) );
  INV_X1 U8284 ( .A(n9582), .ZN(n8926) );
  OAI222_X1 U8285 ( .A1(n9349), .A2(n6575), .B1(n8117), .B2(n6576), .C1(
        P1_U3084), .C2(n8926), .ZN(P1_U3338) );
  INV_X1 U8286 ( .A(n7425), .ZN(n7436) );
  OAI222_X1 U8287 ( .A1(n4267), .A2(n6577), .B1(n7519), .B2(n6576), .C1(
        P2_U3152), .C2(n7436), .ZN(P2_U3343) );
  AND2_X1 U8288 ( .A1(n6579), .A2(n6715), .ZN(n6581) );
  NAND2_X1 U8289 ( .A1(n6580), .A2(n6581), .ZN(n6774) );
  OAI21_X1 U8290 ( .B1(n6580), .B2(n6581), .A(n6774), .ZN(n6582) );
  INV_X1 U8291 ( .A(n6582), .ZN(n6684) );
  OR2_X1 U8292 ( .A1(n6583), .A2(n5676), .ZN(n6585) );
  NAND3_X1 U8293 ( .A1(n7815), .A2(n6099), .A3(n7809), .ZN(n6584) );
  AND2_X1 U8294 ( .A1(n6585), .A2(n6584), .ZN(n9664) );
  NAND2_X1 U8295 ( .A1(n9664), .A2(n9456), .ZN(n9681) );
  INV_X1 U8296 ( .A(n9455), .ZN(n9652) );
  OAI21_X1 U8297 ( .B1(n6586), .B2(n7773), .A(n6980), .ZN(n6587) );
  OR2_X1 U8298 ( .A1(n9679), .A2(n6587), .ZN(n6687) );
  OAI21_X1 U8299 ( .B1(n9652), .B2(n7773), .A(n6687), .ZN(n6591) );
  OR2_X1 U8300 ( .A1(n7765), .A2(n4269), .ZN(n9435) );
  XNOR2_X1 U8301 ( .A(n6580), .B(n6782), .ZN(n6590) );
  NAND2_X1 U8302 ( .A1(n7768), .A2(n9157), .ZN(n6589) );
  OR2_X1 U8303 ( .A1(n7647), .A2(n7771), .ZN(n6588) );
  OAI222_X1 U8304 ( .A1(n9437), .A2(n6775), .B1(n9435), .B2(n6615), .C1(n6590), 
        .C2(n9433), .ZN(n6689) );
  AOI211_X1 U8305 ( .C1(n6684), .C2(n9681), .A(n6591), .B(n6689), .ZN(n9637)
         );
  NAND2_X1 U8306 ( .A1(n9693), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6592) );
  OAI21_X1 U8307 ( .B1(n9637), .B2(n9693), .A(n6592), .ZN(P1_U3524) );
  INV_X1 U8308 ( .A(n6593), .ZN(n6638) );
  AOI22_X1 U8309 ( .A1(n9605), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7485), .ZN(n6594) );
  OAI21_X1 U8310 ( .B1(n6638), .B2(n8117), .A(n6594), .ZN(P1_U3336) );
  INV_X1 U8311 ( .A(n6661), .ZN(n6612) );
  NOR2_X1 U8312 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6595), .ZN(n6604) );
  NAND2_X1 U8313 ( .A1(n6606), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U8314 ( .A1(n6597), .A2(n6596), .ZN(n6598) );
  INV_X1 U8315 ( .A(n6598), .ZN(n6602) );
  INV_X1 U8316 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7108) );
  MUX2_X1 U8317 ( .A(n7108), .B(P2_REG1_REG_10__SCAN_IN), .S(n6661), .Z(n6601)
         );
  MUX2_X1 U8318 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7108), .S(n6661), .Z(n6599)
         );
  NAND2_X1 U8319 ( .A1(n6599), .A2(n6598), .ZN(n6651) );
  INV_X1 U8320 ( .A(n6651), .ZN(n6600) );
  AOI211_X1 U8321 ( .C1(n6602), .C2(n6601), .A(n6600), .B(n9699), .ZN(n6603)
         );
  AOI211_X1 U8322 ( .C1(n9960), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n6604), .B(
        n6603), .ZN(n6611) );
  XNOR2_X1 U8323 ( .A(n6661), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n6607) );
  AOI211_X1 U8324 ( .C1(n6608), .C2(n6607), .A(n6660), .B(n9951), .ZN(n6609)
         );
  INV_X1 U8325 ( .A(n6609), .ZN(n6610) );
  OAI211_X1 U8326 ( .C1(n9964), .C2(n6612), .A(n6611), .B(n6610), .ZN(P2_U3255) );
  NOR2_X1 U8327 ( .A1(n6613), .A2(n6614), .ZN(n7521) );
  AOI21_X1 U8328 ( .B1(n6614), .B2(n6613), .A(n7521), .ZN(n6619) );
  NOR2_X1 U8329 ( .A1(n8813), .A2(n7773), .ZN(n6617) );
  OAI22_X1 U8330 ( .A1(n8864), .A2(n6615), .B1(n6775), .B2(n8850), .ZN(n6616)
         );
  AOI211_X1 U8331 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n7529), .A(n6617), .B(
        n6616), .ZN(n6618) );
  OAI21_X1 U8332 ( .B1(n6619), .B2(n8868), .A(n6618), .ZN(P1_U3220) );
  INV_X1 U8333 ( .A(n6621), .ZN(n6622) );
  AOI21_X1 U8334 ( .B1(n6620), .B2(n6623), .A(n6622), .ZN(n6627) );
  AOI22_X1 U8335 ( .A1(n8312), .A2(n8267), .B1(n8228), .B2(n8314), .ZN(n6646)
         );
  AOI22_X1 U8336 ( .A1(n4262), .A2(n6644), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n6624) );
  OAI21_X1 U8337 ( .B1(n8269), .B2(n6646), .A(n6624), .ZN(n6625) );
  AOI21_X1 U8338 ( .B1(n6841), .B2(n8271), .A(n6625), .ZN(n6626) );
  OAI21_X1 U8339 ( .B1(n6627), .B2(n8289), .A(n6626), .ZN(P2_U3232) );
  XOR2_X1 U8340 ( .A(n6629), .B(n6628), .Z(n6636) );
  INV_X1 U8341 ( .A(n6630), .ZN(n6818) );
  AOI22_X1 U8342 ( .A1(n4262), .A2(n6821), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6634) );
  OR2_X1 U8343 ( .A1(n5023), .A2(n8264), .ZN(n6632) );
  NAND2_X1 U8344 ( .A1(n8311), .A2(n8267), .ZN(n6631) );
  NAND2_X1 U8345 ( .A1(n6632), .A2(n6631), .ZN(n6816) );
  NAND2_X1 U8346 ( .A1(n8281), .A2(n6816), .ZN(n6633) );
  OAI211_X1 U8347 ( .C1(n8285), .C2(n6818), .A(n6634), .B(n6633), .ZN(n6635)
         );
  AOI21_X1 U8348 ( .B1(n6636), .B2(n8239), .A(n6635), .ZN(n6637) );
  INV_X1 U8349 ( .A(n6637), .ZN(P2_U3229) );
  INV_X1 U8350 ( .A(n8337), .ZN(n8333) );
  OAI222_X1 U8351 ( .A1(n4267), .A2(n6639), .B1(n7519), .B2(n6638), .C1(n8333), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  OAI21_X1 U8352 ( .B1(n6641), .B2(n8070), .A(n6640), .ZN(n6846) );
  INV_X1 U8353 ( .A(n6822), .ZN(n6642) );
  AOI211_X1 U8354 ( .C1(n6644), .C2(n6643), .A(n9752), .B(n6642), .ZN(n6840)
         );
  XNOR2_X1 U8355 ( .A(n6645), .B(n8070), .ZN(n6647) );
  INV_X1 U8356 ( .A(n8585), .ZN(n8531) );
  OAI21_X1 U8357 ( .B1(n6647), .B2(n8531), .A(n6646), .ZN(n6839) );
  AOI211_X1 U8358 ( .C1(n9746), .C2(n6846), .A(n6840), .B(n6839), .ZN(n6722)
         );
  OAI22_X1 U8359 ( .A1(n8667), .A2(n6844), .B1(n8676), .B2(n6293), .ZN(n6648)
         );
  INV_X1 U8360 ( .A(n6648), .ZN(n6649) );
  OAI21_X1 U8361 ( .B1(n6722), .B2(n9767), .A(n6649), .ZN(P2_U3524) );
  INV_X1 U8362 ( .A(n6895), .ZN(n6668) );
  NOR2_X1 U8363 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5117), .ZN(n6659) );
  NAND2_X1 U8364 ( .A1(n6661), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U8365 ( .A1(n6651), .A2(n6650), .ZN(n6654) );
  INV_X1 U8366 ( .A(n6654), .ZN(n6657) );
  INV_X1 U8367 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6652) );
  MUX2_X1 U8368 ( .A(n6652), .B(P2_REG1_REG_11__SCAN_IN), .S(n6895), .Z(n6656)
         );
  MUX2_X1 U8369 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6652), .S(n6895), .Z(n6653)
         );
  NAND2_X1 U8370 ( .A1(n6654), .A2(n6653), .ZN(n6897) );
  INV_X1 U8371 ( .A(n6897), .ZN(n6655) );
  AOI211_X1 U8372 ( .C1(n6657), .C2(n6656), .A(n6655), .B(n9699), .ZN(n6658)
         );
  AOI211_X1 U8373 ( .C1(n9960), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n6659), .B(
        n6658), .ZN(n6667) );
  AOI21_X1 U8374 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n6661), .A(n6660), .ZN(
        n6664) );
  NOR2_X1 U8375 ( .A1(n6895), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6662) );
  AOI21_X1 U8376 ( .B1(n6895), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6662), .ZN(
        n6663) );
  NAND2_X1 U8377 ( .A1(n6664), .A2(n6663), .ZN(n6891) );
  OAI21_X1 U8378 ( .B1(n6664), .B2(n6663), .A(n6891), .ZN(n6665) );
  NAND2_X1 U8379 ( .A1(n9697), .A2(n6665), .ZN(n6666) );
  OAI211_X1 U8380 ( .C1(n9964), .C2(n6668), .A(n6667), .B(n6666), .ZN(P2_U3256) );
  NAND2_X1 U8381 ( .A1(n5840), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U8382 ( .A1(n4266), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6674) );
  INV_X1 U8383 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U8384 ( .A1(n6670), .A2(n6669), .ZN(n6671) );
  NAND2_X1 U8385 ( .A1(n4270), .A2(n9022), .ZN(n6673) );
  NAND2_X1 U8386 ( .A1(n4273), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U8387 ( .A1(n8870), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6676) );
  OAI21_X1 U8388 ( .B1(n9044), .B2(n8870), .A(n6676), .ZN(P1_U3583) );
  NAND2_X1 U8389 ( .A1(n8317), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6677) );
  OAI21_X1 U8390 ( .B1(n8182), .B2(n8317), .A(n6677), .ZN(P2_U3578) );
  NAND2_X1 U8391 ( .A1(n7647), .A2(n7812), .ZN(n6678) );
  NAND2_X1 U8392 ( .A1(n7812), .A2(n6679), .ZN(n6680) );
  NOR2_X1 U8393 ( .A1(n6681), .A2(n6680), .ZN(n6682) );
  NAND2_X1 U8394 ( .A1(n6683), .A2(n6682), .ZN(n6966) );
  NAND2_X2 U8395 ( .A1(n9419), .A2(n6966), .ZN(n9424) );
  AND2_X1 U8396 ( .A1(n5676), .A2(n9157), .ZN(n6938) );
  INV_X1 U8397 ( .A(n9664), .ZN(n9438) );
  OAI21_X1 U8398 ( .B1(n6938), .B2(n9438), .A(n6684), .ZN(n6686) );
  NAND2_X1 U8399 ( .A1(n9439), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6685) );
  OAI211_X1 U8400 ( .C1(n9157), .C2(n6687), .A(n6686), .B(n6685), .ZN(n6688)
         );
  OAI21_X1 U8401 ( .B1(n6689), .B2(n6688), .A(n9424), .ZN(n6693) );
  INV_X1 U8402 ( .A(n6690), .ZN(n6691) );
  NAND2_X1 U8403 ( .A1(n9424), .A2(n6691), .ZN(n9418) );
  INV_X1 U8404 ( .A(n7773), .ZN(n6783) );
  NAND2_X1 U8405 ( .A1(n9441), .A2(n6783), .ZN(n6692) );
  OAI211_X1 U8406 ( .C1(n6481), .C2(n9424), .A(n6693), .B(n6692), .ZN(P1_U3290) );
  INV_X1 U8407 ( .A(n6694), .ZN(n6698) );
  NOR2_X1 U8408 ( .A1(n6696), .A2(n6695), .ZN(n6697) );
  NAND2_X1 U8409 ( .A1(n6698), .A2(n6697), .ZN(n6739) );
  OR2_X1 U8410 ( .A1(n6699), .A2(n8357), .ZN(n6921) );
  NAND2_X1 U8411 ( .A1(n7170), .A2(n6921), .ZN(n6700) );
  NOR2_X1 U8412 ( .A1(n5430), .A2(n6701), .ZN(n6702) );
  AOI22_X1 U8413 ( .A1(n6703), .A2(n8582), .B1(n8581), .B2(n7938), .ZN(n6707)
         );
  NOR2_X1 U8414 ( .A1(n6739), .A2(n7909), .ZN(n8593) );
  OAI22_X1 U8415 ( .A1(n8567), .A2(n6272), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8587), .ZN(n6704) );
  AOI21_X1 U8416 ( .B1(n8593), .B2(n6705), .A(n6704), .ZN(n6706) );
  OAI211_X1 U8417 ( .C1(n6708), .C2(n8462), .A(n6707), .B(n6706), .ZN(P2_U3293) );
  INV_X1 U8418 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6718) );
  INV_X1 U8419 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6710) );
  OAI21_X1 U8420 ( .B1(n6710), .B2(n9419), .A(n6709), .ZN(n6711) );
  NAND2_X1 U8421 ( .A1(n6711), .A2(n9424), .ZN(n6717) );
  NOR2_X1 U8422 ( .A1(n6713), .A2(n6712), .ZN(n6714) );
  OAI21_X1 U8423 ( .B1(n9441), .B2(n9446), .A(n6715), .ZN(n6716) );
  OAI211_X1 U8424 ( .C1(n6718), .C2(n9424), .A(n6717), .B(n6716), .ZN(P1_U3291) );
  INV_X1 U8425 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6719) );
  OAI22_X1 U8426 ( .A1(n8711), .A2(n6844), .B1(n9759), .B2(n6719), .ZN(n6720)
         );
  INV_X1 U8427 ( .A(n6720), .ZN(n6721) );
  OAI21_X1 U8428 ( .B1(n6722), .B2(n9758), .A(n6721), .ZN(P2_U3463) );
  OAI21_X1 U8429 ( .B1(n6725), .B2(n6724), .A(n6723), .ZN(n6732) );
  NOR2_X1 U8430 ( .A1(n8285), .A2(n6878), .ZN(n6731) );
  OR2_X1 U8431 ( .A1(n6726), .A2(n8264), .ZN(n6727) );
  OAI21_X1 U8432 ( .B1(n6851), .B2(n8242), .A(n6727), .ZN(n6884) );
  NAND2_X1 U8433 ( .A1(n8281), .A2(n6884), .ZN(n6729) );
  OAI211_X1 U8434 ( .C1(n8274), .C2(n9743), .A(n6729), .B(n6728), .ZN(n6730)
         );
  AOI211_X1 U8435 ( .C1(n6732), .C2(n8239), .A(n6731), .B(n6730), .ZN(n6733)
         );
  INV_X1 U8436 ( .A(n6733), .ZN(P2_U3241) );
  XNOR2_X1 U8437 ( .A(n6734), .B(n8076), .ZN(n6736) );
  INV_X1 U8438 ( .A(n8309), .ZN(n7952) );
  OAI22_X1 U8439 ( .A1(n6735), .A2(n8264), .B1(n7952), .B2(n8242), .ZN(n6761)
         );
  AOI21_X1 U8440 ( .B1(n6736), .B2(n8585), .A(n6761), .ZN(n6792) );
  XOR2_X1 U8441 ( .A(n6737), .B(n8076), .Z(n6793) );
  OR2_X1 U8442 ( .A1(n6793), .A2(n8559), .ZN(n6745) );
  INV_X1 U8443 ( .A(n6762), .ZN(n6738) );
  OAI22_X1 U8444 ( .A1(n8567), .A2(n6323), .B1(n6738), .B2(n8587), .ZN(n6742)
         );
  OAI211_X1 U8445 ( .C1(n6876), .C2(n6797), .A(n8670), .B(n6930), .ZN(n6791)
         );
  INV_X1 U8446 ( .A(n6739), .ZN(n6740) );
  NAND2_X1 U8447 ( .A1(n6740), .A2(n8357), .ZN(n8370) );
  NOR2_X1 U8448 ( .A1(n6791), .A2(n8370), .ZN(n6741) );
  AOI211_X1 U8449 ( .C1(n8581), .C2(n6743), .A(n6742), .B(n6741), .ZN(n6744)
         );
  OAI211_X1 U8450 ( .C1(n8462), .C2(n6792), .A(n6745), .B(n6744), .ZN(P2_U3289) );
  INV_X1 U8451 ( .A(n6746), .ZN(n6748) );
  NOR2_X1 U8452 ( .A1(n6748), .A2(n6747), .ZN(n6749) );
  XNOR2_X1 U8453 ( .A(n6750), .B(n6749), .ZN(n6756) );
  AOI21_X1 U8454 ( .B1(n8860), .B2(n8882), .A(n6751), .ZN(n6753) );
  NAND2_X1 U8455 ( .A1(n8848), .A2(n8884), .ZN(n6752) );
  OAI211_X1 U8456 ( .C1(n9644), .C2(n8813), .A(n6753), .B(n6752), .ZN(n6754)
         );
  AOI21_X1 U8457 ( .B1(n6779), .B2(n8861), .A(n6754), .ZN(n6755) );
  OAI21_X1 U8458 ( .B1(n6756), .B2(n8868), .A(n6755), .ZN(P1_U3216) );
  XNOR2_X1 U8459 ( .A(n6758), .B(n6757), .ZN(n6765) );
  NOR2_X1 U8460 ( .A1(n8274), .A2(n6797), .ZN(n6759) );
  AOI211_X1 U8461 ( .C1(n8281), .C2(n6761), .A(n6760), .B(n6759), .ZN(n6764)
         );
  NAND2_X1 U8462 ( .A1(n8271), .A2(n6762), .ZN(n6763) );
  OAI211_X1 U8463 ( .C1(n6765), .C2(n8289), .A(n6764), .B(n6763), .ZN(P2_U3215) );
  INV_X1 U8464 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6767) );
  INV_X1 U8465 ( .A(n6766), .ZN(n6768) );
  INV_X1 U8466 ( .A(n9620), .ZN(n8931) );
  OAI222_X1 U8467 ( .A1(n9349), .A2(n6767), .B1(n8117), .B2(n6768), .C1(
        P1_U3084), .C2(n8931), .ZN(P1_U3335) );
  INV_X1 U8468 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6769) );
  INV_X1 U8469 ( .A(n8342), .ZN(n8351) );
  OAI222_X1 U8470 ( .A1(n4267), .A2(n6769), .B1(n7519), .B2(n6768), .C1(
        P2_U3152), .C2(n8351), .ZN(P2_U3340) );
  NAND2_X1 U8471 ( .A1(n8317), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6770) );
  OAI21_X1 U8472 ( .B1(n6771), .B2(n8317), .A(n6770), .ZN(P2_U3581) );
  AND2_X1 U8473 ( .A1(n7818), .A2(n4268), .ZN(n6772) );
  NAND2_X1 U8474 ( .A1(n9424), .A2(n6772), .ZN(n9217) );
  INV_X1 U8475 ( .A(n9217), .ZN(n7853) );
  NAND2_X1 U8476 ( .A1(n8885), .A2(n6783), .ZN(n6773) );
  NAND2_X1 U8477 ( .A1(n8884), .A2(n9639), .ZN(n7778) );
  NAND2_X1 U8478 ( .A1(n6775), .A2(n6984), .ZN(n7777) );
  NAND2_X1 U8479 ( .A1(n6775), .A2(n9639), .ZN(n6776) );
  NAND2_X1 U8480 ( .A1(n6978), .A2(n6776), .ZN(n6778) );
  NAND2_X1 U8481 ( .A1(n6777), .A2(n6780), .ZN(n7780) );
  NAND2_X1 U8482 ( .A1(n8883), .A2(n9644), .ZN(n7579) );
  NAND2_X1 U8483 ( .A1(n6778), .A2(n6859), .ZN(n6857) );
  OAI21_X1 U8484 ( .B1(n6778), .B2(n6859), .A(n6857), .ZN(n9648) );
  INV_X1 U8485 ( .A(n9446), .ZN(n9200) );
  OAI21_X1 U8486 ( .B1(n6982), .B2(n9644), .A(n6866), .ZN(n9645) );
  AOI22_X1 U8487 ( .A1(n9441), .A2(n6780), .B1(n9439), .B2(n6779), .ZN(n6781)
         );
  OAI21_X1 U8488 ( .B1(n9200), .B2(n9645), .A(n6781), .ZN(n6789) );
  INV_X1 U8489 ( .A(n6580), .ZN(n7625) );
  NAND2_X1 U8490 ( .A1(n7526), .A2(n6783), .ZN(n6784) );
  NAND2_X1 U8491 ( .A1(n6974), .A2(n7626), .ZN(n6786) );
  XNOR2_X1 U8492 ( .A(n6859), .B(n7582), .ZN(n6787) );
  OAI222_X1 U8493 ( .A1(n9437), .A2(n7839), .B1(n9435), .B2(n6775), .C1(n6787), 
        .C2(n9433), .ZN(n9646) );
  MUX2_X1 U8494 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9646), .S(n9424), .Z(n6788)
         );
  AOI211_X1 U8495 ( .C1(n7853), .C2(n9648), .A(n6789), .B(n6788), .ZN(n6790)
         );
  INV_X1 U8496 ( .A(n6790), .ZN(P1_U3288) );
  OAI211_X1 U8497 ( .C1(n6793), .C2(n8674), .A(n6792), .B(n6791), .ZN(n6799)
         );
  OAI22_X1 U8498 ( .A1(n8667), .A2(n6797), .B1(n8676), .B2(n6329), .ZN(n6794)
         );
  AOI21_X1 U8499 ( .B1(n6799), .B2(n8676), .A(n6794), .ZN(n6795) );
  INV_X1 U8500 ( .A(n6795), .ZN(P2_U3527) );
  INV_X1 U8501 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6796) );
  OAI22_X1 U8502 ( .A1(n8711), .A2(n6797), .B1(n9759), .B2(n6796), .ZN(n6798)
         );
  AOI21_X1 U8503 ( .B1(n6799), .B2(n9759), .A(n6798), .ZN(n6800) );
  INV_X1 U8504 ( .A(n6800), .ZN(P2_U3472) );
  NAND2_X1 U8505 ( .A1(n8583), .A2(n7924), .ZN(n9717) );
  INV_X1 U8506 ( .A(n9717), .ZN(n6807) );
  NAND2_X1 U8507 ( .A1(n9717), .A2(n8585), .ZN(n6802) );
  AND2_X1 U8508 ( .A1(n6802), .A2(n6801), .ZN(n9719) );
  INV_X1 U8509 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6803) );
  OAI22_X1 U8510 ( .A1(n8462), .A2(n9719), .B1(n6803), .B2(n8587), .ZN(n6804)
         );
  AOI21_X1 U8511 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n8462), .A(n6804), .ZN(
        n6806) );
  OAI21_X1 U8512 ( .B1(n8581), .B2(n8593), .A(n9715), .ZN(n6805) );
  OAI211_X1 U8513 ( .C1(n6807), .C2(n8559), .A(n6806), .B(n6805), .ZN(P2_U3296) );
  INV_X1 U8514 ( .A(n6808), .ZN(n6810) );
  OAI222_X1 U8515 ( .A1(n4267), .A2(n6809), .B1(n7519), .B2(n6810), .C1(
        P2_U3152), .C2(n8357), .ZN(P2_U3339) );
  OAI222_X1 U8516 ( .A1(n9349), .A2(n6811), .B1(n8117), .B2(n6810), .C1(n4434), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  XNOR2_X1 U8517 ( .A(n6812), .B(n8073), .ZN(n9739) );
  NAND2_X1 U8518 ( .A1(n6813), .A2(n6814), .ZN(n6815) );
  XNOR2_X1 U8519 ( .A(n6815), .B(n8073), .ZN(n6817) );
  AOI21_X1 U8520 ( .B1(n6817), .B2(n8585), .A(n6816), .ZN(n9736) );
  INV_X1 U8521 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6819) );
  OAI22_X1 U8522 ( .A1(n8567), .A2(n6819), .B1(n6818), .B2(n8587), .ZN(n6820)
         );
  AOI21_X1 U8523 ( .B1(n8581), .B2(n6821), .A(n6820), .ZN(n6827) );
  NAND2_X1 U8524 ( .A1(n6822), .A2(n6821), .ZN(n6823) );
  NAND2_X1 U8525 ( .A1(n6823), .A2(n8670), .ZN(n6824) );
  OR2_X1 U8526 ( .A1(n6875), .A2(n6824), .ZN(n9735) );
  INV_X1 U8527 ( .A(n9735), .ZN(n6825) );
  NAND2_X1 U8528 ( .A1(n8572), .A2(n6825), .ZN(n6826) );
  OAI211_X1 U8529 ( .C1(n9736), .C2(n8462), .A(n6827), .B(n6826), .ZN(n6828)
         );
  AOI21_X1 U8530 ( .B1(n8582), .B2(n9739), .A(n6828), .ZN(n6829) );
  INV_X1 U8531 ( .A(n6829), .ZN(P2_U3291) );
  OAI21_X1 U8532 ( .B1(n6832), .B2(n6831), .A(n6830), .ZN(n6833) );
  NAND2_X1 U8533 ( .A1(n6833), .A2(n8806), .ZN(n6838) );
  AND2_X1 U8534 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9531) );
  AOI21_X1 U8535 ( .B1(n8848), .B2(n8883), .A(n9531), .ZN(n6835) );
  OR2_X1 U8536 ( .A1(n8813), .A2(n6957), .ZN(n6834) );
  OAI211_X1 U8537 ( .C1(n6950), .C2(n8850), .A(n6835), .B(n6834), .ZN(n6836)
         );
  AOI21_X1 U8538 ( .B1(n6940), .B2(n8861), .A(n6836), .ZN(n6837) );
  NAND2_X1 U8539 ( .A1(n6838), .A2(n6837), .ZN(P1_U3228) );
  INV_X1 U8540 ( .A(n6839), .ZN(n6848) );
  NAND2_X1 U8541 ( .A1(n6840), .A2(n8572), .ZN(n6843) );
  INV_X1 U8542 ( .A(n8587), .ZN(n8566) );
  AOI22_X1 U8543 ( .A1(n8462), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n6841), .B2(
        n8566), .ZN(n6842) );
  OAI211_X1 U8544 ( .C1(n8556), .C2(n6844), .A(n6843), .B(n6842), .ZN(n6845)
         );
  AOI21_X1 U8545 ( .B1(n6846), .B2(n8582), .A(n6845), .ZN(n6847) );
  OAI21_X1 U8546 ( .B1(n6848), .B2(n8462), .A(n6847), .ZN(P2_U3292) );
  XNOR2_X1 U8547 ( .A(n6850), .B(n6849), .ZN(n6855) );
  OAI22_X1 U8548 ( .A1(n6851), .A2(n8264), .B1(n7015), .B2(n8242), .ZN(n6924)
         );
  AOI22_X1 U8549 ( .A1(n8281), .A2(n6924), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n6852) );
  OAI21_X1 U8550 ( .B1(n6927), .B2(n8285), .A(n6852), .ZN(n6853) );
  AOI21_X1 U8551 ( .B1(n6935), .B2(n4262), .A(n6853), .ZN(n6854) );
  OAI21_X1 U8552 ( .B1(n6855), .B2(n8289), .A(n6854), .ZN(P2_U3223) );
  NAND2_X1 U8553 ( .A1(n6777), .A2(n9644), .ZN(n6856) );
  NAND2_X1 U8554 ( .A1(n6857), .A2(n6856), .ZN(n6858) );
  NAND2_X1 U8555 ( .A1(n7839), .A2(n6867), .ZN(n7657) );
  NAND2_X1 U8556 ( .A1(n7657), .A2(n7583), .ZN(n6862) );
  OAI21_X1 U8557 ( .B1(n6858), .B2(n6862), .A(n6959), .ZN(n6944) );
  INV_X1 U8558 ( .A(n6944), .ZN(n6869) );
  OAI22_X1 U8559 ( .A1(n9437), .A2(n6950), .B1(n6777), .B2(n9435), .ZN(n6865)
         );
  INV_X1 U8560 ( .A(n6859), .ZN(n6860) );
  NAND2_X1 U8561 ( .A1(n7582), .A2(n6860), .ZN(n6861) );
  XNOR2_X1 U8562 ( .A(n6862), .B(n6947), .ZN(n6863) );
  NOR2_X1 U8563 ( .A1(n6863), .A2(n9433), .ZN(n6864) );
  AOI211_X1 U8564 ( .C1(n9438), .C2(n6944), .A(n6865), .B(n6864), .ZN(n6946)
         );
  INV_X1 U8565 ( .A(n6965), .ZN(n7837) );
  AOI21_X1 U8566 ( .B1(n6867), .B2(n6866), .A(n7837), .ZN(n6939) );
  AOI22_X1 U8567 ( .A1(n6939), .A2(n9661), .B1(n9455), .B2(n6867), .ZN(n6868)
         );
  OAI211_X1 U8568 ( .C1(n6869), .C2(n9456), .A(n6946), .B(n6868), .ZN(n6871)
         );
  NAND2_X1 U8569 ( .A1(n6871), .A2(n9696), .ZN(n6870) );
  OAI21_X1 U8570 ( .B1(n9696), .B2(n6198), .A(n6870), .ZN(P1_U3527) );
  INV_X1 U8571 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U8572 ( .A1(n6871), .A2(n9685), .ZN(n6872) );
  OAI21_X1 U8573 ( .B1(n9685), .B2(n6873), .A(n6872), .ZN(P1_U3466) );
  XNOR2_X1 U8574 ( .A(n6874), .B(n4712), .ZN(n9745) );
  INV_X1 U8575 ( .A(n9745), .ZN(n6890) );
  OAI21_X1 U8576 ( .B1(n6875), .B2(n9743), .A(n8670), .ZN(n6877) );
  OR2_X1 U8577 ( .A1(n6877), .A2(n6876), .ZN(n9741) );
  NOR2_X1 U8578 ( .A1(n8587), .A2(n6878), .ZN(n6879) );
  AOI21_X1 U8579 ( .B1(n8462), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6879), .ZN(
        n6880) );
  OAI21_X1 U8580 ( .B1(n8370), .B2(n9741), .A(n6880), .ZN(n6887) );
  OAI21_X1 U8581 ( .B1(n6883), .B2(n6881), .A(n6882), .ZN(n6885) );
  AOI21_X1 U8582 ( .B1(n6885), .B2(n8585), .A(n6884), .ZN(n9742) );
  NOR2_X1 U8583 ( .A1(n9742), .A2(n8462), .ZN(n6886) );
  AOI211_X1 U8584 ( .C1(n8581), .C2(n6888), .A(n6887), .B(n6886), .ZN(n6889)
         );
  OAI21_X1 U8585 ( .B1(n6890), .B2(n8559), .A(n6889), .ZN(P2_U3290) );
  INV_X1 U8586 ( .A(n6996), .ZN(n6907) );
  XNOR2_X1 U8587 ( .A(n6996), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n6893) );
  AOI211_X1 U8588 ( .C1(n6893), .C2(n6892), .A(n6995), .B(n9951), .ZN(n6894)
         );
  INV_X1 U8589 ( .A(n6894), .ZN(n6906) );
  NAND2_X1 U8590 ( .A1(n6895), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6896) );
  AND2_X1 U8591 ( .A1(n6897), .A2(n6896), .ZN(n6899) );
  INV_X1 U8592 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7315) );
  MUX2_X1 U8593 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7315), .S(n6996), .Z(n6898)
         );
  NAND2_X1 U8594 ( .A1(n6899), .A2(n6898), .ZN(n6993) );
  OAI21_X1 U8595 ( .B1(n6899), .B2(n6898), .A(n6993), .ZN(n6904) );
  NOR2_X1 U8596 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6900), .ZN(n6903) );
  INV_X1 U8597 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6901) );
  NOR2_X1 U8598 ( .A1(n8362), .A2(n6901), .ZN(n6902) );
  AOI211_X1 U8599 ( .C1(n9956), .C2(n6904), .A(n6903), .B(n6902), .ZN(n6905)
         );
  OAI211_X1 U8600 ( .C1(n9964), .C2(n6907), .A(n6906), .B(n6905), .ZN(P2_U3257) );
  XNOR2_X1 U8601 ( .A(n6909), .B(n6908), .ZN(n6910) );
  XNOR2_X1 U8602 ( .A(n6911), .B(n6910), .ZN(n6917) );
  AOI21_X1 U8603 ( .B1(n8860), .B2(n8880), .A(n6912), .ZN(n6914) );
  NAND2_X1 U8604 ( .A1(n8848), .A2(n8882), .ZN(n6913) );
  OAI211_X1 U8605 ( .C1(n9653), .C2(n8813), .A(n6914), .B(n6913), .ZN(n6915)
         );
  AOI21_X1 U8606 ( .B1(n7846), .B2(n8861), .A(n6915), .ZN(n6916) );
  OAI21_X1 U8607 ( .B1(n6917), .B2(n8868), .A(n6916), .ZN(P1_U3225) );
  NAND2_X1 U8608 ( .A1(n6918), .A2(n8075), .ZN(n6919) );
  NAND2_X1 U8609 ( .A1(n6920), .A2(n6919), .ZN(n9749) );
  INV_X1 U8610 ( .A(n6921), .ZN(n6922) );
  NAND2_X1 U8611 ( .A1(n8567), .A2(n6922), .ZN(n7180) );
  XNOR2_X1 U8612 ( .A(n6923), .B(n5085), .ZN(n6925) );
  AOI21_X1 U8613 ( .B1(n6925), .B2(n8585), .A(n6924), .ZN(n6926) );
  OAI21_X1 U8614 ( .B1(n9749), .B2(n7170), .A(n6926), .ZN(n9754) );
  NAND2_X1 U8615 ( .A1(n9754), .A2(n8567), .ZN(n6937) );
  OAI22_X1 U8616 ( .A1(n8567), .A2(n6928), .B1(n6927), .B2(n8587), .ZN(n6934)
         );
  INV_X1 U8617 ( .A(n6929), .ZN(n7176) );
  NAND2_X1 U8618 ( .A1(n6930), .A2(n6935), .ZN(n6931) );
  NAND2_X1 U8619 ( .A1(n7176), .A2(n6931), .ZN(n9753) );
  INV_X1 U8620 ( .A(n8593), .ZN(n6932) );
  NOR2_X1 U8621 ( .A1(n9753), .A2(n6932), .ZN(n6933) );
  AOI211_X1 U8622 ( .C1(n8581), .C2(n6935), .A(n6934), .B(n6933), .ZN(n6936)
         );
  OAI211_X1 U8623 ( .C1(n9749), .C2(n7180), .A(n6937), .B(n6936), .ZN(P2_U3288) );
  NAND2_X1 U8624 ( .A1(n9424), .A2(n6938), .ZN(n9233) );
  INV_X1 U8625 ( .A(n9233), .ZN(n9447) );
  NAND2_X1 U8626 ( .A1(n6939), .A2(n9446), .ZN(n6942) );
  AOI22_X1 U8627 ( .A1(n9451), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n6940), .B2(
        n9439), .ZN(n6941) );
  OAI211_X1 U8628 ( .C1(n6957), .C2(n9418), .A(n6942), .B(n6941), .ZN(n6943)
         );
  AOI21_X1 U8629 ( .B1(n6944), .B2(n9447), .A(n6943), .ZN(n6945) );
  OAI21_X1 U8630 ( .B1(n6946), .B2(n9451), .A(n6945), .ZN(P1_U3287) );
  NAND2_X1 U8631 ( .A1(n7840), .A2(n7824), .ZN(n7662) );
  NAND2_X1 U8632 ( .A1(n8880), .A2(n7825), .ZN(n7660) );
  INV_X1 U8633 ( .A(n6950), .ZN(n8881) );
  NAND2_X1 U8634 ( .A1(n8881), .A2(n9653), .ZN(n7659) );
  NAND2_X1 U8635 ( .A1(n7660), .A2(n7659), .ZN(n6948) );
  NAND2_X1 U8636 ( .A1(n6950), .A2(n7852), .ZN(n6960) );
  NAND2_X1 U8637 ( .A1(n7662), .A2(n6960), .ZN(n7585) );
  INV_X1 U8638 ( .A(n7657), .ZN(n6951) );
  OR2_X1 U8639 ( .A1(n7585), .A2(n6951), .ZN(n6952) );
  NAND2_X1 U8640 ( .A1(n6952), .A2(n6949), .ZN(n7785) );
  NAND2_X1 U8641 ( .A1(n6954), .A2(n7785), .ZN(n6953) );
  NAND2_X1 U8642 ( .A1(n7132), .A2(n7226), .ZN(n7661) );
  INV_X1 U8643 ( .A(n7132), .ZN(n8879) );
  NAND2_X1 U8644 ( .A1(n8879), .A2(n7114), .ZN(n7664) );
  NAND2_X1 U8645 ( .A1(n7661), .A2(n7664), .ZN(n6963) );
  INV_X1 U8646 ( .A(n6963), .ZN(n7629) );
  NAND3_X1 U8647 ( .A1(n6954), .A2(n7785), .A3(n6963), .ZN(n6955) );
  NAND2_X1 U8648 ( .A1(n7119), .A2(n6955), .ZN(n6956) );
  INV_X1 U8649 ( .A(n9435), .ZN(n9136) );
  AOI222_X1 U8650 ( .A1(n9414), .A2(n6956), .B1(n8880), .B2(n9136), .C1(n8878), 
        .C2(n9188), .ZN(n9672) );
  NAND2_X1 U8651 ( .A1(n7839), .A2(n6957), .ZN(n6958) );
  NAND2_X1 U8652 ( .A1(n8881), .A2(n7852), .ZN(n6962) );
  NAND2_X1 U8653 ( .A1(n7851), .A2(n6962), .ZN(n7822) );
  OAI21_X1 U8654 ( .B1(n6964), .B2(n6963), .A(n7116), .ZN(n9674) );
  NAND2_X1 U8655 ( .A1(n9674), .A2(n7853), .ZN(n6971) );
  NAND2_X1 U8656 ( .A1(n7823), .A2(n7114), .ZN(n7141) );
  OAI211_X1 U8657 ( .C1(n7823), .C2(n7114), .A(n7141), .B(n9661), .ZN(n9670)
         );
  INV_X1 U8658 ( .A(n9670), .ZN(n6969) );
  NOR2_X1 U8659 ( .A1(n6966), .A2(n9157), .ZN(n9210) );
  AOI22_X1 U8660 ( .A1(n9451), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7228), .B2(
        n9439), .ZN(n6967) );
  OAI21_X1 U8661 ( .B1(n7114), .B2(n9418), .A(n6967), .ZN(n6968) );
  AOI21_X1 U8662 ( .B1(n6969), .B2(n9210), .A(n6968), .ZN(n6970) );
  OAI211_X1 U8663 ( .C1(n9672), .C2(n9451), .A(n6971), .B(n6970), .ZN(P1_U3284) );
  INV_X1 U8664 ( .A(n6972), .ZN(n7511) );
  OAI222_X1 U8665 ( .A1(n8117), .A2(n7511), .B1(P1_U3084), .B2(n7771), .C1(
        n6973), .C2(n9349), .ZN(P1_U3333) );
  XNOR2_X1 U8666 ( .A(n6974), .B(n7626), .ZN(n6975) );
  NAND2_X1 U8667 ( .A1(n6975), .A2(n9414), .ZN(n6977) );
  AOI22_X1 U8668 ( .A1(n8883), .A2(n9188), .B1(n9136), .B2(n8885), .ZN(n6976)
         );
  NAND2_X1 U8669 ( .A1(n6977), .A2(n6976), .ZN(n9640) );
  INV_X1 U8670 ( .A(n9640), .ZN(n6989) );
  OAI21_X1 U8671 ( .B1(n6979), .B2(n6785), .A(n6978), .ZN(n9642) );
  INV_X1 U8672 ( .A(n9210), .ZN(n7339) );
  NAND2_X1 U8673 ( .A1(n6980), .A2(n6984), .ZN(n6981) );
  NAND2_X1 U8674 ( .A1(n9661), .A2(n6981), .ZN(n6983) );
  OR2_X1 U8675 ( .A1(n6983), .A2(n6982), .ZN(n9638) );
  AOI22_X1 U8676 ( .A1(n9451), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9439), .ZN(n6986) );
  NAND2_X1 U8677 ( .A1(n9441), .A2(n6984), .ZN(n6985) );
  OAI211_X1 U8678 ( .C1(n7339), .C2(n9638), .A(n6986), .B(n6985), .ZN(n6987)
         );
  AOI21_X1 U8679 ( .B1(n9642), .B2(n7853), .A(n6987), .ZN(n6988) );
  OAI21_X1 U8680 ( .B1(n6989), .B2(n9451), .A(n6988), .ZN(P1_U3289) );
  INV_X1 U8681 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6990) );
  MUX2_X1 U8682 ( .A(n6990), .B(P2_REG1_REG_13__SCAN_IN), .S(n7046), .Z(n6991)
         );
  OR2_X1 U8683 ( .A1(n6996), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6992) );
  AND2_X1 U8684 ( .A1(n6991), .A2(n6992), .ZN(n6994) );
  AOI21_X1 U8685 ( .B1(n6993), .B2(n6992), .A(n6991), .ZN(n7040) );
  AOI21_X1 U8686 ( .B1(n6994), .B2(n6993), .A(n7040), .ZN(n7004) );
  NOR2_X1 U8687 ( .A1(n7046), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6997) );
  AOI21_X1 U8688 ( .B1(n7046), .B2(P2_REG2_REG_13__SCAN_IN), .A(n6997), .ZN(
        n6998) );
  OAI21_X1 U8689 ( .B1(n6999), .B2(n6998), .A(n7045), .ZN(n7000) );
  NAND2_X1 U8690 ( .A1(n7000), .A2(n9697), .ZN(n7003) );
  NOR2_X1 U8691 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5143), .ZN(n7220) );
  NOR2_X1 U8692 ( .A1(n9964), .A2(n7041), .ZN(n7001) );
  AOI211_X1 U8693 ( .C1(n9960), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n7220), .B(
        n7001), .ZN(n7002) );
  OAI211_X1 U8694 ( .C1(n7004), .C2(n9699), .A(n7003), .B(n7002), .ZN(P2_U3258) );
  INV_X1 U8695 ( .A(n7005), .ZN(n7008) );
  OAI222_X1 U8696 ( .A1(n8117), .A2(n7008), .B1(P1_U3084), .B2(n7647), .C1(
        n7006), .C2(n9349), .ZN(P1_U3332) );
  OAI222_X1 U8697 ( .A1(n4267), .A2(n7009), .B1(n7519), .B2(n7008), .C1(n8099), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NAND2_X1 U8698 ( .A1(n7010), .A2(n7011), .ZN(n7013) );
  XNOR2_X1 U8699 ( .A(n7013), .B(n7012), .ZN(n7019) );
  INV_X1 U8700 ( .A(n7014), .ZN(n7093) );
  OAI22_X1 U8701 ( .A1(n7015), .A2(n8264), .B1(n7075), .B2(n8242), .ZN(n7085)
         );
  AOI22_X1 U8702 ( .A1(n8281), .A2(n7085), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7016) );
  OAI21_X1 U8703 ( .B1(n7093), .B2(n8285), .A(n7016), .ZN(n7017) );
  AOI21_X1 U8704 ( .B1(n7103), .B2(n4262), .A(n7017), .ZN(n7018) );
  OAI21_X1 U8705 ( .B1(n7019), .B2(n8289), .A(n7018), .ZN(P2_U3219) );
  INV_X1 U8706 ( .A(n7010), .ZN(n7021) );
  AOI21_X1 U8707 ( .B1(n7020), .B2(n7022), .A(n7021), .ZN(n7030) );
  INV_X1 U8708 ( .A(n7177), .ZN(n7027) );
  OR2_X1 U8709 ( .A1(n7033), .A2(n8242), .ZN(n7024) );
  NAND2_X1 U8710 ( .A1(n8309), .A2(n8228), .ZN(n7023) );
  NAND2_X1 U8711 ( .A1(n7024), .A2(n7023), .ZN(n7172) );
  NAND2_X1 U8712 ( .A1(n8281), .A2(n7172), .ZN(n7026) );
  OAI211_X1 U8713 ( .C1(n8285), .C2(n7027), .A(n7026), .B(n7025), .ZN(n7028)
         );
  AOI21_X1 U8714 ( .B1(n7360), .B2(n4262), .A(n7028), .ZN(n7029) );
  OAI21_X1 U8715 ( .B1(n7030), .B2(n8289), .A(n7029), .ZN(P2_U3233) );
  XNOR2_X1 U8716 ( .A(n7031), .B(n7032), .ZN(n7039) );
  NAND2_X1 U8717 ( .A1(n8271), .A2(n7155), .ZN(n7036) );
  OR2_X1 U8718 ( .A1(n7033), .A2(n8264), .ZN(n7034) );
  OAI21_X1 U8719 ( .B1(n7218), .B2(n8242), .A(n7034), .ZN(n7161) );
  NAND2_X1 U8720 ( .A1(n8281), .A2(n7161), .ZN(n7035) );
  OAI211_X1 U8721 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5117), .A(n7036), .B(n7035), .ZN(n7037) );
  AOI21_X1 U8722 ( .B1(n8669), .B2(n4262), .A(n7037), .ZN(n7038) );
  OAI21_X1 U8723 ( .B1(n7039), .B2(n8289), .A(n7038), .ZN(P2_U3238) );
  AOI21_X1 U8724 ( .B1(n7041), .B2(n6990), .A(n7040), .ZN(n7043) );
  INV_X1 U8725 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7450) );
  AOI22_X1 U8726 ( .A1(n7258), .A2(n7450), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7262), .ZN(n7042) );
  NOR2_X1 U8727 ( .A1(n7043), .A2(n7042), .ZN(n7261) );
  AOI21_X1 U8728 ( .B1(n7043), .B2(n7042), .A(n7261), .ZN(n7054) );
  INV_X1 U8729 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7044) );
  AOI22_X1 U8730 ( .A1(n7258), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7044), .B2(
        n7262), .ZN(n7048) );
  OAI21_X1 U8731 ( .B1(n7046), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7045), .ZN(
        n7047) );
  NAND2_X1 U8732 ( .A1(n7048), .A2(n7047), .ZN(n7257) );
  OAI21_X1 U8733 ( .B1(n7048), .B2(n7047), .A(n7257), .ZN(n7049) );
  NAND2_X1 U8734 ( .A1(n7049), .A2(n9697), .ZN(n7053) );
  INV_X1 U8735 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7050) );
  NAND2_X1 U8736 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7417) );
  OAI21_X1 U8737 ( .B1(n8362), .B2(n7050), .A(n7417), .ZN(n7051) );
  AOI21_X1 U8738 ( .B1(n9359), .B2(n7258), .A(n7051), .ZN(n7052) );
  OAI211_X1 U8739 ( .C1(n7054), .C2(n9699), .A(n7053), .B(n7052), .ZN(P2_U3259) );
  INV_X1 U8740 ( .A(n7055), .ZN(n7057) );
  OAI222_X1 U8741 ( .A1(n9349), .A2(n9862), .B1(n8117), .B2(n7057), .C1(n7815), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  OAI222_X1 U8742 ( .A1(n4267), .A2(n7058), .B1(n7519), .B2(n7057), .C1(
        P2_U3152), .C2(n7056), .ZN(P2_U3336) );
  NAND2_X1 U8743 ( .A1(n9455), .A2(n7824), .ZN(n9657) );
  INV_X1 U8744 ( .A(n7059), .ZN(n7063) );
  XNOR2_X1 U8745 ( .A(n7061), .B(n7060), .ZN(n7062) );
  XNOR2_X1 U8746 ( .A(n7063), .B(n7062), .ZN(n7064) );
  NAND2_X1 U8747 ( .A1(n7064), .A2(n8806), .ZN(n7071) );
  AOI21_X1 U8748 ( .B1(n8848), .B2(n8881), .A(n7065), .ZN(n7068) );
  NAND2_X1 U8749 ( .A1(n8861), .A2(n7066), .ZN(n7067) );
  OAI211_X1 U8750 ( .C1(n7132), .C2(n8850), .A(n7068), .B(n7067), .ZN(n7069)
         );
  INV_X1 U8751 ( .A(n7069), .ZN(n7070) );
  OAI211_X1 U8752 ( .C1(n8851), .C2(n9657), .A(n7071), .B(n7070), .ZN(P1_U3237) );
  NAND2_X1 U8753 ( .A1(n7073), .A2(n7957), .ZN(n7074) );
  XNOR2_X1 U8754 ( .A(n7074), .B(n8083), .ZN(n7077) );
  OR2_X1 U8755 ( .A1(n7075), .A2(n8264), .ZN(n7076) );
  OAI21_X1 U8756 ( .B1(n7277), .B2(n8242), .A(n7076), .ZN(n7206) );
  AOI21_X1 U8757 ( .B1(n7077), .B2(n8585), .A(n7206), .ZN(n7308) );
  XNOR2_X1 U8758 ( .A(n7078), .B(n8083), .ZN(n7311) );
  NAND2_X1 U8759 ( .A1(n7311), .A2(n8582), .ZN(n7083) );
  INV_X1 U8760 ( .A(n4798), .ZN(n7079) );
  AOI211_X1 U8761 ( .C1(n7210), .C2(n7152), .A(n9752), .B(n7079), .ZN(n7310)
         );
  INV_X1 U8762 ( .A(n7210), .ZN(n7317) );
  AOI22_X1 U8763 ( .A1(n8462), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7205), .B2(
        n8566), .ZN(n7080) );
  OAI21_X1 U8764 ( .B1(n8556), .B2(n7317), .A(n7080), .ZN(n7081) );
  AOI21_X1 U8765 ( .B1(n7310), .B2(n8572), .A(n7081), .ZN(n7082) );
  OAI211_X1 U8766 ( .C1(n8462), .C2(n7308), .A(n7083), .B(n7082), .ZN(P2_U3284) );
  XOR2_X1 U8767 ( .A(n7084), .B(n8079), .Z(n7086) );
  AOI21_X1 U8768 ( .B1(n7086), .B2(n8585), .A(n7085), .ZN(n7105) );
  OR2_X1 U8769 ( .A1(n7169), .A2(n8077), .ZN(n7167) );
  AND2_X1 U8770 ( .A1(n7167), .A2(n7087), .ZN(n7090) );
  NAND2_X1 U8771 ( .A1(n7167), .A2(n7088), .ZN(n7089) );
  OAI21_X1 U8772 ( .B1(n7090), .B2(n8079), .A(n7089), .ZN(n7106) );
  INV_X1 U8773 ( .A(n7106), .ZN(n7098) );
  INV_X1 U8774 ( .A(n7091), .ZN(n7154) );
  AOI21_X1 U8775 ( .B1(n7174), .B2(n7103), .A(n9752), .ZN(n7092) );
  NAND2_X1 U8776 ( .A1(n7154), .A2(n7092), .ZN(n7104) );
  INV_X1 U8777 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7094) );
  OAI22_X1 U8778 ( .A1(n8567), .A2(n7094), .B1(n7093), .B2(n8587), .ZN(n7095)
         );
  AOI21_X1 U8779 ( .B1(n8581), .B2(n7103), .A(n7095), .ZN(n7096) );
  OAI21_X1 U8780 ( .B1(n7104), .B2(n8370), .A(n7096), .ZN(n7097) );
  AOI21_X1 U8781 ( .B1(n7098), .B2(n8582), .A(n7097), .ZN(n7099) );
  OAI21_X1 U8782 ( .B1(n8462), .B2(n7105), .A(n7099), .ZN(P2_U3286) );
  INV_X1 U8783 ( .A(n7146), .ZN(n7102) );
  AND2_X1 U8784 ( .A1(n7100), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7814) );
  AOI21_X1 U8785 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n7485), .A(n7814), .ZN(
        n7101) );
  OAI21_X1 U8786 ( .B1(n7102), .B2(n8117), .A(n7101), .ZN(P1_U3330) );
  INV_X1 U8787 ( .A(n7103), .ZN(n7113) );
  OAI211_X1 U8788 ( .C1(n7106), .C2(n8674), .A(n7105), .B(n7104), .ZN(n7107)
         );
  INV_X1 U8789 ( .A(n7107), .ZN(n7110) );
  MUX2_X1 U8790 ( .A(n7108), .B(n7110), .S(n8676), .Z(n7109) );
  OAI21_X1 U8791 ( .B1(n7113), .B2(n8667), .A(n7109), .ZN(P2_U3530) );
  INV_X1 U8792 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7111) );
  MUX2_X1 U8793 ( .A(n7111), .B(n7110), .S(n9759), .Z(n7112) );
  OAI21_X1 U8794 ( .B1(n7113), .B2(n8711), .A(n7112), .ZN(P2_U3481) );
  NAND2_X1 U8795 ( .A1(n7132), .A2(n7114), .ZN(n7115) );
  NAND2_X1 U8796 ( .A1(n7231), .A2(n7287), .ZN(n7668) );
  INV_X1 U8797 ( .A(n7287), .ZN(n7373) );
  NAND2_X1 U8798 ( .A1(n7373), .A2(n8878), .ZN(n7184) );
  NAND2_X1 U8799 ( .A1(n7287), .A2(n8878), .ZN(n7118) );
  INV_X1 U8800 ( .A(n8877), .ZN(n7133) );
  OR2_X1 U8801 ( .A1(n7344), .A2(n7133), .ZN(n7670) );
  NAND2_X1 U8802 ( .A1(n7344), .A2(n7133), .ZN(n7669) );
  NAND2_X1 U8803 ( .A1(n7670), .A2(n7669), .ZN(n7632) );
  XOR2_X1 U8804 ( .A(n7325), .B(n7632), .Z(n9682) );
  INV_X1 U8805 ( .A(n7668), .ZN(n7678) );
  NAND2_X1 U8806 ( .A1(n7185), .A2(n7184), .ZN(n7120) );
  XNOR2_X1 U8807 ( .A(n7120), .B(n7632), .ZN(n7122) );
  OAI22_X1 U8808 ( .A1(n9437), .A2(n9434), .B1(n7231), .B2(n9435), .ZN(n7121)
         );
  AOI21_X1 U8809 ( .B1(n7122), .B2(n9414), .A(n7121), .ZN(n9677) );
  NOR2_X1 U8810 ( .A1(n9677), .A2(n9451), .ZN(n7129) );
  AND2_X1 U8811 ( .A1(n7140), .A2(n7344), .ZN(n7123) );
  OR2_X1 U8812 ( .A1(n7123), .A2(n7192), .ZN(n9678) );
  INV_X1 U8813 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7125) );
  INV_X1 U8814 ( .A(n7354), .ZN(n7124) );
  OAI22_X1 U8815 ( .A1(n9424), .A2(n7125), .B1(n7124), .B2(n9419), .ZN(n7126)
         );
  AOI21_X1 U8816 ( .B1(n9441), .B2(n7344), .A(n7126), .ZN(n7127) );
  OAI21_X1 U8817 ( .B1(n9678), .B2(n9200), .A(n7127), .ZN(n7128) );
  AOI211_X1 U8818 ( .C1(n9682), .C2(n7853), .A(n7129), .B(n7128), .ZN(n7130)
         );
  INV_X1 U8819 ( .A(n7130), .ZN(P1_U3282) );
  XNOR2_X1 U8820 ( .A(n7131), .B(n7631), .ZN(n7139) );
  OAI22_X1 U8821 ( .A1(n9437), .A2(n7133), .B1(n7132), .B2(n9435), .ZN(n7138)
         );
  NAND2_X1 U8822 ( .A1(n7135), .A2(n7631), .ZN(n7136) );
  NAND2_X1 U8823 ( .A1(n7134), .A2(n7136), .ZN(n7291) );
  NOR2_X1 U8824 ( .A1(n7291), .A2(n9664), .ZN(n7137) );
  AOI211_X1 U8825 ( .C1(n7139), .C2(n9414), .A(n7138), .B(n7137), .ZN(n7290)
         );
  AOI21_X1 U8826 ( .B1(n7287), .B2(n7141), .A(n4548), .ZN(n7288) );
  AOI22_X1 U8827 ( .A1(n9451), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7375), .B2(
        n9439), .ZN(n7142) );
  OAI21_X1 U8828 ( .B1(n7373), .B2(n9418), .A(n7142), .ZN(n7144) );
  NOR2_X1 U8829 ( .A1(n7291), .A2(n9233), .ZN(n7143) );
  AOI211_X1 U8830 ( .C1(n7288), .C2(n9446), .A(n7144), .B(n7143), .ZN(n7145)
         );
  OAI21_X1 U8831 ( .B1(n7290), .B2(n9451), .A(n7145), .ZN(P1_U3283) );
  NAND2_X1 U8832 ( .A1(n7146), .A2(n8721), .ZN(n7147) );
  OAI211_X1 U8833 ( .C1(n7148), .C2(n4267), .A(n7147), .B(n8111), .ZN(P2_U3335) );
  AND2_X1 U8834 ( .A1(n7150), .A2(n7149), .ZN(n7151) );
  XNOR2_X1 U8835 ( .A(n7151), .B(n7159), .ZN(n8675) );
  INV_X1 U8836 ( .A(n7152), .ZN(n7153) );
  AOI21_X1 U8837 ( .B1(n8669), .B2(n7154), .A(n7153), .ZN(n8671) );
  AOI22_X1 U8838 ( .A1(n8462), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7155), .B2(
        n8566), .ZN(n7156) );
  OAI21_X1 U8839 ( .B1(n8556), .B2(n7157), .A(n7156), .ZN(n7164) );
  NAND3_X1 U8840 ( .A1(n7158), .A2(n7159), .A3(n7962), .ZN(n7160) );
  AOI21_X1 U8841 ( .B1(n7073), .B2(n7160), .A(n8531), .ZN(n7162) );
  NOR2_X1 U8842 ( .A1(n7162), .A2(n7161), .ZN(n8673) );
  NOR2_X1 U8843 ( .A1(n8673), .A2(n8462), .ZN(n7163) );
  AOI211_X1 U8844 ( .C1(n8671), .C2(n8593), .A(n7164), .B(n7163), .ZN(n7165)
         );
  OAI21_X1 U8845 ( .B1(n8559), .B2(n8675), .A(n7165), .ZN(P2_U3285) );
  XNOR2_X1 U8846 ( .A(n7166), .B(n8077), .ZN(n7173) );
  INV_X1 U8847 ( .A(n7167), .ZN(n7168) );
  AOI21_X1 U8848 ( .B1(n8077), .B2(n7169), .A(n7168), .ZN(n7364) );
  NOR2_X1 U8849 ( .A1(n7364), .A2(n7170), .ZN(n7171) );
  AOI211_X1 U8850 ( .C1(n7173), .C2(n8585), .A(n7172), .B(n7171), .ZN(n7363)
         );
  INV_X1 U8851 ( .A(n7174), .ZN(n7175) );
  AOI21_X1 U8852 ( .B1(n7360), .B2(n7176), .A(n7175), .ZN(n7361) );
  INV_X1 U8853 ( .A(n7360), .ZN(n7179) );
  AOI22_X1 U8854 ( .A1(n8462), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7177), .B2(
        n8566), .ZN(n7178) );
  OAI21_X1 U8855 ( .B1(n8556), .B2(n7179), .A(n7178), .ZN(n7182) );
  NOR2_X1 U8856 ( .A1(n7364), .A2(n7180), .ZN(n7181) );
  AOI211_X1 U8857 ( .C1(n7361), .C2(n8593), .A(n7182), .B(n7181), .ZN(n7183)
         );
  OAI21_X1 U8858 ( .B1(n7363), .B2(n8462), .A(n7183), .ZN(P2_U3287) );
  AND2_X1 U8859 ( .A1(n7670), .A2(n7184), .ZN(n7677) );
  NAND2_X1 U8860 ( .A1(n7185), .A2(n7677), .ZN(n7319) );
  NAND2_X1 U8861 ( .A1(n7319), .A2(n7669), .ZN(n7186) );
  OR2_X1 U8862 ( .A1(n7322), .A2(n9434), .ZN(n7681) );
  NAND2_X1 U8863 ( .A1(n7322), .A2(n9434), .ZN(n7674) );
  XNOR2_X1 U8864 ( .A(n7186), .B(n7637), .ZN(n7187) );
  AOI222_X1 U8865 ( .A1(n9414), .A2(n7187), .B1(n8875), .B2(n9188), .C1(n8877), 
        .C2(n9136), .ZN(n9367) );
  OR2_X1 U8866 ( .A1(n7344), .A2(n8877), .ZN(n7323) );
  NAND2_X1 U8867 ( .A1(n7325), .A2(n7323), .ZN(n7188) );
  NAND2_X1 U8868 ( .A1(n7344), .A2(n8877), .ZN(n7328) );
  AND2_X1 U8869 ( .A1(n7188), .A2(n7328), .ZN(n7190) );
  INV_X1 U8870 ( .A(n7637), .ZN(n7327) );
  NAND2_X1 U8871 ( .A1(n7190), .A2(n7327), .ZN(n7189) );
  OAI21_X1 U8872 ( .B1(n7190), .B2(n7327), .A(n7189), .ZN(n9370) );
  NAND2_X1 U8873 ( .A1(n9370), .A2(n7853), .ZN(n7197) );
  INV_X1 U8874 ( .A(n7322), .ZN(n9368) );
  INV_X1 U8875 ( .A(n9444), .ZN(n7191) );
  OAI211_X1 U8876 ( .C1(n9368), .C2(n7192), .A(n7191), .B(n9661), .ZN(n9366)
         );
  INV_X1 U8877 ( .A(n9366), .ZN(n7195) );
  AOI22_X1 U8878 ( .A1(n9451), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7301), .B2(
        n9439), .ZN(n7193) );
  OAI21_X1 U8879 ( .B1(n9368), .B2(n9418), .A(n7193), .ZN(n7194) );
  AOI21_X1 U8880 ( .B1(n7195), .B2(n9210), .A(n7194), .ZN(n7196) );
  OAI211_X1 U8881 ( .C1(n9451), .C2(n9367), .A(n7197), .B(n7196), .ZN(P1_U3281) );
  INV_X1 U8882 ( .A(n7198), .ZN(n7214) );
  OAI222_X1 U8883 ( .A1(n8117), .A2(n7214), .B1(P1_U3084), .B2(n7200), .C1(
        n7199), .C2(n9349), .ZN(P1_U3329) );
  INV_X1 U8884 ( .A(n7202), .ZN(n7203) );
  AOI21_X1 U8885 ( .B1(n7201), .B2(n7204), .A(n7203), .ZN(n7212) );
  INV_X1 U8886 ( .A(n7205), .ZN(n7208) );
  AOI22_X1 U8887 ( .A1(n8281), .A2(n7206), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n7207) );
  OAI21_X1 U8888 ( .B1(n7208), .B2(n8285), .A(n7207), .ZN(n7209) );
  AOI21_X1 U8889 ( .B1(n7210), .B2(n4262), .A(n7209), .ZN(n7211) );
  OAI21_X1 U8890 ( .B1(n7212), .B2(n8289), .A(n7211), .ZN(P2_U3226) );
  OAI222_X1 U8891 ( .A1(n7215), .A2(P2_U3152), .B1(n7519), .B2(n7214), .C1(
        n7213), .C2(n4267), .ZN(P2_U3334) );
  XNOR2_X1 U8892 ( .A(n7217), .B(n7216), .ZN(n7225) );
  INV_X1 U8893 ( .A(n7251), .ZN(n7222) );
  OR2_X1 U8894 ( .A1(n7218), .A2(n8264), .ZN(n7219) );
  OAI21_X1 U8895 ( .B1(n7388), .B2(n8242), .A(n7219), .ZN(n7245) );
  AOI21_X1 U8896 ( .B1(n8281), .B2(n7245), .A(n7220), .ZN(n7221) );
  OAI21_X1 U8897 ( .B1(n7222), .B2(n8285), .A(n7221), .ZN(n7223) );
  AOI21_X1 U8898 ( .B1(n7250), .B2(n4262), .A(n7223), .ZN(n7224) );
  OAI21_X1 U8899 ( .B1(n7225), .B2(n8289), .A(n7224), .ZN(P2_U3236) );
  AND2_X1 U8900 ( .A1(n9455), .A2(n7226), .ZN(n9669) );
  AOI21_X1 U8901 ( .B1(n8848), .B2(n8880), .A(n7227), .ZN(n7230) );
  NAND2_X1 U8902 ( .A1(n8861), .A2(n7228), .ZN(n7229) );
  OAI211_X1 U8903 ( .C1(n7231), .C2(n8850), .A(n7230), .B(n7229), .ZN(n7239)
         );
  INV_X1 U8904 ( .A(n7232), .ZN(n7237) );
  AOI21_X1 U8905 ( .B1(n7236), .B2(n7234), .A(n7233), .ZN(n7235) );
  AOI211_X1 U8906 ( .C1(n7237), .C2(n7236), .A(n8868), .B(n7235), .ZN(n7238)
         );
  AOI211_X1 U8907 ( .C1(n7240), .C2(n9669), .A(n7239), .B(n7238), .ZN(n7241)
         );
  INV_X1 U8908 ( .A(n7241), .ZN(P1_U3211) );
  NAND2_X1 U8909 ( .A1(n7243), .A2(n4458), .ZN(n7244) );
  AOI21_X1 U8910 ( .B1(n7274), .B2(n7244), .A(n8531), .ZN(n7246) );
  OR2_X1 U8911 ( .A1(n7246), .A2(n7245), .ZN(n7405) );
  INV_X1 U8912 ( .A(n7405), .ZN(n7256) );
  INV_X1 U8913 ( .A(n7247), .ZN(n7248) );
  AOI21_X1 U8914 ( .B1(n8084), .B2(n7249), .A(n7248), .ZN(n7407) );
  NAND2_X1 U8915 ( .A1(n7407), .A2(n8582), .ZN(n7255) );
  AOI211_X1 U8916 ( .C1(n7250), .C2(n4798), .A(n9752), .B(n7280), .ZN(n7406)
         );
  INV_X1 U8917 ( .A(n7250), .ZN(n7412) );
  AOI22_X1 U8918 ( .A1(n8462), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7251), .B2(
        n8566), .ZN(n7252) );
  OAI21_X1 U8919 ( .B1(n7412), .B2(n8556), .A(n7252), .ZN(n7253) );
  AOI21_X1 U8920 ( .B1(n7406), .B2(n8572), .A(n7253), .ZN(n7254) );
  OAI211_X1 U8921 ( .C1(n8462), .C2(n7256), .A(n7255), .B(n7254), .ZN(P2_U3283) );
  OAI21_X1 U8922 ( .B1(n7258), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7257), .ZN(
        n7435) );
  XNOR2_X1 U8923 ( .A(n7435), .B(n7425), .ZN(n7260) );
  INV_X1 U8924 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7259) );
  OAI21_X1 U8925 ( .B1(n7260), .B2(n7259), .A(n7437), .ZN(n7268) );
  AOI21_X1 U8926 ( .B1(n7262), .B2(n7450), .A(n7261), .ZN(n7424) );
  XNOR2_X1 U8927 ( .A(n7424), .B(n7436), .ZN(n7263) );
  NAND2_X1 U8928 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7263), .ZN(n7426) );
  OAI211_X1 U8929 ( .C1(n7263), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9956), .B(
        n7426), .ZN(n7266) );
  NAND2_X1 U8930 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8282) );
  INV_X1 U8931 ( .A(n8282), .ZN(n7264) );
  AOI21_X1 U8932 ( .B1(n9960), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7264), .ZN(
        n7265) );
  OAI211_X1 U8933 ( .C1(n9964), .C2(n7436), .A(n7266), .B(n7265), .ZN(n7267)
         );
  AOI21_X1 U8934 ( .B1(n9697), .B2(n7268), .A(n7267), .ZN(n7269) );
  INV_X1 U8935 ( .A(n7269), .ZN(P2_U3260) );
  XNOR2_X1 U8936 ( .A(n7270), .B(n7272), .ZN(n7446) );
  INV_X1 U8937 ( .A(n7446), .ZN(n7286) );
  INV_X1 U8938 ( .A(n7271), .ZN(n7276) );
  AOI21_X1 U8939 ( .B1(n7274), .B2(n7273), .A(n7272), .ZN(n7275) );
  NOR3_X1 U8940 ( .A1(n7276), .A2(n7275), .A3(n8531), .ZN(n7279) );
  OR2_X1 U8941 ( .A1(n7277), .A2(n8264), .ZN(n7278) );
  OAI21_X1 U8942 ( .B1(n7466), .B2(n8242), .A(n7278), .ZN(n7416) );
  OR2_X1 U8943 ( .A1(n7279), .A2(n7416), .ZN(n7444) );
  INV_X1 U8944 ( .A(n7280), .ZN(n7281) );
  AOI211_X1 U8945 ( .C1(n7421), .C2(n7281), .A(n9752), .B(n7391), .ZN(n7445)
         );
  NAND2_X1 U8946 ( .A1(n7445), .A2(n8572), .ZN(n7283) );
  AOI22_X1 U8947 ( .A1(n8462), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7415), .B2(
        n8566), .ZN(n7282) );
  OAI211_X1 U8948 ( .C1(n7452), .C2(n8556), .A(n7283), .B(n7282), .ZN(n7284)
         );
  AOI21_X1 U8949 ( .B1(n7444), .B2(n8567), .A(n7284), .ZN(n7285) );
  OAI21_X1 U8950 ( .B1(n7286), .B2(n8559), .A(n7285), .ZN(P2_U3282) );
  AOI22_X1 U8951 ( .A1(n7288), .A2(n9661), .B1(n9455), .B2(n7287), .ZN(n7289)
         );
  OAI211_X1 U8952 ( .C1(n9456), .C2(n7291), .A(n7290), .B(n7289), .ZN(n7293)
         );
  NAND2_X1 U8953 ( .A1(n7293), .A2(n9696), .ZN(n7292) );
  OAI21_X1 U8954 ( .B1(n9696), .B2(n6205), .A(n7292), .ZN(P1_U3531) );
  INV_X1 U8955 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7295) );
  NAND2_X1 U8956 ( .A1(n7293), .A2(n9685), .ZN(n7294) );
  OAI21_X1 U8957 ( .B1(n9685), .B2(n7295), .A(n7294), .ZN(P1_U3478) );
  XNOR2_X1 U8958 ( .A(n7297), .B(n7296), .ZN(n7298) );
  XNOR2_X1 U8959 ( .A(n7299), .B(n7298), .ZN(n7306) );
  NOR2_X1 U8960 ( .A1(n9368), .A2(n8813), .ZN(n7305) );
  AOI21_X1 U8961 ( .B1(n8848), .B2(n8877), .A(n7300), .ZN(n7303) );
  NAND2_X1 U8962 ( .A1(n8861), .A2(n7301), .ZN(n7302) );
  OAI211_X1 U8963 ( .C1(n7320), .C2(n8850), .A(n7303), .B(n7302), .ZN(n7304)
         );
  AOI211_X1 U8964 ( .C1(n7306), .C2(n8806), .A(n7305), .B(n7304), .ZN(n7307)
         );
  INV_X1 U8965 ( .A(n7307), .ZN(P1_U3215) );
  INV_X1 U8966 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7312) );
  INV_X1 U8967 ( .A(n7308), .ZN(n7309) );
  AOI211_X1 U8968 ( .C1(n7311), .C2(n9746), .A(n7310), .B(n7309), .ZN(n7314)
         );
  MUX2_X1 U8969 ( .A(n7312), .B(n7314), .S(n9759), .Z(n7313) );
  OAI21_X1 U8970 ( .B1(n7317), .B2(n8711), .A(n7313), .ZN(P2_U3487) );
  MUX2_X1 U8971 ( .A(n7315), .B(n7314), .S(n9770), .Z(n7316) );
  OAI21_X1 U8972 ( .B1(n7317), .B2(n8667), .A(n7316), .ZN(P2_U3532) );
  NAND2_X1 U8973 ( .A1(n8771), .A2(n9436), .ZN(n7687) );
  INV_X1 U8974 ( .A(n7681), .ZN(n7318) );
  NAND2_X1 U8975 ( .A1(n7674), .A2(n7669), .ZN(n7679) );
  NAND2_X1 U8976 ( .A1(n7679), .A2(n7681), .ZN(n7575) );
  AND2_X1 U8977 ( .A1(n9442), .A2(n7320), .ZN(n7574) );
  OR2_X1 U8978 ( .A1(n9442), .A2(n7320), .ZN(n7590) );
  XOR2_X1 U8979 ( .A(n7638), .B(n7456), .Z(n7321) );
  AOI222_X1 U8980 ( .A1(n9414), .A2(n7321), .B1(n8873), .B2(n9188), .C1(n8875), 
        .C2(n9136), .ZN(n9464) );
  OR2_X1 U8981 ( .A1(n7322), .A2(n8876), .ZN(n7326) );
  AND2_X1 U8982 ( .A1(n7323), .A2(n7326), .ZN(n7324) );
  NAND2_X1 U8983 ( .A1(n7325), .A2(n7324), .ZN(n9428) );
  NAND2_X1 U8984 ( .A1(n9442), .A2(n8875), .ZN(n7634) );
  INV_X1 U8985 ( .A(n7326), .ZN(n7330) );
  AND2_X1 U8986 ( .A1(n7328), .A2(n7327), .ZN(n7329) );
  AND2_X1 U8987 ( .A1(n7634), .A2(n9427), .ZN(n7331) );
  NAND2_X1 U8988 ( .A1(n9428), .A2(n7331), .ZN(n7334) );
  OR2_X1 U8989 ( .A1(n9442), .A2(n8875), .ZN(n7635) );
  NAND2_X1 U8990 ( .A1(n7334), .A2(n7635), .ZN(n7336) );
  INV_X1 U8991 ( .A(n7638), .ZN(n7332) );
  AND2_X1 U8992 ( .A1(n7332), .A2(n7635), .ZN(n7333) );
  NAND2_X1 U8993 ( .A1(n7334), .A2(n7333), .ZN(n7454) );
  INV_X1 U8994 ( .A(n7454), .ZN(n7335) );
  AOI21_X1 U8995 ( .B1(n7638), .B2(n7336), .A(n7335), .ZN(n9467) );
  NAND2_X1 U8996 ( .A1(n9467), .A2(n7853), .ZN(n7343) );
  INV_X1 U8997 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7338) );
  OAI22_X1 U8998 ( .A1(n9424), .A2(n7338), .B1(n7337), .B2(n9419), .ZN(n7341)
         );
  INV_X1 U8999 ( .A(n8771), .ZN(n9465) );
  OAI211_X1 U9000 ( .C1(n4549), .C2(n9465), .A(n9661), .B(n9405), .ZN(n9463)
         );
  NOR2_X1 U9001 ( .A1(n9463), .A2(n7339), .ZN(n7340) );
  AOI211_X1 U9002 ( .C1(n9441), .C2(n8771), .A(n7341), .B(n7340), .ZN(n7342)
         );
  OAI211_X1 U9003 ( .C1(n9451), .C2(n9464), .A(n7343), .B(n7342), .ZN(P1_U3279) );
  NAND2_X1 U9004 ( .A1(n7344), .A2(n9455), .ZN(n9676) );
  NOR2_X1 U9005 ( .A1(n7346), .A2(n7345), .ZN(n7368) );
  NAND2_X1 U9006 ( .A1(n7346), .A2(n7345), .ZN(n7369) );
  OAI21_X1 U9007 ( .B1(n7368), .B2(n7347), .A(n7369), .ZN(n7351) );
  XNOR2_X1 U9008 ( .A(n7349), .B(n7348), .ZN(n7350) );
  XNOR2_X1 U9009 ( .A(n7351), .B(n7350), .ZN(n7352) );
  NAND2_X1 U9010 ( .A1(n7352), .A2(n8806), .ZN(n7359) );
  AOI21_X1 U9011 ( .B1(n8848), .B2(n8878), .A(n7353), .ZN(n7356) );
  NAND2_X1 U9012 ( .A1(n8861), .A2(n7354), .ZN(n7355) );
  OAI211_X1 U9013 ( .C1(n9434), .C2(n8850), .A(n7356), .B(n7355), .ZN(n7357)
         );
  INV_X1 U9014 ( .A(n7357), .ZN(n7358) );
  OAI211_X1 U9015 ( .C1(n8851), .C2(n9676), .A(n7359), .B(n7358), .ZN(P1_U3229) );
  AOI22_X1 U9016 ( .A1(n7361), .A2(n8670), .B1(n9722), .B2(n7360), .ZN(n7362)
         );
  OAI211_X1 U9017 ( .C1(n7364), .C2(n9748), .A(n7363), .B(n7362), .ZN(n7366)
         );
  NAND2_X1 U9018 ( .A1(n7366), .A2(n8676), .ZN(n7365) );
  OAI21_X1 U9019 ( .B1(n8676), .B2(n6463), .A(n7365), .ZN(P2_U3529) );
  INV_X1 U9020 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U9021 ( .A1(n7366), .A2(n9759), .ZN(n7367) );
  OAI21_X1 U9022 ( .B1(n9759), .B2(n9848), .A(n7367), .ZN(P2_U3478) );
  INV_X1 U9023 ( .A(n7368), .ZN(n7370) );
  NAND2_X1 U9024 ( .A1(n7370), .A2(n7369), .ZN(n7372) );
  XNOR2_X1 U9025 ( .A(n7372), .B(n7371), .ZN(n7381) );
  NOR2_X1 U9026 ( .A1(n8813), .A2(n7373), .ZN(n7380) );
  INV_X1 U9027 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7374) );
  NOR2_X1 U9028 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7374), .ZN(n8891) );
  AOI21_X1 U9029 ( .B1(n8860), .B2(n8877), .A(n8891), .ZN(n7378) );
  NAND2_X1 U9030 ( .A1(n8861), .A2(n7375), .ZN(n7377) );
  NAND2_X1 U9031 ( .A1(n8848), .A2(n8879), .ZN(n7376) );
  NAND3_X1 U9032 ( .A1(n7378), .A2(n7377), .A3(n7376), .ZN(n7379) );
  AOI211_X1 U9033 ( .C1(n7381), .C2(n8806), .A(n7380), .B(n7379), .ZN(n7382)
         );
  INV_X1 U9034 ( .A(n7382), .ZN(P1_U3219) );
  OAI21_X1 U9035 ( .B1(n7384), .B2(n8086), .A(n7383), .ZN(n7489) );
  INV_X1 U9036 ( .A(n7489), .ZN(n7398) );
  OAI211_X1 U9037 ( .C1(n7386), .C2(n7978), .A(n7385), .B(n8585), .ZN(n7390)
         );
  OR2_X1 U9038 ( .A1(n8206), .A2(n8242), .ZN(n7387) );
  OAI21_X1 U9039 ( .B1(n7388), .B2(n8264), .A(n7387), .ZN(n8280) );
  INV_X1 U9040 ( .A(n8280), .ZN(n7389) );
  NAND2_X1 U9041 ( .A1(n7390), .A2(n7389), .ZN(n7487) );
  INV_X1 U9042 ( .A(n7391), .ZN(n7393) );
  INV_X1 U9043 ( .A(n7472), .ZN(n7392) );
  AOI211_X1 U9044 ( .C1(n8287), .C2(n7393), .A(n9752), .B(n7392), .ZN(n7488)
         );
  NAND2_X1 U9045 ( .A1(n7488), .A2(n8572), .ZN(n7395) );
  AOI22_X1 U9046 ( .A1(n8462), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8279), .B2(
        n8566), .ZN(n7394) );
  OAI211_X1 U9047 ( .C1(n7495), .C2(n8556), .A(n7395), .B(n7394), .ZN(n7396)
         );
  AOI21_X1 U9048 ( .B1(n7487), .B2(n8567), .A(n7396), .ZN(n7397) );
  OAI21_X1 U9049 ( .B1(n7398), .B2(n8559), .A(n7397), .ZN(P2_U3281) );
  INV_X1 U9050 ( .A(n7399), .ZN(n7403) );
  OAI222_X1 U9051 ( .A1(n4267), .A2(n7401), .B1(n7519), .B2(n7403), .C1(n7400), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9052 ( .A1(n9349), .A2(n7404), .B1(n8117), .B2(n7403), .C1(n7402), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9053 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7408) );
  AOI211_X1 U9054 ( .C1(n7407), .C2(n9746), .A(n7406), .B(n7405), .ZN(n7410)
         );
  MUX2_X1 U9055 ( .A(n7408), .B(n7410), .S(n9759), .Z(n7409) );
  OAI21_X1 U9056 ( .B1(n7412), .B2(n8711), .A(n7409), .ZN(P2_U3490) );
  MUX2_X1 U9057 ( .A(n6990), .B(n7410), .S(n9770), .Z(n7411) );
  OAI21_X1 U9058 ( .B1(n7412), .B2(n8667), .A(n7411), .ZN(P2_U3533) );
  AOI21_X1 U9059 ( .B1(n7414), .B2(n7413), .A(n4335), .ZN(n7423) );
  INV_X1 U9060 ( .A(n7415), .ZN(n7419) );
  NAND2_X1 U9061 ( .A1(n8281), .A2(n7416), .ZN(n7418) );
  OAI211_X1 U9062 ( .C1(n8285), .C2(n7419), .A(n7418), .B(n7417), .ZN(n7420)
         );
  AOI21_X1 U9063 ( .B1(n7421), .B2(n4262), .A(n7420), .ZN(n7422) );
  OAI21_X1 U9064 ( .B1(n7423), .B2(n8289), .A(n7422), .ZN(P2_U3217) );
  NAND2_X1 U9065 ( .A1(n7425), .A2(n7424), .ZN(n7427) );
  NAND2_X1 U9066 ( .A1(n7427), .A2(n7426), .ZN(n7429) );
  XNOR2_X1 U9067 ( .A(n8322), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7428) );
  NOR2_X1 U9068 ( .A1(n7428), .A2(n7429), .ZN(n8323) );
  AOI21_X1 U9069 ( .B1(n7429), .B2(n7428), .A(n8323), .ZN(n7434) );
  NOR2_X1 U9070 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7430), .ZN(n7431) );
  AOI21_X1 U9071 ( .B1(n9960), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7431), .ZN(
        n7433) );
  NAND2_X1 U9072 ( .A1(n9359), .A2(n8322), .ZN(n7432) );
  OAI211_X1 U9073 ( .C1(n7434), .C2(n9699), .A(n7433), .B(n7432), .ZN(n7443)
         );
  NAND2_X1 U9074 ( .A1(n7436), .A2(n7435), .ZN(n7438) );
  NAND2_X1 U9075 ( .A1(n8322), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7439) );
  OAI21_X1 U9076 ( .B1(n8322), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7439), .ZN(
        n7440) );
  AOI211_X1 U9077 ( .C1(n7441), .C2(n7440), .A(n8318), .B(n9951), .ZN(n7442)
         );
  OR2_X1 U9078 ( .A1(n7443), .A2(n7442), .ZN(P2_U3261) );
  INV_X1 U9079 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7447) );
  AOI211_X1 U9080 ( .C1(n7446), .C2(n9746), .A(n7445), .B(n7444), .ZN(n7449)
         );
  MUX2_X1 U9081 ( .A(n7447), .B(n7449), .S(n9759), .Z(n7448) );
  OAI21_X1 U9082 ( .B1(n7452), .B2(n8711), .A(n7448), .ZN(P2_U3493) );
  MUX2_X1 U9083 ( .A(n7450), .B(n7449), .S(n9770), .Z(n7451) );
  OAI21_X1 U9084 ( .B1(n7452), .B2(n8667), .A(n7451), .ZN(P2_U3534) );
  INV_X1 U9085 ( .A(n9436), .ZN(n8874) );
  NAND2_X1 U9086 ( .A1(n8771), .A2(n8874), .ZN(n7453) );
  NAND2_X1 U9087 ( .A1(n7454), .A2(n7453), .ZN(n9403) );
  XNOR2_X1 U9088 ( .A(n9322), .B(n9412), .ZN(n7640) );
  XNOR2_X1 U9089 ( .A(n7503), .B(n7640), .ZN(n9325) );
  INV_X1 U9090 ( .A(n8871), .ZN(n8780) );
  INV_X1 U9091 ( .A(n7688), .ZN(n7455) );
  OR2_X1 U9092 ( .A1(n8822), .A2(n8769), .ZN(n7680) );
  NAND2_X1 U9093 ( .A1(n8822), .A2(n8769), .ZN(n7693) );
  NAND2_X1 U9094 ( .A1(n9409), .A2(n7693), .ZN(n7504) );
  XNOR2_X1 U9095 ( .A(n7504), .B(n7640), .ZN(n7457) );
  OAI222_X1 U9096 ( .A1(n9437), .A2(n8780), .B1(n9435), .B2(n8769), .C1(n9433), 
        .C2(n7457), .ZN(n9320) );
  AOI211_X1 U9097 ( .C1(n9322), .C2(n9406), .A(n9679), .B(n9226), .ZN(n9321)
         );
  NAND2_X1 U9098 ( .A1(n9321), .A2(n9210), .ZN(n7459) );
  AOI22_X1 U9099 ( .A1(n9451), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8729), .B2(
        n9439), .ZN(n7458) );
  OAI211_X1 U9100 ( .C1(n7460), .C2(n9418), .A(n7459), .B(n7458), .ZN(n7461)
         );
  AOI21_X1 U9101 ( .B1(n9320), .B2(n9424), .A(n7461), .ZN(n7462) );
  OAI21_X1 U9102 ( .B1(n9325), .B2(n9217), .A(n7462), .ZN(P1_U3277) );
  NAND2_X1 U9103 ( .A1(n7463), .A2(n8087), .ZN(n7464) );
  NAND2_X1 U9104 ( .A1(n7465), .A2(n7464), .ZN(n7468) );
  OR2_X1 U9105 ( .A1(n7466), .A2(n8264), .ZN(n7467) );
  OAI21_X1 U9106 ( .B1(n8253), .B2(n8242), .A(n7467), .ZN(n8198) );
  AOI21_X1 U9107 ( .B1(n7468), .B2(n8585), .A(n8198), .ZN(n8662) );
  AND2_X1 U9108 ( .A1(n7469), .A2(n7983), .ZN(n7470) );
  NOR2_X1 U9109 ( .A1(n7471), .A2(n7470), .ZN(n8664) );
  NAND2_X1 U9110 ( .A1(n8664), .A2(n8582), .ZN(n7478) );
  AOI21_X1 U9111 ( .B1(n7472), .B2(n8715), .A(n9752), .ZN(n7473) );
  NAND2_X1 U9112 ( .A1(n7473), .A2(n8551), .ZN(n8661) );
  INV_X1 U9113 ( .A(n8661), .ZN(n7476) );
  INV_X1 U9114 ( .A(n8715), .ZN(n8668) );
  AOI22_X1 U9115 ( .A1(n8462), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8199), .B2(
        n8566), .ZN(n7474) );
  OAI21_X1 U9116 ( .B1(n8668), .B2(n8556), .A(n7474), .ZN(n7475) );
  AOI21_X1 U9117 ( .B1(n7476), .B2(n8572), .A(n7475), .ZN(n7477) );
  OAI211_X1 U9118 ( .C1(n8462), .C2(n8662), .A(n7478), .B(n7477), .ZN(P2_U3280) );
  INV_X1 U9119 ( .A(n7479), .ZN(n7482) );
  OAI222_X1 U9120 ( .A1(n4267), .A2(n9806), .B1(n7519), .B2(n7482), .C1(n7480), 
        .C2(P2_U3152), .ZN(P2_U3332) );
  OAI222_X1 U9121 ( .A1(n9349), .A2(n7483), .B1(n8117), .B2(n7482), .C1(n7481), 
        .C2(P1_U3084), .ZN(P1_U3327) );
  INV_X1 U9122 ( .A(n7560), .ZN(n7496) );
  AOI21_X1 U9123 ( .B1(n7485), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7484), .ZN(
        n7486) );
  OAI21_X1 U9124 ( .B1(n7496), .B2(n8117), .A(n7486), .ZN(P1_U3326) );
  INV_X1 U9125 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7490) );
  AOI211_X1 U9126 ( .C1(n7489), .C2(n9746), .A(n7488), .B(n7487), .ZN(n7492)
         );
  MUX2_X1 U9127 ( .A(n7490), .B(n7492), .S(n9759), .Z(n7491) );
  OAI21_X1 U9128 ( .B1(n7495), .B2(n8711), .A(n7491), .ZN(P2_U3496) );
  INV_X1 U9129 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7493) );
  MUX2_X1 U9130 ( .A(n7493), .B(n7492), .S(n9770), .Z(n7494) );
  OAI21_X1 U9131 ( .B1(n7495), .B2(n8667), .A(n7494), .ZN(P2_U3535) );
  OAI222_X1 U9132 ( .A1(n4267), .A2(n9869), .B1(n7519), .B2(n7496), .C1(
        P2_U3152), .C2(n5394), .ZN(P2_U3331) );
  NAND2_X1 U9133 ( .A1(n7555), .A2(n8721), .ZN(n7498) );
  OAI211_X1 U9134 ( .C1(n4267), .C2(n7499), .A(n7498), .B(n7497), .ZN(P2_U3330) );
  INV_X1 U9135 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7556) );
  NAND2_X1 U9136 ( .A1(n7555), .A2(n9344), .ZN(n7500) );
  OAI211_X1 U9137 ( .C1(n9349), .C2(n7556), .A(n7500), .B(n9484), .ZN(P1_U3325) );
  AND2_X1 U9138 ( .A1(n9322), .A2(n8872), .ZN(n7502) );
  OR2_X1 U9139 ( .A1(n9312), .A2(n9220), .ZN(n7706) );
  NAND2_X1 U9140 ( .A1(n9312), .A2(n9220), .ZN(n9179) );
  NAND2_X1 U9141 ( .A1(n7706), .A2(n9179), .ZN(n8956) );
  XNOR2_X1 U9142 ( .A(n8957), .B(n8956), .ZN(n9314) );
  OR2_X1 U9143 ( .A1(n9322), .A2(n9412), .ZN(n7700) );
  AND2_X1 U9144 ( .A1(n9232), .A2(n8871), .ZN(n7624) );
  NAND2_X1 U9145 ( .A1(n9315), .A2(n8780), .ZN(n8980) );
  NAND2_X1 U9146 ( .A1(n8981), .A2(n8980), .ZN(n9178) );
  XNOR2_X1 U9147 ( .A(n9178), .B(n8956), .ZN(n7505) );
  OAI222_X1 U9148 ( .A1(n9437), .A2(n9190), .B1(n9435), .B2(n8780), .C1(n7505), 
        .C2(n9433), .ZN(n9310) );
  INV_X1 U9149 ( .A(n9312), .ZN(n8785) );
  INV_X1 U9150 ( .A(n9209), .ZN(n7506) );
  AOI211_X1 U9151 ( .C1(n9312), .C2(n9227), .A(n9679), .B(n7506), .ZN(n9311)
         );
  NAND2_X1 U9152 ( .A1(n9311), .A2(n9210), .ZN(n7508) );
  AOI22_X1 U9153 ( .A1(n9451), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8782), .B2(
        n9439), .ZN(n7507) );
  OAI211_X1 U9154 ( .C1(n8785), .C2(n9418), .A(n7508), .B(n7507), .ZN(n7509)
         );
  AOI21_X1 U9155 ( .B1(n9310), .B2(n9424), .A(n7509), .ZN(n7510) );
  OAI21_X1 U9156 ( .B1(n9314), .B2(n9217), .A(n7510), .ZN(P1_U3275) );
  OAI222_X1 U9157 ( .A1(n4267), .A2(n7512), .B1(n7519), .B2(n7511), .C1(n5430), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  INV_X1 U9158 ( .A(SI_29_), .ZN(n7513) );
  AND2_X1 U9159 ( .A1(n7514), .A2(n7513), .ZN(n7517) );
  INV_X1 U9160 ( .A(n7514), .ZN(n7515) );
  NAND2_X1 U9161 ( .A1(n7515), .A2(SI_29_), .ZN(n7516) );
  MUX2_X1 U9162 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7538), .Z(n7534) );
  INV_X1 U9163 ( .A(n7891), .ZN(n8116) );
  INV_X1 U9164 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7892) );
  OAI222_X1 U9165 ( .A1(P2_U3152), .A2(n7520), .B1(n7519), .B2(n8116), .C1(
        n7892), .C2(n4267), .ZN(P2_U3328) );
  NOR2_X1 U9166 ( .A1(n7522), .A2(n7521), .ZN(n7525) );
  AOI21_X1 U9167 ( .B1(n7525), .B2(n7524), .A(n7523), .ZN(n7531) );
  NOR2_X1 U9168 ( .A1(n8813), .A2(n9639), .ZN(n7528) );
  OAI22_X1 U9169 ( .A1(n8864), .A2(n7526), .B1(n6777), .B2(n8850), .ZN(n7527)
         );
  AOI211_X1 U9170 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n7529), .A(n7528), .B(
        n7527), .ZN(n7530) );
  OAI21_X1 U9171 ( .B1(n7531), .B2(n8868), .A(n7530), .ZN(P1_U3235) );
  INV_X1 U9172 ( .A(n7532), .ZN(n7533) );
  NAND2_X1 U9173 ( .A1(n7533), .A2(SI_30_), .ZN(n7537) );
  NAND2_X1 U9174 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  NAND2_X1 U9175 ( .A1(n7537), .A2(n7536), .ZN(n7541) );
  MUX2_X1 U9176 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7538), .Z(n7539) );
  XNOR2_X1 U9177 ( .A(n7539), .B(SI_31_), .ZN(n7540) );
  NOR2_X1 U9178 ( .A1(n7562), .A2(n6266), .ZN(n7542) );
  INV_X1 U9179 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8118) );
  OR2_X1 U9180 ( .A1(n7562), .A2(n8118), .ZN(n7543) );
  NAND2_X1 U9181 ( .A1(n4266), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7546) );
  NAND2_X1 U9182 ( .A1(n5840), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7545) );
  NAND2_X1 U9183 ( .A1(n4273), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7544) );
  AND3_X1 U9184 ( .A1(n7546), .A2(n7545), .A3(n7544), .ZN(n9005) );
  OR2_X1 U9185 ( .A1(n8949), .A2(n7802), .ZN(n7547) );
  NAND2_X1 U9186 ( .A1(n9237), .A2(n8947), .ZN(n7806) );
  NAND2_X1 U9187 ( .A1(n7547), .A2(n7806), .ZN(n7758) );
  INV_X1 U9188 ( .A(n7758), .ZN(n7618) );
  NAND2_X1 U9189 ( .A1(n8113), .A2(n5779), .ZN(n7549) );
  OR2_X1 U9190 ( .A1(n7562), .A2(n9350), .ZN(n7548) );
  NAND2_X1 U9191 ( .A1(n5840), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7554) );
  NAND2_X1 U9192 ( .A1(n4266), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7553) );
  INV_X1 U9193 ( .A(n7550), .ZN(n9011) );
  NAND2_X1 U9194 ( .A1(n4271), .A2(n9011), .ZN(n7552) );
  NAND2_X1 U9195 ( .A1(n4273), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7551) );
  NAND4_X1 U9196 ( .A1(n7554), .A2(n7553), .A3(n7552), .A4(n7551), .ZN(n9027)
         );
  INV_X1 U9197 ( .A(n9027), .ZN(n7750) );
  OR2_X1 U9198 ( .A1(n9242), .A2(n7750), .ZN(n7559) );
  NAND2_X1 U9199 ( .A1(n7555), .A2(n5779), .ZN(n7558) );
  OR2_X1 U9200 ( .A1(n7562), .A2(n7556), .ZN(n7557) );
  NAND2_X1 U9201 ( .A1(n7559), .A2(n9001), .ZN(n7800) );
  NAND2_X1 U9202 ( .A1(n7560), .A2(n5779), .ZN(n7564) );
  OR2_X1 U9203 ( .A1(n7562), .A2(n7561), .ZN(n7563) );
  AND2_X1 U9204 ( .A1(n8997), .A2(n7728), .ZN(n7798) );
  OR2_X1 U9205 ( .A1(n9140), .A2(n9154), .ZN(n7721) );
  INV_X1 U9206 ( .A(n9137), .ZN(n9166) );
  AND2_X1 U9207 ( .A1(n9290), .A2(n9166), .ZN(n8987) );
  NAND2_X1 U9208 ( .A1(n7721), .A2(n8987), .ZN(n7565) );
  NAND2_X1 U9209 ( .A1(n9140), .A2(n9154), .ZN(n8989) );
  NAND2_X1 U9210 ( .A1(n7565), .A2(n8989), .ZN(n7566) );
  NOR2_X1 U9211 ( .A1(n8990), .A2(n7566), .ZN(n7722) );
  INV_X1 U9212 ( .A(n9187), .ZN(n9153) );
  NAND2_X1 U9213 ( .A1(n9295), .A2(n9153), .ZN(n8985) );
  NAND2_X1 U9214 ( .A1(n7567), .A2(n9208), .ZN(n8984) );
  AND2_X1 U9215 ( .A1(n8985), .A2(n8984), .ZN(n7713) );
  INV_X1 U9216 ( .A(n7713), .ZN(n7569) );
  INV_X1 U9217 ( .A(n9290), .ZN(n8961) );
  AND2_X1 U9218 ( .A1(n8961), .A2(n9137), .ZN(n9132) );
  OR2_X1 U9219 ( .A1(n9295), .A2(n9153), .ZN(n7709) );
  INV_X1 U9220 ( .A(n7709), .ZN(n7568) );
  NOR2_X1 U9221 ( .A1(n9132), .A2(n7568), .ZN(n7716) );
  OAI211_X1 U9222 ( .C1(n8982), .C2(n7569), .A(n7716), .B(n7721), .ZN(n7571)
         );
  INV_X1 U9223 ( .A(n8991), .ZN(n7570) );
  AOI21_X1 U9224 ( .B1(n7722), .B2(n7571), .A(n7570), .ZN(n7794) );
  NOR2_X1 U9225 ( .A1(n4503), .A2(n4636), .ZN(n7791) );
  AND2_X1 U9226 ( .A1(n9307), .A2(n9190), .ZN(n9181) );
  INV_X1 U9227 ( .A(n9181), .ZN(n8977) );
  AND2_X1 U9228 ( .A1(n8984), .A2(n8977), .ZN(n7656) );
  INV_X1 U9229 ( .A(n7656), .ZN(n7573) );
  INV_X1 U9230 ( .A(n9179), .ZN(n7572) );
  OR2_X1 U9231 ( .A1(n7573), .A2(n7572), .ZN(n7601) );
  NAND2_X1 U9232 ( .A1(n9322), .A2(n9412), .ZN(n7697) );
  AND2_X1 U9233 ( .A1(n7697), .A2(n7693), .ZN(n7597) );
  INV_X1 U9234 ( .A(n7574), .ZN(n7686) );
  NAND3_X1 U9235 ( .A1(n7687), .A2(n7686), .A3(n7575), .ZN(n7594) );
  NAND2_X1 U9236 ( .A1(n7668), .A2(n7661), .ZN(n7576) );
  NOR2_X1 U9237 ( .A1(n7594), .A2(n7576), .ZN(n7577) );
  NAND3_X1 U9238 ( .A1(n8980), .A2(n7597), .A3(n7577), .ZN(n7578) );
  OR2_X1 U9239 ( .A1(n7601), .A2(n7578), .ZN(n7789) );
  NAND2_X1 U9240 ( .A1(n7583), .A2(n7579), .ZN(n7580) );
  NOR2_X1 U9241 ( .A1(n7581), .A2(n7580), .ZN(n7782) );
  NAND2_X1 U9242 ( .A1(n7582), .A2(n7782), .ZN(n7589) );
  INV_X1 U9243 ( .A(n7583), .ZN(n7584) );
  OAI21_X1 U9244 ( .B1(n7584), .B2(n7780), .A(n7657), .ZN(n7586) );
  AOI21_X1 U9245 ( .B1(n7586), .B2(n7659), .A(n7585), .ZN(n7630) );
  INV_X1 U9246 ( .A(n7630), .ZN(n7587) );
  NAND2_X1 U9247 ( .A1(n7587), .A2(n7660), .ZN(n7588) );
  INV_X1 U9248 ( .A(n7664), .ZN(n7784) );
  AOI21_X1 U9249 ( .B1(n7589), .B2(n7588), .A(n7784), .ZN(n7602) );
  AND2_X1 U9250 ( .A1(n7681), .A2(n7677), .ZN(n7595) );
  NAND2_X1 U9251 ( .A1(n7688), .A2(n7590), .ZN(n7591) );
  NAND2_X1 U9252 ( .A1(n7591), .A2(n7687), .ZN(n7592) );
  NAND2_X1 U9253 ( .A1(n7680), .A2(n7592), .ZN(n7694) );
  INV_X1 U9254 ( .A(n7694), .ZN(n7593) );
  OAI21_X1 U9255 ( .B1(n7595), .B2(n7594), .A(n7593), .ZN(n7596) );
  AOI21_X1 U9256 ( .B1(n7597), .B2(n7596), .A(n4377), .ZN(n7598) );
  INV_X1 U9257 ( .A(n8980), .ZN(n7623) );
  INV_X1 U9258 ( .A(n7624), .ZN(n7703) );
  OAI211_X1 U9259 ( .C1(n7598), .C2(n7623), .A(n7706), .B(n7703), .ZN(n7599)
         );
  INV_X1 U9260 ( .A(n7599), .ZN(n7600) );
  OR2_X1 U9261 ( .A1(n7601), .A2(n7600), .ZN(n7787) );
  OAI21_X1 U9262 ( .B1(n7789), .B2(n7602), .A(n7787), .ZN(n7603) );
  NAND2_X1 U9263 ( .A1(n7791), .A2(n7603), .ZN(n7604) );
  NAND2_X1 U9264 ( .A1(n9273), .A2(n9089), .ZN(n7622) );
  INV_X1 U9265 ( .A(n7622), .ZN(n7650) );
  AOI21_X1 U9266 ( .B1(n7794), .B2(n7604), .A(n7650), .ZN(n7607) );
  INV_X1 U9267 ( .A(n9109), .ZN(n8969) );
  NAND2_X1 U9268 ( .A1(n8966), .A2(n8969), .ZN(n7792) );
  NAND2_X1 U9269 ( .A1(n9103), .A2(n9123), .ZN(n8992) );
  NAND2_X1 U9270 ( .A1(n7792), .A2(n8992), .ZN(n7606) );
  NAND2_X1 U9271 ( .A1(n9069), .A2(n9088), .ZN(n7731) );
  NAND2_X1 U9272 ( .A1(n8967), .A2(n9109), .ZN(n8995) );
  NAND2_X1 U9273 ( .A1(n7731), .A2(n8995), .ZN(n7652) );
  INV_X1 U9274 ( .A(n7652), .ZN(n7605) );
  OAI21_X1 U9275 ( .B1(n7607), .B2(n7606), .A(n7605), .ZN(n7608) );
  NAND3_X1 U9276 ( .A1(n8999), .A2(n7798), .A3(n7608), .ZN(n7616) );
  NAND2_X1 U9277 ( .A1(n4397), .A2(n7609), .ZN(n7610) );
  NAND2_X1 U9278 ( .A1(n9454), .A2(n7610), .ZN(n7759) );
  NAND2_X1 U9279 ( .A1(n9247), .A2(n9044), .ZN(n7742) );
  NAND2_X1 U9280 ( .A1(n9252), .A2(n9058), .ZN(n7738) );
  NAND2_X1 U9281 ( .A1(n9257), .A2(n9073), .ZN(n7621) );
  NAND2_X1 U9282 ( .A1(n7738), .A2(n7621), .ZN(n7611) );
  NAND2_X1 U9283 ( .A1(n7611), .A2(n8999), .ZN(n7612) );
  AND2_X1 U9284 ( .A1(n7742), .A2(n7612), .ZN(n7613) );
  OR2_X1 U9285 ( .A1(n7800), .A2(n7613), .ZN(n7615) );
  NAND2_X1 U9286 ( .A1(n9242), .A2(n7750), .ZN(n7614) );
  AND2_X1 U9287 ( .A1(n7615), .A2(n7614), .ZN(n7801) );
  OAI211_X1 U9288 ( .C1(n7800), .C2(n7616), .A(n7759), .B(n7801), .ZN(n7617)
         );
  NAND2_X1 U9289 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  AND2_X1 U9290 ( .A1(n7747), .A2(n6099), .ZN(n7767) );
  NAND2_X1 U9291 ( .A1(n7619), .A2(n7767), .ZN(n7649) );
  NAND2_X1 U9292 ( .A1(n9454), .A2(n9005), .ZN(n7620) );
  INV_X1 U9293 ( .A(n9025), .ZN(n7740) );
  INV_X1 U9294 ( .A(n9042), .ZN(n9033) );
  XNOR2_X1 U9295 ( .A(n8967), .B(n9109), .ZN(n9086) );
  INV_X1 U9296 ( .A(n8956), .ZN(n9177) );
  AND3_X1 U9297 ( .A1(n7627), .A2(n7626), .A3(n7625), .ZN(n7628) );
  NAND4_X1 U9298 ( .A1(n7630), .A2(n7782), .A3(n7629), .A4(n7628), .ZN(n7633)
         );
  NOR3_X1 U9299 ( .A1(n7633), .A2(n7632), .A3(n7117), .ZN(n7636) );
  NAND2_X1 U9300 ( .A1(n7635), .A2(n7634), .ZN(n9431) );
  NAND4_X1 U9301 ( .A1(n7638), .A2(n7637), .A3(n7636), .A4(n9431), .ZN(n7639)
         );
  NOR4_X1 U9302 ( .A1(n9218), .A2(n7640), .A3(n4355), .A4(n7639), .ZN(n7641)
         );
  AND4_X1 U9303 ( .A1(n9184), .A2(n9177), .A3(n9206), .A4(n7641), .ZN(n7642)
         );
  NAND2_X1 U9304 ( .A1(n9164), .A2(n7642), .ZN(n7643) );
  NOR3_X1 U9305 ( .A1(n9131), .A2(n9150), .A3(n7643), .ZN(n7644) );
  NAND3_X1 U9306 ( .A1(n9105), .A2(n9121), .A3(n7644), .ZN(n7645) );
  NOR4_X1 U9307 ( .A1(n9056), .A2(n9065), .A3(n9086), .A4(n7645), .ZN(n7646)
         );
  NAND4_X1 U9308 ( .A1(n4790), .A2(n7802), .A3(n7806), .A4(n4795), .ZN(n7648)
         );
  NAND2_X1 U9309 ( .A1(n7648), .A2(n7647), .ZN(n7764) );
  AND2_X1 U9310 ( .A1(n7649), .A2(n7764), .ZN(n7766) );
  AND2_X1 U9311 ( .A1(n7792), .A2(n7650), .ZN(n7651) );
  NOR2_X1 U9312 ( .A1(n7652), .A2(n7651), .ZN(n7796) );
  INV_X1 U9313 ( .A(n8995), .ZN(n7653) );
  OAI211_X1 U9314 ( .C1(n7653), .C2(n8992), .A(n7728), .B(n7792), .ZN(n7654)
         );
  INV_X1 U9315 ( .A(n7654), .ZN(n7655) );
  MUX2_X1 U9316 ( .A(n7796), .B(n7655), .S(n7752), .Z(n7727) );
  INV_X1 U9317 ( .A(n7752), .ZN(n7753) );
  MUX2_X1 U9318 ( .A(n8982), .B(n7656), .S(n7753), .Z(n7708) );
  INV_X1 U9319 ( .A(n7660), .ZN(n7663) );
  NAND2_X1 U9320 ( .A1(n7665), .A2(n7664), .ZN(n7667) );
  INV_X1 U9321 ( .A(n7667), .ZN(n7666) );
  INV_X1 U9322 ( .A(n7677), .ZN(n7673) );
  NAND2_X1 U9323 ( .A1(n7669), .A2(n7668), .ZN(n7671) );
  NAND2_X1 U9324 ( .A1(n7671), .A2(n7670), .ZN(n7672) );
  AND4_X1 U9325 ( .A1(n7687), .A2(n7674), .A3(n7752), .A4(n9431), .ZN(n7675)
         );
  NAND3_X1 U9326 ( .A1(n7697), .A2(n7675), .A3(n7693), .ZN(n7676) );
  INV_X1 U9327 ( .A(n7679), .ZN(n7684) );
  NAND2_X1 U9328 ( .A1(n7700), .A2(n7680), .ZN(n7685) );
  NAND4_X1 U9329 ( .A1(n7688), .A2(n7753), .A3(n7681), .A4(n9431), .ZN(n7682)
         );
  OR2_X1 U9330 ( .A1(n7685), .A2(n7682), .ZN(n7683) );
  INV_X1 U9331 ( .A(n7685), .ZN(n7692) );
  NAND2_X1 U9332 ( .A1(n7687), .A2(n7686), .ZN(n7689) );
  NAND2_X1 U9333 ( .A1(n7689), .A2(n7688), .ZN(n7690) );
  AOI21_X1 U9334 ( .B1(n7693), .B2(n7690), .A(n7752), .ZN(n7691) );
  NAND2_X1 U9335 ( .A1(n7692), .A2(n7691), .ZN(n7699) );
  NAND3_X1 U9336 ( .A1(n7694), .A2(n7693), .A3(n7752), .ZN(n7695) );
  NAND2_X1 U9337 ( .A1(n7695), .A2(n7697), .ZN(n7696) );
  OAI21_X1 U9338 ( .B1(n7753), .B2(n7697), .A(n7696), .ZN(n7698) );
  OAI211_X1 U9339 ( .C1(n7753), .C2(n7700), .A(n7699), .B(n7698), .ZN(n7701)
         );
  INV_X1 U9340 ( .A(n9218), .ZN(n9221) );
  NAND2_X1 U9341 ( .A1(n7702), .A2(n9221), .ZN(n7705) );
  MUX2_X1 U9342 ( .A(n8980), .B(n7703), .S(n7752), .Z(n7704) );
  MUX2_X1 U9343 ( .A(n7706), .B(n9179), .S(n7752), .Z(n7707) );
  INV_X1 U9344 ( .A(n8987), .ZN(n7711) );
  NAND3_X1 U9345 ( .A1(n7712), .A2(n7711), .A3(n8985), .ZN(n7718) );
  NAND2_X1 U9346 ( .A1(n7714), .A2(n7713), .ZN(n7715) );
  NAND2_X1 U9347 ( .A1(n7716), .A2(n7715), .ZN(n7717) );
  MUX2_X1 U9348 ( .A(n7718), .B(n7717), .S(n7752), .Z(n7724) );
  INV_X1 U9349 ( .A(n9132), .ZN(n7719) );
  NAND2_X1 U9350 ( .A1(n8991), .A2(n7721), .ZN(n7720) );
  INV_X1 U9351 ( .A(n7721), .ZN(n7723) );
  MUX2_X1 U9352 ( .A(n8995), .B(n7792), .S(n7753), .Z(n7725) );
  NAND2_X1 U9353 ( .A1(n7727), .A2(n7726), .ZN(n7736) );
  AOI21_X1 U9354 ( .B1(n9055), .B2(n8996), .A(n8973), .ZN(n7729) );
  MUX2_X1 U9355 ( .A(n9055), .B(n7729), .S(n7753), .Z(n7730) );
  OAI21_X1 U9356 ( .B1(n8996), .B2(n9055), .A(n7738), .ZN(n7734) );
  NAND2_X1 U9357 ( .A1(n7731), .A2(n8973), .ZN(n7732) );
  NAND2_X1 U9358 ( .A1(n8999), .A2(n7732), .ZN(n7733) );
  MUX2_X1 U9359 ( .A(n7734), .B(n7733), .S(n7752), .Z(n7735) );
  OAI21_X1 U9360 ( .B1(n7736), .B2(n9042), .A(n7735), .ZN(n7737) );
  MUX2_X1 U9361 ( .A(n8999), .B(n7738), .S(n7752), .Z(n7739) );
  NAND3_X1 U9362 ( .A1(n7741), .A2(n7740), .A3(n7739), .ZN(n7744) );
  MUX2_X1 U9363 ( .A(n7742), .B(n9001), .S(n7752), .Z(n7743) );
  AND2_X1 U9364 ( .A1(n7744), .A2(n7743), .ZN(n7749) );
  MUX2_X1 U9365 ( .A(n9027), .B(n9242), .S(n7752), .Z(n7745) );
  NAND3_X1 U9366 ( .A1(n7759), .A2(n7749), .A3(n7745), .ZN(n7746) );
  MUX2_X1 U9367 ( .A(n7746), .B(n7752), .S(n7758), .Z(n7748) );
  NAND2_X1 U9368 ( .A1(n7748), .A2(n7747), .ZN(n7763) );
  AND2_X1 U9369 ( .A1(n7806), .A2(n7752), .ZN(n7761) );
  INV_X1 U9370 ( .A(n7749), .ZN(n7751) );
  INV_X1 U9371 ( .A(n9242), .ZN(n9014) );
  NAND3_X1 U9372 ( .A1(n7751), .A2(n9014), .A3(n7750), .ZN(n7756) );
  NAND2_X1 U9373 ( .A1(n9027), .A2(n7752), .ZN(n7755) );
  NAND2_X1 U9374 ( .A1(n9242), .A2(n7753), .ZN(n7754) );
  NAND3_X1 U9375 ( .A1(n7756), .A2(n7755), .A3(n7754), .ZN(n7757) );
  NOR2_X1 U9376 ( .A1(n7758), .A2(n7757), .ZN(n7760) );
  MUX2_X1 U9377 ( .A(n7761), .B(n7760), .S(n7759), .Z(n7762) );
  INV_X1 U9378 ( .A(n7767), .ZN(n7769) );
  NOR2_X1 U9379 ( .A1(n7769), .A2(n7768), .ZN(n7770) );
  INV_X1 U9380 ( .A(n7772), .ZN(n7775) );
  NAND2_X1 U9381 ( .A1(n8885), .A2(n7773), .ZN(n7774) );
  NAND3_X1 U9382 ( .A1(n7775), .A2(n6099), .A3(n7774), .ZN(n7776) );
  NAND2_X1 U9383 ( .A1(n7777), .A2(n7776), .ZN(n7779) );
  OAI21_X1 U9384 ( .B1(n6974), .B2(n7779), .A(n7778), .ZN(n7781) );
  NAND2_X1 U9385 ( .A1(n7781), .A2(n7780), .ZN(n7783) );
  NAND2_X1 U9386 ( .A1(n7783), .A2(n7782), .ZN(n7786) );
  AOI21_X1 U9387 ( .B1(n7786), .B2(n7785), .A(n7784), .ZN(n7788) );
  OAI21_X1 U9388 ( .B1(n7789), .B2(n7788), .A(n7787), .ZN(n7790) );
  NAND2_X1 U9389 ( .A1(n7791), .A2(n7790), .ZN(n7793) );
  NAND4_X1 U9390 ( .A1(n7794), .A2(n7793), .A3(n7792), .A4(n8992), .ZN(n7795)
         );
  NAND2_X1 U9391 ( .A1(n7796), .A2(n7795), .ZN(n7797) );
  NAND3_X1 U9392 ( .A1(n9033), .A2(n7798), .A3(n7797), .ZN(n7799) );
  NOR2_X1 U9393 ( .A1(n7800), .A2(n7799), .ZN(n7804) );
  INV_X1 U9394 ( .A(n7801), .ZN(n7803) );
  OAI21_X1 U9395 ( .B1(n7804), .B2(n7803), .A(n7802), .ZN(n7805) );
  NAND2_X1 U9396 ( .A1(n4790), .A2(n7805), .ZN(n7807) );
  NAND2_X1 U9397 ( .A1(n7807), .A2(n7806), .ZN(n7810) );
  NAND2_X1 U9398 ( .A1(n7810), .A2(n7809), .ZN(n7811) );
  NAND2_X1 U9399 ( .A1(n7811), .A2(n7814), .ZN(n7820) );
  NAND3_X1 U9400 ( .A1(n7812), .A2(n9490), .A3(n9491), .ZN(n7817) );
  INV_X1 U9401 ( .A(P1_B_REG_SCAN_IN), .ZN(n7813) );
  AOI21_X1 U9402 ( .B1(n7815), .B2(n7814), .A(n7813), .ZN(n7816) );
  OAI21_X1 U9403 ( .B1(n7818), .B2(n7817), .A(n7816), .ZN(n7819) );
  OAI21_X1 U9404 ( .B1(n7821), .B2(n7820), .A(n7819), .ZN(P1_U3240) );
  XOR2_X1 U9405 ( .A(n7830), .B(n7822), .Z(n9663) );
  AOI21_X1 U9406 ( .B1(n7824), .B2(n7836), .A(n7823), .ZN(n9660) );
  NOR2_X1 U9407 ( .A1(n9418), .A2(n7825), .ZN(n7828) );
  OAI22_X1 U9408 ( .A1(n9424), .A2(n6184), .B1(n7826), .B2(n9419), .ZN(n7827)
         );
  AOI211_X1 U9409 ( .C1(n9660), .C2(n9446), .A(n7828), .B(n7827), .ZN(n7835)
         );
  NAND2_X1 U9410 ( .A1(n7831), .A2(n7830), .ZN(n7829) );
  OAI211_X1 U9411 ( .C1(n7831), .C2(n7830), .A(n7829), .B(n9414), .ZN(n7833)
         );
  AOI22_X1 U9412 ( .A1(n9136), .A2(n8881), .B1(n8879), .B2(n9188), .ZN(n7832)
         );
  NAND2_X1 U9413 ( .A1(n7833), .A2(n7832), .ZN(n9658) );
  NAND2_X1 U9414 ( .A1(n9658), .A2(n9424), .ZN(n7834) );
  OAI211_X1 U9415 ( .C1(n9663), .C2(n9217), .A(n7835), .B(n7834), .ZN(P1_U3285) );
  OAI211_X1 U9416 ( .C1(n7837), .C2(n9653), .A(n9661), .B(n7836), .ZN(n9650)
         );
  NOR2_X1 U9417 ( .A1(n9650), .A2(n9157), .ZN(n7845) );
  AOI21_X1 U9418 ( .B1(n7838), .B2(n6961), .A(n9433), .ZN(n7843) );
  OAI22_X1 U9419 ( .A1(n9437), .A2(n7840), .B1(n7839), .B2(n9435), .ZN(n7841)
         );
  AOI21_X1 U9420 ( .B1(n7843), .B2(n7842), .A(n7841), .ZN(n9651) );
  INV_X1 U9421 ( .A(n9651), .ZN(n7844) );
  AOI211_X1 U9422 ( .C1(n9439), .C2(n7846), .A(n7845), .B(n7844), .ZN(n7847)
         );
  MUX2_X1 U9423 ( .A(n7848), .B(n7847), .S(n9424), .Z(n7855) );
  NAND2_X1 U9424 ( .A1(n7849), .A2(n4523), .ZN(n7850) );
  AND2_X1 U9425 ( .A1(n7851), .A2(n7850), .ZN(n9655) );
  AOI22_X1 U9426 ( .A1(n9655), .A2(n7853), .B1(n9441), .B2(n7852), .ZN(n7854)
         );
  NAND2_X1 U9427 ( .A1(n7855), .A2(n7854), .ZN(P1_U3286) );
  NAND2_X1 U9428 ( .A1(n7857), .A2(n7856), .ZN(n7862) );
  INV_X1 U9429 ( .A(n7862), .ZN(n7859) );
  NAND3_X1 U9430 ( .A1(n7860), .A2(n8735), .A3(n7861), .ZN(n7867) );
  INV_X1 U9431 ( .A(n7861), .ZN(n7865) );
  AND2_X1 U9432 ( .A1(n7863), .A2(n7862), .ZN(n7864) );
  NAND2_X1 U9433 ( .A1(n9252), .A2(n5986), .ZN(n7870) );
  OR2_X1 U9434 ( .A1(n9058), .A2(n7868), .ZN(n7869) );
  NAND2_X1 U9435 ( .A1(n7870), .A2(n7869), .ZN(n7871) );
  XNOR2_X1 U9436 ( .A(n7871), .B(n4268), .ZN(n8133) );
  NOR2_X1 U9437 ( .A1(n9058), .A2(n8128), .ZN(n7872) );
  AOI21_X1 U9438 ( .B1(n9252), .B2(n4274), .A(n7872), .ZN(n8119) );
  XNOR2_X1 U9439 ( .A(n8133), .B(n8119), .ZN(n7873) );
  XNOR2_X1 U9440 ( .A(n8121), .B(n7873), .ZN(n7878) );
  AOI22_X1 U9441 ( .A1(n8848), .A2(n8973), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n7874) );
  OAI21_X1 U9442 ( .B1(n9044), .B2(n8850), .A(n7874), .ZN(n7876) );
  NOR2_X1 U9443 ( .A1(n9040), .A2(n8813), .ZN(n7875) );
  AOI211_X1 U9444 ( .C1(n9038), .C2(n8861), .A(n7876), .B(n7875), .ZN(n7877)
         );
  OAI21_X1 U9445 ( .B1(n7878), .B2(n8868), .A(n7877), .ZN(P1_U3212) );
  NAND2_X1 U9446 ( .A1(n7879), .A2(n8582), .ZN(n7887) );
  INV_X1 U9447 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7880) );
  OAI22_X1 U9448 ( .A1(n7881), .A2(n8587), .B1(n7880), .B2(n8567), .ZN(n7884)
         );
  NOR2_X1 U9449 ( .A1(n7882), .A2(n8370), .ZN(n7883) );
  AOI211_X1 U9450 ( .C1(n8581), .C2(n7885), .A(n7884), .B(n7883), .ZN(n7886)
         );
  OAI211_X1 U9451 ( .C1(n7888), .C2(n8462), .A(n7887), .B(n7886), .ZN(P2_U3267) );
  INV_X1 U9452 ( .A(n8047), .ZN(n8052) );
  NAND2_X1 U9453 ( .A1(n7891), .A2(n7898), .ZN(n7894) );
  OR2_X1 U9454 ( .A1(n7899), .A2(n7892), .ZN(n7893) );
  NAND2_X1 U9455 ( .A1(n7896), .A2(n7895), .ZN(n7903) );
  OR2_X1 U9456 ( .A1(n7899), .A2(n6440), .ZN(n7900) );
  INV_X1 U9457 ( .A(n8291), .ZN(n7902) );
  NAND2_X1 U9458 ( .A1(n8373), .A2(n7902), .ZN(n8059) );
  NAND2_X1 U9459 ( .A1(n8063), .A2(n8059), .ZN(n8066) );
  NAND3_X1 U9460 ( .A1(n7904), .A2(n7903), .A3(n8096), .ZN(n7906) );
  NAND2_X1 U9461 ( .A1(n8679), .A2(n7905), .ZN(n8058) );
  NAND2_X1 U9462 ( .A1(n7906), .A2(n8058), .ZN(n7907) );
  XNOR2_X1 U9463 ( .A(n7907), .B(n8417), .ZN(n8105) );
  NAND2_X1 U9464 ( .A1(n7909), .A2(n7908), .ZN(n8104) );
  NOR2_X1 U9465 ( .A1(n8109), .A2(n8099), .ZN(n7910) );
  INV_X1 U9466 ( .A(n7911), .ZN(n7959) );
  NAND2_X1 U9467 ( .A1(n7914), .A2(n7913), .ZN(n7917) );
  INV_X1 U9468 ( .A(n7946), .ZN(n7915) );
  AOI211_X1 U9469 ( .C1(n7941), .C2(n7917), .A(n7916), .B(n7915), .ZN(n7935)
         );
  INV_X1 U9470 ( .A(n7924), .ZN(n7920) );
  INV_X1 U9471 ( .A(n7927), .ZN(n7918) );
  AOI21_X1 U9472 ( .B1(n7920), .B2(n7919), .A(n7918), .ZN(n7922) );
  INV_X1 U9473 ( .A(n7928), .ZN(n7921) );
  OAI21_X1 U9474 ( .B1(n7922), .B2(n7921), .A(n7926), .ZN(n7932) );
  AOI21_X1 U9475 ( .B1(n7925), .B2(n7924), .A(n7923), .ZN(n7930) );
  NAND2_X1 U9476 ( .A1(n7927), .A2(n7926), .ZN(n7929) );
  OAI21_X1 U9477 ( .B1(n7930), .B2(n7929), .A(n7928), .ZN(n7931) );
  MUX2_X1 U9478 ( .A(n7932), .B(n7931), .S(n8045), .Z(n7933) );
  NAND3_X1 U9479 ( .A1(n7933), .A2(n7941), .A3(n6548), .ZN(n7934) );
  OAI21_X1 U9480 ( .B1(n7935), .B2(n4478), .A(n7934), .ZN(n7945) );
  OAI21_X1 U9481 ( .B1(n7939), .B2(n7938), .A(n7937), .ZN(n7940) );
  AOI21_X1 U9482 ( .B1(n7942), .B2(n7944), .A(n8045), .ZN(n7943) );
  AOI21_X1 U9483 ( .B1(n7945), .B2(n7944), .A(n7943), .ZN(n7951) );
  OAI21_X1 U9484 ( .B1(n7946), .B2(n8045), .A(n8076), .ZN(n7950) );
  MUX2_X1 U9485 ( .A(n7948), .B(n7947), .S(n8045), .Z(n7949) );
  OAI211_X1 U9486 ( .C1(n7951), .C2(n7950), .A(n8075), .B(n7949), .ZN(n7956)
         );
  NAND2_X1 U9487 ( .A1(n7952), .A2(n4478), .ZN(n7954) );
  NAND2_X1 U9488 ( .A1(n8309), .A2(n8045), .ZN(n7953) );
  MUX2_X1 U9489 ( .A(n7954), .B(n7953), .S(n9751), .Z(n7955) );
  NAND3_X1 U9490 ( .A1(n7956), .A2(n7960), .A3(n7955), .ZN(n7961) );
  NAND3_X1 U9491 ( .A1(n7961), .A2(n7965), .A3(n7963), .ZN(n7958) );
  NAND2_X1 U9492 ( .A1(n7961), .A2(n7960), .ZN(n7964) );
  NAND3_X1 U9493 ( .A1(n8083), .A2(n7966), .A3(n7965), .ZN(n7970) );
  INV_X1 U9494 ( .A(n7967), .ZN(n7969) );
  INV_X1 U9495 ( .A(n7971), .ZN(n7973) );
  MUX2_X1 U9496 ( .A(n7973), .B(n7972), .S(n8045), .Z(n7974) );
  MUX2_X1 U9497 ( .A(n7976), .B(n7975), .S(n8045), .Z(n7977) );
  OAI211_X1 U9498 ( .C1(n7979), .C2(n5168), .A(n7978), .B(n7977), .ZN(n7984)
         );
  MUX2_X1 U9499 ( .A(n7981), .B(n7980), .S(n8045), .Z(n7982) );
  NAND3_X1 U9500 ( .A1(n7984), .A2(n7983), .A3(n7982), .ZN(n7988) );
  MUX2_X1 U9501 ( .A(n7986), .B(n7985), .S(n8045), .Z(n7987) );
  NAND3_X1 U9502 ( .A1(n7988), .A2(n5380), .A3(n7987), .ZN(n7992) );
  AND2_X1 U9503 ( .A1(n7997), .A2(n7989), .ZN(n7990) );
  MUX2_X1 U9504 ( .A(n7990), .B(n8527), .S(n8045), .Z(n7991) );
  NAND3_X1 U9505 ( .A1(n7992), .A2(n7993), .A3(n7991), .ZN(n7999) );
  NAND2_X1 U9506 ( .A1(n7999), .A2(n7993), .ZN(n7996) );
  INV_X1 U9507 ( .A(n8008), .ZN(n7995) );
  INV_X1 U9508 ( .A(n8001), .ZN(n7994) );
  AOI211_X1 U9509 ( .C1(n7996), .C2(n7998), .A(n7995), .B(n7994), .ZN(n8004)
         );
  NAND3_X1 U9510 ( .A1(n7999), .A2(n7998), .A3(n7997), .ZN(n8002) );
  INV_X1 U9511 ( .A(n8005), .ZN(n8000) );
  AOI21_X1 U9512 ( .B1(n8002), .B2(n8001), .A(n8000), .ZN(n8003) );
  MUX2_X1 U9513 ( .A(n8004), .B(n8003), .S(n8045), .Z(n8013) );
  NAND2_X1 U9514 ( .A1(n8010), .A2(n8005), .ZN(n8006) );
  NAND2_X1 U9515 ( .A1(n8696), .A2(n8297), .ZN(n8009) );
  OAI211_X1 U9516 ( .C1(n8013), .C2(n8006), .A(n8015), .B(n8009), .ZN(n8007)
         );
  NAND2_X1 U9517 ( .A1(n8009), .A2(n8008), .ZN(n8012) );
  OAI211_X1 U9518 ( .C1(n8013), .C2(n8012), .A(n8011), .B(n8010), .ZN(n8014)
         );
  NAND3_X1 U9519 ( .A1(n8016), .A2(n8015), .A3(n8014), .ZN(n8018) );
  INV_X1 U9520 ( .A(n8019), .ZN(n8027) );
  NAND2_X1 U9521 ( .A1(n8021), .A2(n8020), .ZN(n8022) );
  INV_X1 U9522 ( .A(n8034), .ZN(n8032) );
  NAND2_X1 U9523 ( .A1(n8035), .A2(n8028), .ZN(n8029) );
  MUX2_X1 U9524 ( .A(n8030), .B(n8029), .S(n8045), .Z(n8031) );
  NOR3_X1 U9525 ( .A1(n8033), .A2(n8032), .A3(n8031), .ZN(n8039) );
  MUX2_X1 U9526 ( .A(n8035), .B(n8034), .S(n8045), .Z(n8036) );
  NAND2_X1 U9527 ( .A1(n8391), .A2(n8036), .ZN(n8038) );
  OAI21_X1 U9528 ( .B1(n8039), .B2(n8038), .A(n8037), .ZN(n8050) );
  NAND2_X1 U9529 ( .A1(n8041), .A2(n8040), .ZN(n8043) );
  NOR2_X1 U9530 ( .A1(n8403), .A2(n8293), .ZN(n8042) );
  MUX2_X1 U9531 ( .A(n8043), .B(n8042), .S(n8045), .Z(n8049) );
  MUX2_X1 U9532 ( .A(n8045), .B(n8149), .S(n8044), .Z(n8046) );
  OAI22_X1 U9533 ( .A1(n8047), .A2(n8046), .B1(n4478), .B2(n8292), .ZN(n8048)
         );
  OAI21_X1 U9534 ( .B1(n8050), .B2(n8049), .A(n8048), .ZN(n8055) );
  INV_X1 U9535 ( .A(n8060), .ZN(n8051) );
  AOI22_X1 U9536 ( .A1(n8056), .A2(n8059), .B1(n4478), .B2(n8066), .ZN(n8062)
         );
  NAND2_X1 U9537 ( .A1(n8058), .A2(n7895), .ZN(n8067) );
  AOI21_X1 U9538 ( .B1(n8060), .B2(n8059), .A(n8067), .ZN(n8061) );
  INV_X1 U9539 ( .A(n8064), .ZN(n8098) );
  INV_X1 U9540 ( .A(n8066), .ZN(n8096) );
  INV_X1 U9541 ( .A(n8067), .ZN(n8095) );
  INV_X1 U9542 ( .A(n8391), .ZN(n8388) );
  INV_X1 U9543 ( .A(n8068), .ZN(n8407) );
  INV_X1 U9544 ( .A(n8524), .ZN(n8528) );
  NOR2_X1 U9545 ( .A1(n9717), .A2(n8069), .ZN(n8072) );
  NOR2_X1 U9546 ( .A1(n5371), .A2(n5430), .ZN(n8071) );
  NAND4_X1 U9547 ( .A1(n8072), .A2(n8071), .A3(n4567), .A4(n6548), .ZN(n8074)
         );
  NOR3_X1 U9548 ( .A1(n8074), .A2(n8073), .A3(n4712), .ZN(n8078) );
  NAND4_X1 U9549 ( .A1(n8078), .A2(n8077), .A3(n8076), .A4(n8075), .ZN(n8080)
         );
  NOR2_X1 U9550 ( .A1(n8080), .A2(n8079), .ZN(n8081) );
  NAND4_X1 U9551 ( .A1(n8084), .A2(n8083), .A3(n8082), .A4(n8081), .ZN(n8085)
         );
  NOR4_X1 U9552 ( .A1(n8087), .A2(n8086), .A3(n5168), .A4(n8085), .ZN(n8088)
         );
  NAND4_X1 U9553 ( .A1(n8512), .A2(n5380), .A3(n8528), .A4(n8088), .ZN(n8089)
         );
  NOR4_X1 U9554 ( .A1(n8463), .A2(n8480), .A3(n8497), .A4(n8089), .ZN(n8090)
         );
  NAND4_X1 U9555 ( .A1(n8435), .A2(n8407), .A3(n8090), .A4(n4574), .ZN(n8091)
         );
  NOR4_X1 U9556 ( .A1(n8388), .A2(n8092), .A3(n8091), .A4(n8422), .ZN(n8093)
         );
  NAND4_X1 U9557 ( .A1(n8096), .A2(n8095), .A3(n8094), .A4(n8093), .ZN(n8097)
         );
  XNOR2_X1 U9558 ( .A(n8097), .B(n8417), .ZN(n8100) );
  AOI22_X1 U9559 ( .A1(n8100), .A2(n8099), .B1(n8098), .B2(n5430), .ZN(n8101)
         );
  AOI21_X1 U9560 ( .B1(n8105), .B2(n8104), .A(n8103), .ZN(n8112) );
  NAND4_X1 U9561 ( .A1(n8107), .A2(n8106), .A3(n9706), .A4(n8228), .ZN(n8108)
         );
  OAI211_X1 U9562 ( .C1(n8109), .C2(n8111), .A(n8108), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8110) );
  OAI21_X1 U9563 ( .B1(n8112), .B2(n8111), .A(n8110), .ZN(P2_U3244) );
  INV_X1 U9564 ( .A(n8113), .ZN(n9352) );
  OAI222_X1 U9565 ( .A1(n8114), .A2(P2_U3152), .B1(n7519), .B2(n9352), .C1(
        n9866), .C2(n4267), .ZN(P2_U3329) );
  OAI222_X1 U9566 ( .A1(n9349), .A2(n8118), .B1(n8117), .B2(n8116), .C1(
        P1_U3084), .C2(n8115), .ZN(P1_U3323) );
  INV_X1 U9567 ( .A(n8119), .ZN(n8132) );
  NAND2_X1 U9568 ( .A1(n9247), .A2(n5986), .ZN(n8124) );
  OR2_X1 U9569 ( .A1(n9044), .A2(n8122), .ZN(n8123) );
  NAND2_X1 U9570 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  XNOR2_X1 U9571 ( .A(n8125), .B(n5719), .ZN(n8130) );
  NAND2_X1 U9572 ( .A1(n9247), .A2(n4274), .ZN(n8127) );
  OAI21_X1 U9573 ( .B1(n9044), .B2(n8128), .A(n8127), .ZN(n8129) );
  XNOR2_X1 U9574 ( .A(n8130), .B(n8129), .ZN(n8137) );
  INV_X1 U9575 ( .A(n8137), .ZN(n8131) );
  NAND2_X1 U9576 ( .A1(n8131), .A2(n8806), .ZN(n8142) );
  NAND2_X1 U9577 ( .A1(n8133), .A2(n8132), .ZN(n8136) );
  NAND4_X1 U9578 ( .A1(n8143), .A2(n8806), .A3(n8137), .A4(n8136), .ZN(n8141)
         );
  AOI22_X1 U9579 ( .A1(n8860), .A2(n9027), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8135) );
  NAND2_X1 U9580 ( .A1(n8861), .A2(n9022), .ZN(n8134) );
  OAI211_X1 U9581 ( .C1(n9058), .C2(n8864), .A(n8135), .B(n8134), .ZN(n8139)
         );
  NOR3_X1 U9582 ( .A1(n8137), .A2(n8868), .A3(n8136), .ZN(n8138) );
  AOI211_X1 U9583 ( .C1(n8866), .C2(n9247), .A(n8139), .B(n8138), .ZN(n8140)
         );
  OAI211_X1 U9584 ( .C1(n8143), .C2(n8142), .A(n8141), .B(n8140), .ZN(P1_U3218) );
  INV_X1 U9585 ( .A(n8144), .ZN(n8148) );
  AOI21_X1 U9586 ( .B1(n8146), .B2(n8145), .A(n8289), .ZN(n8147) );
  NAND2_X1 U9587 ( .A1(n8148), .A2(n8147), .ZN(n8154) );
  OR2_X1 U9588 ( .A1(n8149), .A2(n8242), .ZN(n8151) );
  OR2_X1 U9589 ( .A1(n8182), .A2(n8264), .ZN(n8150) );
  NAND2_X1 U9590 ( .A1(n8151), .A2(n8150), .ZN(n8393) );
  OAI22_X1 U9591 ( .A1(n8399), .A2(n8285), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9934), .ZN(n8152) );
  AOI21_X1 U9592 ( .B1(n8393), .B2(n8281), .A(n8152), .ZN(n8153) );
  OAI211_X1 U9593 ( .C1(n8403), .C2(n8274), .A(n8154), .B(n8153), .ZN(P2_U3216) );
  XNOR2_X1 U9594 ( .A(n8155), .B(n4331), .ZN(n8162) );
  INV_X1 U9595 ( .A(n8455), .ZN(n8159) );
  OAI22_X1 U9596 ( .A1(n8157), .A2(n8242), .B1(n8156), .B2(n8264), .ZN(n8450)
         );
  AOI22_X1 U9597 ( .A1(n8450), .A2(n8281), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8158) );
  OAI21_X1 U9598 ( .B1(n8159), .B2(n8285), .A(n8158), .ZN(n8160) );
  AOI21_X1 U9599 ( .B1(n8626), .B2(n4262), .A(n8160), .ZN(n8161) );
  OAI21_X1 U9600 ( .B1(n8162), .B2(n8289), .A(n8161), .ZN(P2_U3218) );
  OAI21_X1 U9601 ( .B1(n4339), .B2(n8164), .A(n8163), .ZN(n8165) );
  NAND2_X1 U9602 ( .A1(n8165), .A2(n8239), .ZN(n8170) );
  OAI22_X1 U9603 ( .A1(n8173), .A2(n8242), .B1(n8166), .B2(n8264), .ZN(n8167)
         );
  INV_X1 U9604 ( .A(n8167), .ZN(n8513) );
  NAND2_X1 U9605 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8360) );
  OAI21_X1 U9606 ( .B1(n8269), .B2(n8513), .A(n8360), .ZN(n8168) );
  AOI21_X1 U9607 ( .B1(n8518), .B2(n8271), .A(n8168), .ZN(n8169) );
  OAI211_X1 U9608 ( .C1(n8703), .C2(n8274), .A(n8170), .B(n8169), .ZN(P2_U3221) );
  XNOR2_X1 U9609 ( .A(n8172), .B(n8171), .ZN(n8178) );
  NOR2_X1 U9610 ( .A1(n8173), .A2(n8264), .ZN(n8174) );
  AOI21_X1 U9611 ( .B1(n8296), .B2(n8267), .A(n8174), .ZN(n8483) );
  OAI22_X1 U9612 ( .A1(n8269), .A2(n8483), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9845), .ZN(n8176) );
  NOR2_X1 U9613 ( .A1(n8696), .A2(n8274), .ZN(n8175) );
  AOI211_X1 U9614 ( .C1(n8271), .C2(n8488), .A(n8176), .B(n8175), .ZN(n8177)
         );
  OAI21_X1 U9615 ( .B1(n8178), .B2(n8289), .A(n8177), .ZN(P2_U3225) );
  XNOR2_X1 U9616 ( .A(n5581), .B(n8179), .ZN(n8180) );
  XNOR2_X1 U9617 ( .A(n8181), .B(n8180), .ZN(n8189) );
  OR2_X1 U9618 ( .A1(n8182), .A2(n8242), .ZN(n8184) );
  NAND2_X1 U9619 ( .A1(n8295), .A2(n8228), .ZN(n8183) );
  AND2_X1 U9620 ( .A1(n8184), .A2(n8183), .ZN(n8425) );
  OAI22_X1 U9621 ( .A1(n8425), .A2(n8269), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8185), .ZN(n8186) );
  AOI21_X1 U9622 ( .B1(n8428), .B2(n8271), .A(n8186), .ZN(n8188) );
  NAND2_X1 U9623 ( .A1(n8616), .A2(n4262), .ZN(n8187) );
  OAI211_X1 U9624 ( .C1(n8189), .C2(n8289), .A(n8188), .B(n8187), .ZN(P2_U3227) );
  NAND2_X1 U9625 ( .A1(n4700), .A2(n8191), .ZN(n8192) );
  OAI21_X1 U9626 ( .B1(n4700), .B2(n8191), .A(n8192), .ZN(n8277) );
  NOR2_X1 U9627 ( .A1(n8277), .A2(n8278), .ZN(n8276) );
  INV_X1 U9628 ( .A(n8192), .ZN(n8194) );
  NOR3_X1 U9629 ( .A1(n8276), .A2(n8194), .A3(n8193), .ZN(n8197) );
  INV_X1 U9630 ( .A(n8195), .ZN(n8196) );
  OAI21_X1 U9631 ( .B1(n8197), .B2(n8196), .A(n8239), .ZN(n8203) );
  AOI22_X1 U9632 ( .A1(n8281), .A2(n8198), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n8202) );
  NAND2_X1 U9633 ( .A1(n8715), .A2(n4262), .ZN(n8201) );
  NAND2_X1 U9634 ( .A1(n8271), .A2(n8199), .ZN(n8200) );
  NAND4_X1 U9635 ( .A1(n8203), .A2(n8202), .A3(n8201), .A4(n8200), .ZN(
        P2_U3228) );
  XNOR2_X1 U9636 ( .A(n8205), .B(n8204), .ZN(n8213) );
  INV_X1 U9637 ( .A(n8553), .ZN(n8210) );
  OR2_X1 U9638 ( .A1(n8206), .A2(n8264), .ZN(n8208) );
  NAND2_X1 U9639 ( .A1(n8300), .A2(n8267), .ZN(n8207) );
  NAND2_X1 U9640 ( .A1(n8208), .A2(n8207), .ZN(n8547) );
  AOI22_X1 U9641 ( .A1(n8281), .A2(n8547), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8209) );
  OAI21_X1 U9642 ( .B1(n8210), .B2(n8285), .A(n8209), .ZN(n8211) );
  AOI21_X1 U9643 ( .B1(n8552), .B2(n4262), .A(n8211), .ZN(n8212) );
  OAI21_X1 U9644 ( .B1(n8213), .B2(n8289), .A(n8212), .ZN(P2_U3230) );
  AOI21_X1 U9645 ( .B1(n4331), .B2(n8155), .A(n8214), .ZN(n8218) );
  XNOR2_X1 U9646 ( .A(n8216), .B(n8215), .ZN(n8217) );
  XNOR2_X1 U9647 ( .A(n8218), .B(n8217), .ZN(n8225) );
  OR2_X1 U9648 ( .A1(n8265), .A2(n8242), .ZN(n8220) );
  OR2_X1 U9649 ( .A1(n8243), .A2(n8264), .ZN(n8219) );
  NAND2_X1 U9650 ( .A1(n8220), .A2(n8219), .ZN(n8444) );
  AOI22_X1 U9651 ( .A1(n8444), .A2(n8281), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8221) );
  OAI21_X1 U9652 ( .B1(n8437), .B2(n8285), .A(n8221), .ZN(n8222) );
  AOI21_X1 U9653 ( .B1(n8620), .B2(n4262), .A(n8222), .ZN(n8224) );
  OAI21_X1 U9654 ( .B1(n8225), .B2(n8289), .A(n8224), .ZN(P2_U3231) );
  XNOR2_X1 U9655 ( .A(n8227), .B(n8226), .ZN(n8235) );
  OR2_X1 U9656 ( .A1(n8244), .A2(n8242), .ZN(n8230) );
  NAND2_X1 U9657 ( .A1(n8299), .A2(n8228), .ZN(n8229) );
  AND2_X1 U9658 ( .A1(n8230), .A2(n8229), .ZN(n8499) );
  OAI22_X1 U9659 ( .A1(n8269), .A2(n8499), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8231), .ZN(n8233) );
  NOR2_X1 U9660 ( .A1(n4447), .A2(n8274), .ZN(n8232) );
  AOI211_X1 U9661 ( .C1(n8271), .C2(n8504), .A(n8233), .B(n8232), .ZN(n8234)
         );
  OAI21_X1 U9662 ( .B1(n8235), .B2(n8289), .A(n8234), .ZN(P2_U3235) );
  OAI21_X1 U9663 ( .B1(n8238), .B2(n8237), .A(n8236), .ZN(n8240) );
  NAND2_X1 U9664 ( .A1(n8240), .A2(n8239), .ZN(n8250) );
  INV_X1 U9665 ( .A(n8241), .ZN(n8472) );
  OR2_X1 U9666 ( .A1(n8243), .A2(n8242), .ZN(n8246) );
  OR2_X1 U9667 ( .A1(n8244), .A2(n8264), .ZN(n8245) );
  AND2_X1 U9668 ( .A1(n8246), .A2(n8245), .ZN(n8468) );
  OAI22_X1 U9669 ( .A1(n8468), .A2(n8269), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8247), .ZN(n8248) );
  AOI21_X1 U9670 ( .B1(n8472), .B2(n8271), .A(n8248), .ZN(n8249) );
  OAI211_X1 U9671 ( .C1(n8692), .C2(n8274), .A(n8250), .B(n8249), .ZN(P2_U3237) );
  XNOR2_X1 U9672 ( .A(n8252), .B(n8251), .ZN(n8259) );
  OR2_X1 U9673 ( .A1(n8253), .A2(n8264), .ZN(n8255) );
  NAND2_X1 U9674 ( .A1(n8299), .A2(n8267), .ZN(n8254) );
  AND2_X1 U9675 ( .A1(n8255), .A2(n8254), .ZN(n8530) );
  NAND2_X1 U9676 ( .A1(n8271), .A2(n8536), .ZN(n8256) );
  NAND2_X1 U9677 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8340) );
  OAI211_X1 U9678 ( .C1(n8269), .C2(n8530), .A(n8256), .B(n8340), .ZN(n8257)
         );
  AOI21_X1 U9679 ( .B1(n8535), .B2(n4262), .A(n8257), .ZN(n8258) );
  OAI21_X1 U9680 ( .B1(n8259), .B2(n8289), .A(n8258), .ZN(P2_U3240) );
  AOI211_X1 U9681 ( .C1(n8262), .C2(n8261), .A(n8289), .B(n8260), .ZN(n8263)
         );
  INV_X1 U9682 ( .A(n8263), .ZN(n8273) );
  NOR2_X1 U9683 ( .A1(n8265), .A2(n8264), .ZN(n8266) );
  AOI21_X1 U9684 ( .B1(n8293), .B2(n8267), .A(n8266), .ZN(n8411) );
  OAI22_X1 U9685 ( .A1(n8411), .A2(n8269), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8268), .ZN(n8270) );
  AOI21_X1 U9686 ( .B1(n8415), .B2(n8271), .A(n8270), .ZN(n8272) );
  OAI211_X1 U9687 ( .C1(n8275), .C2(n8274), .A(n8273), .B(n8272), .ZN(P2_U3242) );
  AOI21_X1 U9688 ( .B1(n8278), .B2(n8277), .A(n8276), .ZN(n8290) );
  INV_X1 U9689 ( .A(n8279), .ZN(n8284) );
  NAND2_X1 U9690 ( .A1(n8281), .A2(n8280), .ZN(n8283) );
  OAI211_X1 U9691 ( .C1(n8285), .C2(n8284), .A(n8283), .B(n8282), .ZN(n8286)
         );
  AOI21_X1 U9692 ( .B1(n8287), .B2(n4262), .A(n8286), .ZN(n8288) );
  OAI21_X1 U9693 ( .B1(n8290), .B2(n8289), .A(n8288), .ZN(P2_U3243) );
  MUX2_X1 U9694 ( .A(n8291), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8317), .Z(
        P2_U3582) );
  MUX2_X1 U9695 ( .A(n8292), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8317), .Z(
        P2_U3580) );
  MUX2_X1 U9696 ( .A(n8293), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8317), .Z(
        P2_U3579) );
  MUX2_X1 U9697 ( .A(n8294), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8317), .Z(
        P2_U3577) );
  MUX2_X1 U9698 ( .A(n8295), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8317), .Z(
        P2_U3576) );
  MUX2_X1 U9699 ( .A(n8296), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8317), .Z(
        P2_U3574) );
  MUX2_X1 U9700 ( .A(n8297), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8317), .Z(
        P2_U3573) );
  MUX2_X1 U9701 ( .A(n8298), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8317), .Z(
        P2_U3572) );
  MUX2_X1 U9702 ( .A(n8299), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8317), .Z(
        P2_U3571) );
  MUX2_X1 U9703 ( .A(n8300), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8317), .Z(
        P2_U3570) );
  MUX2_X1 U9704 ( .A(n8301), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8317), .Z(
        P2_U3569) );
  MUX2_X1 U9705 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8302), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9706 ( .A(n8303), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8317), .Z(
        P2_U3566) );
  MUX2_X1 U9707 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8304), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9708 ( .A(n8305), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8317), .Z(
        P2_U3564) );
  MUX2_X1 U9709 ( .A(n8306), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8317), .Z(
        P2_U3563) );
  MUX2_X1 U9710 ( .A(n8307), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8317), .Z(
        P2_U3562) );
  MUX2_X1 U9711 ( .A(n8308), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8317), .Z(
        P2_U3561) );
  MUX2_X1 U9712 ( .A(n8309), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8317), .Z(
        P2_U3560) );
  MUX2_X1 U9713 ( .A(n8310), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8317), .Z(
        P2_U3559) );
  MUX2_X1 U9714 ( .A(n8311), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8317), .Z(
        P2_U3558) );
  MUX2_X1 U9715 ( .A(n8312), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8317), .Z(
        P2_U3557) );
  MUX2_X1 U9716 ( .A(n8313), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8317), .Z(
        P2_U3556) );
  MUX2_X1 U9717 ( .A(n8314), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8317), .Z(
        P2_U3555) );
  MUX2_X1 U9718 ( .A(n8315), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8317), .Z(
        P2_U3554) );
  MUX2_X1 U9719 ( .A(n8316), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8317), .Z(
        P2_U3553) );
  MUX2_X1 U9720 ( .A(n5369), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8317), .Z(
        P2_U3552) );
  NAND2_X1 U9721 ( .A1(n8337), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8319) );
  OAI21_X1 U9722 ( .B1(n8337), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8319), .ZN(
        n8320) );
  NOR2_X1 U9723 ( .A1(n8321), .A2(n8320), .ZN(n8336) );
  AOI211_X1 U9724 ( .C1(n8321), .C2(n8320), .A(n8336), .B(n9951), .ZN(n8331)
         );
  INV_X1 U9725 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8659) );
  XNOR2_X1 U9726 ( .A(n8337), .B(n8659), .ZN(n8326) );
  INV_X1 U9727 ( .A(n8322), .ZN(n8324) );
  INV_X1 U9728 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8665) );
  AOI21_X1 U9729 ( .B1(n8324), .B2(n8665), .A(n8323), .ZN(n8325) );
  NAND2_X1 U9730 ( .A1(n8326), .A2(n8325), .ZN(n8332) );
  OAI211_X1 U9731 ( .C1(n8326), .C2(n8325), .A(n9956), .B(n8332), .ZN(n8329)
         );
  AND2_X1 U9732 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8327) );
  AOI21_X1 U9733 ( .B1(n9960), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8327), .ZN(
        n8328) );
  OAI211_X1 U9734 ( .C1(n9964), .C2(n8333), .A(n8329), .B(n8328), .ZN(n8330)
         );
  OR2_X1 U9735 ( .A1(n8331), .A2(n8330), .ZN(P2_U3262) );
  OAI21_X1 U9736 ( .B1(n8659), .B2(n8333), .A(n8332), .ZN(n8335) );
  INV_X1 U9737 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8654) );
  AOI22_X1 U9738 ( .A1(n8342), .A2(n8654), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8351), .ZN(n8334) );
  NOR2_X1 U9739 ( .A1(n8335), .A2(n8334), .ZN(n8350) );
  AOI21_X1 U9740 ( .B1(n8335), .B2(n8334), .A(n8350), .ZN(n8345) );
  INV_X1 U9741 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9895) );
  OAI21_X1 U9742 ( .B1(n8338), .B2(n9895), .A(n8347), .ZN(n8339) );
  NAND2_X1 U9743 ( .A1(n8339), .A2(n9697), .ZN(n8344) );
  INV_X1 U9744 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9978) );
  OAI21_X1 U9745 ( .B1(n8362), .B2(n9978), .A(n8340), .ZN(n8341) );
  AOI21_X1 U9746 ( .B1(n9359), .B2(n8342), .A(n8341), .ZN(n8343) );
  OAI211_X1 U9747 ( .C1(n8345), .C2(n9699), .A(n8344), .B(n8343), .ZN(P2_U3263) );
  NAND2_X1 U9748 ( .A1(n8346), .A2(n8351), .ZN(n8348) );
  XNOR2_X1 U9749 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8349), .ZN(n8356) );
  INV_X1 U9750 ( .A(n8356), .ZN(n8354) );
  INV_X1 U9751 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8649) );
  AOI21_X1 U9752 ( .B1(n8351), .B2(n8654), .A(n8350), .ZN(n8352) );
  XNOR2_X1 U9753 ( .A(n8649), .B(n8352), .ZN(n8355) );
  OAI21_X1 U9754 ( .B1(n8355), .B2(n9699), .A(n9964), .ZN(n8353) );
  AOI21_X1 U9755 ( .B1(n8354), .B2(n9697), .A(n8353), .ZN(n8359) );
  AOI22_X1 U9756 ( .A1(n8356), .A2(n9697), .B1(n9956), .B2(n8355), .ZN(n8358)
         );
  MUX2_X1 U9757 ( .A(n8359), .B(n8358), .S(n8357), .Z(n8361) );
  OAI211_X1 U9758 ( .C1(n8363), .C2(n8362), .A(n8361), .B(n8360), .ZN(P2_U3264) );
  XNOR2_X1 U9759 ( .A(n8679), .B(n8371), .ZN(n8365) );
  OR2_X1 U9760 ( .A1(n8365), .A2(n9752), .ZN(n8597) );
  NAND2_X1 U9761 ( .A1(n8367), .A2(n8366), .ZN(n8600) );
  NOR2_X1 U9762 ( .A1(n8462), .A2(n8600), .ZN(n8375) );
  AOI21_X1 U9763 ( .B1(n8462), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8375), .ZN(
        n8369) );
  NAND2_X1 U9764 ( .A1(n8679), .A2(n8581), .ZN(n8368) );
  OAI211_X1 U9765 ( .C1(n8597), .C2(n8370), .A(n8369), .B(n8368), .ZN(P2_U3265) );
  INV_X1 U9766 ( .A(n8371), .ZN(n8372) );
  AOI211_X1 U9767 ( .C1(n8374), .C2(n8373), .A(n9752), .B(n8372), .ZN(n8602)
         );
  NAND2_X1 U9768 ( .A1(n8602), .A2(n8572), .ZN(n8377) );
  AOI21_X1 U9769 ( .B1(n8462), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8375), .ZN(
        n8376) );
  OAI211_X1 U9770 ( .C1(n8364), .C2(n8556), .A(n8377), .B(n8376), .ZN(P2_U3266) );
  INV_X1 U9771 ( .A(n8378), .ZN(n8387) );
  NAND2_X1 U9772 ( .A1(n8379), .A2(n8582), .ZN(n8386) );
  AOI22_X1 U9773 ( .A1(n8380), .A2(n8566), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8462), .ZN(n8381) );
  OAI21_X1 U9774 ( .B1(n8382), .B2(n8556), .A(n8381), .ZN(n8383) );
  AOI21_X1 U9775 ( .B1(n8384), .B2(n8572), .A(n8383), .ZN(n8385) );
  OAI211_X1 U9776 ( .C1(n8387), .C2(n8462), .A(n8386), .B(n8385), .ZN(P2_U3268) );
  XNOR2_X1 U9777 ( .A(n8389), .B(n8388), .ZN(n8608) );
  OAI211_X1 U9778 ( .C1(n8392), .C2(n8391), .A(n8390), .B(n8585), .ZN(n8395)
         );
  INV_X1 U9779 ( .A(n8393), .ZN(n8394) );
  NAND2_X1 U9780 ( .A1(n8395), .A2(n8394), .ZN(n8604) );
  INV_X1 U9781 ( .A(n8413), .ZN(n8398) );
  INV_X1 U9782 ( .A(n8396), .ZN(n8397) );
  AOI211_X1 U9783 ( .C1(n8606), .C2(n8398), .A(n9752), .B(n8397), .ZN(n8605)
         );
  NAND2_X1 U9784 ( .A1(n8605), .A2(n8572), .ZN(n8402) );
  INV_X1 U9785 ( .A(n8399), .ZN(n8400) );
  AOI22_X1 U9786 ( .A1(n8400), .A2(n8566), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8462), .ZN(n8401) );
  OAI211_X1 U9787 ( .C1(n8403), .C2(n8556), .A(n8402), .B(n8401), .ZN(n8404)
         );
  AOI21_X1 U9788 ( .B1(n8604), .B2(n8567), .A(n8404), .ZN(n8405) );
  OAI21_X1 U9789 ( .B1(n8608), .B2(n8559), .A(n8405), .ZN(P2_U3269) );
  XNOR2_X1 U9790 ( .A(n8406), .B(n8407), .ZN(n8613) );
  AOI22_X1 U9791 ( .A1(n8611), .A2(n8581), .B1(n8462), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8421) );
  AOI21_X1 U9792 ( .B1(n4730), .B2(n8408), .A(n8407), .ZN(n8409) );
  OAI21_X1 U9793 ( .B1(n8410), .B2(n8409), .A(n8585), .ZN(n8412) );
  NAND2_X1 U9794 ( .A1(n8412), .A2(n8411), .ZN(n8609) );
  INV_X1 U9795 ( .A(n8427), .ZN(n8414) );
  AOI211_X1 U9796 ( .C1(n8611), .C2(n8414), .A(n9752), .B(n8413), .ZN(n8610)
         );
  INV_X1 U9797 ( .A(n8610), .ZN(n8418) );
  INV_X1 U9798 ( .A(n8415), .ZN(n8416) );
  OAI22_X1 U9799 ( .A1(n8418), .A2(n8417), .B1(n8587), .B2(n8416), .ZN(n8419)
         );
  OAI21_X1 U9800 ( .B1(n8609), .B2(n8419), .A(n8567), .ZN(n8420) );
  OAI211_X1 U9801 ( .C1(n8613), .C2(n8559), .A(n8421), .B(n8420), .ZN(P2_U3270) );
  XNOR2_X1 U9802 ( .A(n8423), .B(n8422), .ZN(n8618) );
  OAI211_X1 U9803 ( .C1(n8424), .C2(n4319), .A(n4730), .B(n8585), .ZN(n8426)
         );
  NAND2_X1 U9804 ( .A1(n8426), .A2(n8425), .ZN(n8614) );
  INV_X1 U9805 ( .A(n8616), .ZN(n8431) );
  AOI211_X1 U9806 ( .C1(n8616), .C2(n8436), .A(n9752), .B(n8427), .ZN(n8615)
         );
  NAND2_X1 U9807 ( .A1(n8615), .A2(n8572), .ZN(n8430) );
  AOI22_X1 U9808 ( .A1(n8462), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8428), .B2(
        n8566), .ZN(n8429) );
  OAI211_X1 U9809 ( .C1(n8431), .C2(n8556), .A(n8430), .B(n8429), .ZN(n8432)
         );
  AOI21_X1 U9810 ( .B1(n8614), .B2(n8567), .A(n8432), .ZN(n8433) );
  OAI21_X1 U9811 ( .B1(n8618), .B2(n8559), .A(n8433), .ZN(P2_U3271) );
  AOI21_X1 U9812 ( .B1(n8435), .B2(n8434), .A(n4309), .ZN(n8623) );
  AOI211_X1 U9813 ( .C1(n8620), .C2(n8454), .A(n9752), .B(n5402), .ZN(n8619)
         );
  INV_X1 U9814 ( .A(n8437), .ZN(n8438) );
  AOI22_X1 U9815 ( .A1(n8462), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8438), .B2(
        n8566), .ZN(n8439) );
  OAI21_X1 U9816 ( .B1(n8440), .B2(n8556), .A(n8439), .ZN(n8447) );
  AOI211_X1 U9817 ( .C1(n8443), .C2(n8442), .A(n8531), .B(n8441), .ZN(n8445)
         );
  NOR2_X1 U9818 ( .A1(n8445), .A2(n8444), .ZN(n8622) );
  NOR2_X1 U9819 ( .A1(n8622), .A2(n8462), .ZN(n8446) );
  AOI211_X1 U9820 ( .C1(n8619), .C2(n8572), .A(n8447), .B(n8446), .ZN(n8448)
         );
  OAI21_X1 U9821 ( .B1(n8623), .B2(n8559), .A(n8448), .ZN(P2_U3272) );
  XNOR2_X1 U9822 ( .A(n8449), .B(n8452), .ZN(n8451) );
  AOI21_X1 U9823 ( .B1(n8451), .B2(n8585), .A(n8450), .ZN(n8629) );
  OR2_X1 U9824 ( .A1(n8453), .A2(n8452), .ZN(n8625) );
  NAND3_X1 U9825 ( .A1(n8625), .A2(n8624), .A3(n8582), .ZN(n8461) );
  OAI211_X1 U9826 ( .C1(n8470), .C2(n8457), .A(n8454), .B(n8670), .ZN(n8628)
         );
  INV_X1 U9827 ( .A(n8628), .ZN(n8459) );
  AOI22_X1 U9828 ( .A1(n8462), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8455), .B2(
        n8566), .ZN(n8456) );
  OAI21_X1 U9829 ( .B1(n8457), .B2(n8556), .A(n8456), .ZN(n8458) );
  AOI21_X1 U9830 ( .B1(n8459), .B2(n8572), .A(n8458), .ZN(n8460) );
  OAI211_X1 U9831 ( .C1(n8462), .C2(n8629), .A(n8461), .B(n8460), .ZN(P2_U3273) );
  XNOR2_X1 U9832 ( .A(n8464), .B(n8463), .ZN(n8633) );
  INV_X1 U9833 ( .A(n8633), .ZN(n8477) );
  OAI211_X1 U9834 ( .C1(n8467), .C2(n8466), .A(n8465), .B(n8585), .ZN(n8469)
         );
  NAND2_X1 U9835 ( .A1(n8469), .A2(n8468), .ZN(n8631) );
  AOI211_X1 U9836 ( .C1(n8471), .C2(n8485), .A(n9752), .B(n8470), .ZN(n8632)
         );
  NAND2_X1 U9837 ( .A1(n8632), .A2(n8572), .ZN(n8474) );
  AOI22_X1 U9838 ( .A1(n8462), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8472), .B2(
        n8566), .ZN(n8473) );
  OAI211_X1 U9839 ( .C1(n8692), .C2(n8556), .A(n8474), .B(n8473), .ZN(n8475)
         );
  AOI21_X1 U9840 ( .B1(n8631), .B2(n8567), .A(n8475), .ZN(n8476) );
  OAI21_X1 U9841 ( .B1(n8477), .B2(n8559), .A(n8476), .ZN(P2_U3274) );
  XNOR2_X1 U9842 ( .A(n8479), .B(n8480), .ZN(n8638) );
  INV_X1 U9843 ( .A(n8638), .ZN(n8493) );
  XNOR2_X1 U9844 ( .A(n8481), .B(n8480), .ZN(n8482) );
  NAND2_X1 U9845 ( .A1(n8482), .A2(n8585), .ZN(n8484) );
  NAND2_X1 U9846 ( .A1(n8484), .A2(n8483), .ZN(n8636) );
  INV_X1 U9847 ( .A(n8485), .ZN(n8486) );
  AOI211_X1 U9848 ( .C1(n8487), .C2(n8501), .A(n9752), .B(n8486), .ZN(n8637)
         );
  NAND2_X1 U9849 ( .A1(n8637), .A2(n8572), .ZN(n8490) );
  AOI22_X1 U9850 ( .A1(n8462), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8488), .B2(
        n8566), .ZN(n8489) );
  OAI211_X1 U9851 ( .C1(n8696), .C2(n8556), .A(n8490), .B(n8489), .ZN(n8491)
         );
  AOI21_X1 U9852 ( .B1(n8636), .B2(n8567), .A(n8491), .ZN(n8492) );
  OAI21_X1 U9853 ( .B1(n8493), .B2(n8559), .A(n8492), .ZN(P2_U3275) );
  XOR2_X1 U9854 ( .A(n8494), .B(n8497), .Z(n8643) );
  INV_X1 U9855 ( .A(n8643), .ZN(n8509) );
  NAND2_X1 U9856 ( .A1(n8496), .A2(n8497), .ZN(n8498) );
  NAND3_X1 U9857 ( .A1(n8495), .A2(n8585), .A3(n8498), .ZN(n8500) );
  NAND2_X1 U9858 ( .A1(n8500), .A2(n8499), .ZN(n8641) );
  INV_X1 U9859 ( .A(n8501), .ZN(n8502) );
  AOI211_X1 U9860 ( .C1(n8503), .C2(n8515), .A(n9752), .B(n8502), .ZN(n8642)
         );
  NAND2_X1 U9861 ( .A1(n8642), .A2(n8572), .ZN(n8506) );
  AOI22_X1 U9862 ( .A1(n8462), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8504), .B2(
        n8566), .ZN(n8505) );
  OAI211_X1 U9863 ( .C1(n4447), .C2(n8556), .A(n8506), .B(n8505), .ZN(n8507)
         );
  AOI21_X1 U9864 ( .B1(n8641), .B2(n8567), .A(n8507), .ZN(n8508) );
  OAI21_X1 U9865 ( .B1(n8509), .B2(n8559), .A(n8508), .ZN(P2_U3276) );
  XNOR2_X1 U9866 ( .A(n8510), .B(n8512), .ZN(n8648) );
  INV_X1 U9867 ( .A(n8648), .ZN(n8523) );
  XOR2_X1 U9868 ( .A(n8511), .B(n8512), .Z(n8514) );
  OAI21_X1 U9869 ( .B1(n8514), .B2(n8531), .A(n8513), .ZN(n8646) );
  INV_X1 U9870 ( .A(n8533), .ZN(n8516) );
  AOI211_X1 U9871 ( .C1(n8517), .C2(n8516), .A(n9752), .B(n4448), .ZN(n8647)
         );
  NAND2_X1 U9872 ( .A1(n8647), .A2(n8572), .ZN(n8520) );
  AOI22_X1 U9873 ( .A1(n8462), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8518), .B2(
        n8566), .ZN(n8519) );
  OAI211_X1 U9874 ( .C1(n8703), .C2(n8556), .A(n8520), .B(n8519), .ZN(n8521)
         );
  AOI21_X1 U9875 ( .B1(n8646), .B2(n8567), .A(n8521), .ZN(n8522) );
  OAI21_X1 U9876 ( .B1(n8523), .B2(n8559), .A(n8522), .ZN(P2_U3277) );
  XNOR2_X1 U9877 ( .A(n8525), .B(n8524), .ZN(n8653) );
  INV_X1 U9878 ( .A(n8653), .ZN(n8541) );
  NAND2_X1 U9879 ( .A1(n8526), .A2(n8527), .ZN(n8529) );
  XNOR2_X1 U9880 ( .A(n8529), .B(n8528), .ZN(n8532) );
  OAI21_X1 U9881 ( .B1(n8532), .B2(n8531), .A(n8530), .ZN(n8651) );
  INV_X1 U9882 ( .A(n8550), .ZN(n8534) );
  AOI211_X1 U9883 ( .C1(n8535), .C2(n8534), .A(n9752), .B(n8533), .ZN(n8652)
         );
  NAND2_X1 U9884 ( .A1(n8652), .A2(n8572), .ZN(n8538) );
  AOI22_X1 U9885 ( .A1(n8462), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8536), .B2(
        n8566), .ZN(n8537) );
  OAI211_X1 U9886 ( .C1(n8707), .C2(n8556), .A(n8538), .B(n8537), .ZN(n8539)
         );
  AOI21_X1 U9887 ( .B1(n8651), .B2(n8567), .A(n8539), .ZN(n8540) );
  OAI21_X1 U9888 ( .B1(n8541), .B2(n8559), .A(n8540), .ZN(P2_U3278) );
  OAI21_X1 U9889 ( .B1(n8543), .B2(n8544), .A(n8542), .ZN(n8658) );
  INV_X1 U9890 ( .A(n8658), .ZN(n8560) );
  NAND2_X1 U9891 ( .A1(n8545), .A2(n8544), .ZN(n8546) );
  NAND3_X1 U9892 ( .A1(n8526), .A2(n8585), .A3(n8546), .ZN(n8549) );
  INV_X1 U9893 ( .A(n8547), .ZN(n8548) );
  NAND2_X1 U9894 ( .A1(n8549), .A2(n8548), .ZN(n8656) );
  AOI211_X1 U9895 ( .C1(n8552), .C2(n8551), .A(n9752), .B(n8550), .ZN(n8657)
         );
  NAND2_X1 U9896 ( .A1(n8657), .A2(n8572), .ZN(n8555) );
  AOI22_X1 U9897 ( .A1(n8462), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8553), .B2(
        n8566), .ZN(n8554) );
  OAI211_X1 U9898 ( .C1(n5201), .C2(n8556), .A(n8555), .B(n8554), .ZN(n8557)
         );
  AOI21_X1 U9899 ( .B1(n8656), .B2(n8567), .A(n8557), .ZN(n8558) );
  OAI21_X1 U9900 ( .B1(n8560), .B2(n8559), .A(n8558), .ZN(P2_U3279) );
  NAND2_X1 U9901 ( .A1(n8562), .A2(n5371), .ZN(n8563) );
  NAND2_X1 U9902 ( .A1(n8561), .A2(n8563), .ZN(n8565) );
  AOI21_X1 U9903 ( .B1(n8565), .B2(n8585), .A(n8564), .ZN(n9730) );
  INV_X1 U9904 ( .A(n9730), .ZN(n8568) );
  AOI22_X1 U9905 ( .A1(n8568), .A2(n8567), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8566), .ZN(n8578) );
  INV_X1 U9906 ( .A(n8592), .ZN(n8570) );
  OAI211_X1 U9907 ( .C1(n9731), .C2(n8570), .A(n8569), .B(n8670), .ZN(n9729)
         );
  INV_X1 U9908 ( .A(n9729), .ZN(n8571) );
  AOI22_X1 U9909 ( .A1(n8572), .A2(n8571), .B1(n8462), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n8577) );
  OAI21_X1 U9910 ( .B1(n8574), .B2(n5371), .A(n8573), .ZN(n9733) );
  AOI22_X1 U9911 ( .A1(n8582), .A2(n9733), .B1(n8581), .B2(n8575), .ZN(n8576)
         );
  NAND3_X1 U9912 ( .A1(n8578), .A2(n8577), .A3(n8576), .ZN(P2_U3294) );
  OAI21_X1 U9913 ( .B1(n8069), .B2(n8580), .A(n8579), .ZN(n9727) );
  AOI22_X1 U9914 ( .A1(n8582), .A2(n9727), .B1(n8581), .B2(n8590), .ZN(n8596)
         );
  XNOR2_X1 U9915 ( .A(n8069), .B(n8583), .ZN(n8586) );
  AOI21_X1 U9916 ( .B1(n8586), .B2(n8585), .A(n8584), .ZN(n9724) );
  OAI22_X1 U9917 ( .A1(n8462), .A2(n9724), .B1(n8588), .B2(n8587), .ZN(n8589)
         );
  INV_X1 U9918 ( .A(n8589), .ZN(n8595) );
  NAND2_X1 U9919 ( .A1(n8590), .A2(n9715), .ZN(n8591) );
  AND2_X1 U9920 ( .A1(n8592), .A2(n8591), .ZN(n9721) );
  AOI22_X1 U9921 ( .A1(n8593), .A2(n9721), .B1(n8462), .B2(
        P2_REG2_REG_1__SCAN_IN), .ZN(n8594) );
  NAND3_X1 U9922 ( .A1(n8596), .A2(n8595), .A3(n8594), .ZN(P2_U3295) );
  NAND2_X1 U9923 ( .A1(n8597), .A2(n8600), .ZN(n8677) );
  MUX2_X1 U9924 ( .A(n8677), .B(P2_REG1_REG_31__SCAN_IN), .S(n9767), .Z(n8598)
         );
  AOI21_X1 U9925 ( .B1(n5451), .B2(n8679), .A(n8598), .ZN(n8599) );
  INV_X1 U9926 ( .A(n8599), .ZN(P2_U3551) );
  INV_X1 U9927 ( .A(n8600), .ZN(n8601) );
  NOR2_X1 U9928 ( .A1(n8602), .A2(n8601), .ZN(n8681) );
  MUX2_X1 U9929 ( .A(n9830), .B(n8681), .S(n8676), .Z(n8603) );
  OAI21_X1 U9930 ( .B1(n8364), .B2(n8667), .A(n8603), .ZN(P2_U3550) );
  OAI21_X1 U9931 ( .B1(n8608), .B2(n8674), .A(n8607), .ZN(n8684) );
  MUX2_X1 U9932 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8684), .S(n9770), .Z(
        P2_U3547) );
  OAI21_X1 U9933 ( .B1(n8613), .B2(n8674), .A(n8612), .ZN(n8685) );
  MUX2_X1 U9934 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8685), .S(n9770), .Z(
        P2_U3546) );
  OAI21_X1 U9935 ( .B1(n8618), .B2(n8674), .A(n8617), .ZN(n8686) );
  MUX2_X1 U9936 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8686), .S(n9770), .Z(
        P2_U3545) );
  AOI21_X1 U9937 ( .B1(n9722), .B2(n8620), .A(n8619), .ZN(n8621) );
  OAI211_X1 U9938 ( .C1(n8623), .C2(n8674), .A(n8622), .B(n8621), .ZN(n8687)
         );
  MUX2_X1 U9939 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8687), .S(n8676), .Z(
        P2_U3544) );
  NAND3_X1 U9940 ( .A1(n8625), .A2(n8624), .A3(n9746), .ZN(n8630) );
  NAND2_X1 U9941 ( .A1(n8626), .A2(n9722), .ZN(n8627) );
  NAND4_X1 U9942 ( .A1(n8630), .A2(n8629), .A3(n8628), .A4(n8627), .ZN(n8688)
         );
  MUX2_X1 U9943 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8688), .S(n8676), .Z(
        P2_U3543) );
  INV_X1 U9944 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8634) );
  AOI211_X1 U9945 ( .C1(n8633), .C2(n9746), .A(n8632), .B(n8631), .ZN(n8689)
         );
  MUX2_X1 U9946 ( .A(n8634), .B(n8689), .S(n9770), .Z(n8635) );
  OAI21_X1 U9947 ( .B1(n8692), .B2(n8667), .A(n8635), .ZN(P2_U3542) );
  INV_X1 U9948 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8639) );
  AOI211_X1 U9949 ( .C1(n8638), .C2(n9746), .A(n8637), .B(n8636), .ZN(n8693)
         );
  MUX2_X1 U9950 ( .A(n8639), .B(n8693), .S(n9770), .Z(n8640) );
  OAI21_X1 U9951 ( .B1(n8696), .B2(n8667), .A(n8640), .ZN(P2_U3541) );
  INV_X1 U9952 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8644) );
  AOI211_X1 U9953 ( .C1(n8643), .C2(n9746), .A(n8642), .B(n8641), .ZN(n8697)
         );
  MUX2_X1 U9954 ( .A(n8644), .B(n8697), .S(n8676), .Z(n8645) );
  OAI21_X1 U9955 ( .B1(n4447), .B2(n8667), .A(n8645), .ZN(P2_U3540) );
  AOI211_X1 U9956 ( .C1(n8648), .C2(n9746), .A(n8647), .B(n8646), .ZN(n8700)
         );
  MUX2_X1 U9957 ( .A(n8649), .B(n8700), .S(n9770), .Z(n8650) );
  OAI21_X1 U9958 ( .B1(n8703), .B2(n8667), .A(n8650), .ZN(P2_U3539) );
  AOI211_X1 U9959 ( .C1(n8653), .C2(n9746), .A(n8652), .B(n8651), .ZN(n8704)
         );
  MUX2_X1 U9960 ( .A(n8654), .B(n8704), .S(n9770), .Z(n8655) );
  OAI21_X1 U9961 ( .B1(n8707), .B2(n8667), .A(n8655), .ZN(P2_U3538) );
  AOI211_X1 U9962 ( .C1(n8658), .C2(n9746), .A(n8657), .B(n8656), .ZN(n8708)
         );
  MUX2_X1 U9963 ( .A(n8659), .B(n8708), .S(n9770), .Z(n8660) );
  OAI21_X1 U9964 ( .B1(n5201), .B2(n8667), .A(n8660), .ZN(P2_U3537) );
  NAND2_X1 U9965 ( .A1(n8662), .A2(n8661), .ZN(n8663) );
  AOI21_X1 U9966 ( .B1(n8664), .B2(n9746), .A(n8663), .ZN(n8712) );
  MUX2_X1 U9967 ( .A(n8665), .B(n8712), .S(n9770), .Z(n8666) );
  OAI21_X1 U9968 ( .B1(n8668), .B2(n8667), .A(n8666), .ZN(P2_U3536) );
  AOI22_X1 U9969 ( .A1(n8671), .A2(n8670), .B1(n9722), .B2(n8669), .ZN(n8672)
         );
  OAI211_X1 U9970 ( .C1(n8675), .C2(n8674), .A(n8673), .B(n8672), .ZN(n8718)
         );
  MUX2_X1 U9971 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8718), .S(n8676), .Z(
        P2_U3531) );
  MUX2_X1 U9972 ( .A(n8677), .B(P2_REG0_REG_31__SCAN_IN), .S(n9758), .Z(n8678)
         );
  AOI21_X1 U9973 ( .B1(n8714), .B2(n8679), .A(n8678), .ZN(n8680) );
  INV_X1 U9974 ( .A(n8680), .ZN(P2_U3519) );
  INV_X1 U9975 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8682) );
  MUX2_X1 U9976 ( .A(n8682), .B(n8681), .S(n9759), .Z(n8683) );
  OAI21_X1 U9977 ( .B1(n8364), .B2(n8711), .A(n8683), .ZN(P2_U3518) );
  MUX2_X1 U9978 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8684), .S(n9759), .Z(
        P2_U3515) );
  MUX2_X1 U9979 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8685), .S(n9759), .Z(
        P2_U3514) );
  MUX2_X1 U9980 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8686), .S(n9759), .Z(
        P2_U3513) );
  MUX2_X1 U9981 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8687), .S(n9759), .Z(
        P2_U3512) );
  MUX2_X1 U9982 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8688), .S(n9759), .Z(
        P2_U3511) );
  INV_X1 U9983 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8690) );
  MUX2_X1 U9984 ( .A(n8690), .B(n8689), .S(n9759), .Z(n8691) );
  OAI21_X1 U9985 ( .B1(n8692), .B2(n8711), .A(n8691), .ZN(P2_U3510) );
  INV_X1 U9986 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8694) );
  MUX2_X1 U9987 ( .A(n8694), .B(n8693), .S(n9759), .Z(n8695) );
  OAI21_X1 U9988 ( .B1(n8696), .B2(n8711), .A(n8695), .ZN(P2_U3509) );
  INV_X1 U9989 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8698) );
  MUX2_X1 U9990 ( .A(n8698), .B(n8697), .S(n9759), .Z(n8699) );
  OAI21_X1 U9991 ( .B1(n4447), .B2(n8711), .A(n8699), .ZN(P2_U3508) );
  INV_X1 U9992 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8701) );
  MUX2_X1 U9993 ( .A(n8701), .B(n8700), .S(n9759), .Z(n8702) );
  OAI21_X1 U9994 ( .B1(n8703), .B2(n8711), .A(n8702), .ZN(P2_U3507) );
  INV_X1 U9995 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8705) );
  MUX2_X1 U9996 ( .A(n8705), .B(n8704), .S(n9759), .Z(n8706) );
  OAI21_X1 U9997 ( .B1(n8707), .B2(n8711), .A(n8706), .ZN(P2_U3505) );
  INV_X1 U9998 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8709) );
  MUX2_X1 U9999 ( .A(n8709), .B(n8708), .S(n9759), .Z(n8710) );
  OAI21_X1 U10000 ( .B1(n5201), .B2(n8711), .A(n8710), .ZN(P2_U3502) );
  INV_X1 U10001 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8713) );
  MUX2_X1 U10002 ( .A(n8713), .B(n8712), .S(n9759), .Z(n8717) );
  NAND2_X1 U10003 ( .A1(n8715), .A2(n8714), .ZN(n8716) );
  NAND2_X1 U10004 ( .A1(n8717), .A2(n8716), .ZN(P2_U3499) );
  MUX2_X1 U10005 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8718), .S(n9759), .Z(
        P2_U3484) );
  NAND3_X1 U10006 ( .A1(n9804), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8719) );
  OAI22_X1 U10007 ( .A1(n4827), .A2(n8719), .B1(n6440), .B2(n4267), .ZN(n8720)
         );
  AOI21_X1 U10008 ( .B1(n7897), .B2(n8721), .A(n8720), .ZN(n8722) );
  INV_X1 U10009 ( .A(n8722), .ZN(P2_U3327) );
  MUX2_X1 U10010 ( .A(n8723), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10011 ( .A(n8725), .B(n8724), .ZN(n8726) );
  XNOR2_X1 U10012 ( .A(n8727), .B(n8726), .ZN(n8734) );
  INV_X1 U10013 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8728) );
  NOR2_X1 U10014 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8728), .ZN(n9569) );
  AOI21_X1 U10015 ( .B1(n8848), .B2(n8873), .A(n9569), .ZN(n8731) );
  NAND2_X1 U10016 ( .A1(n8861), .A2(n8729), .ZN(n8730) );
  OAI211_X1 U10017 ( .C1(n8780), .C2(n8850), .A(n8731), .B(n8730), .ZN(n8732)
         );
  AOI21_X1 U10018 ( .B1(n9322), .B2(n8866), .A(n8732), .ZN(n8733) );
  OAI21_X1 U10019 ( .B1(n8734), .B2(n8868), .A(n8733), .ZN(P1_U3213) );
  NAND2_X1 U10020 ( .A1(n8736), .A2(n8735), .ZN(n8738) );
  XNOR2_X1 U10021 ( .A(n8738), .B(n8737), .ZN(n8743) );
  AOI22_X1 U10022 ( .A1(n8860), .A2(n8969), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8740) );
  NAND2_X1 U10023 ( .A1(n8861), .A2(n9101), .ZN(n8739) );
  OAI211_X1 U10024 ( .C1(n9108), .C2(n8864), .A(n8740), .B(n8739), .ZN(n8741)
         );
  AOI21_X1 U10025 ( .B1(n9273), .B2(n8866), .A(n8741), .ZN(n8742) );
  OAI21_X1 U10026 ( .B1(n8743), .B2(n8868), .A(n8742), .ZN(P1_U3214) );
  INV_X1 U10027 ( .A(n8745), .ZN(n8746) );
  AOI21_X1 U10028 ( .B1(n8747), .B2(n8744), .A(n8746), .ZN(n8753) );
  NOR2_X1 U10029 ( .A1(n8748), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8943) );
  AOI21_X1 U10030 ( .B1(n8860), .B2(n9137), .A(n8943), .ZN(n8750) );
  NAND2_X1 U10031 ( .A1(n8861), .A2(n9170), .ZN(n8749) );
  OAI211_X1 U10032 ( .C1(n9208), .C2(n8864), .A(n8750), .B(n8749), .ZN(n8751)
         );
  AOI21_X1 U10033 ( .B1(n9295), .B2(n8866), .A(n8751), .ZN(n8752) );
  OAI21_X1 U10034 ( .B1(n8753), .B2(n8868), .A(n8752), .ZN(P1_U3217) );
  XOR2_X1 U10035 ( .A(n8755), .B(n8754), .Z(n8760) );
  AOI22_X1 U10036 ( .A1(n8860), .A2(n9138), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8756) );
  OAI21_X1 U10037 ( .B1(n9166), .B2(n8864), .A(n8756), .ZN(n8758) );
  NAND2_X1 U10038 ( .A1(n9140), .A2(n9455), .ZN(n9285) );
  NOR2_X1 U10039 ( .A1(n9285), .A2(n8851), .ZN(n8757) );
  AOI211_X1 U10040 ( .C1(n9142), .C2(n8861), .A(n8758), .B(n8757), .ZN(n8759)
         );
  OAI21_X1 U10041 ( .B1(n8760), .B2(n8868), .A(n8759), .ZN(P1_U3221) );
  NAND2_X1 U10042 ( .A1(n8762), .A2(n8761), .ZN(n8764) );
  XOR2_X1 U10043 ( .A(n8764), .B(n8763), .Z(n8773) );
  INV_X1 U10044 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8765) );
  NOR2_X1 U10045 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8765), .ZN(n9544) );
  AOI21_X1 U10046 ( .B1(n8848), .B2(n8875), .A(n9544), .ZN(n8768) );
  NAND2_X1 U10047 ( .A1(n8861), .A2(n8766), .ZN(n8767) );
  OAI211_X1 U10048 ( .C1(n8769), .C2(n8850), .A(n8768), .B(n8767), .ZN(n8770)
         );
  AOI21_X1 U10049 ( .B1(n8866), .B2(n8771), .A(n8770), .ZN(n8772) );
  OAI21_X1 U10050 ( .B1(n8773), .B2(n8868), .A(n8772), .ZN(P1_U3222) );
  OAI21_X1 U10051 ( .B1(n8776), .B2(n8775), .A(n8774), .ZN(n8777) );
  NAND2_X1 U10052 ( .A1(n8777), .A2(n8806), .ZN(n8784) );
  INV_X1 U10053 ( .A(n9190), .ZN(n8959) );
  NOR2_X1 U10054 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8778), .ZN(n9592) );
  AOI21_X1 U10055 ( .B1(n8860), .B2(n8959), .A(n9592), .ZN(n8779) );
  OAI21_X1 U10056 ( .B1(n8780), .B2(n8864), .A(n8779), .ZN(n8781) );
  AOI21_X1 U10057 ( .B1(n8782), .B2(n8861), .A(n8781), .ZN(n8783) );
  OAI211_X1 U10058 ( .C1(n8785), .C2(n8813), .A(n8784), .B(n8783), .ZN(
        P1_U3224) );
  OAI21_X1 U10059 ( .B1(n8788), .B2(n8786), .A(n8787), .ZN(n8789) );
  NAND2_X1 U10060 ( .A1(n8789), .A2(n8806), .ZN(n8793) );
  INV_X1 U10061 ( .A(n9208), .ZN(n8960) );
  INV_X1 U10062 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9898) );
  NOR2_X1 U10063 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9898), .ZN(n9604) );
  AOI21_X1 U10064 ( .B1(n8860), .B2(n8960), .A(n9604), .ZN(n8790) );
  OAI21_X1 U10065 ( .B1(n9220), .B2(n8864), .A(n8790), .ZN(n8791) );
  AOI21_X1 U10066 ( .B1(n9211), .B2(n8861), .A(n8791), .ZN(n8792) );
  OAI211_X1 U10067 ( .C1(n9214), .C2(n8813), .A(n8793), .B(n8792), .ZN(
        P1_U3226) );
  XNOR2_X1 U10068 ( .A(n8795), .B(n8794), .ZN(n8796) );
  NAND2_X1 U10069 ( .A1(n8796), .A2(n8806), .ZN(n8801) );
  OAI22_X1 U10070 ( .A1(n8850), .A2(n9088), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8797), .ZN(n8799) );
  NOR2_X1 U10071 ( .A1(n8864), .A2(n9089), .ZN(n8798) );
  AOI211_X1 U10072 ( .C1(n9092), .C2(n8861), .A(n8799), .B(n8798), .ZN(n8800)
         );
  OAI211_X1 U10073 ( .C1(n8966), .C2(n8813), .A(n8801), .B(n8800), .ZN(
        P1_U3227) );
  NOR2_X1 U10074 ( .A1(n8802), .A2(n4611), .ZN(n8808) );
  AOI21_X1 U10075 ( .B1(n8805), .B2(n8804), .A(n8803), .ZN(n8807) );
  OAI21_X1 U10076 ( .B1(n8808), .B2(n8807), .A(n8806), .ZN(n8812) );
  AOI22_X1 U10077 ( .A1(n8860), .A2(n9124), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8809) );
  OAI21_X1 U10078 ( .B1(n9153), .B2(n8864), .A(n8809), .ZN(n8810) );
  AOI21_X1 U10079 ( .B1(n9155), .B2(n8861), .A(n8810), .ZN(n8811) );
  OAI211_X1 U10080 ( .C1(n8961), .C2(n8813), .A(n8812), .B(n8811), .ZN(
        P1_U3231) );
  XNOR2_X1 U10081 ( .A(n8815), .B(n8814), .ZN(n8816) );
  XNOR2_X1 U10082 ( .A(n8817), .B(n8816), .ZN(n8824) );
  AND2_X1 U10083 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9556) );
  AOI21_X1 U10084 ( .B1(n8848), .B2(n8874), .A(n9556), .ZN(n8820) );
  NAND2_X1 U10085 ( .A1(n8861), .A2(n8818), .ZN(n8819) );
  OAI211_X1 U10086 ( .C1(n9412), .C2(n8850), .A(n8820), .B(n8819), .ZN(n8821)
         );
  AOI21_X1 U10087 ( .B1(n8822), .B2(n8866), .A(n8821), .ZN(n8823) );
  OAI21_X1 U10088 ( .B1(n8824), .B2(n8868), .A(n8823), .ZN(P1_U3232) );
  NAND2_X1 U10089 ( .A1(n8826), .A2(n8825), .ZN(n8828) );
  XNOR2_X1 U10090 ( .A(n8828), .B(n8827), .ZN(n8833) );
  AOI22_X1 U10091 ( .A1(n8860), .A2(n9123), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8830) );
  NAND2_X1 U10092 ( .A1(n8861), .A2(n9118), .ZN(n8829) );
  OAI211_X1 U10093 ( .C1(n9154), .C2(n8864), .A(n8830), .B(n8829), .ZN(n8831)
         );
  AOI21_X1 U10094 ( .B1(n9278), .B2(n8866), .A(n8831), .ZN(n8832) );
  OAI21_X1 U10095 ( .B1(n8833), .B2(n8868), .A(n8832), .ZN(P1_U3233) );
  INV_X1 U10096 ( .A(n8834), .ZN(n8835) );
  AOI21_X1 U10097 ( .B1(n8848), .B2(n8876), .A(n8835), .ZN(n8837) );
  NAND2_X1 U10098 ( .A1(n8861), .A2(n9440), .ZN(n8836) );
  OAI211_X1 U10099 ( .C1(n9436), .C2(n8850), .A(n8837), .B(n8836), .ZN(n8842)
         );
  XNOR2_X1 U10100 ( .A(n8839), .B(n8838), .ZN(n8840) );
  NOR2_X1 U10101 ( .A1(n8840), .A2(n8868), .ZN(n8841) );
  AOI211_X1 U10102 ( .C1(n8866), .C2(n9442), .A(n8842), .B(n8841), .ZN(n8843)
         );
  INV_X1 U10103 ( .A(n8843), .ZN(P1_U3234) );
  NAND2_X1 U10104 ( .A1(n8845), .A2(n8844), .ZN(n8846) );
  XOR2_X1 U10105 ( .A(n8847), .B(n8846), .Z(n8855) );
  NAND2_X1 U10106 ( .A1(n8848), .A2(n8959), .ZN(n8849) );
  NAND2_X1 U10107 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9612) );
  OAI211_X1 U10108 ( .C1(n9153), .C2(n8850), .A(n8849), .B(n9612), .ZN(n8853)
         );
  NAND2_X1 U10109 ( .A1(n7567), .A2(n9455), .ZN(n9300) );
  NOR2_X1 U10110 ( .A1(n9300), .A2(n8851), .ZN(n8852) );
  AOI211_X1 U10111 ( .C1(n9196), .C2(n8861), .A(n8853), .B(n8852), .ZN(n8854)
         );
  OAI21_X1 U10112 ( .B1(n8855), .B2(n8868), .A(n8854), .ZN(P1_U3236) );
  XOR2_X1 U10113 ( .A(n8857), .B(n8856), .Z(n8858) );
  XNOR2_X1 U10114 ( .A(n8859), .B(n8858), .ZN(n8869) );
  INV_X1 U10115 ( .A(n9220), .ZN(n8955) );
  AND2_X1 U10116 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9581) );
  AOI21_X1 U10117 ( .B1(n8860), .B2(n8955), .A(n9581), .ZN(n8863) );
  NAND2_X1 U10118 ( .A1(n8861), .A2(n9230), .ZN(n8862) );
  OAI211_X1 U10119 ( .C1(n9412), .C2(n8864), .A(n8863), .B(n8862), .ZN(n8865)
         );
  AOI21_X1 U10120 ( .B1(n9315), .B2(n8866), .A(n8865), .ZN(n8867) );
  OAI21_X1 U10121 ( .B1(n8869), .B2(n8868), .A(n8867), .ZN(P1_U3239) );
  MUX2_X1 U10122 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n4397), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10123 ( .A(n9027), .B(P1_DATAO_REG_29__SCAN_IN), .S(n8870), .Z(
        P1_U3584) );
  MUX2_X1 U10124 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n8975), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10125 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n8973), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10126 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n8969), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10127 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9123), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10128 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9138), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10129 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9124), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10130 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9137), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10131 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9187), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10132 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n8960), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10133 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n8959), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10134 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n8955), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10135 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8871), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10136 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8872), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10137 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8873), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10138 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8874), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10139 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8875), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10140 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8876), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10141 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8877), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10142 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8878), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10143 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8879), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10144 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8880), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10145 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8881), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10146 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8882), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10147 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8883), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10148 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8884), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10149 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n8885), .S(P1_U4006), .Z(
        P1_U3556) );
  NAND3_X1 U10150 ( .A1(n9607), .A2(n8901), .A3(P1_REG1_REG_8__SCAN_IN), .ZN(
        n8887) );
  OR3_X1 U10151 ( .A1(n8938), .A2(n6187), .A3(n8892), .ZN(n8886) );
  NAND3_X1 U10152 ( .A1(n8888), .A2(n8887), .A3(n8886), .ZN(n8890) );
  AOI22_X1 U10153 ( .A1(n8890), .A2(n8889), .B1(n9495), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n8905) );
  INV_X1 U10154 ( .A(n8891), .ZN(n8904) );
  INV_X1 U10155 ( .A(n8892), .ZN(n8897) );
  INV_X1 U10156 ( .A(n8893), .ZN(n8894) );
  OAI211_X1 U10157 ( .C1(n8897), .C2(n8896), .A(n8895), .B(n8894), .ZN(n8903)
         );
  INV_X1 U10158 ( .A(n8898), .ZN(n8899) );
  OAI211_X1 U10159 ( .C1(n8901), .C2(n8900), .A(n9607), .B(n8899), .ZN(n8902)
         );
  NAND4_X1 U10160 ( .A1(n8905), .A2(n8904), .A3(n8903), .A4(n8902), .ZN(
        P1_U3249) );
  NAND2_X1 U10161 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9545), .ZN(n8906) );
  OAI21_X1 U10162 ( .B1(n9545), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8906), .ZN(
        n9541) );
  OAI21_X1 U10163 ( .B1(n8908), .B2(P1_REG2_REG_11__SCAN_IN), .A(n8907), .ZN(
        n9542) );
  NAND2_X1 U10164 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9557), .ZN(n8909) );
  OAI21_X1 U10165 ( .B1(n9557), .B2(P1_REG2_REG_13__SCAN_IN), .A(n8909), .ZN(
        n9553) );
  NOR2_X1 U10166 ( .A1(n9554), .A2(n9553), .ZN(n9552) );
  NOR2_X1 U10167 ( .A1(n8910), .A2(n8924), .ZN(n8911) );
  INV_X1 U10168 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9566) );
  NOR2_X1 U10169 ( .A1(n9566), .A2(n9567), .ZN(n9565) );
  NOR2_X1 U10170 ( .A1(n8912), .A2(n8926), .ZN(n8913) );
  INV_X1 U10171 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9578) );
  XNOR2_X1 U10172 ( .A(n8912), .B(n8926), .ZN(n9579) );
  NOR2_X1 U10173 ( .A1(n9578), .A2(n9579), .ZN(n9577) );
  NAND2_X1 U10174 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9593), .ZN(n8914) );
  OAI21_X1 U10175 ( .B1(n9593), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8914), .ZN(
        n9589) );
  NOR2_X1 U10176 ( .A1(n9590), .A2(n9589), .ZN(n9588) );
  NAND2_X1 U10177 ( .A1(n9605), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8915) );
  OAI21_X1 U10178 ( .B1(n9605), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8915), .ZN(
        n9601) );
  NOR2_X1 U10179 ( .A1(n9602), .A2(n9601), .ZN(n9600) );
  AOI21_X1 U10180 ( .B1(n9605), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9600), .ZN(
        n9616) );
  INV_X1 U10181 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8917) );
  NOR2_X1 U10182 ( .A1(n9620), .A2(n8917), .ZN(n8916) );
  AOI21_X1 U10183 ( .B1(n9620), .B2(n8917), .A(n8916), .ZN(n9615) );
  AOI21_X1 U10184 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9620), .A(n9614), .ZN(
        n8918) );
  XNOR2_X1 U10185 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8918), .ZN(n8939) );
  INV_X1 U10186 ( .A(n8939), .ZN(n8935) );
  INV_X1 U10187 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8932) );
  XNOR2_X1 U10188 ( .A(n9620), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9623) );
  INV_X1 U10189 ( .A(n9605), .ZN(n8930) );
  INV_X1 U10190 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8929) );
  XOR2_X1 U10191 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9605), .Z(n9609) );
  INV_X1 U10192 ( .A(n9593), .ZN(n8928) );
  INV_X1 U10193 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9863) );
  XOR2_X1 U10194 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9593), .Z(n9595) );
  INV_X1 U10195 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8923) );
  INV_X1 U10196 ( .A(n9557), .ZN(n8922) );
  INV_X1 U10197 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9462) );
  INV_X1 U10198 ( .A(n9545), .ZN(n8921) );
  INV_X1 U10199 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9468) );
  AOI21_X1 U10200 ( .B1(n8920), .B2(n9474), .A(n8919), .ZN(n9548) );
  MUX2_X1 U10201 ( .A(n9468), .B(P1_REG1_REG_12__SCAN_IN), .S(n9545), .Z(n9547) );
  NOR2_X1 U10202 ( .A1(n9548), .A2(n9547), .ZN(n9546) );
  AOI21_X1 U10203 ( .B1(n8921), .B2(n9468), .A(n9546), .ZN(n9559) );
  MUX2_X1 U10204 ( .A(n9462), .B(P1_REG1_REG_13__SCAN_IN), .S(n9557), .Z(n9560) );
  NOR2_X1 U10205 ( .A1(n9559), .A2(n9560), .ZN(n9558) );
  AOI21_X1 U10206 ( .B1(n8922), .B2(n9462), .A(n9558), .ZN(n9572) );
  MUX2_X1 U10207 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n8923), .S(n8924), .Z(n9573) );
  NOR2_X1 U10208 ( .A1(n9572), .A2(n9573), .ZN(n9571) );
  AOI21_X1 U10209 ( .B1(n8924), .B2(n8923), .A(n9571), .ZN(n8925) );
  NAND2_X1 U10210 ( .A1(n9582), .A2(n8925), .ZN(n8927) );
  XNOR2_X1 U10211 ( .A(n8926), .B(n8925), .ZN(n9584) );
  NAND2_X1 U10212 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9584), .ZN(n9583) );
  NAND2_X1 U10213 ( .A1(n8927), .A2(n9583), .ZN(n9596) );
  NAND2_X1 U10214 ( .A1(n9595), .A2(n9596), .ZN(n9594) );
  OAI21_X1 U10215 ( .B1(n8928), .B2(n9863), .A(n9594), .ZN(n9608) );
  NAND2_X1 U10216 ( .A1(n9609), .A2(n9608), .ZN(n9606) );
  OAI21_X1 U10217 ( .B1(n8930), .B2(n8929), .A(n9606), .ZN(n9622) );
  NOR2_X1 U10218 ( .A1(n9623), .A2(n9622), .ZN(n9621) );
  AOI21_X1 U10219 ( .B1(n8932), .B2(n8931), .A(n9621), .ZN(n8934) );
  INV_X1 U10220 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8933) );
  XOR2_X1 U10221 ( .A(n8934), .B(n8933), .Z(n8936) );
  OAI22_X1 U10222 ( .A1(n8935), .A2(n9613), .B1(n8936), .B2(n9625), .ZN(n8941)
         );
  AOI21_X1 U10223 ( .B1(n8936), .B2(n9607), .A(n9619), .ZN(n8937) );
  OAI21_X1 U10224 ( .B1(n8939), .B2(n8938), .A(n8937), .ZN(n8940) );
  INV_X1 U10225 ( .A(n8944), .ZN(P1_U3260) );
  INV_X1 U10226 ( .A(n9295), .ZN(n9173) );
  NAND2_X1 U10227 ( .A1(n4398), .A2(n9010), .ZN(n8945) );
  XNOR2_X1 U10228 ( .A(n9237), .B(n8945), .ZN(n9239) );
  NAND2_X1 U10229 ( .A1(n9491), .A2(P1_B_REG_SCAN_IN), .ZN(n8946) );
  NAND2_X1 U10230 ( .A1(n9188), .A2(n8946), .ZN(n9006) );
  NOR2_X1 U10231 ( .A1(n9006), .A2(n8947), .ZN(n9453) );
  INV_X1 U10232 ( .A(n9453), .ZN(n8948) );
  NOR2_X1 U10233 ( .A1(n8948), .A2(n9451), .ZN(n8953) );
  NOR2_X1 U10234 ( .A1(n8949), .A2(n9418), .ZN(n8950) );
  AOI211_X1 U10235 ( .C1(n9451), .C2(P1_REG2_REG_31__SCAN_IN), .A(n8953), .B(
        n8950), .ZN(n8951) );
  OAI21_X1 U10236 ( .B1(n9239), .B2(n9200), .A(n8951), .ZN(P1_U3261) );
  NOR2_X1 U10237 ( .A1(n4398), .A2(n9418), .ZN(n8952) );
  AOI211_X1 U10238 ( .C1(n9451), .C2(P1_REG2_REG_30__SCAN_IN), .A(n8953), .B(
        n8952), .ZN(n8954) );
  OAI21_X1 U10239 ( .B1(n9200), .B2(n9452), .A(n8954), .ZN(P1_U3262) );
  INV_X1 U10240 ( .A(n9247), .ZN(n9024) );
  NAND2_X1 U10241 ( .A1(n9116), .A2(n4792), .ZN(n8963) );
  AOI21_X1 U10242 ( .B1(n9089), .B2(n9103), .A(n9098), .ZN(n8965) );
  NAND2_X1 U10243 ( .A1(n8967), .A2(n8969), .ZN(n8968) );
  NAND2_X1 U10244 ( .A1(n9082), .A2(n8968), .ZN(n8971) );
  NAND2_X1 U10245 ( .A1(n9055), .A2(n9073), .ZN(n8974) );
  XNOR2_X1 U10246 ( .A(n8976), .B(n9002), .ZN(n9240) );
  INV_X1 U10247 ( .A(n9240), .ZN(n9017) );
  INV_X1 U10248 ( .A(n8982), .ZN(n8979) );
  AND2_X1 U10249 ( .A1(n8977), .A2(n9179), .ZN(n8978) );
  AND2_X1 U10250 ( .A1(n9177), .A2(n8982), .ZN(n8983) );
  NAND2_X1 U10251 ( .A1(n9163), .A2(n9164), .ZN(n8986) );
  NOR2_X1 U10252 ( .A1(n9131), .A2(n9132), .ZN(n8988) );
  NAND2_X1 U10253 ( .A1(n9111), .A2(n8992), .ZN(n9085) );
  INV_X1 U10254 ( .A(n9085), .ZN(n8994) );
  INV_X1 U10255 ( .A(n9086), .ZN(n8993) );
  INV_X1 U10256 ( .A(n8997), .ZN(n8998) );
  INV_X1 U10257 ( .A(n8999), .ZN(n9000) );
  XNOR2_X1 U10258 ( .A(n9003), .B(n9002), .ZN(n9004) );
  NAND2_X1 U10259 ( .A1(n9004), .A2(n9414), .ZN(n9009) );
  INV_X1 U10260 ( .A(n9007), .ZN(n9008) );
  AOI211_X1 U10261 ( .C1(n9242), .C2(n9020), .A(n9679), .B(n9010), .ZN(n9244)
         );
  NAND2_X1 U10262 ( .A1(n9244), .A2(n9210), .ZN(n9013) );
  AOI22_X1 U10263 ( .A1(n9451), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9011), .B2(
        n9439), .ZN(n9012) );
  OAI211_X1 U10264 ( .C1(n9014), .C2(n9418), .A(n9013), .B(n9012), .ZN(n9015)
         );
  AOI21_X1 U10265 ( .B1(n9241), .B2(n9424), .A(n9015), .ZN(n9016) );
  OAI21_X1 U10266 ( .B1(n9017), .B2(n9217), .A(n9016), .ZN(P1_U3355) );
  INV_X1 U10267 ( .A(n9020), .ZN(n9021) );
  AOI21_X1 U10268 ( .B1(n9247), .B2(n9035), .A(n9021), .ZN(n9248) );
  AOI22_X1 U10269 ( .A1(n9451), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9022), .B2(
        n9439), .ZN(n9023) );
  OAI21_X1 U10270 ( .B1(n9024), .B2(n9418), .A(n9023), .ZN(n9031) );
  NAND2_X1 U10271 ( .A1(n9027), .A2(n9188), .ZN(n9028) );
  AOI211_X1 U10272 ( .C1(n9446), .C2(n9248), .A(n9031), .B(n9030), .ZN(n9032)
         );
  OAI21_X1 U10273 ( .B1(n9251), .B2(n9217), .A(n9032), .ZN(P1_U3263) );
  XNOR2_X1 U10274 ( .A(n9034), .B(n9033), .ZN(n9256) );
  INV_X1 U10275 ( .A(n9051), .ZN(n9037) );
  INV_X1 U10276 ( .A(n9035), .ZN(n9036) );
  AOI21_X1 U10277 ( .B1(n9252), .B2(n9037), .A(n9036), .ZN(n9253) );
  AOI22_X1 U10278 ( .A1(n9451), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9038), .B2(
        n9439), .ZN(n9039) );
  OAI21_X1 U10279 ( .B1(n9040), .B2(n9418), .A(n9039), .ZN(n9048) );
  AOI211_X1 U10280 ( .C1(n9043), .C2(n9042), .A(n9433), .B(n9041), .ZN(n9046)
         );
  OAI22_X1 U10281 ( .A1(n9437), .A2(n9044), .B1(n9073), .B2(n9435), .ZN(n9045)
         );
  NOR2_X1 U10282 ( .A1(n9046), .A2(n9045), .ZN(n9255) );
  NOR2_X1 U10283 ( .A1(n9255), .A2(n9451), .ZN(n9047) );
  AOI211_X1 U10284 ( .C1(n9253), .C2(n9446), .A(n9048), .B(n9047), .ZN(n9049)
         );
  OAI21_X1 U10285 ( .B1(n9256), .B2(n9217), .A(n9049), .ZN(P1_U3264) );
  XNOR2_X1 U10286 ( .A(n9050), .B(n9056), .ZN(n9261) );
  INV_X1 U10287 ( .A(n9072), .ZN(n9052) );
  AOI21_X1 U10288 ( .B1(n9257), .B2(n9052), .A(n9051), .ZN(n9258) );
  AOI22_X1 U10289 ( .A1(n9451), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9053), .B2(
        n9439), .ZN(n9054) );
  OAI21_X1 U10290 ( .B1(n9055), .B2(n9418), .A(n9054), .ZN(n9062) );
  AOI211_X1 U10291 ( .C1(n9057), .C2(n9056), .A(n9433), .B(n4310), .ZN(n9060)
         );
  OAI22_X1 U10292 ( .A1(n9437), .A2(n9058), .B1(n9088), .B2(n9435), .ZN(n9059)
         );
  NOR2_X1 U10293 ( .A1(n9060), .A2(n9059), .ZN(n9260) );
  NOR2_X1 U10294 ( .A1(n9260), .A2(n9451), .ZN(n9061) );
  AOI211_X1 U10295 ( .C1(n9446), .C2(n9258), .A(n9062), .B(n9061), .ZN(n9063)
         );
  OAI21_X1 U10296 ( .B1(n9261), .B2(n9217), .A(n9063), .ZN(P1_U3265) );
  XNOR2_X1 U10297 ( .A(n9064), .B(n9065), .ZN(n9267) );
  INV_X1 U10298 ( .A(n9267), .ZN(n9081) );
  AOI22_X1 U10299 ( .A1(n9069), .A2(n9441), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9451), .ZN(n9080) );
  NAND2_X1 U10300 ( .A1(n9066), .A2(n9065), .ZN(n9067) );
  NAND2_X1 U10301 ( .A1(n9067), .A2(n9414), .ZN(n9068) );
  NOR2_X1 U10302 ( .A1(n4324), .A2(n9068), .ZN(n9266) );
  NAND2_X1 U10303 ( .A1(n9069), .A2(n9090), .ZN(n9070) );
  NAND2_X1 U10304 ( .A1(n9070), .A2(n9661), .ZN(n9071) );
  OR2_X1 U10305 ( .A1(n9072), .A2(n9071), .ZN(n9264) );
  OR2_X1 U10306 ( .A1(n9437), .A2(n9073), .ZN(n9075) );
  OR2_X1 U10307 ( .A1(n9109), .A2(n9435), .ZN(n9074) );
  AND2_X1 U10308 ( .A1(n9075), .A2(n9074), .ZN(n9263) );
  NAND2_X1 U10309 ( .A1(n9439), .A2(n9076), .ZN(n9077) );
  OAI211_X1 U10310 ( .C1(n9264), .C2(n9157), .A(n9263), .B(n9077), .ZN(n9078)
         );
  OAI21_X1 U10311 ( .B1(n9266), .B2(n9078), .A(n9424), .ZN(n9079) );
  OAI211_X1 U10312 ( .C1(n9081), .C2(n9217), .A(n9080), .B(n9079), .ZN(
        P1_U3266) );
  XOR2_X1 U10313 ( .A(n9086), .B(n9082), .Z(n9272) );
  AOI22_X1 U10314 ( .A1(n8967), .A2(n9441), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9451), .ZN(n9097) );
  INV_X1 U10315 ( .A(n9083), .ZN(n9084) );
  AOI21_X1 U10316 ( .B1(n9086), .B2(n9085), .A(n9084), .ZN(n9087) );
  OAI222_X1 U10317 ( .A1(n9435), .A2(n9089), .B1(n9437), .B2(n9088), .C1(n9433), .C2(n9087), .ZN(n9269) );
  INV_X1 U10318 ( .A(n9090), .ZN(n9091) );
  AOI211_X1 U10319 ( .C1(n8967), .C2(n9099), .A(n9679), .B(n9091), .ZN(n9270)
         );
  INV_X1 U10320 ( .A(n9270), .ZN(n9094) );
  INV_X1 U10321 ( .A(n9092), .ZN(n9093) );
  OAI22_X1 U10322 ( .A1(n9094), .A2(n9157), .B1(n9419), .B2(n9093), .ZN(n9095)
         );
  OAI21_X1 U10323 ( .B1(n9269), .B2(n9095), .A(n9424), .ZN(n9096) );
  OAI211_X1 U10324 ( .C1(n9272), .C2(n9217), .A(n9097), .B(n9096), .ZN(
        P1_U3267) );
  XNOR2_X1 U10325 ( .A(n9098), .B(n9105), .ZN(n9277) );
  INV_X1 U10326 ( .A(n9117), .ZN(n9100) );
  AOI21_X1 U10327 ( .B1(n9273), .B2(n9100), .A(n4553), .ZN(n9274) );
  AOI22_X1 U10328 ( .A1(n9451), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9101), .B2(
        n9439), .ZN(n9102) );
  OAI21_X1 U10329 ( .B1(n9103), .B2(n9418), .A(n9102), .ZN(n9114) );
  INV_X1 U10330 ( .A(n9104), .ZN(n9107) );
  INV_X1 U10331 ( .A(n9105), .ZN(n9106) );
  AOI21_X1 U10332 ( .B1(n9107), .B2(n9106), .A(n9433), .ZN(n9112) );
  OAI22_X1 U10333 ( .A1(n9437), .A2(n9109), .B1(n9108), .B2(n9435), .ZN(n9110)
         );
  AOI21_X1 U10334 ( .B1(n9112), .B2(n9111), .A(n9110), .ZN(n9276) );
  NOR2_X1 U10335 ( .A1(n9276), .A2(n9451), .ZN(n9113) );
  AOI211_X1 U10336 ( .C1(n9274), .C2(n9446), .A(n9114), .B(n9113), .ZN(n9115)
         );
  OAI21_X1 U10337 ( .B1(n9277), .B2(n9217), .A(n9115), .ZN(P1_U3268) );
  XNOR2_X1 U10338 ( .A(n9116), .B(n9121), .ZN(n9282) );
  AOI21_X1 U10339 ( .B1(n9278), .B2(n4288), .A(n9117), .ZN(n9279) );
  AOI22_X1 U10340 ( .A1(n9451), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9118), .B2(
        n9439), .ZN(n9119) );
  OAI21_X1 U10341 ( .B1(n9120), .B2(n9418), .A(n9119), .ZN(n9127) );
  XNOR2_X1 U10342 ( .A(n9122), .B(n9121), .ZN(n9125) );
  AOI222_X1 U10343 ( .A1(n9414), .A2(n9125), .B1(n9124), .B2(n9136), .C1(n9123), .C2(n9188), .ZN(n9281) );
  NOR2_X1 U10344 ( .A1(n9281), .A2(n9451), .ZN(n9126) );
  AOI211_X1 U10345 ( .C1(n9279), .C2(n9446), .A(n9127), .B(n9126), .ZN(n9128)
         );
  OAI21_X1 U10346 ( .B1(n9282), .B2(n9217), .A(n9128), .ZN(P1_U3269) );
  XOR2_X1 U10347 ( .A(n9129), .B(n9131), .Z(n9283) );
  INV_X1 U10348 ( .A(n9283), .ZN(n9148) );
  AOI22_X1 U10349 ( .A1(n9140), .A2(n9441), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9451), .ZN(n9147) );
  INV_X1 U10350 ( .A(n9130), .ZN(n9133) );
  OAI21_X1 U10351 ( .B1(n9133), .B2(n9132), .A(n9131), .ZN(n9135) );
  NAND2_X1 U10352 ( .A1(n9135), .A2(n9134), .ZN(n9139) );
  AOI222_X1 U10353 ( .A1(n9414), .A2(n9139), .B1(n9138), .B2(n9188), .C1(n9137), .C2(n9136), .ZN(n9286) );
  INV_X1 U10354 ( .A(n9286), .ZN(n9145) );
  INV_X1 U10355 ( .A(n9140), .ZN(n9141) );
  OAI211_X1 U10356 ( .C1(n9141), .C2(n4333), .A(n4288), .B(n9661), .ZN(n9284)
         );
  INV_X1 U10357 ( .A(n9142), .ZN(n9143) );
  OAI22_X1 U10358 ( .A1(n9284), .A2(n9157), .B1(n9419), .B2(n9143), .ZN(n9144)
         );
  OAI21_X1 U10359 ( .B1(n9145), .B2(n9144), .A(n9424), .ZN(n9146) );
  OAI211_X1 U10360 ( .C1(n9148), .C2(n9217), .A(n9147), .B(n9146), .ZN(
        P1_U3270) );
  XNOR2_X1 U10361 ( .A(n9149), .B(n9150), .ZN(n9292) );
  AOI22_X1 U10362 ( .A1(n9290), .A2(n9441), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n9451), .ZN(n9161) );
  XNOR2_X1 U10363 ( .A(n9151), .B(n9150), .ZN(n9152) );
  OAI222_X1 U10364 ( .A1(n9437), .A2(n9154), .B1(n9435), .B2(n9153), .C1(n9152), .C2(n9433), .ZN(n9288) );
  AOI211_X1 U10365 ( .C1(n9290), .C2(n9167), .A(n9679), .B(n4333), .ZN(n9289)
         );
  INV_X1 U10366 ( .A(n9289), .ZN(n9158) );
  INV_X1 U10367 ( .A(n9155), .ZN(n9156) );
  OAI22_X1 U10368 ( .A1(n9158), .A2(n9157), .B1(n9419), .B2(n9156), .ZN(n9159)
         );
  OAI21_X1 U10369 ( .B1(n9288), .B2(n9159), .A(n9424), .ZN(n9160) );
  OAI211_X1 U10370 ( .C1(n9292), .C2(n9217), .A(n9161), .B(n9160), .ZN(
        P1_U3271) );
  XNOR2_X1 U10371 ( .A(n9162), .B(n9164), .ZN(n9297) );
  XOR2_X1 U10372 ( .A(n9164), .B(n9163), .Z(n9165) );
  OAI222_X1 U10373 ( .A1(n9437), .A2(n9166), .B1(n9435), .B2(n9208), .C1(n9165), .C2(n9433), .ZN(n9293) );
  INV_X1 U10374 ( .A(n9195), .ZN(n9169) );
  INV_X1 U10375 ( .A(n9167), .ZN(n9168) );
  AOI211_X1 U10376 ( .C1(n9295), .C2(n9169), .A(n9679), .B(n9168), .ZN(n9294)
         );
  NAND2_X1 U10377 ( .A1(n9294), .A2(n9210), .ZN(n9172) );
  AOI22_X1 U10378 ( .A1(n9451), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9170), .B2(
        n9439), .ZN(n9171) );
  OAI211_X1 U10379 ( .C1(n9173), .C2(n9418), .A(n9172), .B(n9171), .ZN(n9174)
         );
  AOI21_X1 U10380 ( .B1(n9293), .B2(n9424), .A(n9174), .ZN(n9175) );
  OAI21_X1 U10381 ( .B1(n9297), .B2(n9217), .A(n9175), .ZN(P1_U3272) );
  AND2_X1 U10382 ( .A1(n9176), .A2(n9184), .ZN(n9298) );
  NOR3_X1 U10383 ( .A1(n9299), .A2(n9298), .A3(n9217), .ZN(n9203) );
  NAND2_X1 U10384 ( .A1(n9178), .A2(n9177), .ZN(n9180) );
  NAND2_X1 U10385 ( .A1(n9180), .A2(n9179), .ZN(n9205) );
  OR2_X1 U10386 ( .A1(n9205), .A2(n9181), .ZN(n9183) );
  NAND2_X1 U10387 ( .A1(n9183), .A2(n9182), .ZN(n9186) );
  INV_X1 U10388 ( .A(n9184), .ZN(n9185) );
  XNOR2_X1 U10389 ( .A(n9186), .B(n9185), .ZN(n9192) );
  NAND2_X1 U10390 ( .A1(n9188), .A2(n9187), .ZN(n9189) );
  OAI21_X1 U10391 ( .B1(n9190), .B2(n9435), .A(n9189), .ZN(n9191) );
  AOI21_X1 U10392 ( .B1(n9192), .B2(n9414), .A(n9191), .ZN(n9301) );
  NOR2_X1 U10393 ( .A1(n9301), .A2(n9451), .ZN(n9202) );
  NOR2_X1 U10394 ( .A1(n4332), .A2(n9193), .ZN(n9194) );
  OR2_X1 U10395 ( .A1(n9195), .A2(n9194), .ZN(n9302) );
  INV_X1 U10396 ( .A(n9196), .ZN(n9197) );
  OAI22_X1 U10397 ( .A1(n9424), .A2(n8917), .B1(n9197), .B2(n9419), .ZN(n9198)
         );
  AOI21_X1 U10398 ( .B1(n7567), .B2(n9441), .A(n9198), .ZN(n9199) );
  OAI21_X1 U10399 ( .B1(n9302), .B2(n9200), .A(n9199), .ZN(n9201) );
  OR3_X1 U10400 ( .A1(n9203), .A2(n9202), .A3(n9201), .ZN(P1_U3273) );
  XNOR2_X1 U10401 ( .A(n9204), .B(n9206), .ZN(n9309) );
  XOR2_X1 U10402 ( .A(n9206), .B(n9205), .Z(n9207) );
  OAI222_X1 U10403 ( .A1(n9437), .A2(n9208), .B1(n9435), .B2(n9220), .C1(n9207), .C2(n9433), .ZN(n9305) );
  AOI211_X1 U10404 ( .C1(n9307), .C2(n9209), .A(n9679), .B(n4332), .ZN(n9306)
         );
  NAND2_X1 U10405 ( .A1(n9306), .A2(n9210), .ZN(n9213) );
  AOI22_X1 U10406 ( .A1(n9451), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9211), .B2(
        n9439), .ZN(n9212) );
  OAI211_X1 U10407 ( .C1(n9214), .C2(n9418), .A(n9213), .B(n9212), .ZN(n9215)
         );
  AOI21_X1 U10408 ( .B1(n9305), .B2(n9424), .A(n9215), .ZN(n9216) );
  OAI21_X1 U10409 ( .B1(n9309), .B2(n9217), .A(n9216), .ZN(P1_U3274) );
  XNOR2_X1 U10410 ( .A(n9219), .B(n9218), .ZN(n9225) );
  OAI22_X1 U10411 ( .A1(n9437), .A2(n9220), .B1(n9412), .B2(n9435), .ZN(n9224)
         );
  XNOR2_X1 U10412 ( .A(n9222), .B(n9221), .ZN(n9319) );
  NOR2_X1 U10413 ( .A1(n9319), .A2(n9664), .ZN(n9223) );
  AOI211_X1 U10414 ( .C1(n9414), .C2(n9225), .A(n9224), .B(n9223), .ZN(n9318)
         );
  INV_X1 U10415 ( .A(n9226), .ZN(n9229) );
  INV_X1 U10416 ( .A(n9227), .ZN(n9228) );
  AOI21_X1 U10417 ( .B1(n9315), .B2(n9229), .A(n9228), .ZN(n9316) );
  AOI22_X1 U10418 ( .A1(n9451), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9230), .B2(
        n9439), .ZN(n9231) );
  OAI21_X1 U10419 ( .B1(n9232), .B2(n9418), .A(n9231), .ZN(n9235) );
  NOR2_X1 U10420 ( .A1(n9319), .A2(n9233), .ZN(n9234) );
  AOI211_X1 U10421 ( .C1(n9316), .C2(n9446), .A(n9235), .B(n9234), .ZN(n9236)
         );
  OAI21_X1 U10422 ( .B1(n9318), .B2(n9451), .A(n9236), .ZN(P1_U3276) );
  AOI21_X1 U10423 ( .B1(n9237), .B2(n9455), .A(n9453), .ZN(n9238) );
  OAI21_X1 U10424 ( .B1(n9239), .B2(n9679), .A(n9238), .ZN(n9326) );
  MUX2_X1 U10425 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9326), .S(n9696), .Z(
        P1_U3554) );
  NAND2_X1 U10426 ( .A1(n9240), .A2(n9681), .ZN(n9246) );
  MUX2_X1 U10427 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9327), .S(n9696), .Z(
        P1_U3552) );
  AOI22_X1 U10428 ( .A1(n9248), .A2(n9661), .B1(n9455), .B2(n9247), .ZN(n9249)
         );
  OAI211_X1 U10429 ( .C1(n9251), .C2(n9324), .A(n9250), .B(n9249), .ZN(n9328)
         );
  MUX2_X1 U10430 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9328), .S(n9696), .Z(
        P1_U3551) );
  AOI22_X1 U10431 ( .A1(n9253), .A2(n9661), .B1(n9455), .B2(n9252), .ZN(n9254)
         );
  OAI211_X1 U10432 ( .C1(n9256), .C2(n9324), .A(n9255), .B(n9254), .ZN(n9329)
         );
  MUX2_X1 U10433 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9329), .S(n9696), .Z(
        P1_U3550) );
  AOI22_X1 U10434 ( .A1(n9258), .A2(n9661), .B1(n9455), .B2(n9257), .ZN(n9259)
         );
  OAI211_X1 U10435 ( .C1(n9261), .C2(n9324), .A(n9260), .B(n9259), .ZN(n9330)
         );
  MUX2_X1 U10436 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9330), .S(n9696), .Z(
        P1_U3549) );
  NAND3_X1 U10437 ( .A1(n9264), .A2(n9263), .A3(n9262), .ZN(n9265) );
  AOI211_X1 U10438 ( .C1(n9267), .C2(n9681), .A(n9266), .B(n9265), .ZN(n9268)
         );
  INV_X1 U10439 ( .A(n9268), .ZN(n9331) );
  MUX2_X1 U10440 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9331), .S(n9696), .Z(
        P1_U3548) );
  AOI211_X1 U10441 ( .C1(n9455), .C2(n8967), .A(n9270), .B(n9269), .ZN(n9271)
         );
  OAI21_X1 U10442 ( .B1(n9272), .B2(n9324), .A(n9271), .ZN(n9332) );
  MUX2_X1 U10443 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9332), .S(n9696), .Z(
        P1_U3547) );
  AOI22_X1 U10444 ( .A1(n9274), .A2(n9661), .B1(n9455), .B2(n9273), .ZN(n9275)
         );
  OAI211_X1 U10445 ( .C1(n9277), .C2(n9324), .A(n9276), .B(n9275), .ZN(n9333)
         );
  MUX2_X1 U10446 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9333), .S(n9696), .Z(
        P1_U3546) );
  AOI22_X1 U10447 ( .A1(n9279), .A2(n9661), .B1(n9455), .B2(n9278), .ZN(n9280)
         );
  OAI211_X1 U10448 ( .C1(n9282), .C2(n9324), .A(n9281), .B(n9280), .ZN(n9334)
         );
  MUX2_X1 U10449 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9334), .S(n9696), .Z(
        P1_U3545) );
  NAND2_X1 U10450 ( .A1(n9283), .A2(n9681), .ZN(n9287) );
  NAND4_X1 U10451 ( .A1(n9287), .A2(n9286), .A3(n9285), .A4(n9284), .ZN(n9335)
         );
  MUX2_X1 U10452 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9335), .S(n9696), .Z(
        P1_U3544) );
  AOI211_X1 U10453 ( .C1(n9455), .C2(n9290), .A(n9289), .B(n9288), .ZN(n9291)
         );
  OAI21_X1 U10454 ( .B1(n9292), .B2(n9324), .A(n9291), .ZN(n9336) );
  MUX2_X1 U10455 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9336), .S(n9696), .Z(
        P1_U3543) );
  AOI211_X1 U10456 ( .C1(n9455), .C2(n9295), .A(n9294), .B(n9293), .ZN(n9296)
         );
  OAI21_X1 U10457 ( .B1(n9297), .B2(n9324), .A(n9296), .ZN(n9337) );
  MUX2_X1 U10458 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9337), .S(n9696), .Z(
        P1_U3542) );
  NOR3_X1 U10459 ( .A1(n9299), .A2(n9298), .A3(n9324), .ZN(n9304) );
  OAI211_X1 U10460 ( .C1(n9679), .C2(n9302), .A(n9301), .B(n9300), .ZN(n9303)
         );
  OR2_X1 U10461 ( .A1(n9304), .A2(n9303), .ZN(n9338) );
  MUX2_X1 U10462 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9338), .S(n9696), .Z(
        P1_U3541) );
  AOI211_X1 U10463 ( .C1(n9455), .C2(n9307), .A(n9306), .B(n9305), .ZN(n9308)
         );
  OAI21_X1 U10464 ( .B1(n9309), .B2(n9324), .A(n9308), .ZN(n9339) );
  MUX2_X1 U10465 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9339), .S(n9696), .Z(
        P1_U3540) );
  AOI211_X1 U10466 ( .C1(n9455), .C2(n9312), .A(n9311), .B(n9310), .ZN(n9313)
         );
  OAI21_X1 U10467 ( .B1(n9314), .B2(n9324), .A(n9313), .ZN(n9340) );
  MUX2_X1 U10468 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9340), .S(n9696), .Z(
        P1_U3539) );
  AOI22_X1 U10469 ( .A1(n9316), .A2(n9661), .B1(n9455), .B2(n9315), .ZN(n9317)
         );
  OAI211_X1 U10470 ( .C1(n9319), .C2(n9456), .A(n9318), .B(n9317), .ZN(n9341)
         );
  MUX2_X1 U10471 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9341), .S(n9696), .Z(
        P1_U3538) );
  AOI211_X1 U10472 ( .C1(n9455), .C2(n9322), .A(n9321), .B(n9320), .ZN(n9323)
         );
  OAI21_X1 U10473 ( .B1(n9325), .B2(n9324), .A(n9323), .ZN(n9342) );
  MUX2_X1 U10474 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9342), .S(n9696), .Z(
        P1_U3537) );
  MUX2_X1 U10475 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9326), .S(n9685), .Z(
        P1_U3522) );
  MUX2_X1 U10476 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9327), .S(n9685), .Z(
        P1_U3520) );
  MUX2_X1 U10477 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9328), .S(n9685), .Z(
        P1_U3519) );
  MUX2_X1 U10478 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9329), .S(n9685), .Z(
        P1_U3518) );
  MUX2_X1 U10479 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9330), .S(n9685), .Z(
        P1_U3517) );
  MUX2_X1 U10480 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9331), .S(n9685), .Z(
        P1_U3516) );
  MUX2_X1 U10481 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9332), .S(n9685), .Z(
        P1_U3515) );
  MUX2_X1 U10482 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9333), .S(n9685), .Z(
        P1_U3514) );
  MUX2_X1 U10483 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9334), .S(n9685), .Z(
        P1_U3513) );
  MUX2_X1 U10484 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9335), .S(n9685), .Z(
        P1_U3512) );
  MUX2_X1 U10485 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9336), .S(n9685), .Z(
        P1_U3511) );
  MUX2_X1 U10486 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9337), .S(n9685), .Z(
        P1_U3510) );
  MUX2_X1 U10487 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9338), .S(n9685), .Z(
        P1_U3508) );
  MUX2_X1 U10488 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9339), .S(n9685), .Z(
        P1_U3505) );
  MUX2_X1 U10489 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9340), .S(n9685), .Z(
        P1_U3502) );
  MUX2_X1 U10490 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9341), .S(n9685), .Z(
        P1_U3499) );
  MUX2_X1 U10491 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9342), .S(n9685), .Z(
        P1_U3496) );
  MUX2_X1 U10492 ( .A(n9343), .B(P1_D_REG_0__SCAN_IN), .S(n9635), .Z(P1_U3440)
         );
  NAND2_X1 U10493 ( .A1(n7897), .A2(n9344), .ZN(n9348) );
  NAND4_X1 U10494 ( .A1(n5636), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .A4(n9346), .ZN(n9347) );
  OAI211_X1 U10495 ( .C1(n6266), .C2(n9349), .A(n9348), .B(n9347), .ZN(
        P1_U3322) );
  OAI222_X1 U10496 ( .A1(n8117), .A2(n9352), .B1(n9351), .B2(P1_U3084), .C1(
        n9350), .C2(n9349), .ZN(P1_U3324) );
  MUX2_X1 U10497 ( .A(n9353), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10498 ( .A1(n9960), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9365) );
  AOI211_X1 U10499 ( .C1(n9356), .C2(n9355), .A(n9354), .B(n9951), .ZN(n9357)
         );
  AOI21_X1 U10500 ( .B1(n9359), .B2(n9358), .A(n9357), .ZN(n9364) );
  OAI211_X1 U10501 ( .C1(n9362), .C2(n9361), .A(n9956), .B(n9360), .ZN(n9363)
         );
  NAND3_X1 U10502 ( .A1(n9365), .A2(n9364), .A3(n9363), .ZN(P2_U3247) );
  OAI211_X1 U10503 ( .C1(n9368), .C2(n9652), .A(n9367), .B(n9366), .ZN(n9369)
         );
  AOI21_X1 U10504 ( .B1(n9370), .B2(n9681), .A(n9369), .ZN(n9372) );
  INV_X1 U10505 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9371) );
  AOI22_X1 U10506 ( .A1(n9685), .A2(n9372), .B1(n9371), .B2(n9683), .ZN(
        P1_U3484) );
  AOI22_X1 U10507 ( .A1(n9696), .A2(n9372), .B1(n6397), .B2(n9693), .ZN(
        P1_U3533) );
  NOR2_X1 U10508 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9373) );
  AOI21_X1 U10509 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9373), .ZN(n9777) );
  NOR2_X1 U10510 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9374) );
  AOI21_X1 U10511 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9374), .ZN(n9780) );
  NOR2_X1 U10512 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9375) );
  AOI21_X1 U10513 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9375), .ZN(n9783) );
  NOR2_X1 U10514 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9376) );
  AOI21_X1 U10515 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9376), .ZN(n9786) );
  NOR2_X1 U10516 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9377) );
  AOI21_X1 U10517 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9377), .ZN(n9789) );
  NOR2_X1 U10518 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9384) );
  XNOR2_X1 U10519 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9987) );
  NAND2_X1 U10520 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9382) );
  XOR2_X1 U10521 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n9985) );
  NAND2_X1 U10522 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9380) );
  XOR2_X1 U10523 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n9970) );
  AOI21_X1 U10524 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9771) );
  NAND3_X1 U10525 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9773) );
  OAI21_X1 U10526 ( .B1(n9771), .B2(n9378), .A(n9773), .ZN(n9969) );
  NAND2_X1 U10527 ( .A1(n9970), .A2(n9969), .ZN(n9379) );
  NAND2_X1 U10528 ( .A1(n9380), .A2(n9379), .ZN(n9984) );
  NAND2_X1 U10529 ( .A1(n9985), .A2(n9984), .ZN(n9381) );
  NAND2_X1 U10530 ( .A1(n9382), .A2(n9381), .ZN(n9986) );
  NOR2_X1 U10531 ( .A1(n9987), .A2(n9986), .ZN(n9383) );
  NOR2_X1 U10532 ( .A1(n9384), .A2(n9383), .ZN(n9385) );
  NOR2_X1 U10533 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9385), .ZN(n9973) );
  AND2_X1 U10534 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9385), .ZN(n9974) );
  NOR2_X1 U10535 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9974), .ZN(n9386) );
  NOR2_X1 U10536 ( .A1(n9973), .A2(n9386), .ZN(n9387) );
  NAND2_X1 U10537 ( .A1(n9387), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9389) );
  XOR2_X1 U10538 ( .A(n9387), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n9972) );
  NAND2_X1 U10539 ( .A1(n9972), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9388) );
  NAND2_X1 U10540 ( .A1(n9389), .A2(n9388), .ZN(n9390) );
  NAND2_X1 U10541 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9390), .ZN(n9392) );
  XOR2_X1 U10542 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9390), .Z(n9971) );
  NAND2_X1 U10543 ( .A1(n9971), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9391) );
  NAND2_X1 U10544 ( .A1(n9392), .A2(n9391), .ZN(n9393) );
  NAND2_X1 U10545 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9393), .ZN(n9395) );
  XOR2_X1 U10546 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9393), .Z(n9983) );
  NAND2_X1 U10547 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n9983), .ZN(n9394) );
  NAND2_X1 U10548 ( .A1(n9395), .A2(n9394), .ZN(n9396) );
  AND2_X1 U10549 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9396), .ZN(n9397) );
  XNOR2_X1 U10550 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9396), .ZN(n9981) );
  NOR2_X1 U10551 ( .A1(n9982), .A2(n9981), .ZN(n9980) );
  NAND2_X1 U10552 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9398) );
  OAI21_X1 U10553 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9398), .ZN(n9797) );
  AOI21_X1 U10554 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9796), .ZN(n9795) );
  NAND2_X1 U10555 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9927) );
  OAI21_X1 U10556 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9927), .ZN(n9794) );
  NOR2_X1 U10557 ( .A1(n9795), .A2(n9794), .ZN(n9793) );
  AOI21_X1 U10558 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9793), .ZN(n9792) );
  NOR2_X1 U10559 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_12__SCAN_IN), 
        .ZN(n9399) );
  AOI21_X1 U10560 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9399), .ZN(n9791) );
  NAND2_X1 U10561 ( .A1(n9792), .A2(n9791), .ZN(n9790) );
  OAI21_X1 U10562 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9790), .ZN(n9788) );
  NAND2_X1 U10563 ( .A1(n9789), .A2(n9788), .ZN(n9787) );
  OAI21_X1 U10564 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9787), .ZN(n9785) );
  NAND2_X1 U10565 ( .A1(n9786), .A2(n9785), .ZN(n9784) );
  OAI21_X1 U10566 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9784), .ZN(n9782) );
  NAND2_X1 U10567 ( .A1(n9783), .A2(n9782), .ZN(n9781) );
  OAI21_X1 U10568 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9781), .ZN(n9779) );
  NAND2_X1 U10569 ( .A1(n9780), .A2(n9779), .ZN(n9778) );
  OAI21_X1 U10570 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9778), .ZN(n9776) );
  NAND2_X1 U10571 ( .A1(n9777), .A2(n9776), .ZN(n9775) );
  OAI21_X1 U10572 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9775), .ZN(n9977) );
  NOR2_X1 U10573 ( .A1(n9978), .A2(n9977), .ZN(n9400) );
  NAND2_X1 U10574 ( .A1(n9978), .A2(n9977), .ZN(n9976) );
  OAI21_X1 U10575 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9400), .A(n9976), .ZN(
        n9402) );
  XOR2_X1 U10576 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n9401) );
  XNOR2_X1 U10577 ( .A(n9402), .B(n9401), .ZN(ADD_1071_U4) );
  XNOR2_X1 U10578 ( .A(n9404), .B(n4355), .ZN(n9417) );
  INV_X1 U10579 ( .A(n9417), .ZN(n9461) );
  INV_X1 U10580 ( .A(n9405), .ZN(n9407) );
  OAI21_X1 U10581 ( .B1(n9407), .B2(n9457), .A(n9406), .ZN(n9458) );
  INV_X1 U10582 ( .A(n9458), .ZN(n9408) );
  AOI22_X1 U10583 ( .A1(n9461), .A2(n9447), .B1(n9446), .B2(n9408), .ZN(n9426)
         );
  OAI21_X1 U10584 ( .B1(n9411), .B2(n9410), .A(n9409), .ZN(n9415) );
  OAI22_X1 U10585 ( .A1(n9437), .A2(n9412), .B1(n9436), .B2(n9435), .ZN(n9413)
         );
  AOI21_X1 U10586 ( .B1(n9415), .B2(n9414), .A(n9413), .ZN(n9416) );
  OAI21_X1 U10587 ( .B1(n9417), .B2(n9664), .A(n9416), .ZN(n9459) );
  NOR2_X1 U10588 ( .A1(n9457), .A2(n9418), .ZN(n9423) );
  INV_X1 U10589 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9421) );
  OAI22_X1 U10590 ( .A1(n9424), .A2(n9421), .B1(n9420), .B2(n9419), .ZN(n9422)
         );
  AOI211_X1 U10591 ( .C1(n9459), .C2(n9424), .A(n9423), .B(n9422), .ZN(n9425)
         );
  NAND2_X1 U10592 ( .A1(n9426), .A2(n9425), .ZN(P1_U3278) );
  AND2_X1 U10593 ( .A1(n9428), .A2(n9427), .ZN(n9429) );
  XOR2_X1 U10594 ( .A(n9431), .B(n9429), .Z(n9473) );
  XOR2_X1 U10595 ( .A(n9431), .B(n9430), .Z(n9432) );
  OAI222_X1 U10596 ( .A1(n9437), .A2(n9436), .B1(n9435), .B2(n9434), .C1(n9433), .C2(n9432), .ZN(n9472) );
  AOI21_X1 U10597 ( .B1(n9473), .B2(n9438), .A(n9472), .ZN(n9450) );
  AOI222_X1 U10598 ( .A1(n9442), .A2(n9441), .B1(n9440), .B2(n9439), .C1(
        P1_REG2_REG_11__SCAN_IN), .C2(n9451), .ZN(n9449) );
  OAI21_X1 U10599 ( .B1(n9444), .B2(n9469), .A(n9443), .ZN(n9470) );
  INV_X1 U10600 ( .A(n9470), .ZN(n9445) );
  AOI22_X1 U10601 ( .A1(n9473), .A2(n9447), .B1(n9446), .B2(n9445), .ZN(n9448)
         );
  OAI211_X1 U10602 ( .C1(n9451), .C2(n9450), .A(n9449), .B(n9448), .ZN(
        P1_U3280) );
  INV_X1 U10603 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9892) );
  AOI22_X1 U10604 ( .A1(n9696), .A2(n9475), .B1(n9892), .B2(n9693), .ZN(
        P1_U3553) );
  INV_X1 U10605 ( .A(n9456), .ZN(n9667) );
  OAI22_X1 U10606 ( .A1(n9458), .A2(n9679), .B1(n9457), .B2(n9652), .ZN(n9460)
         );
  AOI211_X1 U10607 ( .C1(n9667), .C2(n9461), .A(n9460), .B(n9459), .ZN(n9477)
         );
  AOI22_X1 U10608 ( .A1(n9696), .A2(n9477), .B1(n9462), .B2(n9693), .ZN(
        P1_U3536) );
  OAI211_X1 U10609 ( .C1(n9465), .C2(n9652), .A(n9464), .B(n9463), .ZN(n9466)
         );
  AOI21_X1 U10610 ( .B1(n9467), .B2(n9681), .A(n9466), .ZN(n9479) );
  AOI22_X1 U10611 ( .A1(n9696), .A2(n9479), .B1(n9468), .B2(n9693), .ZN(
        P1_U3535) );
  OAI22_X1 U10612 ( .A1(n9470), .A2(n9679), .B1(n9469), .B2(n9652), .ZN(n9471)
         );
  AOI211_X1 U10613 ( .C1(n9473), .C2(n9681), .A(n9472), .B(n9471), .ZN(n9481)
         );
  AOI22_X1 U10614 ( .A1(n9696), .A2(n9481), .B1(n9474), .B2(n9693), .ZN(
        P1_U3534) );
  INV_X1 U10615 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9890) );
  INV_X1 U10616 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9476) );
  AOI22_X1 U10617 ( .A1(n9685), .A2(n9477), .B1(n9476), .B2(n9683), .ZN(
        P1_U3493) );
  INV_X1 U10618 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9478) );
  AOI22_X1 U10619 ( .A1(n9685), .A2(n9479), .B1(n9478), .B2(n9683), .ZN(
        P1_U3490) );
  INV_X1 U10620 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9480) );
  AOI22_X1 U10621 ( .A1(n9685), .A2(n9481), .B1(n9480), .B2(n9683), .ZN(
        P1_U3487) );
  XNOR2_X1 U10622 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10623 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X1 U10624 ( .A1(n9488), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9483) );
  INV_X1 U10625 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9843) );
  OR2_X1 U10626 ( .A1(n9843), .A2(P1_U3084), .ZN(n9482) );
  OAI21_X1 U10627 ( .B1(n9484), .B2(n9483), .A(n9482), .ZN(n9503) );
  INV_X1 U10628 ( .A(n9503), .ZN(n9485) );
  NOR2_X1 U10629 ( .A1(n9486), .A2(n9485), .ZN(n9494) );
  NOR2_X1 U10630 ( .A1(n9488), .A2(n9487), .ZN(n9489) );
  NAND2_X1 U10631 ( .A1(n9490), .A2(n9489), .ZN(n9502) );
  INV_X1 U10632 ( .A(n9502), .ZN(n9492) );
  NOR2_X1 U10633 ( .A1(n4269), .A2(n9491), .ZN(n9500) );
  OAI22_X1 U10634 ( .A1(n9492), .A2(n9500), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n9922), .ZN(n9493) );
  AOI22_X1 U10635 ( .A1(n9495), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(n9494), .B2(
        n9493), .ZN(n9497) );
  NAND3_X1 U10636 ( .A1(n9607), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9922), .ZN(
        n9496) );
  OAI211_X1 U10637 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n6710), .A(n9497), .B(
        n9496), .ZN(P1_U3241) );
  INV_X1 U10638 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9889) );
  XNOR2_X1 U10639 ( .A(n9499), .B(n9498), .ZN(n9513) );
  NAND2_X1 U10640 ( .A1(n9501), .A2(n9500), .ZN(n9505) );
  NAND4_X1 U10641 ( .A1(n9505), .A2(n9504), .A3(n9503), .A4(n9502), .ZN(n9537)
         );
  OAI21_X1 U10642 ( .B1(n9508), .B2(n9507), .A(n9506), .ZN(n9509) );
  OAI22_X1 U10643 ( .A1(n9625), .A2(n9509), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n4629), .ZN(n9510) );
  AOI21_X1 U10644 ( .B1(n9511), .B2(n9619), .A(n9510), .ZN(n9512) );
  OAI211_X1 U10645 ( .C1(n9513), .C2(n9613), .A(n9537), .B(n9512), .ZN(n9514)
         );
  INV_X1 U10646 ( .A(n9514), .ZN(n9515) );
  OAI21_X1 U10647 ( .B1(n9628), .B2(n9889), .A(n9515), .ZN(P1_U3243) );
  INV_X1 U10648 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9539) );
  INV_X1 U10649 ( .A(n9516), .ZN(n9519) );
  INV_X1 U10650 ( .A(n9517), .ZN(n9518) );
  NAND2_X1 U10651 ( .A1(n9519), .A2(n9518), .ZN(n9520) );
  AND2_X1 U10652 ( .A1(n9521), .A2(n9520), .ZN(n9535) );
  INV_X1 U10653 ( .A(n9522), .ZN(n9523) );
  NAND2_X1 U10654 ( .A1(n9619), .A2(n9523), .ZN(n9534) );
  NAND2_X1 U10655 ( .A1(n9525), .A2(n9524), .ZN(n9528) );
  INV_X1 U10656 ( .A(n9526), .ZN(n9527) );
  NAND2_X1 U10657 ( .A1(n9528), .A2(n9527), .ZN(n9530) );
  NAND2_X1 U10658 ( .A1(n9530), .A2(n9529), .ZN(n9532) );
  AOI21_X1 U10659 ( .B1(n9607), .B2(n9532), .A(n9531), .ZN(n9533) );
  OAI211_X1 U10660 ( .C1(n9535), .C2(n9613), .A(n9534), .B(n9533), .ZN(n9536)
         );
  INV_X1 U10661 ( .A(n9536), .ZN(n9538) );
  OAI211_X1 U10662 ( .C1(n9539), .C2(n9628), .A(n9538), .B(n9537), .ZN(
        P1_U3245) );
  INV_X1 U10663 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9893) );
  AOI211_X1 U10664 ( .C1(n9542), .C2(n9541), .A(n9540), .B(n9613), .ZN(n9543)
         );
  AOI211_X1 U10665 ( .C1(n9619), .C2(n9545), .A(n9544), .B(n9543), .ZN(n9551)
         );
  AOI21_X1 U10666 ( .B1(n9548), .B2(n9547), .A(n9546), .ZN(n9549) );
  OR2_X1 U10667 ( .A1(n9625), .A2(n9549), .ZN(n9550) );
  OAI211_X1 U10668 ( .C1(n9893), .C2(n9628), .A(n9551), .B(n9550), .ZN(
        P1_U3253) );
  INV_X1 U10669 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9564) );
  AOI211_X1 U10670 ( .C1(n9554), .C2(n9553), .A(n9552), .B(n9613), .ZN(n9555)
         );
  AOI211_X1 U10671 ( .C1(n9619), .C2(n9557), .A(n9556), .B(n9555), .ZN(n9563)
         );
  AOI21_X1 U10672 ( .B1(n9560), .B2(n9559), .A(n9558), .ZN(n9561) );
  OR2_X1 U10673 ( .A1(n9625), .A2(n9561), .ZN(n9562) );
  OAI211_X1 U10674 ( .C1(n9564), .C2(n9628), .A(n9563), .B(n9562), .ZN(
        P1_U3254) );
  INV_X1 U10675 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9906) );
  AOI211_X1 U10676 ( .C1(n9567), .C2(n9566), .A(n9565), .B(n9613), .ZN(n9568)
         );
  AOI211_X1 U10677 ( .C1(n9619), .C2(n9570), .A(n9569), .B(n9568), .ZN(n9576)
         );
  AOI21_X1 U10678 ( .B1(n9573), .B2(n9572), .A(n9571), .ZN(n9574) );
  OR2_X1 U10679 ( .A1(n9625), .A2(n9574), .ZN(n9575) );
  OAI211_X1 U10680 ( .C1(n9906), .C2(n9628), .A(n9576), .B(n9575), .ZN(
        P1_U3255) );
  INV_X1 U10681 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9587) );
  AOI211_X1 U10682 ( .C1(n9579), .C2(n9578), .A(n9577), .B(n9613), .ZN(n9580)
         );
  AOI211_X1 U10683 ( .C1(n9619), .C2(n9582), .A(n9581), .B(n9580), .ZN(n9586)
         );
  OAI211_X1 U10684 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9584), .A(n9607), .B(
        n9583), .ZN(n9585) );
  OAI211_X1 U10685 ( .C1(n9587), .C2(n9628), .A(n9586), .B(n9585), .ZN(
        P1_U3256) );
  INV_X1 U10686 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9599) );
  AOI211_X1 U10687 ( .C1(n9590), .C2(n9589), .A(n9588), .B(n9613), .ZN(n9591)
         );
  AOI211_X1 U10688 ( .C1(n9619), .C2(n9593), .A(n9592), .B(n9591), .ZN(n9598)
         );
  OAI211_X1 U10689 ( .C1(n9596), .C2(n9595), .A(n9607), .B(n9594), .ZN(n9597)
         );
  OAI211_X1 U10690 ( .C1(n9599), .C2(n9628), .A(n9598), .B(n9597), .ZN(
        P1_U3257) );
  INV_X1 U10691 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9924) );
  AOI211_X1 U10692 ( .C1(n9602), .C2(n9601), .A(n9600), .B(n9613), .ZN(n9603)
         );
  AOI211_X1 U10693 ( .C1(n9605), .C2(n9619), .A(n9604), .B(n9603), .ZN(n9611)
         );
  OAI211_X1 U10694 ( .C1(n9609), .C2(n9608), .A(n9607), .B(n9606), .ZN(n9610)
         );
  OAI211_X1 U10695 ( .C1(n9924), .C2(n9628), .A(n9611), .B(n9610), .ZN(
        P1_U3258) );
  INV_X1 U10696 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9629) );
  INV_X1 U10697 ( .A(n9612), .ZN(n9618) );
  AOI211_X1 U10698 ( .C1(n9616), .C2(n9615), .A(n9614), .B(n9613), .ZN(n9617)
         );
  AOI211_X1 U10699 ( .C1(n9620), .C2(n9619), .A(n9618), .B(n9617), .ZN(n9627)
         );
  AOI21_X1 U10700 ( .B1(n9623), .B2(n9622), .A(n9621), .ZN(n9624) );
  OR2_X1 U10701 ( .A1(n9625), .A2(n9624), .ZN(n9626) );
  OAI211_X1 U10702 ( .C1(n9629), .C2(n9628), .A(n9627), .B(n9626), .ZN(
        P1_U3259) );
  NOR2_X1 U10703 ( .A1(n9635), .A2(n9630), .ZN(n9631) );
  AND2_X1 U10704 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9632), .ZN(P1_U3292) );
  AND2_X1 U10705 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9632), .ZN(P1_U3293) );
  AND2_X1 U10706 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9632), .ZN(P1_U3294) );
  AND2_X1 U10707 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9632), .ZN(P1_U3295) );
  AND2_X1 U10708 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9632), .ZN(P1_U3296) );
  AND2_X1 U10709 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9632), .ZN(P1_U3297) );
  AND2_X1 U10710 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9632), .ZN(P1_U3298) );
  AND2_X1 U10711 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9632), .ZN(P1_U3299) );
  AND2_X1 U10712 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9632), .ZN(P1_U3300) );
  AND2_X1 U10713 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9632), .ZN(P1_U3301) );
  AND2_X1 U10714 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9632), .ZN(P1_U3302) );
  AND2_X1 U10715 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9632), .ZN(P1_U3303) );
  INV_X1 U10716 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9868) );
  NOR2_X1 U10717 ( .A1(n9631), .A2(n9868), .ZN(P1_U3304) );
  AND2_X1 U10718 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9632), .ZN(P1_U3305) );
  AND2_X1 U10719 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9632), .ZN(P1_U3306) );
  AND2_X1 U10720 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9632), .ZN(P1_U3307) );
  AND2_X1 U10721 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9632), .ZN(P1_U3308) );
  AND2_X1 U10722 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9632), .ZN(P1_U3309) );
  AND2_X1 U10723 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9632), .ZN(P1_U3310) );
  AND2_X1 U10724 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9632), .ZN(P1_U3311) );
  AND2_X1 U10725 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9632), .ZN(P1_U3312) );
  INV_X1 U10726 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9908) );
  NOR2_X1 U10727 ( .A1(n9631), .A2(n9908), .ZN(P1_U3313) );
  AND2_X1 U10728 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9632), .ZN(P1_U3314) );
  AND2_X1 U10729 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9632), .ZN(P1_U3315) );
  AND2_X1 U10730 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9632), .ZN(P1_U3316) );
  AND2_X1 U10731 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9632), .ZN(P1_U3317) );
  AND2_X1 U10732 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9632), .ZN(P1_U3318) );
  AND2_X1 U10733 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9632), .ZN(P1_U3319) );
  AND2_X1 U10734 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9632), .ZN(P1_U3320) );
  AND2_X1 U10735 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9632), .ZN(P1_U3321) );
  INV_X1 U10736 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9634) );
  AOI21_X1 U10737 ( .B1(n9635), .B2(n9634), .A(n9633), .ZN(P1_U3441) );
  INV_X1 U10738 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9636) );
  AOI22_X1 U10739 ( .A1(n9685), .A2(n9637), .B1(n9636), .B2(n9683), .ZN(
        P1_U3457) );
  OAI21_X1 U10740 ( .B1(n9639), .B2(n9652), .A(n9638), .ZN(n9641) );
  AOI211_X1 U10741 ( .C1(n9681), .C2(n9642), .A(n9641), .B(n9640), .ZN(n9687)
         );
  INV_X1 U10742 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9643) );
  AOI22_X1 U10743 ( .A1(n9685), .A2(n9687), .B1(n9643), .B2(n9683), .ZN(
        P1_U3460) );
  OAI22_X1 U10744 ( .A1(n9645), .A2(n9679), .B1(n9644), .B2(n9652), .ZN(n9647)
         );
  AOI211_X1 U10745 ( .C1(n9681), .C2(n9648), .A(n9647), .B(n9646), .ZN(n9688)
         );
  INV_X1 U10746 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9649) );
  AOI22_X1 U10747 ( .A1(n9685), .A2(n9688), .B1(n9649), .B2(n9683), .ZN(
        P1_U3463) );
  OAI211_X1 U10748 ( .C1(n9653), .C2(n9652), .A(n9651), .B(n9650), .ZN(n9654)
         );
  AOI21_X1 U10749 ( .B1(n9655), .B2(n9681), .A(n9654), .ZN(n9690) );
  INV_X1 U10750 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9656) );
  AOI22_X1 U10751 ( .A1(n9685), .A2(n9690), .B1(n9656), .B2(n9683), .ZN(
        P1_U3469) );
  INV_X1 U10752 ( .A(n9663), .ZN(n9666) );
  INV_X1 U10753 ( .A(n9657), .ZN(n9659) );
  AOI211_X1 U10754 ( .C1(n9661), .C2(n9660), .A(n9659), .B(n9658), .ZN(n9662)
         );
  OAI21_X1 U10755 ( .B1(n9664), .B2(n9663), .A(n9662), .ZN(n9665) );
  AOI21_X1 U10756 ( .B1(n9667), .B2(n9666), .A(n9665), .ZN(n9691) );
  INV_X1 U10757 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9668) );
  AOI22_X1 U10758 ( .A1(n9685), .A2(n9691), .B1(n9668), .B2(n9683), .ZN(
        P1_U3472) );
  INV_X1 U10759 ( .A(n9669), .ZN(n9671) );
  NAND3_X1 U10760 ( .A1(n9672), .A2(n9671), .A3(n9670), .ZN(n9673) );
  AOI21_X1 U10761 ( .B1(n9681), .B2(n9674), .A(n9673), .ZN(n9692) );
  INV_X1 U10762 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9675) );
  AOI22_X1 U10763 ( .A1(n9685), .A2(n9692), .B1(n9675), .B2(n9683), .ZN(
        P1_U3475) );
  OAI211_X1 U10764 ( .C1(n9679), .C2(n9678), .A(n9677), .B(n9676), .ZN(n9680)
         );
  AOI21_X1 U10765 ( .B1(n9682), .B2(n9681), .A(n9680), .ZN(n9695) );
  INV_X1 U10766 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9684) );
  AOI22_X1 U10767 ( .A1(n9685), .A2(n9695), .B1(n9684), .B2(n9683), .ZN(
        P1_U3481) );
  INV_X1 U10768 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9686) );
  AOI22_X1 U10769 ( .A1(n9696), .A2(n9687), .B1(n9686), .B2(n9693), .ZN(
        P1_U3525) );
  AOI22_X1 U10770 ( .A1(n9696), .A2(n9688), .B1(n6192), .B2(n9693), .ZN(
        P1_U3526) );
  INV_X1 U10771 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9689) );
  AOI22_X1 U10772 ( .A1(n9696), .A2(n9690), .B1(n9689), .B2(n9693), .ZN(
        P1_U3528) );
  AOI22_X1 U10773 ( .A1(n9696), .A2(n9691), .B1(n6201), .B2(n9693), .ZN(
        P1_U3529) );
  AOI22_X1 U10774 ( .A1(n9696), .A2(n9692), .B1(n6203), .B2(n9693), .ZN(
        P1_U3530) );
  AOI22_X1 U10775 ( .A1(n9696), .A2(n9695), .B1(n9694), .B2(n9693), .ZN(
        P1_U3532) );
  AOI22_X1 U10776 ( .A1(n9697), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n9956), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U10777 ( .A1(n9697), .A2(n9933), .ZN(n9698) );
  OAI211_X1 U10778 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9699), .A(n9698), .B(
        n9964), .ZN(n9700) );
  INV_X1 U10779 ( .A(n9700), .ZN(n9703) );
  AOI22_X1 U10780 ( .A1(n9960), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9702) );
  OAI221_X1 U10781 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9704), .C1(n9878), .C2(
        n9703), .A(n9702), .ZN(P2_U3245) );
  NAND2_X1 U10782 ( .A1(n9706), .A2(n9705), .ZN(n9707) );
  AND2_X1 U10783 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9707), .ZN(P2_U3297) );
  AND2_X1 U10784 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9707), .ZN(P2_U3298) );
  AND2_X1 U10785 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9707), .ZN(P2_U3299) );
  AND2_X1 U10786 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9707), .ZN(P2_U3300) );
  AND2_X1 U10787 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9707), .ZN(P2_U3301) );
  AND2_X1 U10788 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9707), .ZN(P2_U3302) );
  AND2_X1 U10789 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9707), .ZN(P2_U3303) );
  AND2_X1 U10790 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9707), .ZN(P2_U3304) );
  AND2_X1 U10791 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9707), .ZN(P2_U3305) );
  AND2_X1 U10792 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9707), .ZN(P2_U3306) );
  AND2_X1 U10793 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9707), .ZN(P2_U3307) );
  AND2_X1 U10794 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9707), .ZN(P2_U3308) );
  AND2_X1 U10795 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9707), .ZN(P2_U3309) );
  AND2_X1 U10796 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9707), .ZN(P2_U3310) );
  INV_X1 U10797 ( .A(n9707), .ZN(n9711) );
  INV_X1 U10798 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9860) );
  NOR2_X1 U10799 ( .A1(n9711), .A2(n9860), .ZN(P2_U3311) );
  AND2_X1 U10800 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9707), .ZN(P2_U3312) );
  AND2_X1 U10801 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9707), .ZN(P2_U3313) );
  AND2_X1 U10802 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9707), .ZN(P2_U3314) );
  INV_X1 U10803 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9818) );
  NOR2_X1 U10804 ( .A1(n9711), .A2(n9818), .ZN(P2_U3315) );
  AND2_X1 U10805 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9707), .ZN(P2_U3316) );
  AND2_X1 U10806 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9707), .ZN(P2_U3317) );
  AND2_X1 U10807 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9707), .ZN(P2_U3318) );
  INV_X1 U10808 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9865) );
  NOR2_X1 U10809 ( .A1(n9711), .A2(n9865), .ZN(P2_U3319) );
  AND2_X1 U10810 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9707), .ZN(P2_U3320) );
  AND2_X1 U10811 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9707), .ZN(P2_U3321) );
  AND2_X1 U10812 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9707), .ZN(P2_U3322) );
  AND2_X1 U10813 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9707), .ZN(P2_U3323) );
  AND2_X1 U10814 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9707), .ZN(P2_U3324) );
  AND2_X1 U10815 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9707), .ZN(P2_U3325) );
  INV_X1 U10816 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9807) );
  NOR2_X1 U10817 ( .A1(n9711), .A2(n9807), .ZN(P2_U3326) );
  INV_X1 U10818 ( .A(n9708), .ZN(n9712) );
  OAI22_X1 U10819 ( .A1(n9709), .A2(n9712), .B1(P2_D_REG_0__SCAN_IN), .B2(
        n9711), .ZN(n9710) );
  INV_X1 U10820 ( .A(n9710), .ZN(P2_U3437) );
  OAI22_X1 U10821 ( .A1(n9713), .A2(n9712), .B1(P2_D_REG_1__SCAN_IN), .B2(
        n9711), .ZN(n9714) );
  INV_X1 U10822 ( .A(n9714), .ZN(P2_U3438) );
  AOI22_X1 U10823 ( .A1(n9717), .A2(n9746), .B1(n9716), .B2(n9715), .ZN(n9718)
         );
  AND2_X1 U10824 ( .A1(n9719), .A2(n9718), .ZN(n9761) );
  INV_X1 U10825 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9720) );
  AOI22_X1 U10826 ( .A1(n9759), .A2(n9761), .B1(n9720), .B2(n9758), .ZN(
        P2_U3451) );
  INV_X1 U10827 ( .A(n9721), .ZN(n9723) );
  INV_X1 U10828 ( .A(n9722), .ZN(n9750) );
  OAI22_X1 U10829 ( .A1(n9723), .A2(n9752), .B1(n4979), .B2(n9750), .ZN(n9726)
         );
  INV_X1 U10830 ( .A(n9724), .ZN(n9725) );
  AOI211_X1 U10831 ( .C1(n9746), .C2(n9727), .A(n9726), .B(n9725), .ZN(n9763)
         );
  INV_X1 U10832 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9728) );
  AOI22_X1 U10833 ( .A1(n9759), .A2(n9763), .B1(n9728), .B2(n9758), .ZN(
        P2_U3454) );
  OAI211_X1 U10834 ( .C1(n9731), .C2(n9750), .A(n9730), .B(n9729), .ZN(n9732)
         );
  AOI21_X1 U10835 ( .B1(n9746), .B2(n9733), .A(n9732), .ZN(n9764) );
  INV_X1 U10836 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9734) );
  AOI22_X1 U10837 ( .A1(n9759), .A2(n9764), .B1(n9734), .B2(n9758), .ZN(
        P2_U3457) );
  OAI211_X1 U10838 ( .C1(n9737), .C2(n9750), .A(n9736), .B(n9735), .ZN(n9738)
         );
  AOI21_X1 U10839 ( .B1(n9746), .B2(n9739), .A(n9738), .ZN(n9765) );
  INV_X1 U10840 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9740) );
  AOI22_X1 U10841 ( .A1(n9759), .A2(n9765), .B1(n9740), .B2(n9758), .ZN(
        P2_U3466) );
  OAI211_X1 U10842 ( .C1(n9743), .C2(n9750), .A(n9742), .B(n9741), .ZN(n9744)
         );
  AOI21_X1 U10843 ( .B1(n9746), .B2(n9745), .A(n9744), .ZN(n9766) );
  INV_X1 U10844 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9747) );
  AOI22_X1 U10845 ( .A1(n9759), .A2(n9766), .B1(n9747), .B2(n9758), .ZN(
        P2_U3469) );
  INV_X1 U10846 ( .A(n9748), .ZN(n9757) );
  INV_X1 U10847 ( .A(n9749), .ZN(n9756) );
  OAI22_X1 U10848 ( .A1(n9753), .A2(n9752), .B1(n9751), .B2(n9750), .ZN(n9755)
         );
  AOI211_X1 U10849 ( .C1(n9757), .C2(n9756), .A(n9755), .B(n9754), .ZN(n9769)
         );
  INV_X1 U10850 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9814) );
  AOI22_X1 U10851 ( .A1(n9759), .A2(n9769), .B1(n9814), .B2(n9758), .ZN(
        P2_U3475) );
  INV_X1 U10852 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9760) );
  AOI22_X1 U10853 ( .A1(n9770), .A2(n9761), .B1(n9760), .B2(n9767), .ZN(
        P2_U3520) );
  INV_X1 U10854 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9762) );
  AOI22_X1 U10855 ( .A1(n9770), .A2(n9763), .B1(n9762), .B2(n9767), .ZN(
        P2_U3521) );
  AOI22_X1 U10856 ( .A1(n9770), .A2(n9764), .B1(n6294), .B2(n9767), .ZN(
        P2_U3522) );
  AOI22_X1 U10857 ( .A1(n9770), .A2(n9765), .B1(n6291), .B2(n9767), .ZN(
        P2_U3525) );
  AOI22_X1 U10858 ( .A1(n9770), .A2(n9766), .B1(n6300), .B2(n9767), .ZN(
        P2_U3526) );
  AOI22_X1 U10859 ( .A1(n9770), .A2(n9769), .B1(n9768), .B2(n9767), .ZN(
        P2_U3528) );
  INV_X1 U10860 ( .A(n9771), .ZN(n9772) );
  NAND2_X1 U10861 ( .A1(n9773), .A2(n9772), .ZN(n9774) );
  XNOR2_X1 U10862 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9774), .ZN(ADD_1071_U5) );
  XOR2_X1 U10863 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10864 ( .B1(n9777), .B2(n9776), .A(n9775), .ZN(ADD_1071_U56) );
  OAI21_X1 U10865 ( .B1(n9780), .B2(n9779), .A(n9778), .ZN(ADD_1071_U57) );
  OAI21_X1 U10866 ( .B1(n9783), .B2(n9782), .A(n9781), .ZN(ADD_1071_U58) );
  OAI21_X1 U10867 ( .B1(n9786), .B2(n9785), .A(n9784), .ZN(ADD_1071_U59) );
  OAI21_X1 U10868 ( .B1(n9789), .B2(n9788), .A(n9787), .ZN(ADD_1071_U60) );
  OAI21_X1 U10869 ( .B1(n9792), .B2(n9791), .A(n9790), .ZN(ADD_1071_U61) );
  AOI21_X1 U10870 ( .B1(n9795), .B2(n9794), .A(n9793), .ZN(ADD_1071_U62) );
  AOI21_X1 U10871 ( .B1(n9798), .B2(n9797), .A(n9796), .ZN(ADD_1071_U63) );
  INV_X1 U10872 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9801) );
  AOI22_X1 U10873 ( .A1(n9801), .A2(keyinput25), .B1(n9800), .B2(keyinput10), 
        .ZN(n9799) );
  OAI221_X1 U10874 ( .B1(n9801), .B2(keyinput25), .C1(n9800), .C2(keyinput10), 
        .A(n9799), .ZN(n9812) );
  INV_X1 U10875 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9804) );
  INV_X1 U10876 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9803) );
  AOI22_X1 U10877 ( .A1(n9804), .A2(keyinput1), .B1(n9803), .B2(keyinput63), 
        .ZN(n9802) );
  OAI221_X1 U10878 ( .B1(n9804), .B2(keyinput1), .C1(n9803), .C2(keyinput63), 
        .A(n9802), .ZN(n9811) );
  AOI22_X1 U10879 ( .A1(n9807), .A2(keyinput52), .B1(n9806), .B2(keyinput6), 
        .ZN(n9805) );
  OAI221_X1 U10880 ( .B1(n9807), .B2(keyinput52), .C1(n9806), .C2(keyinput6), 
        .A(n9805), .ZN(n9810) );
  AOI22_X1 U10881 ( .A1(n5262), .A2(keyinput34), .B1(n9922), .B2(keyinput31), 
        .ZN(n9808) );
  OAI221_X1 U10882 ( .B1(n5262), .B2(keyinput34), .C1(n9922), .C2(keyinput31), 
        .A(n9808), .ZN(n9809) );
  NOR4_X1 U10883 ( .A1(n9812), .A2(n9811), .A3(n9810), .A4(n9809), .ZN(n9858)
         );
  INV_X1 U10884 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9815) );
  AOI22_X1 U10885 ( .A1(n9815), .A2(keyinput23), .B1(keyinput5), .B2(n9814), 
        .ZN(n9813) );
  OAI221_X1 U10886 ( .B1(n9815), .B2(keyinput23), .C1(n9814), .C2(keyinput5), 
        .A(n9813), .ZN(n9828) );
  AOI22_X1 U10887 ( .A1(n9818), .A2(keyinput37), .B1(keyinput48), .B2(n9817), 
        .ZN(n9816) );
  OAI221_X1 U10888 ( .B1(n9818), .B2(keyinput37), .C1(n9817), .C2(keyinput48), 
        .A(n9816), .ZN(n9827) );
  AOI22_X1 U10889 ( .A1(n9821), .A2(keyinput26), .B1(keyinput47), .B2(n9820), 
        .ZN(n9819) );
  OAI221_X1 U10890 ( .B1(n9821), .B2(keyinput26), .C1(n9820), .C2(keyinput47), 
        .A(n9819), .ZN(n9825) );
  XNOR2_X1 U10891 ( .A(n9924), .B(keyinput20), .ZN(n9824) );
  XNOR2_X1 U10892 ( .A(n9822), .B(keyinput54), .ZN(n9823) );
  OR3_X1 U10893 ( .A1(n9825), .A2(n9824), .A3(n9823), .ZN(n9826) );
  NOR3_X1 U10894 ( .A1(n9828), .A2(n9827), .A3(n9826), .ZN(n9857) );
  AOI22_X1 U10895 ( .A1(n9830), .A2(keyinput7), .B1(n5295), .B2(keyinput16), 
        .ZN(n9829) );
  OAI221_X1 U10896 ( .B1(n9830), .B2(keyinput7), .C1(n5295), .C2(keyinput16), 
        .A(n9829), .ZN(n9841) );
  INV_X1 U10897 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9832) );
  AOI22_X1 U10898 ( .A1(n9832), .A2(keyinput59), .B1(keyinput19), .B2(n5421), 
        .ZN(n9831) );
  OAI221_X1 U10899 ( .B1(n9832), .B2(keyinput59), .C1(n5421), .C2(keyinput19), 
        .A(n9831), .ZN(n9840) );
  AOI22_X1 U10900 ( .A1(n9834), .A2(keyinput24), .B1(n9934), .B2(keyinput51), 
        .ZN(n9833) );
  OAI221_X1 U10901 ( .B1(n9834), .B2(keyinput24), .C1(n9934), .C2(keyinput51), 
        .A(n9833), .ZN(n9839) );
  AOI22_X1 U10902 ( .A1(n9837), .A2(keyinput38), .B1(n9836), .B2(keyinput12), 
        .ZN(n9835) );
  OAI221_X1 U10903 ( .B1(n9837), .B2(keyinput38), .C1(n9836), .C2(keyinput12), 
        .A(n9835), .ZN(n9838) );
  NOR4_X1 U10904 ( .A1(n9841), .A2(n9840), .A3(n9839), .A4(n9838), .ZN(n9856)
         );
  AOI22_X1 U10905 ( .A1(n6463), .A2(keyinput57), .B1(n9843), .B2(keyinput61), 
        .ZN(n9842) );
  OAI221_X1 U10906 ( .B1(n6463), .B2(keyinput57), .C1(n9843), .C2(keyinput61), 
        .A(n9842), .ZN(n9854) );
  AOI22_X1 U10907 ( .A1(n9846), .A2(keyinput33), .B1(n9845), .B2(keyinput53), 
        .ZN(n9844) );
  OAI221_X1 U10908 ( .B1(n9846), .B2(keyinput33), .C1(n9845), .C2(keyinput53), 
        .A(n9844), .ZN(n9853) );
  AOI22_X1 U10909 ( .A1(n6710), .A2(keyinput44), .B1(keyinput45), .B2(n9848), 
        .ZN(n9847) );
  OAI221_X1 U10910 ( .B1(n6710), .B2(keyinput44), .C1(n9848), .C2(keyinput45), 
        .A(n9847), .ZN(n9852) );
  INV_X1 U10911 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9850) );
  AOI22_X1 U10912 ( .A1(n6391), .A2(keyinput35), .B1(n9850), .B2(keyinput30), 
        .ZN(n9849) );
  OAI221_X1 U10913 ( .B1(n6391), .B2(keyinput35), .C1(n9850), .C2(keyinput30), 
        .A(n9849), .ZN(n9851) );
  NOR4_X1 U10914 ( .A1(n9854), .A2(n9853), .A3(n9852), .A4(n9851), .ZN(n9855)
         );
  NAND4_X1 U10915 ( .A1(n9858), .A2(n9857), .A3(n9856), .A4(n9855), .ZN(n9921)
         );
  AOI22_X1 U10916 ( .A1(n9933), .A2(keyinput4), .B1(n9860), .B2(keyinput11), 
        .ZN(n9859) );
  OAI221_X1 U10917 ( .B1(n9933), .B2(keyinput4), .C1(n9860), .C2(keyinput11), 
        .A(n9859), .ZN(n9873) );
  AOI22_X1 U10918 ( .A1(n9863), .A2(keyinput15), .B1(n9862), .B2(keyinput55), 
        .ZN(n9861) );
  OAI221_X1 U10919 ( .B1(n9863), .B2(keyinput15), .C1(n9862), .C2(keyinput55), 
        .A(n9861), .ZN(n9872) );
  AOI22_X1 U10920 ( .A1(n9866), .A2(keyinput18), .B1(n9865), .B2(keyinput46), 
        .ZN(n9864) );
  OAI221_X1 U10921 ( .B1(n9866), .B2(keyinput18), .C1(n9865), .C2(keyinput46), 
        .A(n9864), .ZN(n9871) );
  AOI22_X1 U10922 ( .A1(n9869), .A2(keyinput28), .B1(n9868), .B2(keyinput0), 
        .ZN(n9867) );
  OAI221_X1 U10923 ( .B1(n9869), .B2(keyinput28), .C1(n9868), .C2(keyinput0), 
        .A(n9867), .ZN(n9870) );
  NOR4_X1 U10924 ( .A1(n9873), .A2(n9872), .A3(n9871), .A4(n9870), .ZN(n9919)
         );
  INV_X1 U10925 ( .A(SI_0_), .ZN(n9875) );
  AOI22_X1 U10926 ( .A1(n9875), .A2(keyinput56), .B1(keyinput36), .B2(n9978), 
        .ZN(n9874) );
  OAI221_X1 U10927 ( .B1(n9875), .B2(keyinput56), .C1(n9978), .C2(keyinput36), 
        .A(n9874), .ZN(n9887) );
  INV_X1 U10928 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9877) );
  AOI22_X1 U10929 ( .A1(n9878), .A2(keyinput2), .B1(keyinput43), .B2(n9877), 
        .ZN(n9876) );
  OAI221_X1 U10930 ( .B1(n9878), .B2(keyinput2), .C1(n9877), .C2(keyinput43), 
        .A(n9876), .ZN(n9886) );
  INV_X1 U10931 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9880) );
  AOI22_X1 U10932 ( .A1(n9881), .A2(keyinput62), .B1(keyinput60), .B2(n9880), 
        .ZN(n9879) );
  OAI221_X1 U10933 ( .B1(n9881), .B2(keyinput62), .C1(n9880), .C2(keyinput60), 
        .A(n9879), .ZN(n9885) );
  XNOR2_X1 U10934 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput41), .ZN(n9883) );
  XNOR2_X1 U10935 ( .A(keyinput32), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U10936 ( .A1(n9883), .A2(n9882), .ZN(n9884) );
  NOR4_X1 U10937 ( .A1(n9887), .A2(n9886), .A3(n9885), .A4(n9884), .ZN(n9918)
         );
  AOI22_X1 U10938 ( .A1(n9890), .A2(keyinput50), .B1(keyinput49), .B2(n9889), 
        .ZN(n9888) );
  OAI221_X1 U10939 ( .B1(n9890), .B2(keyinput50), .C1(n9889), .C2(keyinput49), 
        .A(n9888), .ZN(n9902) );
  AOI22_X1 U10940 ( .A1(n9893), .A2(keyinput42), .B1(n9892), .B2(keyinput9), 
        .ZN(n9891) );
  OAI221_X1 U10941 ( .B1(n9893), .B2(keyinput42), .C1(n9892), .C2(keyinput9), 
        .A(n9891), .ZN(n9901) );
  AOI22_X1 U10942 ( .A1(n9895), .A2(keyinput3), .B1(n7125), .B2(keyinput39), 
        .ZN(n9894) );
  OAI221_X1 U10943 ( .B1(n9895), .B2(keyinput3), .C1(n7125), .C2(keyinput39), 
        .A(n9894), .ZN(n9900) );
  INV_X1 U10944 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9897) );
  AOI22_X1 U10945 ( .A1(n9898), .A2(keyinput22), .B1(keyinput21), .B2(n9897), 
        .ZN(n9896) );
  OAI221_X1 U10946 ( .B1(n9898), .B2(keyinput22), .C1(n9897), .C2(keyinput21), 
        .A(n9896), .ZN(n9899) );
  NOR4_X1 U10947 ( .A1(n9902), .A2(n9901), .A3(n9900), .A4(n9899), .ZN(n9917)
         );
  INV_X1 U10948 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9904) );
  AOI22_X1 U10949 ( .A1(n6928), .A2(keyinput8), .B1(keyinput58), .B2(n9904), 
        .ZN(n9903) );
  OAI221_X1 U10950 ( .B1(n6928), .B2(keyinput8), .C1(n9904), .C2(keyinput58), 
        .A(n9903), .ZN(n9915) );
  AOI22_X1 U10951 ( .A1(n5143), .A2(keyinput17), .B1(keyinput40), .B2(n9906), 
        .ZN(n9905) );
  OAI221_X1 U10952 ( .B1(n5143), .B2(keyinput17), .C1(n9906), .C2(keyinput40), 
        .A(n9905), .ZN(n9914) );
  INV_X1 U10953 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U10954 ( .A1(n9909), .A2(keyinput29), .B1(n9908), .B2(keyinput14), 
        .ZN(n9907) );
  OAI221_X1 U10955 ( .B1(n9909), .B2(keyinput29), .C1(n9908), .C2(keyinput14), 
        .A(n9907), .ZN(n9913) );
  XNOR2_X1 U10956 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput13), .ZN(n9911) );
  XNOR2_X1 U10957 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput27), .ZN(n9910)
         );
  NAND2_X1 U10958 ( .A1(n9911), .A2(n9910), .ZN(n9912) );
  NOR4_X1 U10959 ( .A1(n9915), .A2(n9914), .A3(n9913), .A4(n9912), .ZN(n9916)
         );
  NAND4_X1 U10960 ( .A1(n9919), .A2(n9918), .A3(n9917), .A4(n9916), .ZN(n9920)
         );
  NOR2_X1 U10961 ( .A1(n9921), .A2(n9920), .ZN(n9950) );
  NOR4_X1 U10962 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .A3(P1_ADDR_REG_2__SCAN_IN), .A4(n9922), .ZN(n9948) );
  INV_X1 U10963 ( .A(n9923), .ZN(n9928) );
  NAND4_X1 U10964 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .A3(P1_ADDR_REG_5__SCAN_IN), .A4(n9924), .ZN(n9926) );
  NAND4_X1 U10965 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .A4(P1_ADDR_REG_12__SCAN_IN), .ZN(n9925) );
  NOR4_X1 U10966 ( .A1(n9928), .A2(n9927), .A3(n9926), .A4(n9925), .ZN(n9947)
         );
  NAND4_X1 U10967 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_REG0_REG_11__SCAN_IN), 
        .A3(P2_REG0_REG_9__SCAN_IN), .A4(P2_REG1_REG_9__SCAN_IN), .ZN(n9932)
         );
  NAND4_X1 U10968 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_REG1_REG_27__SCAN_IN), 
        .A3(P2_REG2_REG_11__SCAN_IN), .A4(P1_REG0_REG_30__SCAN_IN), .ZN(n9931)
         );
  NAND4_X1 U10969 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(P1_REG1_REG_26__SCAN_IN), .A3(P1_REG1_REG_16__SCAN_IN), .A4(P1_REG2_REG_6__SCAN_IN), .ZN(n9930) );
  NAND4_X1 U10970 ( .A1(SI_25_), .A2(P1_REG2_REG_28__SCAN_IN), .A3(
        P2_REG2_REG_25__SCAN_IN), .A4(P2_REG2_REG_22__SCAN_IN), .ZN(n9929) );
  NOR4_X1 U10971 ( .A1(n9932), .A2(n9931), .A3(n9930), .A4(n9929), .ZN(n9946)
         );
  NAND4_X1 U10972 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(n6928), .A3(n9934), .A4(
        n9933), .ZN(n9944) );
  NOR4_X1 U10973 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .A3(P2_REG3_REG_13__SCAN_IN), .A4(P1_DATAO_REG_29__SCAN_IN), .ZN(n9937) );
  NOR4_X1 U10974 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(SI_28_), .A3(
        P2_REG0_REG_24__SCAN_IN), .A4(P2_REG1_REG_30__SCAN_IN), .ZN(n9936) );
  NOR4_X1 U10975 ( .A1(P1_REG0_REG_27__SCAN_IN), .A2(P1_REG1_REG_22__SCAN_IN), 
        .A3(P2_REG0_REG_8__SCAN_IN), .A4(P1_REG1_REG_30__SCAN_IN), .ZN(n9935)
         );
  NAND3_X1 U10976 ( .A1(n9937), .A2(n9936), .A3(n9935), .ZN(n9943) );
  NAND4_X1 U10977 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(SI_23_), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_REG1_REG_28__SCAN_IN), .ZN(n9942) );
  NOR4_X1 U10978 ( .A1(P1_D_REG_19__SCAN_IN), .A2(SI_0_), .A3(
        P1_REG2_REG_9__SCAN_IN), .A4(P1_REG3_REG_0__SCAN_IN), .ZN(n9940) );
  NOR4_X1 U10979 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG0_REG_21__SCAN_IN), 
        .A3(P2_IR_REG_30__SCAN_IN), .A4(P2_REG2_REG_18__SCAN_IN), .ZN(n9938)
         );
  AND3_X1 U10980 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(P1_DATAO_REG_3__SCAN_IN), 
        .A3(n9938), .ZN(n9939) );
  NAND4_X1 U10981 ( .A1(n9940), .A2(P1_DATAO_REG_26__SCAN_IN), .A3(
        P1_DATAO_REG_6__SCAN_IN), .A4(n9939), .ZN(n9941) );
  NOR4_X1 U10982 ( .A1(n9944), .A2(n9943), .A3(n9942), .A4(n9941), .ZN(n9945)
         );
  NAND4_X1 U10983 ( .A1(n9948), .A2(n9947), .A3(n9946), .A4(n9945), .ZN(n9949)
         );
  XNOR2_X1 U10984 ( .A(n9950), .B(n9949), .ZN(n9968) );
  AOI211_X1 U10985 ( .C1(n9954), .C2(n9953), .A(n9952), .B(n9951), .ZN(n9966)
         );
  OAI211_X1 U10986 ( .C1(n9958), .C2(n9957), .A(n9956), .B(n9955), .ZN(n9962)
         );
  AND2_X1 U10987 ( .A1(P2_U3152), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9959) );
  AOI21_X1 U10988 ( .B1(n9960), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n9959), .ZN(
        n9961) );
  OAI211_X1 U10989 ( .C1(n9964), .C2(n9963), .A(n9962), .B(n9961), .ZN(n9965)
         );
  OR2_X1 U10990 ( .A1(n9966), .A2(n9965), .ZN(n9967) );
  XOR2_X1 U10991 ( .A(n9968), .B(n9967), .Z(P2_U3253) );
  XOR2_X1 U10992 ( .A(n9970), .B(n9969), .Z(ADD_1071_U54) );
  XOR2_X1 U10993 ( .A(n9971), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U10994 ( .A(n9972), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U10995 ( .A1(n9974), .A2(n9973), .ZN(n9975) );
  XNOR2_X1 U10996 ( .A(n9975), .B(n6391), .ZN(ADD_1071_U51) );
  OAI21_X1 U10997 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(n9979) );
  XNOR2_X1 U10998 ( .A(n9979), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U10999 ( .B1(n9982), .B2(n9981), .A(n9980), .ZN(ADD_1071_U47) );
  XOR2_X1 U11000 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n9983), .Z(ADD_1071_U48) );
  XOR2_X1 U11001 ( .A(n9985), .B(n9984), .Z(ADD_1071_U53) );
  XNOR2_X1 U11002 ( .A(n9987), .B(n9986), .ZN(ADD_1071_U52) );
  INV_X1 U4775 ( .A(n9157), .ZN(n4434) );
  CLKBUF_X1 U4768 ( .A(n5897), .Z(n5986) );
  CLKBUF_X1 U4785 ( .A(n8126), .Z(n4274) );
  CLKBUF_X2 U4804 ( .A(n5865), .Z(n4268) );
  AND2_X1 U5145 ( .A1(n5699), .A2(n4281), .ZN(n7773) );
  BUF_X4 U5185 ( .A(n5359), .Z(n4264) );
  CLKBUF_X1 U5317 ( .A(n5392), .Z(n6288) );
endmodule

