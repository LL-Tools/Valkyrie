

module b17_C_AntiSAT_k_256_8 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, 
        keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, 
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, 
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, 
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, 
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, 
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, 
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, 
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, 
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, 
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, 
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, 
        keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, 
        keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, 
        keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, 
        keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, 
        keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, 
        keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, 
        keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, 
        keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, 
        keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, 
        keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, 
        keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, 
        keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, 
        keyinput246, keyinput247, keyinput248, keyinput249, keyinput250, 
        keyinput251, keyinput252, keyinput253, keyinput254, keyinput255, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9787, n9788, n9790, n9791, n9792, n9793, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226;

  OR2_X1 U11231 ( .A1(n14621), .A2(n15935), .ZN(n10348) );
  AND2_X1 U11232 ( .A1(n13196), .A2(n13294), .ZN(n20029) );
  INV_X2 U11233 ( .A(n20135), .ZN(n12122) );
  XOR2_X1 U11234 ( .A(n12189), .B(n12188), .Z(n9860) );
  NOR2_X1 U11235 ( .A1(n10532), .A2(n10531), .ZN(n18199) );
  CLKBUF_X2 U11236 ( .A(n10408), .Z(n17157) );
  INV_X1 U11237 ( .A(n12028), .ZN(n13291) );
  AND2_X1 U11238 ( .A1(n12633), .A2(n15567), .ZN(n10975) );
  INV_X1 U11239 ( .A(n10516), .ZN(n16905) );
  INV_X1 U11240 ( .A(n16858), .ZN(n16882) );
  OR2_X1 U11241 ( .A1(n10853), .A2(n10676), .ZN(n12654) );
  INV_X1 U11242 ( .A(n10511), .ZN(n17138) );
  AND2_X1 U11243 ( .A1(n12633), .A2(n10855), .ZN(n10944) );
  AND2_X1 U11244 ( .A1(n9799), .A2(n10859), .ZN(n12660) );
  BUF_X1 U11245 ( .A(n10877), .Z(n12780) );
  INV_X2 U11246 ( .A(n17160), .ZN(n10414) );
  BUF_X1 U11247 ( .A(n10743), .Z(n14310) );
  BUF_X2 U11248 ( .A(n10864), .Z(n10865) );
  AND2_X1 U11249 ( .A1(n11395), .A2(n11734), .ZN(n11739) );
  NAND2_X1 U11250 ( .A1(n10310), .A2(n10724), .ZN(n10771) );
  AND2_X1 U11251 ( .A1(n11825), .A2(n11820), .ZN(n12308) );
  AND2_X4 U11252 ( .A1(n11825), .A2(n13318), .ZN(n11916) );
  NOR2_X1 U11253 ( .A1(n9946), .A2(n10774), .ZN(n10310) );
  AND2_X2 U11254 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14937) );
  NAND2_X1 U11255 ( .A1(n10734), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10735) );
  NAND2_X1 U11256 ( .A1(n10236), .A2(n10235), .ZN(n10754) );
  CLKBUF_X1 U11257 ( .A(n19239), .Z(n9787) );
  NOR2_X1 U11258 ( .A1(n19536), .A2(n19865), .ZN(n19239) );
  AOI222_X1 U11259 ( .A1(n17450), .A2(P3_EAX_REG_15__SCAN_IN), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17465), .C1(BUF2_REG_15__SCAN_IN), 
        .C2(n17464), .ZN(n17466) );
  NOR2_X4 U11260 ( .A1(n17418), .A2(n18665), .ZN(n17450) );
  NOR2_X2 U11261 ( .A1(n17465), .A2(n18813), .ZN(n17464) );
  AND2_X1 U11262 ( .A1(n10895), .A2(n10894), .ZN(n10898) );
  INV_X1 U11263 ( .A(n15588), .ZN(n12571) );
  INV_X1 U11264 ( .A(n12656), .ZN(n12572) );
  INV_X1 U11265 ( .A(n12817), .ZN(n11236) );
  INV_X1 U11266 ( .A(n12654), .ZN(n12570) );
  NAND2_X1 U11267 ( .A1(n10865), .A2(n10676), .ZN(n12656) );
  AND2_X1 U11268 ( .A1(n12632), .A2(n10676), .ZN(n11020) );
  AND2_X1 U11269 ( .A1(n11149), .A2(n13624), .ZN(n13618) );
  AND2_X1 U11270 ( .A1(n12257), .A2(n11986), .ZN(n11915) );
  AND2_X1 U11271 ( .A1(n10344), .A2(n9997), .ZN(n10073) );
  INV_X1 U11272 ( .A(n11289), .ZN(n11539) );
  INV_X1 U11273 ( .A(n16871), .ZN(n17163) );
  INV_X1 U11274 ( .A(n10435), .ZN(n16916) );
  XNOR2_X1 U11275 ( .A(n13180), .B(n12268), .ZN(n13225) );
  INV_X1 U11276 ( .A(n12026), .ZN(n20169) );
  OR2_X1 U11277 ( .A1(n12924), .A2(n12925), .ZN(n15368) );
  NAND2_X1 U11278 ( .A1(n10095), .A2(n9876), .ZN(n10057) );
  INV_X1 U11279 ( .A(n18637), .ZN(n18043) );
  NOR2_X2 U11280 ( .A1(n13669), .A2(n12026), .ZN(n13684) );
  INV_X1 U11281 ( .A(n20002), .ZN(n15809) );
  AND2_X1 U11282 ( .A1(n14501), .A2(n14502), .ZN(n14504) );
  INV_X1 U11283 ( .A(n13669), .ZN(n20152) );
  NAND2_X1 U11284 ( .A1(n10247), .A2(n9864), .ZN(n14701) );
  CLKBUF_X3 U11286 ( .A(n11467), .Z(n19903) );
  INV_X1 U11287 ( .A(n17845), .ZN(n17818) );
  NAND2_X1 U11288 ( .A1(n19951), .A2(n13679), .ZN(n20002) );
  AOI22_X1 U11289 ( .A1(n17834), .A2(n16309), .B1(n17715), .B2(n16308), .ZN(
        n17745) );
  INV_X1 U11290 ( .A(n17837), .ZN(n17829) );
  OR2_X2 U11291 ( .A1(n17810), .A2(n17811), .ZN(n10050) );
  NOR2_X2 U11292 ( .A1(n13971), .A2(n10362), .ZN(n9788) );
  NOR2_X1 U11293 ( .A1(n13971), .A2(n10362), .ZN(n10397) );
  INV_X1 U11294 ( .A(n10397), .ZN(n10435) );
  NAND2_X2 U11295 ( .A1(n11209), .A2(n11208), .ZN(n11199) );
  NAND2_X2 U11296 ( .A1(n11206), .A2(n11257), .ZN(n11209) );
  INV_X2 U11297 ( .A(n12003), .ZN(n20177) );
  NAND2_X2 U11298 ( .A1(n10355), .A2(n10357), .ZN(n12003) );
  INV_X1 U11299 ( .A(n12120), .ZN(n20192) );
  BUF_X4 U11300 ( .A(n11982), .Z(n13191) );
  AOI22_X1 U11301 ( .A1(n15116), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n12438), .B2(n12437), .ZN(n12441) );
  OR2_X4 U11302 ( .A1(n11872), .A2(n11871), .ZN(n11986) );
  NAND2_X2 U11303 ( .A1(n10049), .A2(n10048), .ZN(n16982) );
  INV_X4 U11304 ( .A(n16982), .ZN(n17057) );
  XNOR2_X2 U11305 ( .A(n12740), .B(n12738), .ZN(n14959) );
  NAND2_X2 U11306 ( .A1(n14963), .A2(n12720), .ZN(n12740) );
  NAND4_X4 U11307 ( .A1(n11840), .A2(n11839), .A3(n11838), .A4(n11837), .ZN(
        n12026) );
  AND3_X2 U11308 ( .A1(n10950), .A2(n10949), .A3(n10335), .ZN(n11515) );
  AND4_X2 U11309 ( .A1(n11910), .A2(n11909), .A3(n11908), .A4(n11907), .ZN(
        n11914) );
  INV_X2 U11310 ( .A(n18172), .ZN(n16818) );
  NOR2_X2 U11311 ( .A1(n10542), .A2(n10541), .ZN(n18172) );
  NAND2_X2 U11312 ( .A1(n11034), .A2(n9943), .ZN(n11149) );
  AOI21_X2 U11313 ( .B1(n15232), .B2(n15231), .A(n15181), .ZN(n15223) );
  NOR2_X4 U11314 ( .A1(n15141), .A2(n15332), .ZN(n15129) );
  NAND2_X2 U11315 ( .A1(n13181), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13180) );
  AND2_X4 U11316 ( .A1(n13397), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11820) );
  NOR2_X2 U11317 ( .A1(n15117), .A2(n11069), .ZN(n15315) );
  AND2_X2 U11318 ( .A1(n14504), .A2(n14496), .ZN(n9814) );
  NAND2_X1 U11319 ( .A1(n15477), .A2(n15476), .ZN(n15479) );
  NAND2_X1 U11320 ( .A1(n9951), .A2(n9949), .ZN(n15477) );
  OR2_X1 U11321 ( .A1(n10309), .A2(n9952), .ZN(n9951) );
  INV_X1 U11322 ( .A(n9803), .ZN(n13782) );
  OR2_X1 U11323 ( .A1(n11149), .A2(n13624), .ZN(n11040) );
  NAND3_X1 U11324 ( .A1(n9959), .A2(n11003), .A3(n11033), .ZN(n11063) );
  XNOR2_X1 U11325 ( .A(n10981), .B(n11526), .ZN(n10983) );
  INV_X1 U11326 ( .A(n9945), .ZN(n11003) );
  NAND2_X1 U11327 ( .A1(n10133), .A2(n10131), .ZN(n16164) );
  NAND2_X1 U11328 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17842), .ZN(n17696) );
  INV_X2 U11329 ( .A(n17759), .ZN(n17715) );
  BUF_X1 U11330 ( .A(n14919), .Z(n9821) );
  XNOR2_X1 U11331 ( .A(n13210), .B(n13209), .ZN(n14919) );
  CLKBUF_X1 U11332 ( .A(n20650), .Z(n9939) );
  NOR2_X2 U11333 ( .A1(n16819), .A2(n16418), .ZN(n17834) );
  NOR2_X1 U11334 ( .A1(n17286), .A2(n17292), .ZN(n17285) );
  OR2_X1 U11335 ( .A1(n11779), .A2(n11747), .ZN(n15443) );
  NOR2_X2 U11336 ( .A1(n16819), .A2(n18076), .ZN(n18066) );
  NAND2_X2 U11337 ( .A1(n18052), .A2(n18043), .ZN(n18076) );
  NOR2_X2 U11338 ( .A1(n17417), .A2(n12462), .ZN(n16417) );
  NAND3_X2 U11339 ( .A1(n18181), .A2(n18199), .A3(n18190), .ZN(n10594) );
  CLKBUF_X2 U11340 ( .A(n11528), .Z(n11713) );
  INV_X1 U11341 ( .A(n11681), .ZN(n11495) );
  BUF_X1 U11342 ( .A(n11992), .Z(n14933) );
  CLKBUF_X2 U11343 ( .A(n11160), .Z(n11289) );
  OR2_X1 U11344 ( .A1(n13093), .A2(n13171), .ZN(n12429) );
  INV_X4 U11345 ( .A(n19903), .ZN(n15614) );
  NAND2_X1 U11346 ( .A1(n20192), .A2(n12256), .ZN(n12426) );
  NAND2_X1 U11347 ( .A1(n20169), .A2(n13669), .ZN(n20821) );
  BUF_X1 U11348 ( .A(n10767), .Z(n15640) );
  NOR2_X1 U11349 ( .A1(n12256), .A2(n12120), .ZN(n13193) );
  INV_X4 U11351 ( .A(n16231), .ZN(n11443) );
  CLKBUF_X1 U11352 ( .A(n10755), .Z(n11732) );
  INV_X4 U11353 ( .A(n12653), .ZN(n12569) );
  NAND2_X1 U11354 ( .A1(n20096), .A2(n20145), .ZN(n20212) );
  BUF_X2 U11355 ( .A(n13734), .Z(n9820) );
  INV_X2 U11356 ( .A(n9796), .ZN(n9790) );
  CLKBUF_X2 U11357 ( .A(n10416), .Z(n17144) );
  CLKBUF_X2 U11358 ( .A(n11877), .Z(n14053) );
  CLKBUF_X2 U11359 ( .A(n12308), .Z(n12281) );
  BUF_X4 U11360 ( .A(n13734), .Z(n9791) );
  BUF_X4 U11361 ( .A(n10417), .Z(n9792) );
  CLKBUF_X2 U11362 ( .A(n11865), .Z(n14199) );
  NAND2_X2 U11363 ( .A1(n18796), .A2(n18775), .ZN(n10360) );
  INV_X1 U11364 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n9801) );
  XNOR2_X1 U11365 ( .A(n11778), .B(n11777), .ZN(n12845) );
  AOI21_X1 U11366 ( .B1(n9967), .B2(n9966), .A(n9964), .ZN(n9963) );
  AOI21_X1 U11367 ( .B1(n9967), .B2(n15127), .A(n15126), .ZN(n15128) );
  OR2_X1 U11368 ( .A1(n12839), .A2(n16199), .ZN(n11781) );
  AND2_X1 U11369 ( .A1(n12799), .A2(n12798), .ZN(n14304) );
  NOR2_X1 U11370 ( .A1(n15130), .A2(n10303), .ZN(n12435) );
  AOI211_X1 U11371 ( .C1(n15847), .C2(n14633), .A(n14632), .B(n14631), .ZN(
        n14634) );
  XNOR2_X1 U11372 ( .A(n9858), .B(n14289), .ZN(n14367) );
  INV_X1 U11373 ( .A(n14957), .ZN(n10234) );
  INV_X1 U11374 ( .A(n9814), .ZN(n14495) );
  NAND2_X1 U11375 ( .A1(n14701), .A2(n14700), .ZN(n14699) );
  OR2_X1 U11376 ( .A1(n12719), .A2(n12718), .ZN(n12720) );
  NAND2_X1 U11377 ( .A1(n10093), .A2(n17507), .ZN(n17504) );
  INV_X1 U11378 ( .A(n17506), .ZN(n10093) );
  NAND2_X1 U11379 ( .A1(n13960), .A2(n13959), .ZN(n13961) );
  NOR2_X2 U11380 ( .A1(n13893), .A2(n13895), .ZN(n13960) );
  AND2_X1 U11381 ( .A1(n12403), .A2(n9886), .ZN(n9994) );
  NAND2_X1 U11382 ( .A1(n9802), .A2(n13752), .ZN(n13893) );
  AND2_X1 U11383 ( .A1(n12376), .A2(n15861), .ZN(n9810) );
  NOR2_X1 U11384 ( .A1(n14739), .A2(n14738), .ZN(n14723) );
  AND2_X1 U11385 ( .A1(n11041), .A2(n11040), .ZN(n11036) );
  INV_X1 U11386 ( .A(n11040), .ZN(n13620) );
  AND2_X1 U11387 ( .A1(n15852), .A2(n12399), .ZN(n13800) );
  INV_X1 U11388 ( .A(n11156), .ZN(n11041) );
  NAND2_X1 U11389 ( .A1(n11064), .A2(n11067), .ZN(n11065) );
  OAI21_X1 U11390 ( .B1(n11149), .B2(n11289), .A(n19020), .ZN(n11150) );
  AND2_X1 U11391 ( .A1(n12373), .A2(n12372), .ZN(n15867) );
  NAND2_X1 U11392 ( .A1(n10041), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10040) );
  NAND2_X1 U11393 ( .A1(n10305), .A2(n10304), .ZN(n10303) );
  NAND2_X1 U11394 ( .A1(n11063), .A2(n9961), .ZN(n11156) );
  OR2_X1 U11395 ( .A1(n11063), .A2(n11539), .ZN(n11067) );
  XNOR2_X1 U11396 ( .A(n12394), .B(n12381), .ZN(n13649) );
  NAND2_X1 U11397 ( .A1(n13402), .A2(n13401), .ZN(n13520) );
  NOR2_X1 U11398 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16465), .ZN(n16477) );
  AND2_X1 U11399 ( .A1(n10063), .A2(n17963), .ZN(n10061) );
  NOR2_X1 U11400 ( .A1(n13522), .A2(n13521), .ZN(n13523) );
  NAND2_X1 U11401 ( .A1(n13389), .A2(n13388), .ZN(n13402) );
  AND2_X1 U11402 ( .A1(n10064), .A2(n10094), .ZN(n10063) );
  NOR2_X1 U11403 ( .A1(n16535), .A2(n16469), .ZN(n16498) );
  OR2_X1 U11404 ( .A1(n9834), .A2(n17978), .ZN(n10064) );
  NOR2_X1 U11405 ( .A1(n13126), .A2(n15654), .ZN(n13204) );
  XNOR2_X1 U11406 ( .A(n13167), .B(n13166), .ZN(n19846) );
  INV_X1 U11407 ( .A(n16174), .ZN(n10133) );
  OR2_X1 U11408 ( .A1(n11014), .A2(n11013), .ZN(n11033) );
  XNOR2_X1 U11409 ( .A(n12271), .B(n21116), .ZN(n13278) );
  INV_X1 U11410 ( .A(n10057), .ZN(n10472) );
  NAND2_X1 U11411 ( .A1(n10057), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18036) );
  NAND2_X1 U11412 ( .A1(n16190), .A2(n15509), .ZN(n16174) );
  NOR2_X1 U11413 ( .A1(n10007), .A2(n10006), .ZN(n18860) );
  AND4_X1 U11414 ( .A1(n10849), .A2(n10848), .A3(n10847), .A4(n10846), .ZN(
        n10850) );
  NAND2_X1 U11415 ( .A1(n17327), .A2(n17838), .ZN(n17759) );
  NOR2_X2 U11416 ( .A1(n16191), .A2(n15520), .ZN(n16190) );
  NAND2_X1 U11417 ( .A1(n13226), .A2(n12270), .ZN(n12271) );
  NAND2_X1 U11418 ( .A1(n15522), .A2(n15521), .ZN(n15520) );
  NOR3_X1 U11419 ( .A1(n11199), .A2(n11197), .A3(n11200), .ZN(n11218) );
  OAI21_X2 U11420 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18808), .A(n16418), 
        .ZN(n17845) );
  OR2_X1 U11421 ( .A1(n13134), .A2(n13133), .ZN(n13135) );
  AND2_X1 U11422 ( .A1(n12499), .A2(n12498), .ZN(n13072) );
  INV_X1 U11423 ( .A(n14926), .ZN(n14927) );
  NAND2_X1 U11424 ( .A1(n12249), .A2(n12248), .ZN(n12273) );
  AND2_X1 U11425 ( .A1(n10843), .A2(n10842), .ZN(n10988) );
  NAND2_X1 U11426 ( .A1(n12509), .A2(n12508), .ZN(n13134) );
  AND2_X1 U11427 ( .A1(n12296), .A2(n12295), .ZN(n14926) );
  AND2_X1 U11428 ( .A1(n10833), .A2(n10840), .ZN(n13565) );
  AND2_X1 U11429 ( .A1(n10843), .A2(n10840), .ZN(n10997) );
  NAND2_X1 U11430 ( .A1(n20029), .A2(n11986), .ZN(n14529) );
  NAND2_X1 U11431 ( .A1(n12261), .A2(n12260), .ZN(n12268) );
  XNOR2_X1 U11432 ( .A(n12247), .B(n12245), .ZN(n13207) );
  OAI21_X1 U11433 ( .B1(n13175), .B2(n12391), .A(n12267), .ZN(n13181) );
  NAND2_X1 U11434 ( .A1(n12221), .A2(n12392), .ZN(n12247) );
  INV_X1 U11435 ( .A(n18066), .ZN(n18611) );
  AND2_X1 U11436 ( .A1(n10082), .A2(n10084), .ZN(n13208) );
  NOR2_X1 U11437 ( .A1(n12489), .A2(n12485), .ZN(n10842) );
  NAND2_X1 U11438 ( .A1(n10083), .A2(n20223), .ZN(n10082) );
  NAND2_X1 U11439 ( .A1(n12493), .A2(n12492), .ZN(n13047) );
  AND2_X1 U11440 ( .A1(n12489), .A2(n9968), .ZN(n10839) );
  INV_X2 U11441 ( .A(n19172), .ZN(n19201) );
  NAND2_X1 U11442 ( .A1(n12241), .A2(n12240), .ZN(n20223) );
  INV_X2 U11443 ( .A(n17385), .ZN(n17402) );
  INV_X2 U11444 ( .A(n17193), .ZN(n9793) );
  NAND2_X1 U11445 ( .A1(n10828), .A2(n10827), .ZN(n9969) );
  OAI21_X1 U11446 ( .B1(n10821), .B2(n16211), .A(n10804), .ZN(n10822) );
  NAND2_X1 U11447 ( .A1(n10790), .A2(n10789), .ZN(n10827) );
  NOR2_X2 U11448 ( .A1(n17327), .A2(n16318), .ZN(n17754) );
  NOR2_X1 U11449 ( .A1(n10134), .A2(n10132), .ZN(n10131) );
  INV_X1 U11450 ( .A(n11300), .ZN(n10820) );
  NOR2_X1 U11451 ( .A1(n17417), .A2(n13972), .ZN(n16436) );
  NAND2_X1 U11452 ( .A1(n11435), .A2(n11416), .ZN(n12826) );
  INV_X1 U11453 ( .A(n16166), .ZN(n10132) );
  INV_X1 U11454 ( .A(n11109), .ZN(n11085) );
  NOR2_X1 U11455 ( .A1(n13092), .A2(n12018), .ZN(n12154) );
  MUX2_X1 U11456 ( .A(n11521), .B(n11093), .S(n11084), .Z(n11109) );
  NOR2_X1 U11457 ( .A1(n17344), .A2(n10621), .ZN(n10618) );
  NAND2_X1 U11458 ( .A1(n10091), .A2(n10330), .ZN(n10090) );
  INV_X1 U11459 ( .A(n20821), .ZN(n12397) );
  AND2_X1 U11460 ( .A1(n11031), .A2(n11030), .ZN(n11535) );
  AND2_X1 U11461 ( .A1(n11995), .A2(n11994), .ZN(n11996) );
  NOR2_X1 U11462 ( .A1(n12219), .A2(n20824), .ZN(n12220) );
  INV_X2 U11463 ( .A(n13654), .ZN(n14287) );
  NAND2_X1 U11464 ( .A1(n10329), .A2(n10334), .ZN(n17844) );
  OR2_X1 U11465 ( .A1(n12426), .A2(n14382), .ZN(n12017) );
  OR2_X1 U11466 ( .A1(n10980), .A2(n10979), .ZN(n11526) );
  AOI21_X1 U11467 ( .B1(n11438), .B2(n11732), .A(n12830), .ZN(n10218) );
  AND2_X1 U11468 ( .A1(n10776), .A2(n11740), .ZN(n10724) );
  INV_X2 U11469 ( .A(U212), .ZN(n16369) );
  NOR2_X2 U11470 ( .A1(n10494), .A2(n10493), .ZN(n18813) );
  AOI211_X1 U11471 ( .C1(n17164), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n10550), .B(n10549), .ZN(n10551) );
  OR3_X2 U11472 ( .A1(n10424), .A2(n10423), .A3(n10422), .ZN(n17352) );
  OR2_X1 U11473 ( .A1(n12213), .A2(n12212), .ZN(n12265) );
  OR2_X2 U11474 ( .A1(n11860), .A2(n11859), .ZN(n12250) );
  NAND4_X2 U11475 ( .A1(n11903), .A2(n11902), .A3(n11901), .A4(n11900), .ZN(
        n12120) );
  NAND4_X2 U11476 ( .A1(n11936), .A2(n11935), .A3(n11934), .A4(n11933), .ZN(
        n13669) );
  OR2_X1 U11477 ( .A1(n12202), .A2(n12201), .ZN(n12396) );
  NAND2_X1 U11478 ( .A1(n10237), .A2(n10238), .ZN(n10753) );
  AND4_X1 U11479 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11901) );
  AND4_X1 U11480 ( .A1(n11928), .A2(n11927), .A3(n11926), .A4(n11925), .ZN(
        n11934) );
  AND4_X1 U11481 ( .A1(n11819), .A2(n11818), .A3(n11817), .A4(n11816), .ZN(
        n11840) );
  INV_X4 U11482 ( .A(n11631), .ZN(n12667) );
  AND4_X1 U11483 ( .A1(n11836), .A2(n11835), .A3(n11834), .A4(n11833), .ZN(
        n11837) );
  AND4_X1 U11484 ( .A1(n11920), .A2(n11919), .A3(n11918), .A4(n11917), .ZN(
        n11936) );
  AND4_X1 U11485 ( .A1(n11932), .A2(n11931), .A3(n11930), .A4(n11929), .ZN(
        n11933) );
  AND4_X1 U11486 ( .A1(n11824), .A2(n11823), .A3(n11822), .A4(n11821), .ZN(
        n11839) );
  AND4_X1 U11487 ( .A1(n11924), .A2(n11923), .A3(n11922), .A4(n11921), .ZN(
        n11935) );
  AND4_X1 U11488 ( .A1(n11830), .A2(n11829), .A3(n11828), .A4(n11827), .ZN(
        n11838) );
  AND4_X1 U11489 ( .A1(n11887), .A2(n11886), .A3(n11885), .A4(n11884), .ZN(
        n11903) );
  AND2_X1 U11490 ( .A1(n11912), .A2(n11911), .ZN(n11913) );
  AND4_X1 U11491 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n11900) );
  AND4_X1 U11492 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11902) );
  NAND2_X1 U11493 ( .A1(n9865), .A2(n10672), .ZN(n10238) );
  NAND2_X1 U11494 ( .A1(n10729), .A2(n10676), .ZN(n10736) );
  NAND2_X1 U11495 ( .A1(n10661), .A2(n10336), .ZN(n10236) );
  NAND2_X2 U11496 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19840), .ZN(n19833) );
  NAND2_X2 U11497 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20795), .ZN(n20798) );
  BUF_X2 U11498 ( .A(n10396), .Z(n17089) );
  NAND2_X2 U11499 ( .A1(n19840), .A2(n19786), .ZN(n19832) );
  BUF_X2 U11500 ( .A(n10416), .Z(n10565) );
  AND2_X1 U11501 ( .A1(n10674), .A2(n10673), .ZN(n10679) );
  INV_X2 U11502 ( .A(n20768), .ZN(n20771) );
  AND3_X1 U11503 ( .A1(n10671), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10670), .ZN(n10672) );
  INV_X2 U11504 ( .A(n16404), .ZN(U215) );
  NAND2_X1 U11505 ( .A1(n10865), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11629) );
  NAND2_X2 U11506 ( .A1(n18754), .A2(n18699), .ZN(n18752) );
  INV_X2 U11507 ( .A(n16406), .ZN(n16408) );
  NAND2_X2 U11508 ( .A1(n18754), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18757) );
  BUF_X4 U11509 ( .A(n10447), .Z(n9795) );
  NOR2_X1 U11510 ( .A1(n10359), .A2(n10363), .ZN(n10398) );
  INV_X2 U11511 ( .A(n16272), .ZN(n9796) );
  AND2_X2 U11512 ( .A1(n11831), .A2(n14937), .ZN(n12306) );
  AND2_X2 U11513 ( .A1(n11825), .A2(n11826), .ZN(n14149) );
  AND2_X1 U11514 ( .A1(n10241), .A2(n11826), .ZN(n11877) );
  OR2_X1 U11515 ( .A1(n18633), .A2(n10359), .ZN(n10328) );
  BUF_X4 U11516 ( .A(n10387), .Z(n9797) );
  BUF_X2 U11517 ( .A(n10851), .Z(n10852) );
  CLKBUF_X1 U11518 ( .A(n10879), .Z(n15567) );
  NAND2_X1 U11519 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n10497), .ZN(
        n18632) );
  NAND2_X1 U11520 ( .A1(n10495), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n18633) );
  NAND2_X1 U11521 ( .A1(n10497), .A2(n10495), .ZN(n10363) );
  AND2_X2 U11522 ( .A1(n11826), .A2(n11832), .ZN(n11866) );
  AND2_X2 U11523 ( .A1(n14937), .A2(n13318), .ZN(n12309) );
  INV_X2 U11524 ( .A(n19898), .ZN(n9798) );
  AND2_X2 U11525 ( .A1(n10879), .A2(n16211), .ZN(n12639) );
  AND2_X2 U11526 ( .A1(n13233), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11831) );
  INV_X1 U11527 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18775) );
  AND2_X1 U11528 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18619) );
  AND2_X1 U11529 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10858) );
  CLKBUF_X1 U11530 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n18641) );
  NOR2_X2 U11531 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11826) );
  INV_X1 U11532 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13233) );
  INV_X1 U11533 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13397) );
  NAND4_X1 U11534 ( .A1(n10767), .A2(n12830), .A3(n10753), .A4(n13457), .ZN(
        n10778) );
  NAND2_X1 U11535 ( .A1(n10754), .A2(n10759), .ZN(n11438) );
  AND3_X1 U11536 ( .A1(n10754), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10766), 
        .ZN(n12758) );
  AOI21_X2 U11537 ( .B1(n14950), .B2(n14945), .A(n14947), .ZN(n12799) );
  NOR2_X2 U11538 ( .A1(n14994), .A2(n10226), .ZN(n10225) );
  OR2_X1 U11539 ( .A1(n13046), .A2(n13047), .ZN(n12499) );
  XNOR2_X1 U11540 ( .A(n12305), .B(n14927), .ZN(n20146) );
  NAND2_X1 U11541 ( .A1(n9985), .A2(n12376), .ZN(n15860) );
  AND2_X1 U11542 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9799) );
  INV_X1 U11543 ( .A(n11182), .ZN(n9800) );
  NAND2_X1 U11544 ( .A1(n11188), .A2(n11257), .ZN(n11186) );
  OR2_X2 U11545 ( .A1(n11300), .A2(n9801), .ZN(n10811) );
  NOR2_X2 U11546 ( .A1(n12305), .A2(n14926), .ZN(n12332) );
  AND2_X1 U11547 ( .A1(n10271), .A2(n13751), .ZN(n9802) );
  NAND2_X1 U11548 ( .A1(n13752), .A2(n13751), .ZN(n9803) );
  INV_X1 U11549 ( .A(n15117), .ZN(n9804) );
  AND2_X2 U11550 ( .A1(n11746), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9805) );
  NAND2_X2 U11551 ( .A1(n15129), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15117) );
  AND2_X1 U11552 ( .A1(n11746), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10816) );
  OAI21_X2 U11553 ( .B1(n15151), .B2(n15342), .A(n11251), .ZN(n9957) );
  XNOR2_X2 U11554 ( .A(n10800), .B(n10802), .ZN(n10825) );
  AOI21_X2 U11555 ( .B1(n14707), .B2(n14856), .A(n12410), .ZN(n14857) );
  NOR2_X2 U11556 ( .A1(n13970), .A2(n13969), .ZN(n16434) );
  NOR2_X4 U11557 ( .A1(n18664), .A2(n16459), .ZN(n16790) );
  OR2_X2 U11558 ( .A1(n16231), .A2(n10766), .ZN(n10313) );
  NAND2_X2 U11559 ( .A1(n10841), .A2(n10840), .ZN(n19374) );
  NOR2_X2 U11560 ( .A1(n15069), .A2(n15060), .ZN(n15062) );
  CLKBUF_X1 U11561 ( .A(n12271), .Z(n9806) );
  NAND2_X1 U11562 ( .A1(n9985), .A2(n9810), .ZN(n9807) );
  AND2_X2 U11563 ( .A1(n9807), .A2(n9808), .ZN(n13799) );
  OR2_X1 U11564 ( .A1(n9809), .A2(n15862), .ZN(n9808) );
  INV_X1 U11565 ( .A(n15861), .ZN(n9809) );
  NAND2_X1 U11566 ( .A1(n10087), .A2(n10086), .ZN(n9811) );
  NAND2_X1 U11567 ( .A1(n10087), .A2(n10086), .ZN(n12419) );
  AND3_X2 U11568 ( .A1(n10952), .A2(n10888), .A3(n9915), .ZN(n10985) );
  XNOR2_X1 U11569 ( .A(n10823), .B(n10822), .ZN(n10824) );
  NAND2_X2 U11570 ( .A1(n10797), .A2(n10796), .ZN(n11464) );
  NAND2_X2 U11571 ( .A1(n15559), .A2(n11734), .ZN(n10786) );
  XNOR2_X1 U11572 ( .A(n9860), .B(n12273), .ZN(n13229) );
  AND2_X1 U11573 ( .A1(n14416), .A2(n10262), .ZN(n9812) );
  AND2_X1 U11574 ( .A1(n9814), .A2(n10262), .ZN(n14415) );
  CLKBUF_X1 U11575 ( .A(n13279), .Z(n9813) );
  NAND2_X1 U11576 ( .A1(n13278), .A2(n13277), .ZN(n13279) );
  OR2_X1 U11577 ( .A1(n12247), .A2(n12246), .ZN(n12248) );
  INV_X2 U11578 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10795) );
  NAND2_X2 U11579 ( .A1(n10313), .A2(n11071), .ZN(n11731) );
  NOR2_X1 U11580 ( .A1(n12435), .A2(n12434), .ZN(n12436) );
  NAND2_X1 U11581 ( .A1(n13524), .A2(n13523), .ZN(n13644) );
  NAND2_X2 U11582 ( .A1(n16119), .A2(n11068), .ZN(n15262) );
  XNOR2_X2 U11583 ( .A(n12151), .B(n12150), .ZN(n20277) );
  CLKBUF_X1 U11584 ( .A(n13226), .Z(n9815) );
  NAND2_X1 U11585 ( .A1(n12390), .A2(n15861), .ZN(n9816) );
  NAND2_X1 U11586 ( .A1(n10247), .A2(n9819), .ZN(n9817) );
  AND2_X2 U11587 ( .A1(n9817), .A2(n9818), .ZN(n10087) );
  OR2_X1 U11588 ( .A1(n10332), .A2(n14700), .ZN(n9818) );
  AND2_X1 U11589 ( .A1(n9864), .A2(n15852), .ZN(n9819) );
  NAND2_X1 U11590 ( .A1(n13225), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13226) );
  AOI21_X1 U11591 ( .B1(n12170), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12171), .ZN(n12176) );
  NAND2_X1 U11592 ( .A1(n10247), .A2(n9877), .ZN(n14685) );
  NOR2_X2 U11593 ( .A1(n15216), .A2(n15404), .ZN(n15204) );
  AND2_X1 U11594 ( .A1(n12192), .A2(n12190), .ZN(n12239) );
  NAND2_X1 U11595 ( .A1(n12153), .A2(n12152), .ZN(n12192) );
  AND2_X1 U11596 ( .A1(n10825), .A2(n12485), .ZN(n10844) );
  NAND2_X2 U11597 ( .A1(n9812), .A2(n9814), .ZN(n14406) );
  AOI21_X1 U11598 ( .B1(n10078), .B2(n15872), .A(n9880), .ZN(n9986) );
  AND2_X2 U11599 ( .A1(n12009), .A2(n11998), .ZN(n12142) );
  AND2_X1 U11600 ( .A1(n14359), .A2(n10838), .ZN(n10833) );
  NOR2_X1 U11601 ( .A1(n10838), .A2(n12503), .ZN(n10845) );
  XNOR2_X2 U11602 ( .A(n9857), .B(n10962), .ZN(n13547) );
  NAND2_X2 U11603 ( .A1(n12150), .A2(n12146), .ZN(n12170) );
  NAND2_X2 U11604 ( .A1(n12144), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12150) );
  OR2_X2 U11605 ( .A1(n14406), .A2(n10269), .ZN(n14394) );
  XNOR2_X2 U11606 ( .A(n12303), .B(n20118), .ZN(n13463) );
  NAND2_X2 U11607 ( .A1(n13279), .A2(n12272), .ZN(n12303) );
  NAND2_X2 U11608 ( .A1(n12142), .A2(n20169), .ZN(n12428) );
  NOR2_X2 U11609 ( .A1(n13961), .A2(n10255), .ZN(n14501) );
  AND2_X1 U11610 ( .A1(n11831), .A2(n10241), .ZN(n13734) );
  XNOR2_X2 U11611 ( .A(n12192), .B(n12191), .ZN(n13147) );
  AND2_X2 U11612 ( .A1(n14937), .A2(n13318), .ZN(n9822) );
  NAND2_X1 U11613 ( .A1(n9958), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10821) );
  OAI21_X1 U11614 ( .B1(n10073), .B2(n9825), .A(n10072), .ZN(n9996) );
  INV_X1 U11615 ( .A(n18194), .ZN(n10595) );
  BUF_X1 U11616 ( .A(n11866), .Z(n14186) );
  OAI21_X1 U11617 ( .B1(n12380), .B2(n12323), .A(n12322), .ZN(n12331) );
  INV_X1 U11618 ( .A(n12380), .ZN(n12365) );
  AOI21_X1 U11619 ( .B1(n10778), .B2(n10776), .A(n11443), .ZN(n10777) );
  NOR2_X1 U11620 ( .A1(n17337), .A2(n10628), .ZN(n10613) );
  AND2_X1 U11621 ( .A1(n14443), .A2(n10265), .ZN(n10264) );
  NAND2_X1 U11622 ( .A1(n13935), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14260) );
  NOR2_X1 U11623 ( .A1(n14463), .A2(n14492), .ZN(n10265) );
  NAND2_X1 U11624 ( .A1(n20214), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13654) );
  NAND2_X1 U11625 ( .A1(n12419), .A2(n15852), .ZN(n14654) );
  OR2_X1 U11626 ( .A1(n12099), .A2(n12028), .ZN(n12117) );
  INV_X1 U11627 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10129) );
  INV_X1 U11628 ( .A(n11243), .ZN(n11245) );
  INV_X1 U11629 ( .A(n11147), .ZN(n10143) );
  OR2_X1 U11630 ( .A1(n10838), .A2(n12504), .ZN(n12509) );
  INV_X1 U11631 ( .A(n13422), .ZN(n10125) );
  AND4_X1 U11632 ( .A1(n11047), .A2(n11046), .A3(n11045), .A4(n11044), .ZN(
        n11062) );
  AND4_X1 U11633 ( .A1(n11058), .A2(n11057), .A3(n11056), .A4(n11055), .ZN(
        n11059) );
  NAND2_X1 U11634 ( .A1(n11257), .A2(n9855), .ZN(n11285) );
  NAND2_X1 U11635 ( .A1(n10001), .A2(n11275), .ZN(n10297) );
  INV_X1 U11636 ( .A(n11272), .ZN(n10001) );
  NAND2_X1 U11637 ( .A1(n15151), .A2(n15342), .ZN(n11253) );
  NAND2_X1 U11638 ( .A1(n9945), .A2(n9944), .ZN(n9943) );
  OAI21_X1 U11639 ( .B1(n12503), .B2(n12504), .A(n12502), .ZN(n12510) );
  NAND2_X1 U11640 ( .A1(n10312), .A2(n10776), .ZN(n10311) );
  NAND2_X1 U11641 ( .A1(n10756), .A2(n11443), .ZN(n10312) );
  AND2_X1 U11642 ( .A1(n10774), .A2(n13572), .ZN(n10768) );
  NAND2_X1 U11643 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10362) );
  NOR2_X1 U11644 ( .A1(n16417), .A2(n10597), .ZN(n13972) );
  NAND2_X1 U11645 ( .A1(n9970), .A2(n9874), .ZN(n10639) );
  NOR2_X1 U11646 ( .A1(n18199), .A2(n10591), .ZN(n10592) );
  AND2_X1 U11647 ( .A1(n15726), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13294) );
  OR2_X1 U11648 ( .A1(n14383), .A2(n13053), .ZN(n14363) );
  NAND2_X1 U11649 ( .A1(n14635), .A2(n10349), .ZN(n14604) );
  OAI22_X1 U11650 ( .A1(n19887), .A2(n19885), .B1(n15734), .B2(n11106), .ZN(
        n11463) );
  NAND2_X1 U11651 ( .A1(n12834), .A2(n11432), .ZN(n10279) );
  NAND2_X1 U11652 ( .A1(n12806), .A2(n11719), .ZN(n11787) );
  INV_X1 U11653 ( .A(n12805), .ZN(n10157) );
  INV_X1 U11654 ( .A(n12964), .ZN(n10156) );
  INV_X1 U11655 ( .A(n15281), .ZN(n15283) );
  OR2_X1 U11656 ( .A1(n11234), .A2(n15195), .ZN(n9825) );
  AOI21_X1 U11657 ( .B1(n9950), .B2(n9953), .A(n9923), .ZN(n9949) );
  INV_X1 U11658 ( .A(n10306), .ZN(n9950) );
  NOR2_X1 U11659 ( .A1(n18181), .A2(n10596), .ZN(n12462) );
  INV_X1 U11660 ( .A(n16815), .ZN(n16598) );
  INV_X2 U11661 ( .A(n10544), .ZN(n16885) );
  INV_X1 U11662 ( .A(n10603), .ZN(n10593) );
  INV_X1 U11663 ( .A(n18813), .ZN(n16819) );
  AND2_X1 U11664 ( .A1(n11983), .A2(n11986), .ZN(n12155) );
  NOR2_X1 U11665 ( .A1(n20821), .A2(n20192), .ZN(n12018) );
  AND2_X1 U11666 ( .A1(n13781), .A2(n13866), .ZN(n10274) );
  AND2_X1 U11667 ( .A1(n13781), .A2(n13810), .ZN(n10273) );
  NOR2_X1 U11668 ( .A1(n10337), .A2(n20169), .ZN(n10081) );
  OR2_X1 U11669 ( .A1(n12233), .A2(n12232), .ZN(n12255) );
  AND2_X2 U11670 ( .A1(n20177), .A2(n12250), .ZN(n12257) );
  OR2_X1 U11671 ( .A1(n12294), .A2(n12293), .ZN(n12346) );
  OR2_X1 U11672 ( .A1(n12120), .A2(n20824), .ZN(n12243) );
  OR2_X1 U11673 ( .A1(n13669), .A2(n20824), .ZN(n12222) );
  OR2_X1 U11674 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20143), .ZN(
        n11807) );
  AND2_X1 U11675 ( .A1(n20978), .A2(n13315), .ZN(n10140) );
  INV_X1 U11676 ( .A(n14988), .ZN(n10229) );
  INV_X1 U11677 ( .A(n11032), .ZN(n9960) );
  NAND2_X1 U11678 ( .A1(n10985), .A2(n11526), .ZN(n9945) );
  AOI22_X1 U11679 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19281), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U11680 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n15603), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U11681 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n13565), .B1(
        n10995), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U11682 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19408), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U11683 ( .A1(n10997), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n19436), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U11684 ( .A1(n10742), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10750) );
  NAND2_X1 U11685 ( .A1(n10748), .A2(n10676), .ZN(n10749) );
  AOI21_X1 U11686 ( .B1(n18645), .B2(n18641), .A(n10496), .ZN(n10503) );
  AND2_X1 U11687 ( .A1(n10504), .A2(n10608), .ZN(n10496) );
  AND2_X1 U11688 ( .A1(n13193), .A2(n11984), .ZN(n13059) );
  NAND2_X1 U11689 ( .A1(n12009), .A2(n12008), .ZN(n12163) );
  NOR2_X1 U11690 ( .A1(n12250), .A2(n12003), .ZN(n13192) );
  NAND2_X1 U11691 ( .A1(n14219), .A2(n10270), .ZN(n10269) );
  INV_X1 U11692 ( .A(n14407), .ZN(n10270) );
  INV_X1 U11693 ( .A(n14260), .ZN(n14277) );
  NOR2_X1 U11694 ( .A1(n10258), .A2(n14517), .ZN(n10257) );
  INV_X1 U11695 ( .A(n10259), .ZN(n10258) );
  AOI21_X1 U11696 ( .B1(n15852), .B2(n10089), .A(n14833), .ZN(n10086) );
  INV_X1 U11697 ( .A(n14493), .ZN(n10160) );
  NOR2_X1 U11698 ( .A1(n14499), .A2(n10162), .ZN(n10161) );
  INV_X1 U11699 ( .A(n14505), .ZN(n10162) );
  NOR2_X1 U11700 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10250) );
  NOR2_X1 U11701 ( .A1(n13871), .A2(n10167), .ZN(n10166) );
  INV_X1 U11702 ( .A(n13919), .ZN(n10167) );
  INV_X1 U11703 ( .A(n12401), .ZN(n9992) );
  NAND2_X1 U11704 ( .A1(n10172), .A2(n13708), .ZN(n10171) );
  INV_X1 U11705 ( .A(n10173), .ZN(n10172) );
  INV_X1 U11706 ( .A(n12366), .ZN(n10252) );
  NAND2_X1 U11707 ( .A1(n20185), .A2(n13669), .ZN(n12112) );
  NAND2_X1 U11708 ( .A1(n11940), .A2(n12120), .ZN(n12380) );
  AND2_X1 U11709 ( .A1(n12242), .A2(n20824), .ZN(n10083) );
  NAND2_X1 U11710 ( .A1(n10766), .A2(n16231), .ZN(n11071) );
  INV_X1 U11711 ( .A(n11114), .ZN(n10144) );
  NOR2_X1 U11712 ( .A1(n11114), .A2(n11113), .ZN(n11133) );
  OAI21_X1 U11713 ( .B1(n11085), .B2(n12817), .A(n11110), .ZN(n11114) );
  NAND2_X1 U11714 ( .A1(n12817), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11110) );
  NAND2_X1 U11715 ( .A1(n10813), .A2(n10812), .ZN(n10814) );
  NAND2_X1 U11716 ( .A1(n10066), .A2(n10276), .ZN(n10275) );
  AND2_X1 U11717 ( .A1(n12740), .A2(n12738), .ZN(n12742) );
  NOR2_X1 U11718 ( .A1(n10227), .A2(n10223), .ZN(n10222) );
  NAND2_X1 U11719 ( .A1(n10221), .A2(n10228), .ZN(n10227) );
  INV_X1 U11720 ( .A(n10228), .ZN(n10226) );
  AND2_X1 U11721 ( .A1(n10155), .A2(n10154), .ZN(n10153) );
  INV_X1 U11722 ( .A(n15416), .ZN(n10154) );
  OR2_X1 U11723 ( .A1(n11146), .A2(n11145), .ZN(n11532) );
  NAND2_X1 U11724 ( .A1(n11733), .A2(n10779), .ZN(n10780) );
  OR2_X1 U11725 ( .A1(n15341), .A2(n11769), .ZN(n15281) );
  AND2_X1 U11726 ( .A1(n10294), .A2(n10293), .ZN(n10292) );
  INV_X1 U11727 ( .A(n14978), .ZN(n10293) );
  NOR2_X1 U11728 ( .A1(n12935), .A2(n10295), .ZN(n10294) );
  AND2_X1 U11729 ( .A1(n13759), .A2(n15448), .ZN(n10155) );
  AND2_X1 U11730 ( .A1(n10284), .A2(n10283), .ZN(n10282) );
  INV_X1 U11731 ( .A(n15024), .ZN(n10283) );
  NOR2_X1 U11732 ( .A1(n15033), .A2(n10285), .ZN(n10284) );
  INV_X1 U11733 ( .A(n13605), .ZN(n10285) );
  OR2_X1 U11734 ( .A1(n16175), .A2(n10136), .ZN(n10135) );
  INV_X1 U11735 ( .A(n15501), .ZN(n10136) );
  OR2_X1 U11736 ( .A1(n10135), .A2(n15480), .ZN(n10134) );
  INV_X1 U11737 ( .A(n13200), .ZN(n11321) );
  AND2_X1 U11738 ( .A1(n11172), .A2(n20978), .ZN(n11179) );
  INV_X1 U11739 ( .A(n11451), .ZN(n11455) );
  AND2_X2 U11740 ( .A1(n10751), .A2(n13572), .ZN(n11734) );
  AND2_X1 U11741 ( .A1(n10663), .A2(n10662), .ZN(n10667) );
  INV_X1 U11742 ( .A(n11721), .ZN(n10796) );
  NAND2_X1 U11743 ( .A1(n10068), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9947) );
  NAND2_X1 U11744 ( .A1(n10067), .A2(n10676), .ZN(n9948) );
  INV_X2 U11745 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16211) );
  NOR2_X1 U11746 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18796), .ZN(
        n10504) );
  OAI211_X1 U11747 ( .C1(n16884), .C2(n10404), .A(n10403), .B(n10326), .ZN(
        n10405) );
  NOR2_X1 U11748 ( .A1(n18632), .A2(n10362), .ZN(n10447) );
  INV_X1 U11749 ( .A(n10362), .ZN(n10048) );
  INV_X1 U11750 ( .A(n10363), .ZN(n10049) );
  NAND2_X1 U11751 ( .A1(n18796), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10361) );
  AND2_X1 U11752 ( .A1(n17248), .A2(n10106), .ZN(n10603) );
  INV_X1 U11753 ( .A(n18185), .ZN(n10106) );
  NAND2_X1 U11754 ( .A1(n10029), .A2(n10028), .ZN(n10022) );
  NOR2_X1 U11755 ( .A1(n17709), .A2(n17710), .ZN(n10028) );
  NOR2_X1 U11756 ( .A1(n17746), .A2(n16693), .ZN(n10029) );
  NOR2_X1 U11757 ( .A1(n10060), .A2(n17862), .ZN(n10059) );
  NAND2_X1 U11758 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17760), .ZN(
        n10642) );
  OAI21_X1 U11759 ( .B1(n17787), .B2(n10051), .A(n10052), .ZN(n10470) );
  NAND2_X1 U11760 ( .A1(n17771), .A2(n9862), .ZN(n10052) );
  NAND2_X1 U11761 ( .A1(n10056), .A2(n9862), .ZN(n10051) );
  NOR2_X1 U11762 ( .A1(n17784), .A2(n10633), .ZN(n10635) );
  NOR2_X1 U11763 ( .A1(n10464), .A2(n17337), .ZN(n10466) );
  INV_X1 U11764 ( .A(n17334), .ZN(n10614) );
  NOR2_X1 U11765 ( .A1(n17814), .A2(n10627), .ZN(n10629) );
  INV_X1 U11766 ( .A(n17352), .ZN(n10621) );
  XNOR2_X1 U11767 ( .A(n10090), .B(n17352), .ZN(n10460) );
  NAND2_X1 U11768 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18775), .ZN(
        n10359) );
  INV_X1 U11769 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18645) );
  NAND2_X1 U11770 ( .A1(n13189), .A2(n13291), .ZN(n10181) );
  CLKBUF_X1 U11771 ( .A(n12028), .Z(n14360) );
  OR2_X1 U11772 ( .A1(n15834), .A2(n10352), .ZN(n14035) );
  INV_X1 U11773 ( .A(n13514), .ZN(n14286) );
  NAND2_X1 U11774 ( .A1(n14242), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14281) );
  OR2_X1 U11775 ( .A1(n14180), .A2(n14179), .ZN(n14214) );
  OR2_X1 U11776 ( .A1(n14142), .A2(n14434), .ZN(n14143) );
  AND2_X1 U11777 ( .A1(n10264), .A2(n10263), .ZN(n10262) );
  INV_X1 U11778 ( .A(n14430), .ZN(n10263) );
  OR2_X1 U11779 ( .A1(n14118), .A2(n14117), .ZN(n14138) );
  NOR2_X2 U11780 ( .A1(n13644), .A2(n13643), .ZN(n13656) );
  AOI21_X1 U11781 ( .B1(n13519), .B2(n13951), .A(n13518), .ZN(n13522) );
  AOI21_X1 U11782 ( .B1(n13490), .B2(n13951), .A(n13489), .ZN(n13521) );
  NOR2_X1 U11783 ( .A1(n10179), .A2(n10178), .ZN(n14379) );
  NOR2_X1 U11784 ( .A1(n14431), .A2(n10175), .ZN(n14383) );
  NAND2_X1 U11785 ( .A1(n14405), .A2(n10176), .ZN(n10175) );
  NOR3_X1 U11786 ( .A1(n10177), .A2(n14417), .A3(n10178), .ZN(n10176) );
  NAND2_X1 U11787 ( .A1(n14604), .A2(n15852), .ZN(n12422) );
  OR2_X1 U11788 ( .A1(n14456), .A2(n14433), .ZN(n14431) );
  NAND2_X1 U11789 ( .A1(n14461), .A2(n14454), .ZN(n14456) );
  INV_X1 U11790 ( .A(n14699), .ZN(n12418) );
  NAND2_X1 U11791 ( .A1(n13918), .A2(n10166), .ZN(n13898) );
  AND2_X1 U11792 ( .A1(n9868), .A2(n13830), .ZN(n13918) );
  NAND2_X1 U11793 ( .A1(n9816), .A2(n12401), .ZN(n9995) );
  NAND2_X1 U11794 ( .A1(n20093), .A2(n20092), .ZN(n20091) );
  AND3_X1 U11795 ( .A1(n12035), .A2(n13243), .A3(n10181), .ZN(n13405) );
  NAND2_X1 U11796 ( .A1(n12112), .A2(n12099), .ZN(n14364) );
  AND2_X1 U11797 ( .A1(n12002), .A2(n13294), .ZN(n12425) );
  NAND2_X1 U11798 ( .A1(n9860), .A2(n12274), .ZN(n12305) );
  AND2_X1 U11799 ( .A1(n9821), .A2(n13175), .ZN(n20478) );
  OR2_X1 U11800 ( .A1(n9821), .A2(n20147), .ZN(n20539) );
  AND2_X1 U11801 ( .A1(n9823), .A2(n10128), .ZN(n10127) );
  INV_X1 U11802 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n10128) );
  NOR2_X1 U11803 ( .A1(n10149), .A2(n10147), .ZN(n10146) );
  NAND2_X1 U11804 ( .A1(n10150), .A2(n15007), .ZN(n10149) );
  NAND2_X1 U11805 ( .A1(n10148), .A2(n11208), .ZN(n10147) );
  NAND2_X1 U11806 ( .A1(n9925), .A2(n18880), .ZN(n10200) );
  OAI22_X1 U11807 ( .A1(n12850), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19904), 
        .B2(n12849), .ZN(n10188) );
  INV_X1 U11808 ( .A(n10820), .ZN(n11390) );
  NAND3_X1 U11809 ( .A1(n13136), .A2(n12513), .A3(n13137), .ZN(n10240) );
  INV_X1 U11810 ( .A(n10158), .ZN(n12806) );
  INV_X1 U11811 ( .A(n11438), .ZN(n12804) );
  NOR2_X1 U11812 ( .A1(n11520), .A2(n10125), .ZN(n10121) );
  CLKBUF_X1 U11813 ( .A(n11437), .Z(n19135) );
  NOR2_X1 U11814 ( .A1(n10195), .A2(n9892), .ZN(n10193) );
  INV_X1 U11815 ( .A(n12852), .ZN(n10194) );
  NAND2_X1 U11816 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10195) );
  OR2_X1 U11817 ( .A1(n11065), .A2(n15527), .ZN(n11066) );
  XNOR2_X1 U11818 ( .A(n11067), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16120) );
  NAND2_X1 U11819 ( .A1(n10297), .A2(n10296), .ZN(n10000) );
  NOR2_X1 U11820 ( .A1(n10300), .A2(n11774), .ZN(n10296) );
  INV_X1 U11821 ( .A(n11775), .ZN(n11283) );
  INV_X1 U11822 ( .A(n15106), .ZN(n11282) );
  NOR2_X1 U11823 ( .A1(n10323), .A2(n11374), .ZN(n10322) );
  NAND2_X1 U11824 ( .A1(n10324), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10323) );
  NAND2_X1 U11825 ( .A1(n9804), .A2(n10324), .ZN(n15113) );
  NAND2_X1 U11826 ( .A1(n11253), .A2(n10004), .ZN(n11270) );
  INV_X1 U11827 ( .A(n11192), .ZN(n9998) );
  AND2_X1 U11828 ( .A1(n18860), .A2(n11233), .ZN(n15195) );
  OR2_X1 U11829 ( .A1(n11685), .A2(n16152), .ZN(n11686) );
  AND2_X1 U11830 ( .A1(n10307), .A2(n16113), .ZN(n10306) );
  AND2_X1 U11831 ( .A1(n11170), .A2(n10308), .ZN(n10307) );
  INV_X1 U11832 ( .A(n15259), .ZN(n10308) );
  NAND2_X1 U11833 ( .A1(n11159), .A2(n9831), .ZN(n10309) );
  NAND2_X1 U11834 ( .A1(n10042), .A2(n10040), .ZN(n10045) );
  NAND2_X1 U11835 ( .A1(n10043), .A2(n10982), .ZN(n10042) );
  NAND2_X1 U11836 ( .A1(n10984), .A2(n13623), .ZN(n10043) );
  XNOR2_X1 U11837 ( .A(n12494), .B(n12495), .ZN(n13046) );
  INV_X1 U11838 ( .A(n19134), .ZN(n13032) );
  NAND2_X1 U11839 ( .A1(n19846), .A2(n19078), .ZN(n19441) );
  NAND2_X1 U11840 ( .A1(n19860), .A2(n19868), .ZN(n19502) );
  OR2_X1 U11841 ( .A1(n19846), .A2(n19878), .ZN(n19620) );
  OR2_X1 U11842 ( .A1(n19860), .A2(n19868), .ZN(n19705) );
  NOR2_X1 U11843 ( .A1(n16487), .A2(n16486), .ZN(n16485) );
  OR2_X1 U11844 ( .A1(n16609), .A2(n10012), .ZN(n10010) );
  OR2_X1 U11845 ( .A1(n17627), .A2(n16601), .ZN(n10012) );
  OR2_X1 U11846 ( .A1(n16609), .A2(n17627), .ZN(n10013) );
  NOR2_X1 U11847 ( .A1(n10120), .A2(n17174), .ZN(n10117) );
  NAND2_X1 U11848 ( .A1(n15656), .A2(n10107), .ZN(n16817) );
  NAND2_X1 U11849 ( .A1(n9906), .A2(n10108), .ZN(n10107) );
  INV_X1 U11850 ( .A(n15657), .ZN(n10108) );
  NOR2_X1 U11851 ( .A1(n18669), .A2(n18607), .ZN(n17416) );
  NAND2_X1 U11852 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10014) );
  NOR2_X1 U11853 ( .A1(n9832), .A2(n10033), .ZN(n10031) );
  NAND2_X1 U11854 ( .A1(n17682), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10645) );
  NOR2_X2 U11855 ( .A1(n21007), .A2(n17624), .ZN(n17599) );
  INV_X1 U11856 ( .A(n10022), .ZN(n17677) );
  AND2_X1 U11857 ( .A1(n17636), .A2(n9905), .ZN(n10094) );
  NAND2_X1 U11858 ( .A1(n9973), .A2(n9971), .ZN(n17991) );
  NAND2_X1 U11859 ( .A1(n17752), .A2(n9975), .ZN(n9973) );
  AOI21_X1 U11860 ( .B1(n9975), .B2(n9929), .A(n9972), .ZN(n9971) );
  INV_X1 U11861 ( .A(n17654), .ZN(n9972) );
  NAND2_X1 U11862 ( .A1(n9974), .A2(n9975), .ZN(n18017) );
  OR2_X1 U11863 ( .A1(n17752), .A2(n9929), .ZN(n9974) );
  OR2_X1 U11864 ( .A1(n17752), .A2(n18070), .ZN(n9976) );
  XNOR2_X1 U11865 ( .A(n10635), .B(n10636), .ZN(n17774) );
  OR2_X1 U11866 ( .A1(n17774), .A2(n18091), .ZN(n9970) );
  NOR2_X1 U11867 ( .A1(n17787), .A2(n10055), .ZN(n17772) );
  INV_X1 U11868 ( .A(n10056), .ZN(n10055) );
  OAI21_X1 U11869 ( .B1(n15657), .B2(n10598), .A(n16436), .ZN(n13969) );
  NAND2_X1 U11870 ( .A1(n13052), .A2(n13348), .ZN(n20826) );
  INV_X1 U11871 ( .A(n11986), .ZN(n20214) );
  NAND2_X1 U11872 ( .A1(n14221), .A2(n20145), .ZN(n14591) );
  AND2_X1 U11873 ( .A1(n11721), .A2(n12970), .ZN(n12973) );
  INV_X1 U11874 ( .A(n19062), .ZN(n19047) );
  AND2_X1 U11875 ( .A1(n19205), .A2(n19902), .ZN(n19062) );
  INV_X1 U11876 ( .A(n19868), .ZN(n19342) );
  NAND2_X1 U11877 ( .A1(n9824), .A2(n11433), .ZN(n14329) );
  OR2_X1 U11878 ( .A1(n12832), .A2(n11432), .ZN(n11433) );
  OR2_X1 U11879 ( .A1(n16024), .A2(n14984), .ZN(n12837) );
  NAND2_X1 U11880 ( .A1(n11787), .A2(n11720), .ZN(n14325) );
  OR2_X1 U11881 ( .A1(n12806), .A2(n11719), .ZN(n11720) );
  INV_X1 U11882 ( .A(n19878), .ZN(n19078) );
  OAI21_X1 U11883 ( .B1(n15315), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15113), .ZN(n15295) );
  NAND2_X1 U11884 ( .A1(n15317), .A2(n9787), .ZN(n15125) );
  NAND2_X1 U11885 ( .A1(n12980), .A2(n11417), .ZN(n16150) );
  AOI21_X1 U11886 ( .B1(n19085), .B2(n16192), .A(n11793), .ZN(n11794) );
  NAND2_X1 U11887 ( .A1(n9835), .A2(n10158), .ZN(n16020) );
  NAND2_X1 U11888 ( .A1(n12444), .A2(n12443), .ZN(n15296) );
  AOI21_X1 U11889 ( .B1(n16182), .B2(n15317), .A(n15316), .ZN(n9965) );
  INV_X1 U11890 ( .A(n16194), .ZN(n16182) );
  OR2_X1 U11891 ( .A1(n11779), .A2(n19891), .ZN(n16187) );
  INV_X1 U11892 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19883) );
  NAND2_X1 U11893 ( .A1(n19654), .A2(n19469), .ZN(n15596) );
  INV_X1 U11894 ( .A(n16471), .ZN(n10020) );
  OR2_X1 U11895 ( .A1(n16464), .A2(n10018), .ZN(n10017) );
  OAI21_X1 U11896 ( .B1(n16472), .B2(P3_EBX_REG_30__SCAN_IN), .A(n10019), .ZN(
        n10018) );
  NAND2_X1 U11897 ( .A1(n16767), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n10019) );
  NOR2_X2 U11898 ( .A1(n18515), .A2(n16812), .ZN(n16796) );
  NAND2_X1 U11899 ( .A1(n18638), .A2(n15738), .ZN(n17345) );
  INV_X1 U11900 ( .A(n15738), .ZN(n17349) );
  NAND2_X1 U11901 ( .A1(n10098), .A2(n16265), .ZN(n10047) );
  NAND2_X1 U11902 ( .A1(n16264), .A2(n10099), .ZN(n10105) );
  NOR2_X1 U11903 ( .A1(n16262), .A2(n16265), .ZN(n10099) );
  NAND2_X1 U11904 ( .A1(n10652), .A2(n9863), .ZN(n10653) );
  INV_X1 U11905 ( .A(n17470), .ZN(n17483) );
  NOR2_X2 U11906 ( .A1(n17849), .A2(n17327), .ZN(n17755) );
  INV_X1 U11907 ( .A(n17838), .ZN(n17849) );
  NAND2_X1 U11908 ( .A1(n9981), .A2(n9980), .ZN(n9979) );
  AOI21_X1 U11909 ( .B1(n16301), .B2(n18068), .A(n9920), .ZN(n9980) );
  NAND2_X1 U11910 ( .A1(n16302), .A2(n18066), .ZN(n9981) );
  OAI21_X1 U11911 ( .B1(n10100), .B2(n10484), .A(n12484), .ZN(n10103) );
  NOR2_X1 U11912 ( .A1(n12483), .A2(n12482), .ZN(n12484) );
  OR3_X1 U11913 ( .A1(n16262), .A2(n10104), .A3(n16265), .ZN(n10100) );
  OR2_X1 U11914 ( .A1(n16262), .A2(n10484), .ZN(n10098) );
  NOR2_X1 U11915 ( .A1(n12466), .A2(n18669), .ZN(n18134) );
  CLKBUF_X1 U11916 ( .A(n18134), .Z(n18150) );
  AOI22_X1 U11917 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U11918 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10744) );
  OR2_X1 U11919 ( .A1(n11398), .A2(n11097), .ZN(n11074) );
  NAND2_X1 U11920 ( .A1(n17344), .A2(n9983), .ZN(n10615) );
  NAND2_X1 U11921 ( .A1(n17352), .A2(n17844), .ZN(n9983) );
  OR2_X1 U11922 ( .A1(n10502), .A2(n10503), .ZN(n10498) );
  AND2_X2 U11923 ( .A1(n10159), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11825) );
  NAND2_X1 U11924 ( .A1(n10254), .A2(n12354), .ZN(n12367) );
  AND2_X1 U11925 ( .A1(n13669), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11940) );
  NOR2_X1 U11926 ( .A1(n12187), .A2(n12186), .ZN(n12297) );
  NAND2_X1 U11927 ( .A1(n12017), .A2(n12016), .ZN(n13092) );
  NAND2_X1 U11928 ( .A1(n11986), .A2(n12120), .ZN(n11993) );
  NOR2_X1 U11929 ( .A1(n11213), .A2(n10003), .ZN(n10002) );
  NAND2_X1 U11930 ( .A1(n10823), .A2(n10822), .ZN(n10276) );
  INV_X1 U11931 ( .A(n11735), .ZN(n10779) );
  NAND2_X1 U11932 ( .A1(n11003), .A2(n11002), .ZN(n11034) );
  NAND2_X1 U11933 ( .A1(n10990), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10895) );
  AOI22_X1 U11934 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19408), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10896) );
  NAND2_X1 U11935 ( .A1(n10799), .A2(n9940), .ZN(n10802) );
  NAND2_X1 U11936 ( .A1(n9958), .A2(n9941), .ZN(n9940) );
  AOI21_X1 U11937 ( .B1(n11464), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10798), 
        .ZN(n10799) );
  NOR2_X1 U11938 ( .A1(n10795), .A2(n19904), .ZN(n9941) );
  AOI21_X1 U11939 ( .B1(n10864), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10663) );
  NAND2_X1 U11940 ( .A1(n11438), .A2(n15625), .ZN(n10769) );
  AOI22_X1 U11941 ( .A1(n10864), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12639), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U11942 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10681) );
  NAND2_X1 U11943 ( .A1(n10616), .A2(n10618), .ZN(n10464) );
  INV_X1 U11944 ( .A(n17341), .ZN(n10616) );
  INV_X1 U11945 ( .A(n10615), .ZN(n10617) );
  NOR2_X1 U11946 ( .A1(n11808), .A2(n11807), .ZN(n11969) );
  INV_X1 U11947 ( .A(n12257), .ZN(n13056) );
  OR2_X1 U11948 ( .A1(n10269), .A2(n14396), .ZN(n10268) );
  NOR2_X1 U11949 ( .A1(n10260), .A2(n13962), .ZN(n10259) );
  INV_X1 U11950 ( .A(n14522), .ZN(n10260) );
  AND2_X1 U11951 ( .A1(n10272), .A2(n13868), .ZN(n10271) );
  OR2_X1 U11952 ( .A1(n10273), .A2(n10274), .ZN(n10272) );
  NAND2_X1 U11953 ( .A1(n10332), .A2(n9937), .ZN(n10248) );
  INV_X1 U11954 ( .A(n14708), .ZN(n10251) );
  AND2_X1 U11955 ( .A1(n10166), .A2(n10165), .ZN(n10164) );
  INV_X1 U11956 ( .A(n13897), .ZN(n10165) );
  NOR2_X1 U11957 ( .A1(n15981), .A2(n10168), .ZN(n13784) );
  NAND2_X1 U11958 ( .A1(n10170), .A2(n10169), .ZN(n10168) );
  INV_X1 U11959 ( .A(n15942), .ZN(n10169) );
  INV_X1 U11960 ( .A(n10171), .ZN(n10170) );
  NAND2_X1 U11961 ( .A1(n9881), .A2(n10174), .ZN(n10173) );
  OR2_X1 U11962 ( .A1(n12364), .A2(n12363), .ZN(n12384) );
  INV_X1 U11963 ( .A(n20092), .ZN(n10080) );
  INV_X1 U11964 ( .A(n12330), .ZN(n10078) );
  OR2_X1 U11965 ( .A1(n12321), .A2(n12320), .ZN(n12345) );
  INV_X1 U11966 ( .A(n12117), .ZN(n12105) );
  NAND2_X1 U11967 ( .A1(n13291), .A2(n12099), .ZN(n12109) );
  NAND2_X1 U11968 ( .A1(n10082), .A2(n10081), .ZN(n12261) );
  NAND2_X1 U11969 ( .A1(n11982), .A2(n11986), .ZN(n13171) );
  AND3_X1 U11970 ( .A1(n12012), .A2(n12011), .A3(n12010), .ZN(n13100) );
  AND2_X2 U11971 ( .A1(n11915), .A2(n13059), .ZN(n13118) );
  INV_X1 U11972 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20420) );
  OAI21_X1 U11973 ( .B1(n13662), .B2(n16002), .A(n20805), .ZN(n20150) );
  NAND2_X1 U11974 ( .A1(n12243), .A2(n12222), .ZN(n12377) );
  OR2_X1 U11975 ( .A1(n11808), .A2(n11805), .ZN(n11806) );
  CLKBUF_X1 U11976 ( .A(n11071), .Z(n11084) );
  NOR2_X1 U11977 ( .A1(n11266), .A2(n11263), .ZN(n10145) );
  INV_X1 U11978 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10130) );
  NOR2_X1 U11979 ( .A1(n11237), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11238) );
  INV_X1 U11980 ( .A(n11200), .ZN(n10148) );
  INV_X1 U11981 ( .A(n11197), .ZN(n10150) );
  NAND2_X1 U11982 ( .A1(n11212), .A2(n11195), .ZN(n11205) );
  NAND2_X1 U11983 ( .A1(n9800), .A2(n10002), .ZN(n11216) );
  AND2_X1 U11984 ( .A1(n10140), .A2(n18954), .ZN(n10139) );
  NAND2_X1 U11985 ( .A1(n9800), .A2(n11187), .ZN(n11214) );
  AND2_X1 U11986 ( .A1(n11172), .A2(n10140), .ZN(n11181) );
  INV_X1 U11987 ( .A(n11153), .ZN(n10141) );
  AND4_X1 U11988 ( .A1(n11132), .A2(n10142), .A3(n10144), .A4(n10141), .ZN(
        n11166) );
  NOR2_X1 U11989 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12633) );
  AND2_X1 U11990 ( .A1(n12535), .A2(n13758), .ZN(n10239) );
  NAND2_X1 U11991 ( .A1(n10876), .A2(n10875), .ZN(n10886) );
  INV_X1 U11992 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10196) );
  NOR2_X1 U11993 ( .A1(n11420), .A2(n10212), .ZN(n10211) );
  OR2_X1 U11994 ( .A1(n11419), .A2(n16106), .ZN(n11420) );
  INV_X1 U11995 ( .A(n10214), .ZN(n10212) );
  NOR2_X1 U11996 ( .A1(n15264), .A2(n10215), .ZN(n10214) );
  INV_X1 U11997 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10215) );
  INV_X1 U11998 ( .A(n12856), .ZN(n10213) );
  NOR2_X1 U11999 ( .A1(n13286), .A2(n13199), .ZN(n10281) );
  INV_X1 U12000 ( .A(n13158), .ZN(n11305) );
  AND2_X1 U12001 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10185) );
  INV_X1 U12002 ( .A(n11293), .ZN(n10075) );
  NAND2_X1 U12003 ( .A1(n10760), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10762) );
  XNOR2_X1 U12004 ( .A(n11286), .B(n11279), .ZN(n11280) );
  OAI21_X1 U12005 ( .B1(n10340), .B2(n12434), .A(n15105), .ZN(n10300) );
  NOR2_X1 U12006 ( .A1(n11069), .A2(n15297), .ZN(n10324) );
  INV_X1 U12007 ( .A(n15151), .ZN(n11252) );
  OR2_X1 U12008 ( .A1(n12438), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10343) );
  INV_X1 U12009 ( .A(n15131), .ZN(n10305) );
  NOR2_X1 U12010 ( .A1(n16038), .A2(n11539), .ZN(n11273) );
  NAND2_X1 U12011 ( .A1(n10320), .A2(n10316), .ZN(n15141) );
  NOR2_X1 U12012 ( .A1(n10317), .A2(n15342), .ZN(n10316) );
  INV_X1 U12013 ( .A(n10318), .ZN(n10317) );
  NOR2_X1 U12014 ( .A1(n10319), .A2(n15359), .ZN(n10318) );
  INV_X1 U12015 ( .A(n10321), .ZN(n10319) );
  NOR2_X1 U12016 ( .A1(n20968), .A2(n15372), .ZN(n10321) );
  INV_X1 U12017 ( .A(n9953), .ZN(n9952) );
  AND2_X1 U12018 ( .A1(n11178), .A2(n9954), .ZN(n9953) );
  INV_X1 U12019 ( .A(n15493), .ZN(n9954) );
  INV_X1 U12020 ( .A(n11784), .ZN(n11702) );
  INV_X1 U12021 ( .A(n11380), .ZN(n11314) );
  NAND2_X1 U12022 ( .A1(n11092), .A2(n10327), .ZN(n9942) );
  AND2_X1 U12023 ( .A1(n11305), .A2(n10289), .ZN(n10288) );
  INV_X1 U12024 ( .A(n13076), .ZN(n10289) );
  INV_X1 U12025 ( .A(n13159), .ZN(n10290) );
  NAND2_X1 U12026 ( .A1(n10956), .A2(n11515), .ZN(n10951) );
  AOI22_X1 U12027 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10988), .B1(
        n10987), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10846) );
  AND4_X1 U12028 ( .A1(n10928), .A2(n10927), .A3(n10926), .A4(n10925), .ZN(
        n10929) );
  AND4_X1 U12029 ( .A1(n10715), .A2(n10714), .A3(n10713), .A4(n10712), .ZN(
        n10716) );
  INV_X1 U12030 ( .A(n11409), .ZN(n11415) );
  AND4_X1 U12031 ( .A1(n13457), .A2(n10037), .A3(n15625), .A4(n13572), .ZN(
        n9962) );
  NOR2_X1 U12032 ( .A1(n17183), .A2(n10119), .ZN(n10118) );
  INV_X1 U12033 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n10119) );
  INV_X1 U12034 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16870) );
  OR2_X1 U12035 ( .A1(n10360), .A2(n18632), .ZN(n16871) );
  NOR2_X1 U12036 ( .A1(n10359), .A2(n18632), .ZN(n10417) );
  OR2_X1 U12037 ( .A1(n18633), .A2(n10361), .ZN(n16858) );
  NOR2_X1 U12038 ( .A1(n18633), .A2(n10360), .ZN(n10418) );
  NOR2_X1 U12039 ( .A1(n10363), .A2(n10360), .ZN(n10409) );
  NOR2_X1 U12040 ( .A1(n17477), .A2(n17471), .ZN(n10648) );
  AND2_X1 U12041 ( .A1(n10614), .A2(n10466), .ZN(n10468) );
  NOR2_X1 U12042 ( .A1(n17620), .A2(n10478), .ZN(n17579) );
  INV_X1 U12043 ( .A(n17967), .ZN(n10065) );
  OR2_X1 U12044 ( .A1(n9859), .A2(n17999), .ZN(n9975) );
  NOR2_X1 U12045 ( .A1(n12458), .A2(n18622), .ZN(n13976) );
  NAND2_X1 U12046 ( .A1(n10601), .A2(n10603), .ZN(n12458) );
  OR2_X1 U12047 ( .A1(n10595), .A2(n18621), .ZN(n15657) );
  OAI211_X1 U12048 ( .C1(n12166), .C2(n20169), .A(n12165), .B(n12164), .ZN(
        n12190) );
  NOR2_X1 U12049 ( .A1(n12161), .A2(n12160), .ZN(n12165) );
  AND2_X1 U12050 ( .A1(n14073), .A2(n14072), .ZN(n14496) );
  AND2_X1 U12051 ( .A1(n14052), .A2(n14051), .ZN(n14502) );
  NAND2_X1 U12052 ( .A1(n10256), .A2(n10257), .ZN(n10255) );
  INV_X1 U12053 ( .A(n14510), .ZN(n10256) );
  NAND2_X1 U12054 ( .A1(n10267), .A2(n14378), .ZN(n10266) );
  INV_X1 U12055 ( .A(n10268), .ZN(n10267) );
  NAND2_X1 U12056 ( .A1(n14176), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14180) );
  OAI21_X1 U12057 ( .B1(n10352), .B2(n14640), .A(n14198), .ZN(n14407) );
  OAI21_X1 U12058 ( .B1(n10352), .B2(n14657), .A(n14161), .ZN(n14430) );
  AND2_X1 U12059 ( .A1(n14665), .A2(n14282), .ZN(n14139) );
  NAND2_X1 U12060 ( .A1(n9814), .A2(n10264), .ZN(n14429) );
  NAND2_X1 U12061 ( .A1(n13675), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14118) );
  INV_X1 U12062 ( .A(n14089), .ZN(n13675) );
  OR2_X1 U12063 ( .A1(n14673), .A2(n10352), .ZN(n14120) );
  NAND2_X1 U12064 ( .A1(n9814), .A2(n14092), .ZN(n14462) );
  NAND2_X1 U12065 ( .A1(n13984), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13998) );
  AND2_X1 U12066 ( .A1(n13924), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13984) );
  NAND2_X1 U12067 ( .A1(n13878), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13942) );
  AND2_X1 U12068 ( .A1(n13851), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13878) );
  CLKBUF_X1 U12069 ( .A(n13893), .Z(n13894) );
  INV_X1 U12070 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13836) );
  AND2_X1 U12071 ( .A1(n13776), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13807) );
  OR2_X1 U12072 ( .A1(n13700), .A2(n13674), .ZN(n13733) );
  AND3_X1 U12073 ( .A1(n13704), .A2(n13703), .A3(n13702), .ZN(n13707) );
  CLKBUF_X1 U12074 ( .A(n13752), .Z(n13706) );
  NAND2_X1 U12075 ( .A1(n13650), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13700) );
  AND2_X1 U12076 ( .A1(n13637), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13650) );
  INV_X1 U12077 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13513) );
  NOR2_X1 U12078 ( .A1(n13511), .A2(n13513), .ZN(n13637) );
  INV_X1 U12079 ( .A(n13520), .ZN(n13524) );
  AND2_X1 U12080 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n13390), .ZN(
        n13484) );
  NAND2_X1 U12081 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13391) );
  NAND2_X1 U12082 ( .A1(n13463), .A2(n13462), .ZN(n13461) );
  NAND2_X1 U12083 ( .A1(n13240), .A2(n13239), .ZN(n13389) );
  INV_X1 U12084 ( .A(n13241), .ZN(n13240) );
  INV_X1 U12085 ( .A(n10245), .ZN(n10244) );
  OAI21_X1 U12086 ( .B1(n15852), .B2(n14798), .A(n9936), .ZN(n10245) );
  NOR2_X1 U12087 ( .A1(n14624), .A2(n14798), .ZN(n10076) );
  NOR2_X1 U12088 ( .A1(n14431), .A2(n14417), .ZN(n14418) );
  INV_X1 U12089 ( .A(n14653), .ZN(n9989) );
  INV_X1 U12090 ( .A(n14623), .ZN(n14661) );
  OR2_X1 U12091 ( .A1(n14841), .A2(n12133), .ZN(n14796) );
  AND2_X1 U12092 ( .A1(n14514), .A2(n9844), .ZN(n14461) );
  NAND2_X1 U12093 ( .A1(n14514), .A2(n10161), .ZN(n14497) );
  NAND2_X1 U12094 ( .A1(n14514), .A2(n14505), .ZN(n14506) );
  NAND2_X1 U12095 ( .A1(n12418), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14686) );
  NOR2_X1 U12096 ( .A1(n14520), .A2(n14512), .ZN(n14514) );
  OR2_X1 U12097 ( .A1(n14523), .A2(n14518), .ZN(n14520) );
  OR2_X1 U12098 ( .A1(n14525), .A2(n14526), .ZN(n14523) );
  AND2_X1 U12099 ( .A1(n13918), .A2(n10163), .ZN(n14885) );
  AND2_X1 U12100 ( .A1(n10164), .A2(n14883), .ZN(n10163) );
  AOI21_X1 U12101 ( .B1(n9994), .B2(n9992), .A(n9879), .ZN(n9991) );
  INV_X1 U12102 ( .A(n9994), .ZN(n9993) );
  OR2_X1 U12103 ( .A1(n15981), .A2(n10171), .ZN(n15943) );
  NOR2_X1 U12104 ( .A1(n15981), .A2(n10173), .ZN(n15967) );
  OR2_X1 U12105 ( .A1(n15981), .A2(n15980), .ZN(n15983) );
  NAND2_X1 U12106 ( .A1(n12045), .A2(n12044), .ZN(n15981) );
  INV_X1 U12107 ( .A(n13493), .ZN(n12044) );
  INV_X1 U12108 ( .A(n13494), .ZN(n12045) );
  NOR2_X1 U12109 ( .A1(n14915), .A2(n15930), .ZN(n14892) );
  XNOR2_X1 U12110 ( .A(n12035), .B(n13189), .ZN(n13726) );
  AND2_X1 U12111 ( .A1(n14868), .A2(n14870), .ZN(n15930) );
  NAND2_X1 U12112 ( .A1(n20824), .A2(n20150), .ZN(n20315) );
  NAND2_X1 U12113 ( .A1(n10246), .A2(n14925), .ZN(n20288) );
  INV_X1 U12114 ( .A(n20315), .ZN(n20218) );
  INV_X1 U12115 ( .A(n12250), .ZN(n20185) );
  INV_X1 U12116 ( .A(n20478), .ZN(n20617) );
  AOI21_X1 U12117 ( .B1(n20581), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20315), 
        .ZN(n20667) );
  AND2_X1 U12118 ( .A1(n11409), .A2(n11100), .ZN(n16226) );
  NAND2_X1 U12119 ( .A1(n9925), .A2(n16037), .ZN(n10207) );
  NAND2_X1 U12120 ( .A1(n10206), .A2(n9925), .ZN(n10205) );
  NAND2_X1 U12121 ( .A1(n11245), .A2(n9823), .ZN(n11259) );
  NAND2_X1 U12122 ( .A1(n10190), .A2(n9925), .ZN(n10186) );
  NAND2_X1 U12124 ( .A1(n10192), .A2(n10191), .ZN(n10190) );
  INV_X1 U12125 ( .A(n15163), .ZN(n10191) );
  OR2_X1 U12126 ( .A1(n19041), .A2(n15168), .ZN(n10192) );
  OAI21_X1 U12127 ( .B1(n11238), .B2(n11203), .A(n11239), .ZN(n11243) );
  INV_X1 U12128 ( .A(n11241), .ZN(n11239) );
  NOR2_X1 U12129 ( .A1(n15679), .A2(n15681), .ZN(n15680) );
  INV_X1 U12130 ( .A(n11237), .ZN(n10006) );
  OR2_X1 U12131 ( .A1(n18890), .A2(n19041), .ZN(n10201) );
  INV_X1 U12132 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11419) );
  AND2_X1 U12133 ( .A1(n11132), .A2(n11133), .ZN(n11148) );
  NOR3_X1 U12134 ( .A1(n12948), .A2(n12442), .A3(n9922), .ZN(n12832) );
  NAND2_X1 U12135 ( .A1(n14990), .A2(n10292), .ZN(n14975) );
  NAND2_X1 U12136 ( .A1(n11321), .A2(n11320), .ZN(n13287) );
  INV_X1 U12137 ( .A(n12742), .ZN(n10232) );
  NAND2_X1 U12138 ( .A1(n10231), .A2(n10230), .ZN(n14952) );
  OAI21_X1 U12139 ( .B1(n14957), .B2(n12742), .A(n12760), .ZN(n10230) );
  NAND2_X1 U12140 ( .A1(n10234), .A2(n10233), .ZN(n10231) );
  NOR2_X1 U12141 ( .A1(n12742), .A2(n12760), .ZN(n10233) );
  NAND2_X1 U12142 ( .A1(n14952), .A2(n14951), .ZN(n14950) );
  NAND2_X1 U12143 ( .A1(n14962), .A2(n14964), .ZN(n14963) );
  OAI211_X1 U12144 ( .C1(n10224), .C2(n10221), .A(n10220), .B(n10219), .ZN(
        n14983) );
  NOR2_X1 U12145 ( .A1(n10226), .A2(n10223), .ZN(n10224) );
  NOR2_X1 U12146 ( .A1(n15368), .A2(n15369), .ZN(n15367) );
  AND2_X1 U12147 ( .A1(n10153), .A2(n10152), .ZN(n10151) );
  INV_X1 U12148 ( .A(n15097), .ZN(n10152) );
  NAND2_X1 U12149 ( .A1(n15460), .A2(n10153), .ZN(n15419) );
  NAND2_X1 U12150 ( .A1(n15537), .A2(n10338), .ZN(n15522) );
  NAND2_X1 U12151 ( .A1(n10126), .A2(n10124), .ZN(n10123) );
  NOR2_X1 U12152 ( .A1(n13559), .A2(n10125), .ZN(n10124) );
  INV_X1 U12153 ( .A(n11520), .ZN(n10126) );
  INV_X1 U12154 ( .A(n12816), .ZN(n19101) );
  INV_X1 U12155 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n21083) );
  NAND2_X1 U12156 ( .A1(n12854), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12852) );
  NOR2_X1 U12157 ( .A1(n12856), .A2(n10210), .ZN(n12854) );
  NAND2_X1 U12158 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n10211), .ZN(
        n10210) );
  NOR2_X1 U12159 ( .A1(n12862), .A2(n10183), .ZN(n10182) );
  NAND2_X1 U12160 ( .A1(n10290), .A2(n11305), .ZN(n13161) );
  INV_X1 U12161 ( .A(n10838), .ZN(n13138) );
  NAND2_X1 U12162 ( .A1(n10297), .A2(n10299), .ZN(n11773) );
  INV_X1 U12163 ( .A(n10300), .ZN(n10299) );
  OR3_X1 U12164 ( .A1(n12896), .A2(n11539), .A3(n11386), .ZN(n11775) );
  INV_X1 U12165 ( .A(n10278), .ZN(n12951) );
  AND2_X1 U12166 ( .A1(n10278), .A2(n10277), .ZN(n12835) );
  INV_X1 U12167 ( .A(n12442), .ZN(n10277) );
  NOR2_X1 U12168 ( .A1(n12962), .A2(n11539), .ZN(n12439) );
  AND2_X1 U12169 ( .A1(n14990), .A2(n9927), .ZN(n14966) );
  INV_X1 U12170 ( .A(n14965), .ZN(n10291) );
  NAND2_X1 U12171 ( .A1(n10138), .A2(n10137), .ZN(n15069) );
  INV_X1 U12172 ( .A(n15067), .ZN(n10137) );
  NAND2_X1 U12173 ( .A1(n15367), .A2(n12938), .ZN(n12937) );
  CLKBUF_X1 U12174 ( .A(n15141), .Z(n15142) );
  NAND2_X1 U12175 ( .A1(n14990), .A2(n10294), .ZN(n14977) );
  NAND2_X1 U12176 ( .A1(n10071), .A2(n9825), .ZN(n10070) );
  AND2_X1 U12177 ( .A1(n15385), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15353) );
  NOR2_X1 U12178 ( .A1(n14999), .A2(n12922), .ZN(n14990) );
  OR2_X1 U12179 ( .A1(n14998), .A2(n15001), .ZN(n14999) );
  NAND2_X1 U12180 ( .A1(n15433), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10315) );
  AND2_X1 U12181 ( .A1(n13606), .A2(n9911), .ZN(n15017) );
  NAND2_X1 U12182 ( .A1(n15460), .A2(n10155), .ZN(n15417) );
  AND2_X1 U12183 ( .A1(n15460), .A2(n15448), .ZN(n15450) );
  NAND2_X1 U12184 ( .A1(n13606), .A2(n10284), .ZN(n15031) );
  NOR2_X1 U12185 ( .A1(n13585), .A2(n13586), .ZN(n13606) );
  AND3_X1 U12186 ( .A1(n11684), .A2(n11683), .A3(n11682), .ZN(n16152) );
  NAND2_X1 U12187 ( .A1(n15479), .A2(n11192), .ZN(n15176) );
  OR2_X1 U12188 ( .A1(n13413), .A2(n13468), .ZN(n13475) );
  OR2_X1 U12189 ( .A1(n13475), .A2(n13474), .ZN(n13585) );
  AND3_X1 U12190 ( .A1(n11624), .A2(n11623), .A3(n11622), .ZN(n15480) );
  NOR2_X1 U12191 ( .A1(n16174), .A2(n10134), .ZN(n16165) );
  AND2_X1 U12192 ( .A1(n11321), .A2(n9828), .ZN(n13415) );
  AND2_X1 U12193 ( .A1(n15481), .A2(n13596), .ZN(n15495) );
  OR2_X1 U12194 ( .A1(n11067), .A2(n11488), .ZN(n11068) );
  NOR2_X1 U12195 ( .A1(n13159), .A2(n10286), .ZN(n13142) );
  NAND2_X1 U12196 ( .A1(n10288), .A2(n10287), .ZN(n10286) );
  INV_X1 U12197 ( .A(n13128), .ZN(n10287) );
  NAND2_X1 U12198 ( .A1(n10290), .A2(n10288), .ZN(n13129) );
  AOI21_X1 U12199 ( .B1(n13426), .B2(n11289), .A(n21168), .ZN(n10301) );
  NAND2_X1 U12200 ( .A1(n11126), .A2(n21168), .ZN(n13544) );
  AND2_X1 U12201 ( .A1(n15437), .A2(n15443), .ZN(n15481) );
  NAND2_X1 U12202 ( .A1(n11499), .A2(n11498), .ZN(n13039) );
  XNOR2_X1 U12203 ( .A(n11509), .B(n11510), .ZN(n13081) );
  INV_X2 U12204 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15562) );
  AND2_X1 U12205 ( .A1(n10786), .A2(n12828), .ZN(n15582) );
  AND2_X1 U12206 ( .A1(n13135), .A2(n13163), .ZN(n13167) );
  NAND2_X1 U12207 ( .A1(n13136), .A2(n13137), .ZN(n13166) );
  INV_X1 U12208 ( .A(n15608), .ZN(n15646) );
  OR3_X1 U12209 ( .A1(n13565), .A2(n19270), .A3(n19654), .ZN(n13571) );
  OR2_X1 U12210 ( .A1(n19441), .A2(n19705), .ZN(n19463) );
  INV_X1 U12211 ( .A(n10990), .ZN(n19533) );
  OR2_X1 U12212 ( .A1(n19846), .A2(n19078), .ZN(n19650) );
  NAND2_X2 U12213 ( .A1(n9787), .A2(n19100), .ZN(n15650) );
  NOR2_X1 U12214 ( .A1(n18813), .A2(n16818), .ZN(n10599) );
  INV_X1 U12215 ( .A(n13975), .ZN(n18613) );
  OAI21_X1 U12216 ( .B1(n10509), .B2(n10610), .A(n10611), .ZN(n18607) );
  NOR3_X1 U12217 ( .A1(n16290), .A2(n17841), .A3(n10015), .ZN(n16286) );
  AND2_X1 U12218 ( .A1(n16516), .A2(n10009), .ZN(n16507) );
  NAND2_X1 U12219 ( .A1(n16453), .A2(n16452), .ZN(n16539) );
  INV_X1 U12220 ( .A(n17535), .ZN(n16452) );
  INV_X1 U12221 ( .A(n16541), .ZN(n16453) );
  AND2_X1 U12222 ( .A1(n16586), .A2(n10009), .ZN(n16580) );
  AND3_X1 U12223 ( .A1(n10010), .A2(n10009), .A3(n10011), .ZN(n16588) );
  OR2_X1 U12224 ( .A1(n16588), .A2(n17603), .ZN(n16586) );
  NAND2_X1 U12225 ( .A1(n9890), .A2(n17612), .ZN(n10011) );
  INV_X1 U12226 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n21066) );
  NOR2_X1 U12227 ( .A1(n16933), .A2(n10110), .ZN(n10109) );
  NOR2_X1 U12228 ( .A1(n16821), .A2(n16617), .ZN(n10114) );
  INV_X1 U12229 ( .A(n10405), .ZN(n10091) );
  NOR2_X1 U12230 ( .A1(n10361), .A2(n18632), .ZN(n10408) );
  AOI21_X1 U12231 ( .B1(n13973), .B2(n18665), .A(n18811), .ZN(n17358) );
  NOR2_X1 U12232 ( .A1(n17858), .A2(n12474), .ZN(n16277) );
  NOR2_X1 U12233 ( .A1(n16290), .A2(n17841), .ZN(n16285) );
  NAND2_X1 U12234 ( .A1(n17599), .A2(n10031), .ZN(n17517) );
  NOR2_X1 U12235 ( .A1(n10645), .A2(n10022), .ZN(n10026) );
  NOR2_X1 U12236 ( .A1(n21066), .A2(n17699), .ZN(n17682) );
  NAND2_X1 U12237 ( .A1(n17708), .A2(n17677), .ZN(n17693) );
  INV_X1 U12238 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16693) );
  INV_X1 U12239 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17709) );
  INV_X1 U12240 ( .A(n18036), .ZN(n16308) );
  AND2_X1 U12241 ( .A1(n10027), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17708) );
  INV_X1 U12242 ( .A(n17781), .ZN(n10027) );
  NAND2_X1 U12243 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10008) );
  INV_X1 U12244 ( .A(n16315), .ZN(n10058) );
  OAI221_X1 U12245 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17685), 
        .C1(n17871), .C2(n17526), .A(n17525), .ZN(n17506) );
  NAND2_X1 U12246 ( .A1(n17667), .A2(n9982), .ZN(n17858) );
  AND2_X1 U12247 ( .A1(n12471), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9982) );
  OR2_X1 U12248 ( .A1(n17915), .A2(n17523), .ZN(n17899) );
  NOR2_X1 U12249 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17581), .ZN(
        n17569) );
  NAND2_X1 U12250 ( .A1(n17753), .A2(n17735), .ZN(n17653) );
  OAI21_X1 U12251 ( .B1(n18621), .B2(n13969), .A(n18620), .ZN(n18637) );
  AND2_X1 U12252 ( .A1(n9976), .A2(n9859), .ZN(n18037) );
  AOI21_X1 U12253 ( .B1(n10643), .B2(n10642), .A(n10641), .ZN(n17752) );
  INV_X1 U12254 ( .A(n18609), .ZN(n12467) );
  OR2_X1 U12255 ( .A1(n10639), .A2(n10640), .ZN(n17760) );
  NOR2_X1 U12256 ( .A1(n17796), .A2(n10631), .ZN(n17786) );
  NOR2_X1 U12257 ( .A1(n17786), .A2(n17785), .ZN(n17784) );
  XNOR2_X1 U12258 ( .A(n10629), .B(n10630), .ZN(n17797) );
  NOR2_X1 U12259 ( .A1(n17797), .A2(n17798), .ZN(n17796) );
  INV_X1 U12260 ( .A(n17844), .ZN(n10622) );
  NAND2_X1 U12261 ( .A1(n18825), .A2(n13976), .ZN(n18612) );
  XNOR2_X1 U12262 ( .A(n10460), .B(n10459), .ZN(n17824) );
  NOR2_X1 U12263 ( .A1(n18076), .A2(n12454), .ZN(n18609) );
  NOR2_X1 U12264 ( .A1(n10596), .A2(n10604), .ZN(n13968) );
  INV_X1 U12265 ( .A(n18612), .ZN(n18635) );
  INV_X1 U12266 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18515) );
  NOR2_X1 U12267 ( .A1(n10584), .A2(n10583), .ZN(n18181) );
  NOR2_X1 U12268 ( .A1(n10522), .A2(n10521), .ZN(n18185) );
  INV_X1 U12269 ( .A(n10602), .ZN(n18190) );
  NOR2_X1 U12270 ( .A1(n10563), .A2(n10562), .ZN(n18194) );
  NAND2_X1 U12271 ( .A1(n18671), .A2(n18170), .ZN(n18251) );
  INV_X1 U12272 ( .A(n19101), .ZN(n19100) );
  INV_X1 U12273 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15803) );
  INV_X1 U12274 ( .A(n19947), .ZN(n19965) );
  AND2_X1 U12275 ( .A1(n12035), .A2(n10181), .ZN(n13244) );
  INV_X1 U12276 ( .A(n19988), .ZN(n20012) );
  INV_X1 U12277 ( .A(n19984), .ZN(n19996) );
  OR2_X1 U12278 ( .A1(n20826), .A2(n13666), .ZN(n19951) );
  INV_X1 U12279 ( .A(n19972), .ZN(n15816) );
  INV_X1 U12280 ( .A(n14529), .ZN(n20025) );
  INV_X1 U12281 ( .A(n20029), .ZN(n14527) );
  AND2_X1 U12282 ( .A1(n20029), .A2(n20214), .ZN(n20024) );
  INV_X1 U12283 ( .A(n20024), .ZN(n20015) );
  INV_X1 U12284 ( .A(n14600), .ZN(n14587) );
  AND2_X2 U12285 ( .A1(n13254), .A2(n13294), .ZN(n14600) );
  OR2_X1 U12286 ( .A1(n13253), .A2(n13252), .ZN(n13254) );
  OR2_X1 U12287 ( .A1(n14587), .A2(n13255), .ZN(n14602) );
  NAND2_X1 U12288 ( .A1(n13295), .A2(n13385), .ZN(n13296) );
  XNOR2_X1 U12289 ( .A(n13678), .B(n14371), .ZN(n14300) );
  OR2_X1 U12290 ( .A1(n20097), .A2(n13183), .ZN(n14742) );
  AND2_X1 U12291 ( .A1(n14742), .A2(n13223), .ZN(n15847) );
  INV_X1 U12292 ( .A(n14742), .ZN(n20090) );
  INV_X1 U12293 ( .A(n20097), .ZN(n19922) );
  NAND2_X1 U12294 ( .A1(n14363), .A2(n14362), .ZN(n14366) );
  NAND2_X1 U12295 ( .A1(n14383), .A2(n14384), .ZN(n14362) );
  OR2_X1 U12296 ( .A1(n14383), .A2(n12119), .ZN(n14482) );
  XNOR2_X1 U12297 ( .A(n9987), .B(n14808), .ZN(n14814) );
  NAND2_X1 U12298 ( .A1(n9990), .A2(n9988), .ZN(n9987) );
  OAI21_X1 U12299 ( .B1(n14623), .B2(n9989), .A(n10332), .ZN(n9988) );
  NAND2_X1 U12300 ( .A1(n14655), .A2(n15852), .ZN(n9990) );
  NAND2_X1 U12301 ( .A1(n10085), .A2(n15852), .ZN(n14678) );
  NAND2_X1 U12302 ( .A1(n12418), .A2(n10088), .ZN(n10085) );
  NAND2_X1 U12303 ( .A1(n13918), .A2(n13919), .ZN(n13872) );
  OR3_X1 U12304 ( .A1(n15953), .A2(n15913), .A3(n14872), .ZN(n15915) );
  NAND2_X1 U12305 ( .A1(n9995), .A2(n12403), .ZN(n13825) );
  NAND2_X1 U12306 ( .A1(n15873), .A2(n15872), .ZN(n15871) );
  NAND2_X1 U12307 ( .A1(n20091), .A2(n12330), .ZN(n15873) );
  INV_X1 U12308 ( .A(n15935), .ZN(n20123) );
  AND2_X1 U12309 ( .A1(n15930), .A2(n20132), .ZN(n15952) );
  INV_X1 U12310 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20581) );
  INV_X1 U12311 ( .A(n13208), .ZN(n13209) );
  NAND2_X1 U12312 ( .A1(n13335), .A2(n12177), .ZN(n13091) );
  NOR2_X1 U12313 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15992) );
  NOR2_X2 U12314 ( .A1(n20288), .A2(n20617), .ZN(n20304) );
  AND2_X1 U12315 ( .A1(n20515), .A2(n20478), .ZN(n20535) );
  INV_X1 U12316 ( .A(n20615), .ZN(n20574) );
  INV_X1 U12317 ( .A(n20555), .ZN(n20662) );
  INV_X1 U12318 ( .A(n20561), .ZN(n20682) );
  INV_X1 U12319 ( .A(n20564), .ZN(n20688) );
  INV_X1 U12320 ( .A(n20567), .ZN(n20694) );
  INV_X1 U12321 ( .A(n20570), .ZN(n20702) );
  INV_X1 U12322 ( .A(n20573), .ZN(n20708) );
  INV_X1 U12323 ( .A(n20579), .ZN(n20715) );
  AND2_X1 U12324 ( .A1(n15722), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15726) );
  NAND2_X1 U12325 ( .A1(n13293), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20805) );
  INV_X1 U12326 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19902) );
  OR2_X1 U12327 ( .A1(n16016), .A2(n12961), .ZN(n10202) );
  INV_X1 U12328 ( .A(n10203), .ZN(n12960) );
  AND2_X1 U12329 ( .A1(n10205), .A2(n10204), .ZN(n16026) );
  AND2_X1 U12330 ( .A1(n10207), .A2(n15134), .ZN(n10204) );
  INV_X1 U12331 ( .A(n16037), .ZN(n10208) );
  AND2_X1 U12332 ( .A1(n10198), .A2(n9912), .ZN(n18867) );
  INV_X1 U12333 ( .A(n18869), .ZN(n10197) );
  NOR2_X1 U12334 ( .A1(n19041), .A2(n18918), .ZN(n18903) );
  OR2_X1 U12335 ( .A1(n19895), .A2(n12894), .ZN(n19069) );
  INV_X1 U12336 ( .A(n19035), .ZN(n19080) );
  CLKBUF_X1 U12337 ( .A(n13588), .Z(n13608) );
  NAND2_X1 U12338 ( .A1(n13285), .A2(n12516), .ZN(n13408) );
  INV_X1 U12339 ( .A(n15038), .ZN(n15021) );
  XNOR2_X1 U12340 ( .A(n11787), .B(n11786), .ZN(n19085) );
  AND2_X1 U12341 ( .A1(n13035), .A2(n19100), .ZN(n19090) );
  AND2_X1 U12342 ( .A1(n13035), .A2(n19101), .ZN(n19089) );
  AND2_X1 U12343 ( .A1(n19121), .A2(n9931), .ZN(n19088) );
  NOR2_X1 U12344 ( .A1(n16174), .A2(n16175), .ZN(n15500) );
  NOR2_X1 U12345 ( .A1(n13267), .A2(n11520), .ZN(n13423) );
  OR2_X1 U12346 ( .A1(n19088), .A2(n13035), .ZN(n19123) );
  INV_X1 U12347 ( .A(n19092), .ZN(n19099) );
  INV_X1 U12348 ( .A(n19093), .ZN(n19127) );
  AND2_X1 U12349 ( .A1(n12973), .A2(n12887), .ZN(n19205) );
  AND2_X1 U12350 ( .A1(n12973), .A2(n19903), .ZN(n19231) );
  INV_X1 U12351 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15264) );
  INV_X1 U12352 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15276) );
  AND2_X1 U12353 ( .A1(n16150), .A2(n13018), .ZN(n16143) );
  INV_X1 U12354 ( .A(n9787), .ZN(n16130) );
  XNOR2_X1 U12355 ( .A(n9999), .B(n11291), .ZN(n11782) );
  NAND2_X1 U12356 ( .A1(n10000), .A2(n11284), .ZN(n9999) );
  AOI21_X1 U12357 ( .B1(n12900), .B2(n16192), .A(n10351), .ZN(n11772) );
  NAND2_X1 U12358 ( .A1(n10298), .A2(n11275), .ZN(n15107) );
  NAND2_X1 U12359 ( .A1(n11272), .A2(n10340), .ZN(n10298) );
  AOI21_X1 U12360 ( .B1(n15479), .B2(n10073), .A(n9825), .ZN(n15172) );
  NOR2_X1 U12361 ( .A1(n16163), .A2(n16155), .ZN(n15467) );
  NAND2_X1 U12363 ( .A1(n9955), .A2(n11178), .ZN(n15492) );
  NAND2_X1 U12364 ( .A1(n10309), .A2(n10306), .ZN(n9955) );
  AND2_X1 U12365 ( .A1(n10309), .A2(n10307), .ZN(n16111) );
  NAND2_X1 U12366 ( .A1(n10309), .A2(n11170), .ZN(n15260) );
  OR2_X1 U12367 ( .A1(n11779), .A2(n11724), .ZN(n16177) );
  NAND2_X1 U12368 ( .A1(n10039), .A2(n10040), .ZN(n10038) );
  INV_X1 U12369 ( .A(n16187), .ZN(n16196) );
  OR2_X1 U12370 ( .A1(n11779), .A2(n11466), .ZN(n16194) );
  INV_X1 U12371 ( .A(n16177), .ZN(n16192) );
  OR2_X1 U12372 ( .A1(n12494), .A2(n13037), .ZN(n19878) );
  INV_X1 U12373 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19873) );
  XNOR2_X1 U12374 ( .A(n13071), .B(n13072), .ZN(n19860) );
  XNOR2_X1 U12375 ( .A(n13048), .B(n13047), .ZN(n19868) );
  INV_X1 U12376 ( .A(n19350), .ZN(n19368) );
  INV_X1 U12377 ( .A(n19371), .ZN(n19396) );
  OAI21_X1 U12378 ( .B1(n19488), .B2(n19473), .A(n19707), .ZN(n19490) );
  OAI211_X1 U12379 ( .C1(n19661), .C2(n19660), .A(n19707), .B(n19659), .ZN(
        n19693) );
  NOR2_X2 U12380 ( .A1(n19620), .A2(n19619), .ZN(n19691) );
  INV_X1 U12381 ( .A(n19248), .ZN(n19701) );
  INV_X1 U12382 ( .A(n19251), .ZN(n19714) );
  INV_X1 U12383 ( .A(n19256), .ZN(n19726) );
  INV_X1 U12384 ( .A(n19261), .ZN(n19738) );
  INV_X1 U12385 ( .A(n19264), .ZN(n19744) );
  NOR2_X2 U12386 ( .A1(n19650), .A2(n19705), .ZN(n19755) );
  INV_X1 U12387 ( .A(n19269), .ZN(n19750) );
  AND2_X1 U12388 ( .A1(n12826), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16252) );
  AND2_X1 U12389 ( .A1(n16539), .A2(n10009), .ZN(n16526) );
  AND2_X1 U12390 ( .A1(n16567), .A2(n10009), .ZN(n16557) );
  NOR2_X1 U12391 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16592), .ZN(n16576) );
  AND2_X1 U12392 ( .A1(n10013), .A2(n10009), .ZN(n16600) );
  NAND2_X1 U12393 ( .A1(n10010), .A2(n10011), .ZN(n16599) );
  NOR2_X1 U12394 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16634), .ZN(n16620) );
  AOI21_X1 U12395 ( .B1(n16442), .B2(n16665), .A(n9890), .ZN(n16609) );
  NOR2_X1 U12396 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16655), .ZN(n16641) );
  NAND2_X1 U12397 ( .A1(n16790), .A2(n16466), .ZN(n16664) );
  INV_X1 U12398 ( .A(n16790), .ZN(n16756) );
  NAND2_X1 U12399 ( .A1(n16457), .A2(n18826), .ZN(n16800) );
  INV_X1 U12400 ( .A(n16775), .ZN(n16809) );
  INV_X1 U12401 ( .A(n17248), .ZN(n18206) );
  NOR2_X1 U12402 ( .A1(n21021), .A2(n16930), .ZN(n16929) );
  NAND3_X1 U12403 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n16963), .ZN(n16949) );
  INV_X1 U12404 ( .A(n16949), .ZN(n16955) );
  NAND2_X1 U12405 ( .A1(n16968), .A2(n9854), .ZN(n16960) );
  INV_X1 U12406 ( .A(n16960), .ZN(n16963) );
  NOR2_X1 U12407 ( .A1(n21069), .A2(n16993), .ZN(n16968) );
  AND2_X1 U12408 ( .A1(n17053), .A2(n10111), .ZN(n17005) );
  NOR2_X1 U12409 ( .A1(n17248), .A2(n10113), .ZN(n10111) );
  NAND2_X1 U12410 ( .A1(n17053), .A2(n10112), .ZN(n17017) );
  NAND2_X1 U12411 ( .A1(n17053), .A2(P3_EBX_REG_17__SCAN_IN), .ZN(n17019) );
  NOR2_X1 U12412 ( .A1(n16820), .A2(n17068), .ZN(n17053) );
  AND2_X1 U12413 ( .A1(n17136), .A2(n9852), .ZN(n17069) );
  NAND2_X1 U12414 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17069), .ZN(n17068) );
  NAND2_X1 U12415 ( .A1(n17136), .A2(n9849), .ZN(n17081) );
  NOR2_X1 U12416 ( .A1(n17111), .A2(n16688), .ZN(n10115) );
  NAND2_X1 U12417 ( .A1(n17136), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n17108) );
  INV_X1 U12418 ( .A(n17152), .ZN(n17124) );
  AND2_X1 U12419 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17124), .ZN(n17136) );
  AND2_X1 U12420 ( .A1(n17188), .A2(n10116), .ZN(n17153) );
  AND2_X1 U12421 ( .A1(n9850), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n10116) );
  NAND2_X1 U12422 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17153), .ZN(n17152) );
  NAND2_X1 U12423 ( .A1(n17188), .A2(n9850), .ZN(n17155) );
  NOR2_X1 U12424 ( .A1(n17195), .A2(n17191), .ZN(n17188) );
  NAND2_X1 U12425 ( .A1(n17188), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n17187) );
  INV_X1 U12426 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17195) );
  NAND2_X1 U12427 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17196), .ZN(n17191) );
  NOR2_X1 U12428 ( .A1(n17204), .A2(n17201), .ZN(n17196) );
  NAND2_X1 U12429 ( .A1(n9826), .A2(P3_EBX_REG_0__SCAN_IN), .ZN(n17204) );
  INV_X1 U12430 ( .A(n17214), .ZN(n17209) );
  NAND2_X1 U12431 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17228), .ZN(n17223) );
  NOR2_X1 U12432 ( .A1(n17365), .A2(n17233), .ZN(n17228) );
  NAND2_X1 U12433 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17234), .ZN(n17233) );
  NOR2_X1 U12434 ( .A1(n17248), .A2(n17243), .ZN(n17239) );
  NOR3_X1 U12435 ( .A1(n17281), .A2(n17249), .A3(n15662), .ZN(n17244) );
  INV_X1 U12436 ( .A(n17250), .ZN(n17279) );
  INV_X1 U12437 ( .A(n17254), .ZN(n17280) );
  NAND4_X1 U12438 ( .A1(n17320), .A2(P3_EAX_REG_11__SCAN_IN), .A3(
        P3_EAX_REG_9__SCAN_IN), .A4(n15661), .ZN(n17292) );
  NOR2_X1 U12439 ( .A1(n17349), .A2(n18206), .ZN(n17321) );
  NOR2_X1 U12440 ( .A1(n10382), .A2(n10381), .ZN(n17334) );
  AND3_X1 U12441 ( .A1(n10434), .A2(n10433), .A3(n10432), .ZN(n17337) );
  INV_X1 U12442 ( .A(n10090), .ZN(n17344) );
  INV_X1 U12443 ( .A(n17354), .ZN(n17348) );
  INV_X1 U12444 ( .A(n17321), .ZN(n17350) );
  AOI21_X1 U12445 ( .B1(n15659), .B2(n15658), .A(n18669), .ZN(n15738) );
  NOR2_X1 U12446 ( .A1(n18638), .A2(n17350), .ZN(n17354) );
  NAND2_X1 U12447 ( .A1(n17388), .A2(n17414), .ZN(n17385) );
  CLKBUF_X1 U12448 ( .A(n17456), .Z(n17465) );
  AND2_X1 U12449 ( .A1(n17599), .A2(n9887), .ZN(n17502) );
  INV_X1 U12450 ( .A(n17520), .ZN(n10030) );
  INV_X1 U12451 ( .A(n17988), .ZN(n17547) );
  NAND2_X1 U12452 ( .A1(n17599), .A2(n9827), .ZN(n17589) );
  NAND3_X1 U12453 ( .A1(n10024), .A2(n10023), .A3(n17677), .ZN(n17624) );
  INV_X1 U12454 ( .A(n10645), .ZN(n10024) );
  NOR2_X1 U12455 ( .A1(n17781), .A2(n10025), .ZN(n10023) );
  NAND2_X1 U12456 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n10646), .ZN(
        n10025) );
  NAND2_X1 U12457 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17640) );
  NAND2_X1 U12458 ( .A1(n17667), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17988) );
  INV_X1 U12459 ( .A(n17991), .ZN(n17667) );
  INV_X1 U12460 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17699) );
  INV_X1 U12461 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17710) );
  NOR2_X1 U12462 ( .A1(n10008), .A2(n17804), .ZN(n17783) );
  NAND2_X1 U12463 ( .A1(n17783), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17781) );
  INV_X1 U12464 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17804) );
  BUF_X1 U12465 ( .A(n10649), .Z(n18552) );
  INV_X1 U12466 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18779) );
  INV_X1 U12467 ( .A(n17834), .ZN(n17850) );
  INV_X1 U12468 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18661) );
  NAND2_X1 U12469 ( .A1(n10062), .A2(n10063), .ZN(n17630) );
  NOR2_X1 U12470 ( .A1(n17989), .A2(n17661), .ZN(n17982) );
  INV_X1 U12471 ( .A(n18015), .ZN(n18068) );
  INV_X1 U12472 ( .A(n10095), .ZN(n17766) );
  INV_X1 U12473 ( .A(n9970), .ZN(n17773) );
  INV_X1 U12474 ( .A(n17771), .ZN(n10053) );
  INV_X1 U12475 ( .A(n17772), .ZN(n10054) );
  INV_X1 U12476 ( .A(n10092), .ZN(n17800) );
  INV_X1 U12477 ( .A(n18156), .ZN(n18139) );
  INV_X1 U12478 ( .A(n18154), .ZN(n18141) );
  INV_X1 U12479 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18654) );
  INV_X2 U12480 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18796) );
  AND2_X1 U12481 ( .A1(n12912), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20145)
         );
  OAI21_X1 U12483 ( .B1(n14329), .B2(n19047), .A(n12898), .ZN(n12899) );
  AND2_X1 U12484 ( .A1(n12837), .A2(n12836), .ZN(n12838) );
  OAI21_X1 U12485 ( .B1(n16020), .B2(n19092), .A(n12823), .ZN(n12824) );
  NOR2_X1 U12486 ( .A1(n12844), .A2(n12843), .ZN(n12847) );
  AOI21_X1 U12487 ( .B1(n12450), .B2(n9787), .A(n12449), .ZN(n12451) );
  NOR2_X1 U12488 ( .A1(n15315), .A2(n16145), .ZN(n15127) );
  OAI21_X1 U12489 ( .B1(n15318), .B2(n16187), .A(n9963), .ZN(P2_U3019) );
  INV_X1 U12490 ( .A(n9965), .ZN(n9964) );
  NOR2_X1 U12491 ( .A1(n15315), .A2(n16199), .ZN(n9966) );
  OR2_X1 U12492 ( .A1(n16473), .A2(n9930), .ZN(n10021) );
  NOR2_X1 U12493 ( .A1(n10020), .A2(n10017), .ZN(n10016) );
  AOI211_X1 U12494 ( .C1(n16490), .C2(n16498), .A(n16489), .B(n16488), .ZN(
        n16491) );
  NOR2_X1 U12495 ( .A1(n10654), .A2(n10653), .ZN(n10655) );
  NAND2_X1 U12496 ( .A1(n10105), .A2(n10047), .ZN(n12468) );
  AOI21_X1 U12497 ( .B1(n17484), .B2(n17483), .A(n17482), .ZN(n17486) );
  OAI211_X1 U12498 ( .C1(n16307), .C2(n10104), .A(n9978), .B(n9977), .ZN(
        P3_U2831) );
  AOI21_X1 U12499 ( .B1(n16306), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n16305), .ZN(n9977) );
  NAND2_X1 U12500 ( .A1(n9979), .A2(n18150), .ZN(n9978) );
  NOR2_X1 U12501 ( .A1(n10104), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10097) );
  INV_X1 U12502 ( .A(n10418), .ZN(n10516) );
  AND3_X1 U12503 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n10184), .A3(
        n10185), .ZN(n12861) );
  INV_X1 U12504 ( .A(n10766), .ZN(n11467) );
  NAND2_X1 U12505 ( .A1(n14595), .A2(n10259), .ZN(n14516) );
  NAND2_X1 U12506 ( .A1(n10320), .A2(n10321), .ZN(n15159) );
  INV_X1 U12507 ( .A(n10320), .ZN(n15188) );
  OAI22_X1 U12508 ( .A1(n12959), .A2(n10202), .B1(n9925), .B2(n16016), .ZN(
        n16011) );
  INV_X2 U12509 ( .A(n10188), .ZN(n19041) );
  AND2_X1 U12510 ( .A1(n9847), .A2(n10129), .ZN(n9823) );
  AND2_X1 U12511 ( .A1(n10843), .A2(n10844), .ZN(n10986) );
  NOR2_X1 U12512 ( .A1(n15245), .A2(n11757), .ZN(n15236) );
  OR3_X1 U12513 ( .A1(n12948), .A2(n12442), .A3(n9921), .ZN(n9824) );
  INV_X1 U12514 ( .A(n10409), .ZN(n10544) );
  AND2_X1 U12515 ( .A1(n16817), .A2(n9904), .ZN(n9826) );
  NOR2_X1 U12516 ( .A1(n15188), .A2(n20968), .ZN(n15166) );
  AND2_X1 U12517 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9827) );
  AND2_X1 U12518 ( .A1(n10281), .A2(n13313), .ZN(n9828) );
  AND2_X1 U12519 ( .A1(n10059), .A2(n10058), .ZN(n9829) );
  INV_X1 U12520 ( .A(n15872), .ZN(n10243) );
  AND2_X1 U12521 ( .A1(n13782), .A2(n13781), .ZN(n13867) );
  INV_X1 U12522 ( .A(n10209), .ZN(n16036) );
  XOR2_X1 U12523 ( .A(n11070), .B(n12849), .Z(n9830) );
  AND2_X1 U12524 ( .A1(n10203), .A2(n9925), .ZN(n16015) );
  AND2_X1 U12525 ( .A1(n11158), .A2(n9901), .ZN(n9831) );
  NAND2_X1 U12526 ( .A1(n17567), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9832) );
  AND4_X1 U12527 ( .A1(n11001), .A2(n11000), .A3(n10999), .A4(n10998), .ZN(
        n9833) );
  AND2_X1 U12528 ( .A1(n17735), .A2(n10065), .ZN(n9834) );
  NAND2_X1 U12529 ( .A1(n9883), .A2(n12805), .ZN(n9835) );
  AND3_X1 U12530 ( .A1(n14677), .A2(n9811), .A3(n9936), .ZN(n14622) );
  AND2_X1 U12532 ( .A1(n10002), .A2(n9919), .ZN(n9837) );
  AND2_X1 U12533 ( .A1(n9828), .A2(n13414), .ZN(n9838) );
  AND2_X1 U12534 ( .A1(n9829), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9839) );
  INV_X1 U12535 ( .A(n18078), .ZN(n10104) );
  NAND2_X1 U12536 ( .A1(n10213), .A2(n10214), .ZN(n12855) );
  NAND2_X1 U12537 ( .A1(n10194), .A2(n10193), .ZN(n12867) );
  NAND2_X1 U12538 ( .A1(n13610), .A2(n10239), .ZN(n13757) );
  NAND2_X1 U12539 ( .A1(n10122), .A2(n10121), .ZN(n13424) );
  OR2_X1 U12540 ( .A1(n12852), .A2(n9892), .ZN(n9840) );
  AND2_X1 U12541 ( .A1(n11421), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9841) );
  AND2_X1 U12542 ( .A1(n10161), .A2(n10160), .ZN(n9842) );
  OAI211_X1 U12543 ( .C1(n11039), .C2(n11041), .A(n11037), .B(n11038), .ZN(
        n15531) );
  NOR2_X1 U12544 ( .A1(n15680), .A2(n19041), .ZN(n12933) );
  INV_X1 U12545 ( .A(n10201), .ZN(n18879) );
  AND2_X1 U12546 ( .A1(n9907), .A2(n12516), .ZN(n9843) );
  AND2_X1 U12547 ( .A1(n9842), .A2(n14459), .ZN(n9844) );
  AND2_X1 U12548 ( .A1(n12514), .A2(n12515), .ZN(n9845) );
  AND2_X1 U12549 ( .A1(n9841), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9846) );
  AND2_X1 U12550 ( .A1(n11244), .A2(n10130), .ZN(n9847) );
  AND2_X1 U12551 ( .A1(n12817), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n9848) );
  AND2_X1 U12552 ( .A1(n10115), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n9849) );
  AND2_X1 U12553 ( .A1(n10118), .A2(n10117), .ZN(n9850) );
  AND2_X1 U12554 ( .A1(n11766), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9851) );
  AND2_X1 U12555 ( .A1(n9849), .A2(P3_EBX_REG_14__SCAN_IN), .ZN(n9852) );
  AND2_X1 U12556 ( .A1(n9851), .A2(n9938), .ZN(n9853) );
  AND2_X1 U12557 ( .A1(n10109), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n9854) );
  AND2_X1 U12558 ( .A1(n10845), .A2(n10844), .ZN(n10987) );
  NAND2_X1 U12559 ( .A1(n15262), .A2(n9851), .ZN(n15245) );
  NAND2_X1 U12560 ( .A1(n11245), .A2(n10127), .ZN(n9855) );
  NAND2_X1 U12561 ( .A1(n11984), .A2(n12256), .ZN(n11989) );
  INV_X1 U12562 ( .A(n14404), .ZN(n10179) );
  OR3_X1 U12563 ( .A1(n16290), .A2(n17841), .A3(n10014), .ZN(n9856) );
  AND2_X1 U12564 ( .A1(n10888), .A2(n10887), .ZN(n9857) );
  OR2_X1 U12565 ( .A1(n14406), .A2(n10266), .ZN(n9858) );
  NAND2_X1 U12566 ( .A1(n15262), .A2(n11766), .ZN(n16080) );
  NAND2_X1 U12567 ( .A1(n10185), .A2(n10184), .ZN(n12860) );
  OR2_X1 U12568 ( .A1(n10638), .A2(n10642), .ZN(n9859) );
  NAND2_X1 U12569 ( .A1(n15262), .A2(n11755), .ZN(n15474) );
  NOR2_X1 U12570 ( .A1(n13961), .A2(n13962), .ZN(n13997) );
  AND2_X1 U12571 ( .A1(n10320), .A2(n10318), .ZN(n9861) );
  OR2_X1 U12572 ( .A1(n15245), .A2(n10315), .ZN(n15224) );
  INV_X1 U12573 ( .A(n10398), .ZN(n10511) );
  NAND2_X1 U12574 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10469), .ZN(
        n9862) );
  OR2_X1 U12575 ( .A1(n17496), .A2(n12479), .ZN(n9863) );
  AND2_X1 U12576 ( .A1(n10251), .A2(n10248), .ZN(n9864) );
  AND2_X1 U12577 ( .A1(n9814), .A2(n10265), .ZN(n14442) );
  AND2_X1 U12578 ( .A1(n10669), .A2(n10668), .ZN(n9865) );
  AND2_X1 U12579 ( .A1(n10845), .A2(n10840), .ZN(n10996) );
  OR3_X1 U12580 ( .A1(n12831), .A2(n14304), .A3(n15038), .ZN(n9866) );
  INV_X1 U12581 ( .A(n10471), .ZN(n10096) );
  OR2_X1 U12582 ( .A1(n15295), .A2(n16145), .ZN(n9867) );
  AND2_X1 U12583 ( .A1(n13784), .A2(n12065), .ZN(n9868) );
  NAND2_X1 U12584 ( .A1(n15262), .A2(n9853), .ZN(n15216) );
  NAND2_X1 U12585 ( .A1(n9957), .A2(n11253), .ZN(n15130) );
  NAND2_X1 U12586 ( .A1(n12488), .A2(n12487), .ZN(n12494) );
  AND4_X1 U12587 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(
        n9869) );
  NAND2_X1 U12588 ( .A1(n11245), .A2(n9847), .ZN(n9870) );
  AND2_X1 U12589 ( .A1(n10845), .A2(n10839), .ZN(n10995) );
  NOR2_X1 U12590 ( .A1(n12944), .A2(n19041), .ZN(n12959) );
  OR3_X1 U12591 ( .A1(n12831), .A2(n14304), .A3(n19093), .ZN(n9871) );
  AND4_X1 U12592 ( .A1(n10834), .A2(n10837), .A3(n10835), .A4(n10836), .ZN(
        n9872) );
  AND2_X1 U12593 ( .A1(n11443), .A2(n11467), .ZN(n11395) );
  NAND2_X1 U12594 ( .A1(n10045), .A2(n10044), .ZN(n11039) );
  OR2_X1 U12595 ( .A1(n10463), .A2(n10462), .ZN(n9873) );
  OR2_X1 U12596 ( .A1(n10635), .A2(n10636), .ZN(n9874) );
  AOI21_X1 U12597 ( .B1(n18860), .B2(n11289), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15196) );
  AND2_X1 U12598 ( .A1(n11500), .A2(n10036), .ZN(n9875) );
  NAND2_X1 U12599 ( .A1(n9869), .A2(n9833), .ZN(n11002) );
  INV_X1 U12600 ( .A(n11002), .ZN(n9944) );
  OR2_X1 U12601 ( .A1(n10470), .A2(n10096), .ZN(n9876) );
  NAND2_X1 U12602 ( .A1(n9995), .A2(n9994), .ZN(n14749) );
  INV_X1 U12603 ( .A(n10138), .ZN(n15079) );
  NOR2_X1 U12604 ( .A1(n12937), .A2(n15080), .ZN(n10138) );
  AND2_X1 U12605 ( .A1(n9864), .A2(n10250), .ZN(n9877) );
  AND2_X1 U12606 ( .A1(n17504), .A2(n9829), .ZN(n9878) );
  AND2_X1 U12607 ( .A1(n15852), .A2(n15951), .ZN(n9879) );
  AND2_X1 U12608 ( .A1(n10832), .A2(n12485), .ZN(n10840) );
  INV_X1 U12609 ( .A(n10225), .ZN(n12677) );
  AND2_X1 U12610 ( .A1(n12352), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9880) );
  AND2_X1 U12611 ( .A1(n15965), .A2(n15964), .ZN(n9881) );
  INV_X1 U12612 ( .A(n10033), .ZN(n10032) );
  NAND2_X1 U12613 ( .A1(n9827), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10033) );
  AND2_X1 U12614 ( .A1(n13039), .A2(n13038), .ZN(n11509) );
  INV_X2 U12615 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10676) );
  AND2_X1 U12616 ( .A1(n15640), .A2(n10037), .ZN(n9882) );
  NAND2_X1 U12617 ( .A1(n13782), .A2(n10273), .ZN(n13865) );
  OR2_X1 U12618 ( .A1(n15118), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9967) );
  OR2_X1 U12619 ( .A1(n12952), .A2(n12964), .ZN(n9883) );
  NAND2_X1 U12620 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12862) );
  INV_X1 U12621 ( .A(n12862), .ZN(n10184) );
  AND3_X1 U12622 ( .A1(n10302), .A2(n10305), .A3(n10343), .ZN(n9884) );
  OR2_X1 U12623 ( .A1(n17798), .A2(n10465), .ZN(n9885) );
  OR2_X1 U12624 ( .A1(n15852), .A2(n15951), .ZN(n9886) );
  AND2_X1 U12625 ( .A1(n10031), .A2(n10030), .ZN(n9887) );
  AND2_X1 U12626 ( .A1(n11251), .A2(n15342), .ZN(n9888) );
  NAND2_X1 U12627 ( .A1(n14595), .A2(n10257), .ZN(n10261) );
  NAND2_X1 U12628 ( .A1(n10750), .A2(n10749), .ZN(n10766) );
  AND2_X1 U12629 ( .A1(n17490), .A2(n10483), .ZN(n16262) );
  AND2_X1 U12630 ( .A1(n15129), .A2(n10322), .ZN(n15112) );
  AND2_X1 U12631 ( .A1(n10141), .A2(n11164), .ZN(n9889) );
  INV_X2 U12632 ( .A(n13529), .ZN(n10867) );
  XOR2_X2 U12633 ( .A(n9856), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .Z(n9890)
         );
  INV_X1 U12634 ( .A(n9890), .ZN(n10009) );
  NAND2_X1 U12635 ( .A1(n11468), .A2(n19903), .ZN(n11681) );
  NAND2_X1 U12636 ( .A1(n10026), .A2(n17708), .ZN(n9891) );
  OR2_X1 U12637 ( .A1(n21083), .A2(n10196), .ZN(n9892) );
  AND2_X1 U12638 ( .A1(n17599), .A2(n10032), .ZN(n9893) );
  INV_X1 U12639 ( .A(n10333), .ZN(n10221) );
  OR2_X1 U12640 ( .A1(n16174), .A2(n10135), .ZN(n9894) );
  NAND2_X1 U12641 ( .A1(n13606), .A2(n13605), .ZN(n13604) );
  AND2_X1 U12642 ( .A1(n14514), .A2(n9842), .ZN(n9895) );
  AND2_X1 U12643 ( .A1(n13606), .A2(n10282), .ZN(n9896) );
  NOR2_X1 U12644 ( .A1(n12858), .A2(n15276), .ZN(n12859) );
  NOR2_X1 U12645 ( .A1(n12856), .A2(n15264), .ZN(n12857) );
  NOR2_X1 U12646 ( .A1(n12852), .A2(n21083), .ZN(n12853) );
  AND2_X1 U12647 ( .A1(n16968), .A2(n10109), .ZN(n9897) );
  AND2_X1 U12648 ( .A1(n16968), .A2(P3_EBX_REG_22__SCAN_IN), .ZN(n9898) );
  AND2_X1 U12649 ( .A1(n12155), .A2(n11985), .ZN(n11988) );
  AND2_X1 U12650 ( .A1(n14990), .A2(n14989), .ZN(n9899) );
  AND2_X1 U12651 ( .A1(n17053), .A2(n10114), .ZN(n9900) );
  NOR2_X1 U12652 ( .A1(n16126), .A2(n16123), .ZN(n9901) );
  AND2_X1 U12653 ( .A1(n13610), .A2(n12535), .ZN(n13756) );
  XNOR2_X1 U12654 ( .A(n9824), .B(n11392), .ZN(n11783) );
  INV_X1 U12655 ( .A(n15169), .ZN(n10072) );
  AND2_X1 U12656 ( .A1(n9843), .A2(n12517), .ZN(n9902) );
  INV_X1 U12657 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10495) );
  XNOR2_X1 U12658 ( .A(n12717), .B(n12718), .ZN(n14962) );
  NAND2_X1 U12659 ( .A1(n10213), .A2(n10211), .ZN(n9903) );
  NAND2_X1 U12660 ( .A1(n10038), .A2(n10043), .ZN(n13617) );
  INV_X1 U12661 ( .A(n13426), .ZN(n10074) );
  AND3_X1 U12662 ( .A1(n16819), .A2(n16818), .A3(n18663), .ZN(n9904) );
  OR2_X1 U12663 ( .A1(n11162), .A2(n12817), .ZN(n11257) );
  INV_X1 U12664 ( .A(n13199), .ZN(n11320) );
  OR2_X1 U12665 ( .A1(n17685), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9905) );
  AND3_X1 U12666 ( .A1(n18190), .A2(n18206), .A3(n15663), .ZN(n9906) );
  INV_X1 U12667 ( .A(n14492), .ZN(n14092) );
  INV_X1 U12668 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19904) );
  AND2_X1 U12669 ( .A1(n13312), .A2(n13411), .ZN(n9907) );
  NAND2_X1 U12670 ( .A1(n10961), .A2(n10960), .ZN(n10982) );
  INV_X1 U12671 ( .A(n10982), .ZN(n10039) );
  OR2_X1 U12672 ( .A1(n14329), .A2(n16194), .ZN(n9908) );
  OR2_X1 U12673 ( .A1(n12297), .A2(n12243), .ZN(n9909) );
  AND2_X1 U12674 ( .A1(n10209), .A2(n10208), .ZN(n9910) );
  AND2_X1 U12675 ( .A1(n10282), .A2(n15015), .ZN(n9911) );
  AND2_X1 U12676 ( .A1(n10200), .A2(n10197), .ZN(n9912) );
  AND2_X1 U12677 ( .A1(n10239), .A2(n12568), .ZN(n9913) );
  AND2_X1 U12678 ( .A1(n9902), .A2(n12518), .ZN(n9914) );
  INV_X1 U12679 ( .A(n10337), .ZN(n10084) );
  AND2_X1 U12680 ( .A1(n10951), .A2(n10887), .ZN(n9915) );
  INV_X1 U12681 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19469) );
  INV_X1 U12682 ( .A(n10352), .ZN(n14282) );
  AND3_X1 U12683 ( .A1(n10240), .A2(n13135), .A3(n12514), .ZN(n13075) );
  AND2_X1 U12684 ( .A1(n13285), .A2(n9843), .ZN(n13409) );
  INV_X1 U12685 ( .A(n13267), .ZN(n10122) );
  NOR3_X1 U12686 ( .A1(n12852), .A2(n9892), .A3(n15234), .ZN(n12866) );
  AND2_X1 U12687 ( .A1(n13285), .A2(n9902), .ZN(n13477) );
  NAND2_X1 U12688 ( .A1(n12870), .A2(n9841), .ZN(n12874) );
  NOR2_X1 U12689 ( .A1(n12867), .A2(n15214), .ZN(n12851) );
  NAND2_X1 U12690 ( .A1(n17188), .A2(n10118), .ZN(n9916) );
  INV_X1 U12691 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10216) );
  INV_X1 U12692 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10159) );
  OR2_X1 U12693 ( .A1(n11779), .A2(n19885), .ZN(n16199) );
  INV_X1 U12694 ( .A(n16199), .ZN(n16183) );
  AND2_X1 U12695 ( .A1(n12870), .A2(n11421), .ZN(n12872) );
  AND2_X1 U12696 ( .A1(n13918), .A2(n10164), .ZN(n9917) );
  AND2_X1 U12697 ( .A1(n11321), .A2(n10281), .ZN(n9918) );
  OR2_X1 U12698 ( .A1(n11236), .A2(n11194), .ZN(n9919) );
  INV_X1 U12699 ( .A(n11187), .ZN(n10003) );
  AND4_X1 U12700 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16304), .A3(
        n18778), .A4(n16303), .ZN(n9920) );
  OR2_X1 U12701 ( .A1(n12949), .A2(n10279), .ZN(n9921) );
  OR2_X1 U12702 ( .A1(n12949), .A2(n10280), .ZN(n9922) );
  AND2_X1 U12703 ( .A1(n13118), .A2(n13669), .ZN(n12141) );
  INV_X1 U12704 ( .A(n15003), .ZN(n10223) );
  NAND2_X1 U12705 ( .A1(n11455), .A2(n9942), .ZN(n11722) );
  AND2_X1 U12706 ( .A1(n11185), .A2(n15497), .ZN(n9923) );
  AND2_X1 U12707 ( .A1(n17136), .A2(n10115), .ZN(n9924) );
  INV_X1 U12708 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9984) );
  AND2_X1 U12710 ( .A1(n10054), .A2(n10053), .ZN(n9926) );
  INV_X1 U12711 ( .A(n14405), .ZN(n10180) );
  AND2_X1 U12712 ( .A1(n12851), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12870) );
  INV_X1 U12713 ( .A(n15980), .ZN(n10174) );
  AND2_X1 U12714 ( .A1(n10292), .A2(n10291), .ZN(n9927) );
  AND2_X1 U12715 ( .A1(n10201), .A2(n15227), .ZN(n9928) );
  INV_X1 U12716 ( .A(n10396), .ZN(n16859) );
  INV_X1 U12717 ( .A(n17164), .ZN(n16884) );
  INV_X1 U12718 ( .A(n16145), .ZN(n19241) );
  NAND2_X1 U12719 ( .A1(n12250), .A2(n12026), .ZN(n14382) );
  NOR2_X1 U12721 ( .A1(n12876), .A2(n11422), .ZN(n12445) );
  INV_X1 U12722 ( .A(n14989), .ZN(n10295) );
  AND2_X1 U12723 ( .A1(n12445), .A2(n11423), .ZN(n12840) );
  OR2_X1 U12724 ( .A1(n17999), .A2(n18070), .ZN(n9929) );
  XNOR2_X1 U12725 ( .A(n11425), .B(n11424), .ZN(n12850) );
  OR2_X1 U12726 ( .A1(n16799), .A2(n16474), .ZN(n9930) );
  AND2_X1 U12727 ( .A1(n12817), .A2(n10034), .ZN(n9931) );
  AND3_X1 U12728 ( .A1(n10157), .A2(n12953), .A3(n10156), .ZN(n9932) );
  AND2_X1 U12729 ( .A1(n10145), .A2(n11277), .ZN(n9933) );
  NOR2_X1 U12730 ( .A1(n20545), .A2(n20363), .ZN(n9934) );
  NOR2_X1 U12731 ( .A1(n20545), .A2(n20659), .ZN(n9935) );
  AND2_X1 U12732 ( .A1(n14653), .A2(n14808), .ZN(n9936) );
  INV_X1 U12733 ( .A(n10089), .ZN(n10088) );
  NAND3_X1 U12734 ( .A1(n14860), .A2(n14863), .A3(n15892), .ZN(n9937) );
  AND2_X1 U12735 ( .A1(n10314), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9938) );
  INV_X1 U12736 ( .A(n10113), .ZN(n10112) );
  NAND2_X1 U12737 ( .A1(n10114), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n10113) );
  INV_X1 U12738 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n10120) );
  INV_X1 U12739 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n10110) );
  INV_X1 U12740 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10015) );
  INV_X1 U12741 ( .A(n10315), .ZN(n10314) );
  NOR2_X1 U12742 ( .A1(n14995), .A2(n10229), .ZN(n10228) );
  NOR2_X1 U12743 ( .A1(n14994), .A2(n14995), .ZN(n14987) );
  NOR2_X2 U12744 ( .A1(n19220), .A2(n19536), .ZN(n19745) );
  OAI221_X2 U12745 ( .B1(n19900), .B2(n16252), .C1(n19140), .C2(n16252), .A(
        n19904), .ZN(n19536) );
  OAI22_X2 U12746 ( .A1(n21115), .A2(n20210), .B1(n14590), .B2(n20212), .ZN(
        n20672) );
  OAI22_X2 U12747 ( .A1(n20182), .A2(n20210), .B1(n20181), .B2(n20212), .ZN(
        n20690) );
  OAI22_X2 U12748 ( .A1(n20189), .A2(n20212), .B1(n21006), .B2(n20210), .ZN(
        n20696) );
  NAND2_X1 U12749 ( .A1(n20096), .A2(n20144), .ZN(n20210) );
  OAI22_X2 U12750 ( .A1(n20191), .A2(n20212), .B1(n20190), .B2(n20210), .ZN(
        n20642) );
  NOR3_X2 U12751 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20660), .A3(
        n20659), .ZN(n20651) );
  NOR3_X2 U12752 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18509), .A3(
        n18387), .ZN(n18359) );
  OAI22_X2 U12753 ( .A1(n20184), .A2(n20212), .B1(n20183), .B2(n20210), .ZN(
        n20638) );
  OAI22_X2 U12754 ( .A1(n20149), .A2(n20212), .B1(n20148), .B2(n20210), .ZN(
        n20630) );
  NOR3_X4 U12755 ( .A1(n18650), .A2(n18653), .A3(n18644), .ZN(n18600) );
  NAND2_X2 U12756 ( .A1(n12890), .A2(n12889), .ZN(n19063) );
  NOR2_X2 U12757 ( .A1(n20215), .A2(n20199), .ZN(n20703) );
  NAND2_X1 U12758 ( .A1(n20151), .A2(n20150), .ZN(n20215) );
  AND2_X4 U12759 ( .A1(n10879), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10866) );
  AND2_X2 U12760 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10879) );
  AND2_X4 U12761 ( .A1(n10856), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12632) );
  NOR2_X2 U12762 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10856) );
  NAND3_X1 U12763 ( .A1(n11455), .A2(n9942), .A3(n16231), .ZN(n10783) );
  NAND2_X1 U12764 ( .A1(n10691), .A2(n10690), .ZN(n10755) );
  INV_X2 U12765 ( .A(n10755), .ZN(n13457) );
  NAND2_X1 U12766 ( .A1(n13457), .A2(n10037), .ZN(n9946) );
  NAND2_X2 U12767 ( .A1(n9948), .A2(n9947), .ZN(n10037) );
  INV_X1 U12768 ( .A(n12503), .ZN(n9956) );
  NOR2_X2 U12769 ( .A1(n10838), .A2(n9956), .ZN(n10843) );
  AND2_X2 U12770 ( .A1(n11248), .A2(n10339), .ZN(n15151) );
  OAI211_X1 U12771 ( .C1(n10788), .C2(n9958), .A(P2_STATE2_REG_0__SCAN_IN), 
        .B(n10787), .ZN(n10790) );
  NAND3_X1 U12772 ( .A1(n10783), .A2(n10782), .A3(n11743), .ZN(n9958) );
  NOR2_X1 U12773 ( .A1(n9944), .A2(n9960), .ZN(n9959) );
  NAND2_X1 U12774 ( .A1(n11033), .A2(n11032), .ZN(n11035) );
  NAND2_X1 U12775 ( .A1(n11034), .A2(n11035), .ZN(n9961) );
  NAND2_X4 U12776 ( .A1(n10723), .A2(n10722), .ZN(n13572) );
  NAND2_X2 U12777 ( .A1(n10710), .A2(n10711), .ZN(n15625) );
  AND2_X2 U12778 ( .A1(n9962), .A2(n10756), .ZN(n11451) );
  NAND2_X1 U12779 ( .A1(n10825), .A2(n9969), .ZN(n10046) );
  INV_X1 U12780 ( .A(n9969), .ZN(n10826) );
  INV_X2 U12781 ( .A(n9968), .ZN(n12485) );
  NAND2_X1 U12782 ( .A1(n10831), .A2(n9969), .ZN(n9968) );
  INV_X1 U12783 ( .A(n9976), .ZN(n17751) );
  INV_X2 U12784 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10497) );
  NAND4_X1 U12785 ( .A1(n11984), .A2(n12256), .A3(n12120), .A4(n11986), .ZN(
        n11992) );
  NAND2_X1 U12786 ( .A1(n11992), .A2(n12250), .ZN(n11997) );
  AND2_X4 U12787 ( .A1(n10241), .A2(n13318), .ZN(n11906) );
  AND2_X2 U12788 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13318) );
  AND2_X2 U12789 ( .A1(n9984), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10241) );
  NAND2_X1 U12790 ( .A1(n15866), .A2(n12374), .ZN(n9985) );
  NAND2_X1 U12791 ( .A1(n9986), .A2(n10079), .ZN(n15866) );
  OAI21_X2 U12792 ( .B1(n13799), .B2(n9993), .A(n9991), .ZN(n15851) );
  INV_X1 U12793 ( .A(n9996), .ZN(n10071) );
  NOR2_X1 U12794 ( .A1(n15196), .A2(n9998), .ZN(n9997) );
  NAND4_X1 U12795 ( .A1(n11132), .A2(n10144), .A3(n10142), .A4(n9889), .ZN(
        n11162) );
  AND2_X2 U12796 ( .A1(n11186), .A2(n9837), .ZN(n11212) );
  INV_X1 U12797 ( .A(n10005), .ZN(n10004) );
  OAI21_X1 U12798 ( .B1(n11252), .B2(n15149), .A(n9884), .ZN(n10005) );
  MUX2_X1 U12799 ( .A(n9848), .B(n11236), .S(n11218), .Z(n10007) );
  NOR2_X1 U12800 ( .A1(n10008), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17799) );
  NOR2_X1 U12801 ( .A1(n17841), .A2(n10008), .ZN(n16770) );
  AOI21_X1 U12802 ( .B1(n17803), .B2(n10008), .A(n17818), .ZN(n17812) );
  INV_X1 U12803 ( .A(n10013), .ZN(n16608) );
  INV_X1 U12804 ( .A(n16286), .ZN(n10647) );
  NAND2_X1 U12805 ( .A1(n10021), .A2(n10016), .ZN(P3_U2640) );
  NOR2_X1 U12806 ( .A1(n16485), .A2(n9890), .ZN(n16473) );
  CLKBUF_X1 U12807 ( .A(n10037), .Z(n10034) );
  INV_X2 U12808 ( .A(n10037), .ZN(n12830) );
  CLKBUF_X1 U12809 ( .A(n12830), .Z(n10035) );
  NOR2_X1 U12810 ( .A1(n10035), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11490) );
  AND2_X1 U12811 ( .A1(n10035), .A2(n19469), .ZN(n11487) );
  AND2_X1 U12812 ( .A1(n11732), .A2(n10037), .ZN(n10325) );
  MUX2_X1 U12813 ( .A(n10037), .B(n19883), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11497) );
  NAND2_X1 U12814 ( .A1(n11438), .A2(n10034), .ZN(n11506) );
  MUX2_X1 U12815 ( .A(n10767), .B(n10037), .S(n11732), .Z(n10770) );
  NAND2_X1 U12816 ( .A1(n11440), .A2(n10034), .ZN(n11442) );
  AOI21_X1 U12817 ( .B1(n10035), .B2(P2_EAX_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10036) );
  NAND2_X1 U12818 ( .A1(n11444), .A2(n10034), .ZN(n11445) );
  NAND2_X1 U12819 ( .A1(n15646), .A2(n10034), .ZN(n19269) );
  INV_X1 U12820 ( .A(n10984), .ZN(n10041) );
  INV_X1 U12821 ( .A(n13618), .ZN(n10044) );
  NAND2_X1 U12822 ( .A1(n10982), .A2(n10983), .ZN(n13593) );
  NAND2_X1 U12823 ( .A1(n10039), .A2(n10984), .ZN(n13594) );
  AND2_X2 U12824 ( .A1(n15204), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10320) );
  XNOR2_X2 U12825 ( .A(n10824), .B(n10066), .ZN(n12503) );
  NAND2_X2 U12826 ( .A1(n10046), .A2(n10803), .ZN(n10066) );
  INV_X1 U12827 ( .A(n10050), .ZN(n17809) );
  AND2_X2 U12828 ( .A1(n10050), .A2(n9873), .ZN(n17802) );
  XNOR2_X1 U12829 ( .A(n10463), .B(n10462), .ZN(n17810) );
  NOR2_X1 U12830 ( .A1(n17823), .A2(n10461), .ZN(n10463) );
  NAND2_X1 U12831 ( .A1(n10467), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10056) );
  XNOR2_X1 U12832 ( .A(n10470), .B(n10096), .ZN(n17767) );
  NAND2_X1 U12833 ( .A1(n17504), .A2(n9839), .ZN(n16264) );
  INV_X1 U12834 ( .A(n10481), .ZN(n10060) );
  NAND2_X1 U12835 ( .A1(n17504), .A2(n10059), .ZN(n17491) );
  AND2_X1 U12836 ( .A1(n17504), .A2(n10481), .ZN(n10482) );
  AND2_X1 U12837 ( .A1(n17753), .A2(n9834), .ZN(n17637) );
  NAND2_X1 U12838 ( .A1(n10062), .A2(n10061), .ZN(n17628) );
  OR2_X2 U12839 ( .A1(n17753), .A2(n17978), .ZN(n10062) );
  NAND2_X1 U12840 ( .A1(n9872), .A2(n10850), .ZN(n10888) );
  NAND4_X1 U12841 ( .A1(n10695), .A2(n10694), .A3(n10692), .A4(n10693), .ZN(
        n10067) );
  NAND4_X1 U12842 ( .A1(n10698), .A2(n10699), .A3(n10696), .A4(n10697), .ZN(
        n10068) );
  NAND3_X1 U12843 ( .A1(n10070), .A2(n10069), .A3(n15170), .ZN(n15157) );
  NAND2_X1 U12844 ( .A1(n10071), .A2(n15479), .ZN(n10069) );
  AOI21_X1 U12845 ( .B1(n13547), .B2(n11539), .A(n10074), .ZN(n11126) );
  XNOR2_X2 U12846 ( .A(n11294), .B(n10075), .ZN(n10838) );
  AND2_X2 U12847 ( .A1(n11820), .A2(n10241), .ZN(n12314) );
  AND2_X2 U12848 ( .A1(n14654), .A2(n10076), .ZN(n14635) );
  NAND2_X1 U12849 ( .A1(n20093), .A2(n10077), .ZN(n10079) );
  NOR2_X1 U12850 ( .A1(n10243), .A2(n10080), .ZN(n10077) );
  XNOR2_X2 U12851 ( .A(n12329), .B(n20109), .ZN(n20093) );
  NAND2_X1 U12852 ( .A1(n20223), .A2(n12242), .ZN(n13725) );
  NAND3_X1 U12853 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10089) );
  NOR2_X2 U12854 ( .A1(n17789), .A2(n17788), .ZN(n17787) );
  AND2_X2 U12855 ( .A1(n10092), .A2(n9885), .ZN(n17789) );
  OR2_X2 U12856 ( .A1(n17802), .A2(n17801), .ZN(n10092) );
  OR2_X2 U12857 ( .A1(n17767), .A2(n18085), .ZN(n10095) );
  NAND2_X1 U12858 ( .A1(n10098), .A2(n10097), .ZN(n10101) );
  NAND2_X1 U12859 ( .A1(n10102), .A2(n10101), .ZN(P3_U2832) );
  INV_X1 U12860 ( .A(n10103), .ZN(n10102) );
  NOR2_X2 U12861 ( .A1(n13267), .A2(n10123), .ZN(n13630) );
  NOR2_X1 U12862 ( .A1(n13266), .A2(n13265), .ZN(n13267) );
  NAND2_X1 U12863 ( .A1(n11245), .A2(n11244), .ZN(n11254) );
  NAND2_X1 U12864 ( .A1(n11172), .A2(n10139), .ZN(n11188) );
  NAND3_X1 U12865 ( .A1(n11132), .A2(n10144), .A3(n10142), .ZN(n11154) );
  NOR2_X2 U12866 ( .A1(n11113), .A2(n10143), .ZN(n10142) );
  NAND2_X1 U12867 ( .A1(n11285), .A2(n10145), .ZN(n11276) );
  NAND2_X1 U12868 ( .A1(n11285), .A2(n9933), .ZN(n11286) );
  NAND2_X1 U12869 ( .A1(n11285), .A2(n11262), .ZN(n11267) );
  INV_X1 U12870 ( .A(n11276), .ZN(n11278) );
  NAND2_X1 U12871 ( .A1(n11209), .A2(n10146), .ZN(n11237) );
  OR2_X2 U12872 ( .A1(n11199), .A2(n11200), .ZN(n11202) );
  AND2_X2 U12873 ( .A1(n15460), .A2(n10151), .ZN(n15393) );
  NAND2_X1 U12874 ( .A1(n15062), .A2(n12953), .ZN(n12952) );
  NAND2_X1 U12875 ( .A1(n15062), .A2(n9932), .ZN(n10158) );
  NOR3_X1 U12876 ( .A1(n14431), .A2(n10180), .A3(n14417), .ZN(n14404) );
  INV_X1 U12877 ( .A(n12118), .ZN(n10177) );
  INV_X1 U12878 ( .A(n14226), .ZN(n10178) );
  NAND2_X1 U12879 ( .A1(n13404), .A2(n13405), .ZN(n13494) );
  NAND3_X1 U12880 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10183) );
  NAND2_X1 U12881 ( .A1(n10182), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12858) );
  AOI21_X1 U12882 ( .B1(n15679), .B2(n9925), .A(n10190), .ZN(n10189) );
  NAND2_X1 U12883 ( .A1(n10187), .A2(n10186), .ZN(n16051) );
  NAND2_X1 U12884 ( .A1(n15679), .A2(n10188), .ZN(n10187) );
  NAND2_X1 U12885 ( .A1(n12870), .A2(n9846), .ZN(n12876) );
  INV_X1 U12886 ( .A(n18890), .ZN(n10199) );
  NAND2_X1 U12887 ( .A1(n10198), .A2(n10200), .ZN(n18868) );
  NAND2_X1 U12888 ( .A1(n10199), .A2(n9925), .ZN(n10198) );
  OR2_X1 U12889 ( .A1(n12959), .A2(n12961), .ZN(n10203) );
  NAND2_X1 U12890 ( .A1(n10205), .A2(n10207), .ZN(n16025) );
  INV_X1 U12891 ( .A(n16052), .ZN(n10206) );
  OR2_X1 U12892 ( .A1(n16052), .A2(n19041), .ZN(n10209) );
  NAND2_X2 U12893 ( .A1(n10275), .A2(n10814), .ZN(n11294) );
  NAND2_X1 U12894 ( .A1(n10217), .A2(n10777), .ZN(n10781) );
  NAND2_X1 U12895 ( .A1(n11728), .A2(n15625), .ZN(n10217) );
  NAND2_X1 U12896 ( .A1(n11448), .A2(n10218), .ZN(n11728) );
  NAND2_X1 U12897 ( .A1(n10775), .A2(n13457), .ZN(n11448) );
  NAND2_X1 U12898 ( .A1(n15002), .A2(n15003), .ZN(n14994) );
  NAND2_X1 U12899 ( .A1(n15002), .A2(n10222), .ZN(n10219) );
  OR2_X1 U12900 ( .A1(n15002), .A2(n10221), .ZN(n10220) );
  AOI21_X1 U12901 ( .B1(n10234), .B2(n10232), .A(n12760), .ZN(n12763) );
  INV_X1 U12902 ( .A(n10754), .ZN(n10767) );
  NAND4_X1 U12903 ( .A1(n10236), .A2(n10238), .A3(n10235), .A4(n10237), .ZN(
        n10774) );
  NAND4_X1 U12904 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(
        n10235) );
  NAND2_X1 U12905 ( .A1(n10678), .A2(n10679), .ZN(n10237) );
  NAND2_X1 U12906 ( .A1(n13610), .A2(n9913), .ZN(n15010) );
  NAND2_X1 U12907 ( .A1(n13285), .A2(n9914), .ZN(n13588) );
  NAND3_X1 U12908 ( .A1(n10240), .A2(n13135), .A3(n9845), .ZN(n13126) );
  NAND3_X1 U12909 ( .A1(n13335), .A2(n12177), .A3(n20824), .ZN(n10242) );
  NAND2_X1 U12910 ( .A1(n10242), .A2(n9909), .ZN(n12189) );
  NAND2_X1 U12911 ( .A1(n14677), .A2(n9811), .ZN(n14623) );
  NAND3_X1 U12912 ( .A1(n14677), .A2(n9811), .A3(n10244), .ZN(n14636) );
  INV_X1 U12913 ( .A(n14636), .ZN(n12421) );
  NAND2_X1 U12914 ( .A1(n13229), .A2(n12382), .ZN(n12254) );
  NAND2_X1 U12915 ( .A1(n13229), .A2(n14926), .ZN(n20390) );
  NAND2_X1 U12916 ( .A1(n13229), .A2(n14927), .ZN(n20666) );
  INV_X1 U12917 ( .A(n13229), .ZN(n14925) );
  INV_X1 U12918 ( .A(n20146), .ZN(n10246) );
  OR2_X2 U12919 ( .A1(n15851), .A2(n10249), .ZN(n10247) );
  AND2_X1 U12920 ( .A1(n12411), .A2(n15852), .ZN(n10249) );
  NAND2_X2 U12921 ( .A1(n10253), .A2(n10252), .ZN(n12394) );
  INV_X1 U12922 ( .A(n12367), .ZN(n10253) );
  INV_X1 U12923 ( .A(n12353), .ZN(n10254) );
  INV_X1 U12924 ( .A(n10261), .ZN(n14509) );
  NOR2_X1 U12925 ( .A1(n14406), .A2(n14407), .ZN(n14218) );
  NOR2_X1 U12926 ( .A1(n14406), .A2(n10268), .ZN(n14395) );
  NOR2_X1 U12927 ( .A1(n12948), .A2(n12949), .ZN(n10278) );
  INV_X1 U12928 ( .A(n12834), .ZN(n10280) );
  NAND2_X1 U12929 ( .A1(n11321), .A2(n9838), .ZN(n13413) );
  OAI21_X1 U12930 ( .B1(n13547), .B2(n10074), .A(n10301), .ZN(n13543) );
  INV_X1 U12931 ( .A(n15138), .ZN(n10304) );
  NOR2_X1 U12932 ( .A1(n15138), .A2(n9888), .ZN(n10302) );
  NAND2_X1 U12933 ( .A1(n11159), .A2(n11158), .ZN(n15270) );
  NOR2_X4 U12934 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13531) );
  NAND2_X1 U12935 ( .A1(n10310), .A2(n10765), .ZN(n11092) );
  AND4_X2 U12936 ( .A1(n10325), .A2(n10769), .A3(n11731), .A4(n10311), .ZN(
        n15559) );
  AND2_X2 U12937 ( .A1(n10843), .A2(n10839), .ZN(n10990) );
  NAND2_X1 U12938 ( .A1(n10952), .A2(n10951), .ZN(n10962) );
  NAND2_X1 U12939 ( .A1(n13147), .A2(n20824), .ZN(n12216) );
  INV_X1 U12940 ( .A(n11982), .ZN(n11984) );
  NAND2_X1 U12941 ( .A1(n12216), .A2(n12215), .ZN(n12263) );
  INV_X1 U12942 ( .A(n13285), .ZN(n13202) );
  XNOR2_X1 U12943 ( .A(n12510), .B(n12511), .ZN(n13071) );
  NAND2_X1 U12944 ( .A1(n12510), .A2(n12512), .ZN(n13137) );
  NAND2_X1 U12945 ( .A1(n12485), .A2(n12505), .ZN(n12488) );
  OAI211_X1 U12946 ( .C1(n13654), .C2(n13658), .A(n13653), .B(n13652), .ZN(
        n13655) );
  CLKBUF_X1 U12947 ( .A(n15010), .Z(n15018) );
  NAND2_X1 U12948 ( .A1(n13649), .A2(n13951), .ZN(n13653) );
  INV_X1 U12949 ( .A(n13207), .ZN(n13210) );
  NOR2_X1 U12950 ( .A1(n14304), .A2(n14303), .ZN(n14322) );
  AOI21_X1 U12951 ( .B1(n14367), .B2(n20096), .A(n14301), .ZN(n14302) );
  NAND2_X1 U12952 ( .A1(n11397), .A2(n11734), .ZN(n10785) );
  NAND2_X1 U12953 ( .A1(n10781), .A2(n10780), .ZN(n10782) );
  NAND2_X1 U12954 ( .A1(n10704), .A2(n10676), .ZN(n10711) );
  NAND2_X1 U12955 ( .A1(n10709), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10710) );
  NAND2_X1 U12956 ( .A1(n10716), .A2(n10676), .ZN(n10723) );
  INV_X1 U12957 ( .A(n10983), .ZN(n10984) );
  AND4_X1 U12958 ( .A1(n11729), .A2(n11448), .A3(n11447), .A4(n11446), .ZN(
        n11449) );
  AND3_X1 U12959 ( .A1(n10677), .A2(n10676), .A3(n10675), .ZN(n10678) );
  AOI22_X1 U12960 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U12961 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U12962 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12632), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10708) );
  AND2_X2 U12963 ( .A1(n20058), .A2(n20046), .ZN(n20056) );
  OR2_X1 U12964 ( .A1(n13348), .A2(n12026), .ZN(n13385) );
  INV_X1 U12965 ( .A(n10865), .ZN(n12635) );
  INV_X1 U12966 ( .A(n10857), .ZN(n10968) );
  INV_X1 U12967 ( .A(n10944), .ZN(n11015) );
  AND2_X1 U12968 ( .A1(n17248), .A2(n9826), .ZN(n17193) );
  AND4_X1 U12969 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10326) );
  INV_X1 U12970 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19942) );
  INV_X1 U12971 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19864) );
  AND2_X1 U12972 ( .A1(n13572), .A2(n10766), .ZN(n10327) );
  AND4_X1 U12973 ( .A1(n10453), .A2(n10452), .A3(n10451), .A4(n10450), .ZN(
        n10329) );
  AND2_X1 U12974 ( .A1(n10407), .A2(n10406), .ZN(n10330) );
  NOR4_X1 U12975 ( .A1(n20666), .A2(n20622), .A3(n9821), .A4(n20669), .ZN(
        n10331) );
  NAND2_X1 U12976 ( .A1(n10737), .A2(n11443), .ZN(n11437) );
  AND2_X4 U12977 ( .A1(n12394), .A2(n12393), .ZN(n10332) );
  XOR2_X1 U12978 ( .A(n12675), .B(n12693), .Z(n10333) );
  AND4_X1 U12979 ( .A1(n10457), .A2(n10456), .A3(n10455), .A4(n10454), .ZN(
        n10334) );
  AND4_X1 U12980 ( .A1(n10948), .A2(n10947), .A3(n10946), .A4(n10945), .ZN(
        n10335) );
  AND2_X1 U12981 ( .A1(n10660), .A2(n10659), .ZN(n10336) );
  AND2_X1 U12982 ( .A1(n12244), .A2(n12255), .ZN(n10337) );
  OR2_X1 U12983 ( .A1(n11539), .A2(n11681), .ZN(n10338) );
  OR3_X1 U12984 ( .A1(n12934), .A2(n11539), .A3(n15359), .ZN(n10339) );
  NAND2_X1 U12985 ( .A1(n11271), .A2(n15297), .ZN(n10340) );
  AND2_X1 U12986 ( .A1(n9908), .A2(n11772), .ZN(n10341) );
  OR2_X1 U12987 ( .A1(n19071), .A2(n13015), .ZN(n10342) );
  AND4_X1 U12988 ( .A1(n15185), .A2(n15197), .A3(n15240), .A4(n11217), .ZN(
        n10344) );
  INV_X1 U12989 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10446) );
  INV_X1 U12990 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10459) );
  OR2_X1 U12991 ( .A1(n18947), .A2(n11539), .ZN(n11190) );
  AND2_X1 U12992 ( .A1(n11292), .A2(n15614), .ZN(n19242) );
  NOR2_X1 U12993 ( .A1(n15968), .A2(n15967), .ZN(n10345) );
  INV_X1 U12994 ( .A(n17682), .ZN(n17664) );
  INV_X1 U12995 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12416) );
  INV_X1 U12996 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17663) );
  NOR2_X1 U12997 ( .A1(n20545), .A2(n20511), .ZN(n10346) );
  AND4_X1 U12998 ( .A1(n11554), .A2(n11553), .A3(n11552), .A4(n11551), .ZN(
        n10347) );
  INV_X1 U12999 ( .A(n17574), .ZN(n16448) );
  INV_X1 U13000 ( .A(n11487), .ZN(n11701) );
  AND2_X1 U13001 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10349) );
  INV_X1 U13002 ( .A(n13960), .ZN(n14596) );
  AND2_X1 U13003 ( .A1(n14974), .A2(n12698), .ZN(n10350) );
  NAND2_X1 U13004 ( .A1(n11771), .A2(n12842), .ZN(n10351) );
  BUF_X1 U13005 ( .A(n14149), .Z(n14015) );
  OR2_X1 U13006 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n10352) );
  AND3_X1 U13007 ( .A1(n11556), .A2(n11555), .A3(n10347), .ZN(n13284) );
  INV_X1 U13008 ( .A(n13284), .ZN(n12516) );
  NAND2_X1 U13009 ( .A1(n14983), .A2(n14982), .ZN(n14981) );
  NAND2_X1 U13010 ( .A1(n15393), .A2(n15392), .ZN(n12924) );
  OR2_X1 U13011 ( .A1(n11783), .A2(n16130), .ZN(n10353) );
  AND2_X1 U13012 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10354) );
  OAI21_X1 U13013 ( .B1(n13592), .B2(n13591), .A(n11131), .ZN(n13615) );
  AND4_X1 U13014 ( .A1(n11846), .A2(n11845), .A3(n11844), .A4(n11843), .ZN(
        n10355) );
  AND2_X1 U13015 ( .A1(n11905), .A2(n11904), .ZN(n10356) );
  AND4_X1 U13016 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n10357) );
  NAND2_X1 U13017 ( .A1(n13669), .A2(n12026), .ZN(n12028) );
  OR2_X1 U13018 ( .A1(n11946), .A2(n11945), .ZN(n11951) );
  INV_X1 U13019 ( .A(n12377), .ZN(n11956) );
  OR2_X1 U13020 ( .A1(n12342), .A2(n12341), .ZN(n12368) );
  AND3_X1 U13021 ( .A1(n12238), .A2(n12237), .A3(n12236), .ZN(n12245) );
  NAND2_X1 U13022 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10662) );
  NOR2_X1 U13023 ( .A1(n19894), .A2(n10354), .ZN(n10761) );
  NAND2_X1 U13024 ( .A1(n11079), .A2(n11078), .ZN(n11082) );
  AOI22_X1 U13025 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10739) );
  AND2_X1 U13026 ( .A1(n19894), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10798) );
  OAI21_X1 U13027 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n10497), .A(
        n10498), .ZN(n10499) );
  INV_X1 U13028 ( .A(n11941), .ZN(n11809) );
  INV_X1 U13029 ( .A(n14138), .ZN(n13676) );
  NAND2_X1 U13030 ( .A1(n12332), .A2(n12331), .ZN(n12353) );
  NAND2_X1 U13031 ( .A1(n12019), .A2(n14933), .ZN(n12166) );
  INV_X1 U13032 ( .A(n10773), .ZN(n10756) );
  OR2_X1 U13033 ( .A1(n11792), .A2(n11770), .ZN(n11771) );
  INV_X1 U13034 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11191) );
  AND4_X1 U13035 ( .A1(n11051), .A2(n11050), .A3(n11049), .A4(n11048), .ZN(
        n11061) );
  INV_X1 U13036 ( .A(n13785), .ZN(n12065) );
  NOR2_X1 U13037 ( .A1(n14214), .A2(n14629), .ZN(n14242) );
  NAND2_X1 U13038 ( .A1(n13676), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14142) );
  INV_X1 U13039 ( .A(n14597), .ZN(n13959) );
  INV_X1 U13040 ( .A(n13750), .ZN(n13751) );
  OR2_X1 U13041 ( .A1(n13180), .A2(n12269), .ZN(n12270) );
  INV_X1 U13042 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12415) );
  AND2_X1 U13043 ( .A1(n12064), .A2(n12063), .ZN(n13785) );
  AND2_X1 U13044 ( .A1(n11450), .A2(n11449), .ZN(n11727) );
  INV_X1 U13045 ( .A(n15020), .ZN(n12568) );
  NAND2_X1 U13046 ( .A1(n11190), .A2(n11191), .ZN(n11192) );
  OAI21_X1 U13047 ( .B1(n11156), .B2(n11289), .A(n19009), .ZN(n11157) );
  NAND2_X1 U13048 ( .A1(n11496), .A2(n11495), .ZN(n11499) );
  INV_X1 U13049 ( .A(n16569), .ZN(n16449) );
  INV_X1 U13050 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n21164) );
  AND2_X1 U13051 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n10632), .ZN(
        n10633) );
  NAND2_X1 U13052 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10450) );
  NOR2_X1 U13053 ( .A1(n12380), .A2(n12391), .ZN(n11966) );
  AND2_X1 U13054 ( .A1(n11806), .A2(n11807), .ZN(n11939) );
  AND2_X1 U13055 ( .A1(n14386), .A2(n14282), .ZN(n14283) );
  NOR2_X1 U13056 ( .A1(n13998), .A2(n15784), .ZN(n14030) );
  AND2_X1 U13057 ( .A1(n13869), .A2(n13914), .ZN(n13868) );
  INV_X1 U13058 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13674) );
  AOI21_X1 U13059 ( .B1(n13642), .B2(n13951), .A(n13641), .ZN(n13643) );
  NAND2_X1 U13060 ( .A1(n12416), .A2(n12415), .ZN(n12417) );
  NAND2_X1 U13061 ( .A1(n20421), .A2(n20824), .ZN(n12296) );
  INV_X1 U13062 ( .A(n13175), .ZN(n20147) );
  NAND2_X1 U13063 ( .A1(n11090), .A2(n11089), .ZN(n11409) );
  INV_X1 U13064 ( .A(n13587), .ZN(n12518) );
  INV_X1 U13065 ( .A(n15028), .ZN(n12535) );
  INV_X1 U13066 ( .A(n15495), .ZN(n15440) );
  OR2_X1 U13067 ( .A1(n11779), .A2(n13530), .ZN(n15437) );
  NAND2_X1 U13068 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10419) );
  INV_X1 U13069 ( .A(n17640), .ZN(n10646) );
  NOR2_X1 U13070 ( .A1(n16316), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10483) );
  OAI21_X1 U13071 ( .B1(n10480), .B2(n17860), .A(n17754), .ZN(n10481) );
  OAI21_X1 U13072 ( .B1(n10478), .B2(n17523), .A(n10477), .ZN(n10479) );
  NAND2_X1 U13073 ( .A1(n10468), .A2(n10612), .ZN(n16318) );
  NOR2_X1 U13074 ( .A1(n17825), .A2(n17824), .ZN(n17823) );
  OR2_X1 U13075 ( .A1(n14451), .A2(n14231), .ZN(n14409) );
  AND2_X1 U13076 ( .A1(n14050), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14068) );
  NAND2_X1 U13077 ( .A1(n12280), .A2(n12279), .ZN(n20309) );
  NAND2_X1 U13078 ( .A1(n20826), .A2(n13667), .ZN(n19940) );
  OR2_X1 U13079 ( .A1(n15762), .A2(n10352), .ZN(n14072) );
  INV_X1 U13080 ( .A(n14143), .ZN(n14176) );
  AND2_X1 U13081 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n14030), .ZN(
        n14050) );
  NOR2_X1 U13082 ( .A1(n13942), .A2(n15803), .ZN(n13924) );
  NOR2_X1 U13083 ( .A1(n13835), .A2(n13836), .ZN(n13851) );
  NOR2_X1 U13084 ( .A1(n13733), .A2(n19942), .ZN(n13776) );
  INV_X1 U13085 ( .A(n13706), .ZN(n13749) );
  INV_X1 U13086 ( .A(n13238), .ZN(n13239) );
  INV_X1 U13087 ( .A(n14635), .ZN(n14637) );
  AND2_X1 U13088 ( .A1(n14825), .A2(n12135), .ZN(n14809) );
  AND2_X1 U13089 ( .A1(n12076), .A2(n12075), .ZN(n13897) );
  INV_X1 U13090 ( .A(n13784), .ZN(n15945) );
  XNOR2_X1 U13091 ( .A(n12263), .B(n12262), .ZN(n13175) );
  OR2_X1 U13092 ( .A1(n9821), .A2(n13175), .ZN(n20586) );
  INV_X1 U13093 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20660) );
  AND2_X1 U13094 ( .A1(n16226), .A2(n13032), .ZN(n12970) );
  AND3_X1 U13095 ( .A1(n11531), .A2(n11530), .A3(n11529), .ZN(n13559) );
  OR2_X1 U13096 ( .A1(n15596), .A2(n19902), .ZN(n19865) );
  NOR2_X1 U13097 ( .A1(n12946), .A2(n11539), .ZN(n12438) );
  AND2_X1 U13098 ( .A1(n16189), .A2(n11754), .ZN(n15513) );
  AND2_X1 U13099 ( .A1(n15607), .A2(n15606), .ZN(n15648) );
  AND2_X1 U13100 ( .A1(n19464), .A2(n19651), .ZN(n19467) );
  NAND2_X1 U13101 ( .A1(n19860), .A2(n19342), .ZN(n19847) );
  NAND2_X1 U13102 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19707), .ZN(n15608) );
  NAND2_X2 U13103 ( .A1(n19101), .A2(n9787), .ZN(n15651) );
  NOR2_X1 U13104 ( .A1(n17488), .A2(n16507), .ZN(n16506) );
  NOR2_X1 U13105 ( .A1(n16558), .A2(n16557), .ZN(n16556) );
  NOR2_X1 U13106 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16685), .ZN(n16671) );
  NOR2_X1 U13107 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16730), .ZN(n16717) );
  OR2_X1 U13108 ( .A1(n18826), .A2(n18172), .ZN(n16459) );
  INV_X1 U13109 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17775) );
  NAND2_X1 U13110 ( .A1(n17675), .A2(n17845), .ZN(n17564) );
  OR2_X1 U13111 ( .A1(n15675), .A2(n12479), .ZN(n12481) );
  INV_X1 U13112 ( .A(n17754), .ZN(n17685) );
  INV_X1 U13113 ( .A(n17628), .ZN(n17629) );
  NOR2_X2 U13114 ( .A1(n18623), .A2(n18635), .ZN(n18052) );
  INV_X1 U13115 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18617) );
  NAND2_X1 U13116 ( .A1(n11978), .A2(n11977), .ZN(n13293) );
  NAND2_X1 U13117 ( .A1(n14068), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14089) );
  INV_X1 U13118 ( .A(n19986), .ZN(n19998) );
  AND2_X1 U13119 ( .A1(n14300), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13679) );
  AND2_X1 U13120 ( .A1(n20826), .A2(n13672), .ZN(n19988) );
  INV_X1 U13121 ( .A(n14591), .ZN(n14557) );
  NAND2_X1 U13122 ( .A1(n13807), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13835) );
  NAND2_X1 U13123 ( .A1(n13484), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13511) );
  AND3_X1 U13124 ( .A1(n15707), .A2(n13294), .A3(n13293), .ZN(n20097) );
  INV_X1 U13125 ( .A(n14796), .ZN(n14829) );
  NOR2_X1 U13126 ( .A1(n15890), .A2(n15828), .ZN(n15881) );
  OR2_X1 U13127 ( .A1(n20120), .A2(n14866), .ZN(n15953) );
  OR2_X1 U13128 ( .A1(n12123), .A2(n14910), .ZN(n20120) );
  AND2_X1 U13129 ( .A1(n12425), .A2(n12121), .ZN(n20126) );
  INV_X1 U13130 ( .A(n20288), .ZN(n20276) );
  NOR2_X2 U13131 ( .A1(n20288), .A2(n20586), .ZN(n20271) );
  NOR2_X2 U13132 ( .A1(n20288), .A2(n20509), .ZN(n20332) );
  OAI21_X1 U13133 ( .B1(n9934), .B2(n20316), .A(n20628), .ZN(n20333) );
  INV_X1 U13134 ( .A(n20426), .ZN(n20446) );
  INV_X1 U13135 ( .A(n20539), .ZN(n20419) );
  AND2_X1 U13136 ( .A1(n20515), .A2(n20456), .ZN(n20504) );
  AND2_X1 U13137 ( .A1(n14925), .A2(n20146), .ZN(n20515) );
  INV_X1 U13138 ( .A(n20552), .ZN(n20575) );
  INV_X1 U13139 ( .A(n20623), .ZN(n20652) );
  INV_X1 U13140 ( .A(n20558), .ZN(n20676) );
  INV_X1 U13141 ( .A(n20723), .ZN(n20697) );
  INV_X1 U13142 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n15722) );
  INV_X1 U13143 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20735) );
  AND2_X1 U13144 ( .A1(n16224), .A2(n16226), .ZN(n13025) );
  INV_X1 U13145 ( .A(n19069), .ZN(n19049) );
  AND2_X1 U13146 ( .A1(n19231), .A2(n16249), .ZN(n19064) );
  INV_X1 U13147 ( .A(n19121), .ZN(n19125) );
  NAND2_X1 U13148 ( .A1(n15125), .A2(n15124), .ZN(n15126) );
  INV_X1 U13149 ( .A(n16150), .ZN(n19237) );
  XNOR2_X1 U13150 ( .A(n11247), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15158) );
  NOR2_X1 U13151 ( .A1(n15519), .A2(n16203), .ZN(n16153) );
  INV_X1 U13152 ( .A(n19275), .ZN(n19265) );
  NAND2_X1 U13153 ( .A1(n19846), .A2(n19878), .ZN(n19401) );
  NOR2_X1 U13154 ( .A1(n19705), .A2(n19401), .ZN(n19404) );
  INV_X1 U13155 ( .A(n19463), .ZN(n19489) );
  INV_X1 U13156 ( .A(n19528), .ZN(n19519) );
  OR2_X1 U13157 ( .A1(n19860), .A2(n19342), .ZN(n19619) );
  INV_X1 U13158 ( .A(n19536), .ZN(n19707) );
  INV_X1 U13159 ( .A(n19673), .ZN(n19721) );
  NOR2_X1 U13160 ( .A1(n19620), .A2(n19705), .ZN(n19698) );
  NOR2_X1 U13161 ( .A1(n16575), .A2(n16468), .ZN(n16543) );
  NOR2_X1 U13162 ( .A1(n16607), .A2(n16461), .ZN(n16582) );
  NOR2_X1 U13163 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16616), .ZN(n16602) );
  NOR2_X1 U13164 ( .A1(n16664), .A2(n16460), .ZN(n16639) );
  NOR2_X1 U13165 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16704), .ZN(n16691) );
  NOR2_X1 U13166 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16751), .ZN(n16733) );
  INV_X1 U13167 ( .A(n16800), .ZN(n16812) );
  NAND2_X1 U13168 ( .A1(n17416), .A2(n18606), .ZN(n18826) );
  NOR2_X1 U13169 ( .A1(n17433), .A2(n17223), .ZN(n17218) );
  INV_X1 U13170 ( .A(n17238), .ZN(n17234) );
  NAND2_X1 U13171 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17285), .ZN(n17281) );
  NOR2_X1 U13172 ( .A1(n17349), .A2(n17290), .ZN(n17320) );
  INV_X1 U13173 ( .A(n17345), .ZN(n17353) );
  OR2_X1 U13174 ( .A1(n17481), .A2(n17480), .ZN(n17482) );
  INV_X1 U13175 ( .A(n17696), .ZN(n17604) );
  NOR2_X1 U13176 ( .A1(n17999), .A2(n18036), .ZN(n18016) );
  NAND2_X1 U13177 ( .A1(n12481), .A2(n12480), .ZN(n12482) );
  INV_X1 U13178 ( .A(n17504), .ZN(n17505) );
  INV_X1 U13179 ( .A(n18639), .ZN(n18623) );
  NOR2_X1 U13180 ( .A1(n9790), .A2(n18150), .ZN(n18144) );
  INV_X1 U13181 ( .A(n18669), .ZN(n18663) );
  INV_X1 U13182 ( .A(n18501), .ZN(n18505) );
  OAI22_X1 U13183 ( .A1(n18608), .A2(n12467), .B1(n13975), .B2(n18611), .ZN(
        n18660) );
  INV_X1 U13184 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n16410) );
  NAND3_X1 U13185 ( .A1(n12141), .A2(n13294), .A3(n13293), .ZN(n13348) );
  NAND2_X1 U13186 ( .A1(n19951), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19986) );
  NAND2_X1 U13187 ( .A1(n19951), .A2(n13683), .ZN(n19947) );
  INV_X1 U13188 ( .A(n19982), .ZN(n20004) );
  OR2_X1 U13189 ( .A1(n20058), .A2(n20152), .ZN(n20030) );
  INV_X1 U13190 ( .A(n20056), .ZN(n20045) );
  NAND2_X1 U13191 ( .A1(n13296), .A2(n15718), .ZN(n20058) );
  INV_X1 U13192 ( .A(n20086), .ZN(n13381) );
  INV_X1 U13193 ( .A(n15847), .ZN(n20101) );
  NOR4_X1 U13194 ( .A1(n14767), .A2(n14766), .A3(n14765), .A4(n14764), .ZN(
        n14768) );
  INV_X1 U13195 ( .A(n20126), .ZN(n15936) );
  OR2_X1 U13196 ( .A1(n12432), .A2(n12431), .ZN(n15935) );
  INV_X1 U13197 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20143) );
  INV_X1 U13198 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15995) );
  NAND2_X1 U13199 ( .A1(n20276), .A2(n20419), .ZN(n20248) );
  AOI22_X1 U13200 ( .A1(n20254), .A2(n20251), .B1(n20481), .B2(n20362), .ZN(
        n20275) );
  OR2_X1 U13201 ( .A1(n20390), .A2(n20539), .ZN(n20359) );
  AOI22_X1 U13202 ( .A1(n20367), .A2(n20364), .B1(n20362), .B2(n20544), .ZN(
        n20389) );
  OR2_X1 U13203 ( .A1(n20390), .A2(n20509), .ZN(n20426) );
  NAND2_X1 U13204 ( .A1(n20515), .A2(n20419), .ZN(n20476) );
  AOI22_X1 U13205 ( .A1(n20486), .A2(n20483), .B1(n20481), .B2(n20480), .ZN(
        n20508) );
  NAND2_X1 U13206 ( .A1(n20515), .A2(n20510), .ZN(n20552) );
  OR2_X1 U13207 ( .A1(n20666), .A2(n20539), .ZN(n20615) );
  OR2_X1 U13208 ( .A1(n20666), .A2(n20617), .ZN(n20700) );
  INV_X1 U13209 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20824) );
  INV_X1 U13210 ( .A(n20803), .ZN(n20727) );
  AND2_X1 U13211 ( .A1(n13025), .A2(n13032), .ZN(n19895) );
  AOI21_X1 U13212 ( .B1(n12900), .B2(n19064), .A(n12899), .ZN(n12901) );
  INV_X1 U13213 ( .A(n19064), .ZN(n19053) );
  AND2_X1 U13214 ( .A1(n12829), .A2(n13032), .ZN(n15036) );
  OR2_X1 U13215 ( .A1(n14984), .A2(n12830), .ZN(n15038) );
  NAND2_X1 U13216 ( .A1(n12803), .A2(n12802), .ZN(n19121) );
  NOR2_X1 U13217 ( .A1(n19127), .A2(n19099), .ZN(n19133) );
  INV_X1 U13218 ( .A(n19123), .ZN(n19120) );
  OR2_X1 U13219 ( .A1(n19203), .A2(n19142), .ZN(n19168) );
  NAND2_X1 U13220 ( .A1(n19139), .A2(n19906), .ZN(n19203) );
  INV_X1 U13221 ( .A(n19231), .ZN(n19136) );
  NAND2_X1 U13222 ( .A1(n12845), .A2(n19242), .ZN(n12846) );
  INV_X1 U13223 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19019) );
  INV_X1 U13224 ( .A(n16143), .ZN(n19247) );
  NAND2_X1 U13225 ( .A1(n12845), .A2(n16196), .ZN(n11780) );
  BUF_X1 U13226 ( .A(n12503), .Z(n14359) );
  INV_X1 U13227 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16246) );
  INV_X1 U13228 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16240) );
  AOI21_X1 U13229 ( .B1(n15602), .B2(n15647), .A(n19536), .ZN(n15655) );
  OR2_X1 U13230 ( .A1(n19401), .A2(n19502), .ZN(n19275) );
  AOI211_X2 U13231 ( .C1(n19280), .C2(n19648), .A(n19536), .B(n19279), .ZN(
        n19309) );
  AOI21_X1 U13232 ( .B1(n19315), .B2(n19320), .A(n19314), .ZN(n19341) );
  OR2_X1 U13233 ( .A1(n19401), .A2(n19619), .ZN(n19371) );
  AOI21_X1 U13234 ( .B1(n19376), .B2(n19379), .A(n19375), .ZN(n19400) );
  INV_X1 U13235 ( .A(n19404), .ZN(n19461) );
  OAI22_X1 U13236 ( .A1(n19468), .A2(n19488), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19472), .ZN(n19493) );
  NAND2_X1 U13237 ( .A1(n19462), .A2(n19494), .ZN(n19528) );
  NOR2_X1 U13238 ( .A1(n19537), .A2(n19536), .ZN(n19561) );
  INV_X1 U13239 ( .A(n19578), .ZN(n19572) );
  OR2_X1 U13240 ( .A1(n19650), .A2(n19619), .ZN(n19646) );
  AOI21_X1 U13241 ( .B1(n19656), .B2(n19660), .A(n19655), .ZN(n19697) );
  INV_X1 U13242 ( .A(n19678), .ZN(n19737) );
  INV_X1 U13243 ( .A(n19698), .ZN(n19759) );
  INV_X1 U13244 ( .A(n19845), .ZN(n19768) );
  INV_X1 U13245 ( .A(n19913), .ZN(n19840) );
  NAND2_X1 U13246 ( .A1(n18663), .A2(n18660), .ZN(n16418) );
  NAND2_X1 U13247 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16582), .ZN(n16575) );
  INV_X1 U13248 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n21007) );
  INV_X1 U13249 ( .A(n16796), .ZN(n16798) );
  INV_X1 U13250 ( .A(n16767), .ZN(n16810) );
  INV_X1 U13251 ( .A(n16317), .ZN(n17327) );
  NOR2_X1 U13252 ( .A1(n10393), .A2(n10392), .ZN(n17341) );
  INV_X1 U13253 ( .A(n17383), .ZN(n17382) );
  NAND2_X1 U13254 ( .A1(n17416), .A2(n17358), .ZN(n17414) );
  INV_X1 U13255 ( .A(n17464), .ZN(n17452) );
  INV_X1 U13256 ( .A(n17450), .ZN(n17462) );
  INV_X1 U13257 ( .A(n17755), .ZN(n17733) );
  INV_X1 U13258 ( .A(n10649), .ZN(n18464) );
  INV_X1 U13259 ( .A(n18144), .ZN(n18109) );
  INV_X1 U13260 ( .A(n18134), .ZN(n18142) );
  INV_X1 U13261 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18650) );
  INV_X1 U13262 ( .A(n18754), .ZN(n18822) );
  INV_X1 U13263 ( .A(n16367), .ZN(n16372) );
  NAND2_X1 U13264 ( .A1(n9866), .A2(n12838), .ZN(P2_U2858) );
  NAND2_X1 U13265 ( .A1(n9871), .A2(n12825), .ZN(P2_U2890) );
  OAI211_X1 U13266 ( .C1(n15307), .C2(n12452), .A(n12451), .B(n9867), .ZN(
        P2_U2986) );
  INV_X2 U13267 ( .A(n18619), .ZN(n13971) );
  AOI22_X1 U13268 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16916), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10372) );
  INV_X2 U13269 ( .A(n10511), .ZN(n17156) );
  NOR2_X2 U13270 ( .A1(n18633), .A2(n10362), .ZN(n10416) );
  AOI22_X1 U13271 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10371) );
  NOR2_X2 U13272 ( .A1(n10361), .A2(n10363), .ZN(n10387) );
  NOR2_X2 U13273 ( .A1(n10359), .A2(n13971), .ZN(n10396) );
  AOI22_X1 U13274 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10358) );
  OAI21_X1 U13275 ( .B1(n10516), .B2(n16870), .A(n10358), .ZN(n10369) );
  NOR2_X2 U13276 ( .A1(n10360), .A2(n13971), .ZN(n17164) );
  AOI22_X1 U13277 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U13278 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13279 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16882), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10365) );
  NAND3_X1 U13280 ( .A1(n18796), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n18619), .ZN(n17160) );
  AOI22_X1 U13281 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10364) );
  NAND4_X1 U13282 ( .A1(n10367), .A2(n10366), .A3(n10365), .A4(n10364), .ZN(
        n10368) );
  AOI211_X1 U13283 ( .C1(n9797), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n10369), .B(n10368), .ZN(n10370) );
  NAND3_X1 U13284 ( .A1(n10372), .A2(n10371), .A3(n10370), .ZN(n16317) );
  AOI22_X1 U13285 ( .A1(n10396), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10416), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13286 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10375) );
  AOI22_X1 U13287 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U13288 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10373) );
  NAND4_X1 U13289 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n10382) );
  AOI22_X1 U13290 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13291 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U13292 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16882), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13293 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10377) );
  NAND4_X1 U13294 ( .A1(n10380), .A2(n10379), .A3(n10378), .A4(n10377), .ZN(
        n10381) );
  AOI22_X1 U13295 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13296 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U13297 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16882), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10384) );
  INV_X2 U13298 ( .A(n10516), .ZN(n17162) );
  AOI22_X1 U13299 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10383) );
  NAND4_X1 U13300 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n10393) );
  AOI22_X1 U13301 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10397), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13302 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13303 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13304 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10388) );
  NAND4_X1 U13305 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .ZN(
        n10392) );
  INV_X1 U13306 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10404) );
  INV_X1 U13307 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n21128) );
  AOI22_X1 U13308 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10394) );
  OAI21_X1 U13309 ( .B1(n16982), .B2(n21128), .A(n10394), .ZN(n10395) );
  INV_X1 U13310 ( .A(n10395), .ZN(n10403) );
  AOI22_X1 U13311 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10408), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U13312 ( .A1(n10387), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9792), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10401) );
  AOI22_X1 U13313 ( .A1(n10414), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__2__SCAN_IN), .B2(n10396), .ZN(n10400) );
  AOI22_X1 U13314 ( .A1(n10398), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10397), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U13315 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16882), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U13316 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16885), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U13317 ( .A1(n10408), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n16882), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13318 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10396), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17163), .ZN(n10412) );
  AOI22_X1 U13319 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n9795), .ZN(n10411) );
  AOI22_X1 U13320 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10409), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10410) );
  NAND4_X1 U13321 ( .A1(n10413), .A2(n10412), .A3(n10411), .A4(n10410), .ZN(
        n10424) );
  INV_X1 U13322 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U13323 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10414), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17057), .ZN(n10415) );
  OAI21_X1 U13324 ( .B1(n17200), .B2(n10435), .A(n10415), .ZN(n10423) );
  AOI22_X1 U13325 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17138), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10421) );
  AOI22_X1 U13326 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10418), .B1(
        n9792), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10420) );
  NAND3_X1 U13327 ( .A1(n10421), .A2(n10420), .A3(n10419), .ZN(n10422) );
  AOI22_X1 U13328 ( .A1(n10387), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U13329 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10433) );
  INV_X1 U13330 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n20970) );
  AOI22_X1 U13331 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16916), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10425) );
  OAI21_X1 U13332 ( .B1(n10516), .B2(n20970), .A(n10425), .ZN(n10431) );
  AOI22_X1 U13333 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13334 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16882), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13335 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13336 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10426) );
  NAND4_X1 U13337 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10430) );
  AOI211_X1 U13338 ( .C1(n16885), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n10431), .B(n10430), .ZN(n10432) );
  AOI22_X1 U13339 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13340 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10444) );
  INV_X1 U13341 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n21159) );
  AOI22_X1 U13342 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10436) );
  OAI21_X1 U13343 ( .B1(n10544), .B2(n21159), .A(n10436), .ZN(n10442) );
  AOI22_X1 U13344 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16882), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13345 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9795), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13346 ( .A1(n10396), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U13347 ( .A1(n10387), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10437) );
  NAND4_X1 U13348 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10441) );
  AOI211_X1 U13349 ( .C1(n10397), .C2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n10442), .B(n10441), .ZN(n10443) );
  NAND3_X1 U13350 ( .A1(n10445), .A2(n10444), .A3(n10443), .ZN(n10612) );
  INV_X1 U13351 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17871) );
  INV_X1 U13352 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17978) );
  INV_X1 U13353 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17811) );
  XNOR2_X1 U13354 ( .A(n17352), .B(n10446), .ZN(n17836) );
  INV_X1 U13355 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17207) );
  AOI22_X1 U13356 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10447), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10448) );
  OAI21_X1 U13357 ( .B1(n10435), .B2(n17207), .A(n10448), .ZN(n10449) );
  INV_X1 U13358 ( .A(n10449), .ZN(n10453) );
  AOI22_X1 U13359 ( .A1(n10396), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13360 ( .A1(n10408), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13361 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13362 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13363 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16882), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10455) );
  AOI22_X1 U13364 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10454) );
  NAND2_X1 U13365 ( .A1(n17844), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17843) );
  NOR2_X1 U13366 ( .A1(n17836), .A2(n17843), .ZN(n17835) );
  NOR2_X1 U13367 ( .A1(n17352), .A2(n10446), .ZN(n10458) );
  NOR2_X1 U13368 ( .A1(n17835), .A2(n10458), .ZN(n17825) );
  NOR2_X1 U13369 ( .A1(n10459), .A2(n10460), .ZN(n10461) );
  XOR2_X1 U13370 ( .A(n17341), .B(n10618), .Z(n10462) );
  XNOR2_X1 U13371 ( .A(n17337), .B(n10464), .ZN(n10465) );
  XOR2_X1 U13372 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n10465), .Z(
        n17801) );
  INV_X1 U13373 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17798) );
  XNOR2_X1 U13374 ( .A(n10614), .B(n10466), .ZN(n17788) );
  NAND2_X1 U13375 ( .A1(n17789), .A2(n17788), .ZN(n10467) );
  INV_X1 U13376 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18091) );
  XOR2_X1 U13377 ( .A(n10612), .B(n10468), .Z(n10469) );
  XOR2_X1 U13378 ( .A(n18091), .B(n10469), .Z(n17771) );
  AOI21_X1 U13379 ( .B1(n16318), .B2(n17327), .A(n17754), .ZN(n10471) );
  INV_X1 U13380 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18085) );
  INV_X1 U13381 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18070) );
  NAND2_X2 U13382 ( .A1(n10472), .A2(n18070), .ZN(n17735) );
  NAND2_X1 U13383 ( .A1(n18036), .A2(n17735), .ZN(n17758) );
  INV_X1 U13384 ( .A(n17758), .ZN(n18067) );
  NAND2_X1 U13385 ( .A1(n18067), .A2(n17754), .ZN(n17753) );
  INV_X1 U13386 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17690) );
  INV_X1 U13387 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18006) );
  NOR2_X1 U13388 ( .A1(n17690), .A2(n18006), .ZN(n17654) );
  INV_X1 U13389 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18063) );
  INV_X1 U13390 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17726) );
  NOR2_X1 U13391 ( .A1(n18063), .A2(n17726), .ZN(n18034) );
  NAND2_X1 U13392 ( .A1(n18034), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17702) );
  INV_X1 U13393 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18032) );
  NOR2_X1 U13394 ( .A1(n17702), .A2(n18032), .ZN(n17673) );
  AND2_X1 U13395 ( .A1(n17654), .A2(n17673), .ZN(n17976) );
  NAND2_X1 U13396 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17976), .ZN(
        n17967) );
  NOR4_X1 U13397 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10473) );
  NAND4_X1 U13398 ( .A1(n10473), .A2(n17690), .A3(n18006), .A4(n18032), .ZN(
        n10474) );
  OAI21_X1 U13399 ( .B1(n17735), .B2(n10474), .A(n17685), .ZN(n17636) );
  NAND2_X1 U13400 ( .A1(n17628), .A2(n17685), .ZN(n10475) );
  INV_X1 U13401 ( .A(n10475), .ZN(n17555) );
  INV_X1 U13402 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17963) );
  NOR2_X1 U13403 ( .A1(n17978), .A2(n17963), .ZN(n17962) );
  INV_X1 U13404 ( .A(n17962), .ZN(n17620) );
  INV_X1 U13405 ( .A(n17637), .ZN(n10478) );
  NOR2_X1 U13406 ( .A1(n17555), .A2(n17579), .ZN(n17580) );
  INV_X1 U13407 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17623) );
  NAND2_X1 U13408 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17582) );
  INV_X1 U13409 ( .A(n17582), .ZN(n17938) );
  NAND2_X1 U13410 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17938), .ZN(
        n17920) );
  OR2_X1 U13411 ( .A1(n17623), .A2(n17920), .ZN(n17914) );
  INV_X1 U13412 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17930) );
  NOR2_X1 U13413 ( .A1(n17914), .A2(n17930), .ZN(n16312) );
  INV_X1 U13414 ( .A(n16312), .ZN(n17881) );
  NOR2_X1 U13415 ( .A1(n17580), .A2(n17881), .ZN(n17554) );
  NAND2_X1 U13416 ( .A1(n17962), .A2(n16312), .ZN(n17853) );
  INV_X1 U13417 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17906) );
  OR2_X1 U13418 ( .A1(n17853), .A2(n17906), .ZN(n17523) );
  NAND2_X1 U13419 ( .A1(n17623), .A2(n17685), .ZN(n17617) );
  NOR2_X1 U13420 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17617), .ZN(
        n10476) );
  INV_X1 U13421 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21062) );
  NAND2_X1 U13422 ( .A1(n10476), .A2(n21062), .ZN(n17581) );
  NAND3_X1 U13423 ( .A1(n17569), .A2(n17930), .A3(n17906), .ZN(n10477) );
  AND2_X1 U13424 ( .A1(n10475), .A2(n10479), .ZN(n17533) );
  INV_X1 U13425 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17893) );
  NAND2_X1 U13426 ( .A1(n17533), .A2(n17893), .ZN(n17532) );
  NAND3_X1 U13427 ( .A1(n17554), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17532), .ZN(n10480) );
  INV_X1 U13428 ( .A(n10480), .ZN(n17526) );
  NAND2_X1 U13429 ( .A1(n17685), .A2(n17532), .ZN(n17525) );
  INV_X1 U13430 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17507) );
  NOR2_X1 U13431 ( .A1(n17871), .A2(n17507), .ZN(n12470) );
  INV_X1 U13432 ( .A(n12470), .ZN(n17860) );
  NAND2_X1 U13433 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17754), .ZN(
        n16315) );
  INV_X1 U13434 ( .A(n16264), .ZN(n10484) );
  NOR2_X2 U13435 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n10482), .ZN(
        n17490) );
  INV_X1 U13436 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17467) );
  NAND2_X1 U13437 ( .A1(n17467), .A2(n17685), .ZN(n16316) );
  INV_X1 U13438 ( .A(n16316), .ZN(n15670) );
  INV_X1 U13439 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16265) );
  AOI22_X1 U13440 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16882), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13441 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13442 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n9795), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13443 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10485) );
  NAND4_X1 U13444 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .ZN(
        n10494) );
  AOI22_X1 U13445 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16885), .B1(
        n9792), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13446 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9797), .ZN(n10491) );
  INV_X1 U13447 ( .A(n16884), .ZN(n17143) );
  AOI22_X1 U13448 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13449 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17163), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10489) );
  NAND4_X1 U13450 ( .A1(n10492), .A2(n10491), .A3(n10490), .A4(n10489), .ZN(
        n10493) );
  INV_X1 U13451 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18671) );
  NOR2_X1 U13452 ( .A1(n18671), .A2(n18661), .ZN(n18809) );
  NAND2_X1 U13453 ( .A1(n18779), .A2(n18809), .ZN(n18669) );
  AOI22_X1 U13454 ( .A1(n18641), .A2(n18645), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n10495), .ZN(n10608) );
  OAI22_X1 U13455 ( .A1(n10497), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18650), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10502) );
  OAI22_X1 U13456 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18654), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n10499), .ZN(n10506) );
  NOR2_X1 U13457 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18654), .ZN(
        n10500) );
  NAND2_X1 U13458 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10499), .ZN(
        n10505) );
  AOI22_X1 U13459 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n10506), .B1(
        n10500), .B2(n10505), .ZN(n10607) );
  NAND2_X1 U13460 ( .A1(n10503), .A2(n10502), .ZN(n10501) );
  OAI211_X1 U13461 ( .C1(n10503), .C2(n10502), .A(n10607), .B(n10501), .ZN(
        n10610) );
  AOI21_X1 U13462 ( .B1(n18796), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n10504), .ZN(n10606) );
  INV_X1 U13463 ( .A(n10606), .ZN(n10510) );
  XNOR2_X1 U13464 ( .A(n10608), .B(n10504), .ZN(n10509) );
  AND2_X1 U13465 ( .A1(n10505), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10507) );
  OAI22_X1 U13466 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18617), .B1(
        n10507), .B2(n10506), .ZN(n10508) );
  INV_X1 U13467 ( .A(n10508), .ZN(n10611) );
  INV_X1 U13468 ( .A(n18607), .ZN(n12455) );
  OAI21_X1 U13469 ( .B1(n10610), .B2(n10510), .A(n12455), .ZN(n18608) );
  INV_X4 U13470 ( .A(n10328), .ZN(n17161) );
  AOI22_X1 U13471 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9797), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10515) );
  INV_X1 U13472 ( .A(n10511), .ZN(n16878) );
  AOI22_X1 U13473 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16878), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13474 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13475 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10512) );
  NAND4_X1 U13476 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10522) );
  AOI22_X1 U13477 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16916), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13478 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13479 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13480 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10517) );
  NAND4_X1 U13481 ( .A1(n10520), .A2(n10519), .A3(n10518), .A4(n10517), .ZN(
        n10521) );
  AOI22_X1 U13482 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13483 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U13484 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U13485 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10523) );
  NAND4_X1 U13486 ( .A1(n10526), .A2(n10525), .A3(n10524), .A4(n10523), .ZN(
        n10532) );
  AOI22_X1 U13487 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13488 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13489 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13490 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10527) );
  NAND4_X1 U13491 ( .A1(n10530), .A2(n10529), .A3(n10528), .A4(n10527), .ZN(
        n10531) );
  AOI22_X1 U13492 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13493 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13494 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13495 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10533) );
  NAND4_X1 U13496 ( .A1(n10536), .A2(n10535), .A3(n10534), .A4(n10533), .ZN(
        n10542) );
  AOI22_X1 U13497 ( .A1(n10387), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13498 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13499 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13500 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10537) );
  NAND4_X1 U13501 ( .A1(n10540), .A2(n10539), .A3(n10538), .A4(n10537), .ZN(
        n10541) );
  AOI22_X1 U13502 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13503 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U13504 ( .A1(n10396), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10543) );
  OAI21_X1 U13505 ( .B1(n10328), .B2(n16870), .A(n10543), .ZN(n10550) );
  AOI22_X1 U13506 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9788), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10548) );
  INV_X2 U13507 ( .A(n16858), .ZN(n17158) );
  AOI22_X1 U13508 ( .A1(n16878), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10547) );
  INV_X1 U13509 ( .A(n10544), .ZN(n17145) );
  INV_X2 U13510 ( .A(n16871), .ZN(n17137) );
  AOI22_X1 U13511 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13512 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10545) );
  NAND4_X1 U13513 ( .A1(n10548), .A2(n10547), .A3(n10546), .A4(n10545), .ZN(
        n10549) );
  NAND3_X2 U13514 ( .A1(n10553), .A2(n10552), .A3(n10551), .ZN(n17248) );
  NAND2_X1 U13515 ( .A1(n18172), .A2(n17248), .ZN(n10591) );
  AOI22_X1 U13516 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16885), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13517 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13518 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13519 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10554) );
  NAND4_X1 U13520 ( .A1(n10557), .A2(n10556), .A3(n10555), .A4(n10554), .ZN(
        n10563) );
  AOI22_X1 U13521 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13522 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13523 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13524 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10397), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10558) );
  NAND4_X1 U13525 ( .A1(n10561), .A2(n10560), .A3(n10559), .A4(n10558), .ZN(
        n10562) );
  AOI22_X1 U13526 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13527 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9792), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13528 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10564) );
  OAI21_X1 U13529 ( .B1(n10511), .B2(n21164), .A(n10564), .ZN(n10571) );
  AOI22_X1 U13530 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13531 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13532 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13533 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10566) );
  NAND4_X1 U13534 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n10570) );
  AOI211_X1 U13535 ( .C1(n17161), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n10571), .B(n10570), .ZN(n10572) );
  NAND3_X1 U13536 ( .A1(n10574), .A2(n10573), .A3(n10572), .ZN(n10602) );
  NOR2_X1 U13537 ( .A1(n18194), .A2(n10602), .ZN(n10585) );
  NAND3_X1 U13538 ( .A1(n18185), .A2(n10592), .A3(n10585), .ZN(n10596) );
  AOI22_X1 U13539 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13540 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10577) );
  AOI22_X1 U13541 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9797), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U13542 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10575) );
  NAND4_X1 U13543 ( .A1(n10578), .A2(n10577), .A3(n10576), .A4(n10575), .ZN(
        n10584) );
  AOI22_X1 U13544 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10582) );
  AOI22_X1 U13545 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10581) );
  AOI22_X1 U13546 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10580) );
  AOI22_X1 U13547 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10579) );
  NAND4_X1 U13548 ( .A1(n10582), .A2(n10581), .A3(n10580), .A4(n10579), .ZN(
        n10583) );
  NAND2_X1 U13549 ( .A1(n18181), .A2(n10595), .ZN(n12456) );
  NAND2_X1 U13550 ( .A1(n12456), .A2(n10594), .ZN(n10601) );
  INV_X1 U13551 ( .A(n18199), .ZN(n15663) );
  NOR2_X1 U13552 ( .A1(n18194), .A2(n15663), .ZN(n18638) );
  NOR2_X1 U13553 ( .A1(n18172), .A2(n16819), .ZN(n10600) );
  OAI21_X1 U13554 ( .B1(n18206), .B2(n18638), .A(n10600), .ZN(n12459) );
  OR2_X1 U13555 ( .A1(n12456), .A2(n18199), .ZN(n12457) );
  AOI21_X1 U13556 ( .B1(n10594), .B2(n12457), .A(n16818), .ZN(n10590) );
  NOR2_X1 U13557 ( .A1(n18194), .A2(n18199), .ZN(n10587) );
  NOR2_X1 U13558 ( .A1(n18206), .A2(n10587), .ZN(n10588) );
  INV_X1 U13559 ( .A(n18181), .ZN(n12453) );
  NOR3_X1 U13560 ( .A1(n10599), .A2(n10585), .A3(n12453), .ZN(n10586) );
  OAI22_X1 U13561 ( .A1(n18190), .A2(n10588), .B1(n10587), .B2(n10586), .ZN(
        n10589) );
  AOI211_X1 U13562 ( .C1(n18185), .C2(n10591), .A(n10590), .B(n10589), .ZN(
        n12460) );
  OAI211_X1 U13563 ( .C1(n18185), .C2(n10601), .A(n12459), .B(n12460), .ZN(
        n10604) );
  NAND2_X1 U13564 ( .A1(n18181), .A2(n18185), .ZN(n18621) );
  NAND2_X1 U13565 ( .A1(n18813), .A2(n10592), .ZN(n10598) );
  NOR4_X4 U13566 ( .A1(n18172), .A2(n10595), .A3(n10594), .A4(n10593), .ZN(
        n17417) );
  INV_X1 U13567 ( .A(n10599), .ZN(n10597) );
  NOR2_X2 U13568 ( .A1(n13968), .A2(n13969), .ZN(n18639) );
  NOR2_X1 U13569 ( .A1(n10600), .A2(n10599), .ZN(n18825) );
  NAND2_X1 U13570 ( .A1(n18199), .A2(n10602), .ZN(n18622) );
  NOR2_X1 U13571 ( .A1(n18813), .A2(n10603), .ZN(n10605) );
  AOI21_X1 U13572 ( .B1(n10605), .B2(n16436), .A(n10604), .ZN(n18620) );
  XNOR2_X1 U13573 ( .A(n16819), .B(n12453), .ZN(n12454) );
  NAND3_X1 U13574 ( .A1(n10608), .A2(n10607), .A3(n10606), .ZN(n10609) );
  NAND3_X1 U13575 ( .A1(n10611), .A2(n10610), .A3(n10609), .ZN(n13975) );
  NOR2_X4 U13576 ( .A1(n18813), .A2(n16418), .ZN(n17838) );
  NAND2_X1 U13577 ( .A1(n12468), .A2(n17755), .ZN(n10656) );
  INV_X1 U13578 ( .A(n10612), .ZN(n17330) );
  NAND2_X1 U13579 ( .A1(n10616), .A2(n10615), .ZN(n10628) );
  NAND2_X1 U13580 ( .A1(n10613), .A2(n10614), .ZN(n10634) );
  NOR2_X1 U13581 ( .A1(n17330), .A2(n10634), .ZN(n10637) );
  NAND2_X1 U13582 ( .A1(n10637), .A2(n16317), .ZN(n10638) );
  XOR2_X1 U13583 ( .A(n10614), .B(n10613), .Z(n10632) );
  XNOR2_X1 U13584 ( .A(n10616), .B(n10617), .ZN(n10626) );
  AND2_X1 U13585 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n10626), .ZN(
        n10627) );
  AOI21_X1 U13586 ( .B1(n10618), .B2(n17844), .A(n10617), .ZN(n10619) );
  NOR2_X1 U13587 ( .A1(n10619), .A2(n10459), .ZN(n10625) );
  XOR2_X1 U13588 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10619), .Z(
        n17827) );
  INV_X1 U13589 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21150) );
  NOR2_X1 U13590 ( .A1(n10621), .A2(n21150), .ZN(n10623) );
  NAND3_X1 U13591 ( .A1(n10622), .A2(n10621), .A3(n21150), .ZN(n10620) );
  OAI221_X1 U13592 ( .B1(n10623), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n10622), .C2(n10621), .A(n10620), .ZN(n17826) );
  NOR2_X1 U13593 ( .A1(n17827), .A2(n17826), .ZN(n10624) );
  NOR2_X1 U13594 ( .A1(n10625), .A2(n10624), .ZN(n17816) );
  XOR2_X1 U13595 ( .A(n17811), .B(n10626), .Z(n17815) );
  NOR2_X1 U13596 ( .A1(n17816), .A2(n17815), .ZN(n17814) );
  XNOR2_X1 U13597 ( .A(n17337), .B(n10628), .ZN(n10630) );
  NOR2_X1 U13598 ( .A1(n10629), .A2(n10630), .ZN(n10631) );
  XNOR2_X1 U13599 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n10632), .ZN(
        n17785) );
  XNOR2_X1 U13600 ( .A(n17330), .B(n10634), .ZN(n10636) );
  XOR2_X1 U13601 ( .A(n16317), .B(n10637), .Z(n10640) );
  INV_X1 U13602 ( .A(n10638), .ZN(n10643) );
  NAND2_X1 U13603 ( .A1(n10640), .A2(n10639), .ZN(n17761) );
  OAI21_X1 U13604 ( .B1(n10643), .B2(n10642), .A(n17761), .ZN(n10641) );
  INV_X1 U13605 ( .A(n17673), .ZN(n17999) );
  NAND2_X1 U13606 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17882) );
  INV_X1 U13607 ( .A(n17882), .ZN(n17854) );
  NAND2_X1 U13608 ( .A1(n17854), .A2(n12470), .ZN(n17851) );
  NOR2_X1 U13609 ( .A1(n17853), .A2(n17851), .ZN(n12471) );
  NAND2_X1 U13610 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16295) );
  INV_X1 U13611 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16284) );
  NOR2_X1 U13612 ( .A1(n16295), .A2(n16284), .ZN(n16304) );
  INV_X1 U13613 ( .A(n16304), .ZN(n12474) );
  INV_X1 U13614 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17989) );
  NAND2_X1 U13615 ( .A1(n17654), .A2(n18016), .ZN(n17661) );
  NAND2_X1 U13616 ( .A1(n12471), .A2(n17982), .ZN(n17855) );
  NOR2_X1 U13617 ( .A1(n12474), .A2(n17855), .ZN(n16282) );
  OAI22_X1 U13618 ( .A1(n16277), .A2(n17850), .B1(n16282), .B2(n17759), .ZN(
        n10644) );
  AND2_X1 U13619 ( .A1(n10644), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10654) );
  NAND2_X1 U13620 ( .A1(n18779), .A2(n18515), .ZN(n18824) );
  NAND2_X1 U13621 ( .A1(n18661), .A2(n18515), .ZN(n16413) );
  NAND2_X1 U13622 ( .A1(n18824), .A2(n16413), .ZN(n18159) );
  INV_X1 U13623 ( .A(n18159), .ZN(n18808) );
  INV_X1 U13624 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18812) );
  NOR2_X1 U13625 ( .A1(n18779), .A2(n18812), .ZN(n17803) );
  NOR2_X2 U13626 ( .A1(n17818), .A2(n17803), .ZN(n17842) );
  INV_X1 U13627 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17841) );
  NAND2_X1 U13628 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17746) );
  INV_X1 U13629 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17588) );
  INV_X1 U13630 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n20966) );
  INV_X1 U13631 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17577) );
  NOR2_X1 U13632 ( .A1(n20966), .A2(n17577), .ZN(n17567) );
  NAND2_X1 U13633 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17520) );
  NAND2_X1 U13634 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17502), .ZN(
        n17477) );
  NAND2_X1 U13635 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17471) );
  INV_X1 U13636 ( .A(n10648), .ZN(n16290) );
  INV_X1 U13637 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n21077) );
  AOI22_X1 U13638 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16286), .B1(
        n10647), .B2(n21077), .ZN(n16474) );
  NAND2_X1 U13639 ( .A1(n10648), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10650) );
  NAND2_X1 U13640 ( .A1(n18671), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17846) );
  INV_X1 U13641 ( .A(n17846), .ZN(n17675) );
  NAND2_X1 U13642 ( .A1(n18617), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18781) );
  OAI221_X1 U13643 ( .B1(n18661), .B2(P3_STATE2_REG_1__SCAN_IN), .C1(
        P3_STATE2_REG_2__SCAN_IN), .C2(n18779), .A(n18781), .ZN(n18170) );
  NAND3_X1 U13644 ( .A1(n18661), .A2(n18515), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18512) );
  NOR2_X1 U13645 ( .A1(n18251), .A2(n18512), .ZN(n10649) );
  OAI21_X1 U13646 ( .B1(n17841), .B2(n17564), .A(n18464), .ZN(n17678) );
  INV_X1 U13647 ( .A(n17678), .ZN(n17694) );
  OR2_X1 U13648 ( .A1(n10650), .A2(n17694), .ZN(n16275) );
  NOR2_X1 U13649 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17564), .ZN(
        n16287) );
  NAND2_X1 U13650 ( .A1(n18552), .A2(n10650), .ZN(n16291) );
  OAI211_X1 U13651 ( .C1(n16285), .C2(n17846), .A(n16291), .B(n17845), .ZN(
        n16294) );
  NOR2_X1 U13652 ( .A1(n16287), .A2(n16294), .ZN(n16273) );
  NOR3_X1 U13653 ( .A1(n18824), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n16272) );
  NAND2_X1 U13654 ( .A1(n9790), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n12480) );
  OAI221_X1 U13655 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16275), .C1(
        n21077), .C2(n16273), .A(n12480), .ZN(n10651) );
  AOI21_X1 U13656 ( .B1(n17604), .B2(n16474), .A(n10651), .ZN(n10652) );
  INV_X1 U13657 ( .A(n18037), .ZN(n16309) );
  NOR2_X2 U13658 ( .A1(n17745), .A2(n17967), .ZN(n17633) );
  NAND2_X1 U13659 ( .A1(n12471), .A2(n17633), .ZN(n17496) );
  NAND2_X1 U13660 ( .A1(n16304), .A2(n16265), .ZN(n12479) );
  NAND2_X1 U13661 ( .A1(n10656), .A2(n10655), .ZN(P3_U2800) );
  AND2_X4 U13662 ( .A1(n13531), .A2(n15562), .ZN(n10851) );
  AOI22_X1 U13663 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10658) );
  AND2_X4 U13664 ( .A1(n10858), .A2(n15562), .ZN(n10864) );
  AOI22_X1 U13665 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10657) );
  AND3_X1 U13666 ( .A1(n10658), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10657), .ZN(n10661) );
  AND2_X4 U13667 ( .A1(n13531), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10743) );
  AOI22_X1 U13668 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10660) );
  AND3_X4 U13669 ( .A1(n15562), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n16211), .ZN(n12636) );
  AND3_X4 U13670 ( .A1(n10795), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U13671 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U13672 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13673 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13674 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U13675 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13676 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13677 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U13678 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13679 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13680 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13681 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13682 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13683 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10680) );
  NAND4_X1 U13684 ( .A1(n10683), .A2(n10682), .A3(n10681), .A4(n10680), .ZN(
        n10684) );
  NAND2_X1 U13685 ( .A1(n10684), .A2(n10676), .ZN(n10691) );
  AOI22_X1 U13686 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13687 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13688 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13689 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10685) );
  NAND4_X1 U13690 ( .A1(n10688), .A2(n10687), .A3(n10686), .A4(n10685), .ZN(
        n10689) );
  NAND2_X1 U13691 ( .A1(n10689), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10690) );
  AOI22_X1 U13692 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13693 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13694 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13695 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13696 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13697 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U13698 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13699 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13700 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13701 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13702 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10700) );
  NAND4_X1 U13703 ( .A1(n10703), .A2(n10702), .A3(n10701), .A4(n10700), .ZN(
        n10704) );
  AOI22_X1 U13704 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U13705 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13706 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10705) );
  NAND4_X1 U13707 ( .A1(n10708), .A2(n10707), .A3(n10706), .A4(n10705), .ZN(
        n10709) );
  INV_X1 U13708 ( .A(n15625), .ZN(n10776) );
  AOI22_X1 U13709 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13710 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U13711 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13712 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10851), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13713 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10717) );
  AND2_X1 U13714 ( .A1(n10717), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10721) );
  AOI22_X1 U13715 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13716 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10719) );
  AOI22_X1 U13717 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10851), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10718) );
  NAND4_X1 U13718 ( .A1(n10721), .A2(n10720), .A3(n10719), .A4(n10718), .ZN(
        n10722) );
  INV_X1 U13719 ( .A(n13572), .ZN(n11740) );
  INV_X1 U13720 ( .A(n10771), .ZN(n10737) );
  AOI22_X1 U13721 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U13722 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U13723 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13724 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10725) );
  NAND4_X1 U13725 ( .A1(n10728), .A2(n10727), .A3(n10726), .A4(n10725), .ZN(
        n10729) );
  AOI22_X1 U13726 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U13727 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U13728 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13729 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10730) );
  NAND4_X1 U13730 ( .A1(n10733), .A2(n10732), .A3(n10731), .A4(n10730), .ZN(
        n10734) );
  NAND2_X4 U13731 ( .A1(n10736), .A2(n10735), .ZN(n16231) );
  AOI22_X1 U13732 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U13733 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10738) );
  NAND4_X1 U13734 ( .A1(n10741), .A2(n10740), .A3(n10739), .A4(n10738), .ZN(
        n10742) );
  AOI22_X1 U13735 ( .A1(n10851), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10866), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13736 ( .A1(n12636), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10877), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13737 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10745) );
  NAND4_X1 U13738 ( .A1(n10747), .A2(n10746), .A3(n10745), .A4(n10744), .ZN(
        n10748) );
  INV_X1 U13739 ( .A(n15625), .ZN(n10751) );
  INV_X1 U13740 ( .A(n10753), .ZN(n15635) );
  INV_X4 U13741 ( .A(n15635), .ZN(n12817) );
  NAND3_X1 U13742 ( .A1(n11739), .A2(n12817), .A3(n9882), .ZN(n10752) );
  AND2_X2 U13743 ( .A1(n11437), .A2(n10752), .ZN(n10797) );
  NAND2_X1 U13744 ( .A1(n10753), .A2(n10754), .ZN(n10773) );
  INV_X1 U13745 ( .A(n10753), .ZN(n10759) );
  AND2_X2 U13746 ( .A1(n11451), .A2(n16231), .ZN(n11721) );
  NAND2_X1 U13747 ( .A1(n11721), .A2(n11467), .ZN(n10757) );
  NAND3_X1 U13748 ( .A1(n10797), .A2(n10786), .A3(n10757), .ZN(n10758) );
  AND2_X2 U13749 ( .A1(n10758), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10805) );
  INV_X2 U13750 ( .A(n11071), .ZN(n11397) );
  NOR2_X2 U13751 ( .A1(n10785), .A2(n10778), .ZN(n11746) );
  NAND2_X1 U13752 ( .A1(n9805), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10763) );
  NAND2_X2 U13753 ( .A1(n11721), .A2(n12758), .ZN(n10815) );
  INV_X1 U13754 ( .A(n10815), .ZN(n10760) );
  NOR2_X1 U13755 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19894) );
  INV_X1 U13756 ( .A(n19894), .ZN(n16250) );
  NAND3_X1 U13757 ( .A1(n10763), .A2(n10762), .A3(n10761), .ZN(n10764) );
  AOI21_X1 U13758 ( .B1(n10805), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n10764), .ZN(n10784) );
  AND2_X1 U13759 ( .A1(n13572), .A2(n15625), .ZN(n10765) );
  NAND3_X1 U13760 ( .A1(n10770), .A2(n10769), .A3(n10768), .ZN(n10772) );
  NAND3_X1 U13761 ( .A1(n10772), .A2(n10771), .A3(n11443), .ZN(n11743) );
  NAND2_X1 U13762 ( .A1(n10774), .A2(n10773), .ZN(n11440) );
  INV_X1 U13763 ( .A(n11440), .ZN(n10775) );
  INV_X1 U13764 ( .A(n10778), .ZN(n11738) );
  INV_X1 U13765 ( .A(n11738), .ZN(n11733) );
  NAND2_X1 U13766 ( .A1(n11438), .A2(n11467), .ZN(n11735) );
  NAND2_X1 U13767 ( .A1(n10784), .A2(n10821), .ZN(n10828) );
  NAND2_X1 U13768 ( .A1(n10786), .A2(n10785), .ZN(n10788) );
  INV_X1 U13769 ( .A(n11746), .ZN(n12828) );
  NAND2_X1 U13770 ( .A1(n15582), .A2(n15562), .ZN(n10787) );
  NAND2_X1 U13771 ( .A1(n19894), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10789) );
  INV_X1 U13772 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10793) );
  NAND2_X1 U13773 ( .A1(n10816), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10792) );
  NAND2_X1 U13774 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10791) );
  OAI211_X1 U13775 ( .C1(n10793), .C2(n10815), .A(n10792), .B(n10791), .ZN(
        n10794) );
  AOI21_X2 U13776 ( .B1(n10805), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10794), .ZN(n10800) );
  INV_X1 U13777 ( .A(n10800), .ZN(n10801) );
  OR2_X1 U13778 ( .A1(n10802), .A2(n10801), .ZN(n10803) );
  AOI21_X1 U13779 ( .B1(n19904), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10804) );
  INV_X1 U13780 ( .A(n10805), .ZN(n11300) );
  INV_X1 U13781 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10808) );
  NAND2_X1 U13782 ( .A1(n9805), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10807) );
  NAND2_X1 U13783 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10806) );
  OAI211_X1 U13784 ( .C1(n10808), .C2(n10815), .A(n10807), .B(n10806), .ZN(
        n10809) );
  INV_X1 U13785 ( .A(n10809), .ZN(n10810) );
  NAND2_X2 U13786 ( .A1(n10811), .A2(n10810), .ZN(n10823) );
  INV_X1 U13787 ( .A(n10822), .ZN(n10813) );
  INV_X1 U13788 ( .A(n10823), .ZN(n10812) );
  BUF_X4 U13789 ( .A(n10815), .Z(n11380) );
  BUF_X8 U13790 ( .A(n9805), .Z(n11387) );
  NAND2_X1 U13791 ( .A1(n11387), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10818) );
  NAND2_X1 U13792 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10817) );
  OAI211_X1 U13793 ( .C1(n19789), .C2(n11380), .A(n10818), .B(n10817), .ZN(
        n10819) );
  AOI21_X2 U13794 ( .B1(n10820), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10819), .ZN(n11295) );
  INV_X1 U13795 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19858) );
  OAI22_X1 U13796 ( .A1(n10821), .A2(n10676), .B1(n16250), .B2(n19858), .ZN(
        n11297) );
  XNOR2_X2 U13797 ( .A(n11295), .B(n11297), .ZN(n11293) );
  INV_X1 U13798 ( .A(n10825), .ZN(n10832) );
  XNOR2_X2 U13799 ( .A(n10832), .B(n10826), .ZN(n12489) );
  INV_X1 U13800 ( .A(n10827), .ZN(n10830) );
  INV_X1 U13801 ( .A(n10828), .ZN(n10829) );
  NAND2_X1 U13802 ( .A1(n10830), .A2(n10829), .ZN(n10831) );
  AND2_X2 U13803 ( .A1(n10833), .A2(n10842), .ZN(n15603) );
  AND2_X1 U13804 ( .A1(n10845), .A2(n10842), .ZN(n10989) );
  AND2_X2 U13805 ( .A1(n10833), .A2(n10839), .ZN(n19281) );
  AND2_X2 U13806 ( .A1(n10833), .A2(n10844), .ZN(n19316) );
  AOI22_X1 U13807 ( .A1(n10990), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n19316), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10834) );
  AND2_X2 U13808 ( .A1(n10838), .A2(n9956), .ZN(n10841) );
  AND2_X2 U13809 ( .A1(n10841), .A2(n10839), .ZN(n19408) );
  INV_X1 U13810 ( .A(n19374), .ZN(n11004) );
  AND2_X2 U13811 ( .A1(n10841), .A2(n10842), .ZN(n19346) );
  AOI22_X1 U13812 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11004), .B1(
        n19346), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10848) );
  AND2_X2 U13813 ( .A1(n10841), .A2(n10844), .ZN(n19436) );
  INV_X1 U13814 ( .A(n10852), .ZN(n10853) );
  NAND2_X1 U13815 ( .A1(n12570), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10876) );
  NOR2_X1 U13816 ( .A1(n10795), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10854) );
  AND2_X2 U13817 ( .A1(n12633), .A2(n10854), .ZN(n12661) );
  AND2_X1 U13818 ( .A1(n10795), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10855) );
  AOI22_X1 U13819 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12661), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10863) );
  NAND2_X1 U13820 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10862) );
  AND2_X2 U13821 ( .A1(n14310), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10902) );
  NAND2_X1 U13822 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10861) );
  AND2_X1 U13823 ( .A1(n12633), .A2(n10856), .ZN(n10857) );
  AND2_X1 U13824 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U13825 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10860) );
  NAND4_X1 U13826 ( .A1(n10863), .A2(n10862), .A3(n10861), .A4(n10860), .ZN(
        n10874) );
  INV_X2 U13827 ( .A(n11629), .ZN(n12668) );
  NAND2_X1 U13828 ( .A1(n12668), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10872) );
  INV_X1 U13829 ( .A(n10866), .ZN(n13529) );
  NAND2_X2 U13830 ( .A1(n10867), .A2(n10676), .ZN(n15588) );
  NAND2_X1 U13831 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10871) );
  BUF_X1 U13832 ( .A(n12632), .Z(n10868) );
  INV_X1 U13833 ( .A(n10868), .ZN(n10869) );
  OR2_X2 U13834 ( .A1(n10869), .A2(n10676), .ZN(n12653) );
  NAND2_X1 U13835 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10870) );
  NAND3_X1 U13836 ( .A1(n10872), .A2(n10871), .A3(n10870), .ZN(n10873) );
  NOR2_X1 U13837 ( .A1(n10874), .A2(n10873), .ZN(n10875) );
  AND2_X2 U13838 ( .A1(n12780), .A2(n10676), .ZN(n12666) );
  AND2_X2 U13839 ( .A1(n12780), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10918) );
  AOI22_X1 U13840 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12666), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10884) );
  BUF_X1 U13841 ( .A(n12636), .Z(n10878) );
  AND2_X2 U13842 ( .A1(n10878), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10937) );
  AOI22_X1 U13843 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10883) );
  BUF_X1 U13844 ( .A(n12639), .Z(n10880) );
  NAND2_X2 U13845 ( .A1(n10880), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11631) );
  NAND2_X1 U13846 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10882) );
  NAND2_X1 U13847 ( .A1(n12572), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10881) );
  NAND4_X1 U13848 ( .A1(n10884), .A2(n10883), .A3(n10882), .A4(n10881), .ZN(
        n10885) );
  NOR2_X1 U13849 ( .A1(n10886), .A2(n10885), .ZN(n11521) );
  NAND2_X1 U13850 ( .A1(n19903), .A2(n11521), .ZN(n10887) );
  AOI22_X1 U13851 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19316), .B1(
        n19436), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U13852 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19346), .B1(
        n10997), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U13853 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n13565), .B1(
        n10995), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U13854 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19281), .B1(
        n10988), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10889) );
  AND4_X1 U13855 ( .A1(n10892), .A2(n10891), .A3(n10890), .A4(n10889), .ZN(
        n10901) );
  AOI22_X1 U13856 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n15603), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10899) );
  INV_X1 U13857 ( .A(n19374), .ZN(n10893) );
  AOI21_X1 U13858 ( .B1(n10893), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n19903), .ZN(n10894) );
  AOI22_X1 U13859 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10989), .B1(
        n10987), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10897) );
  AND4_X2 U13860 ( .A1(n10899), .A2(n10898), .A3(n10897), .A4(n10896), .ZN(
        n10900) );
  NAND2_X1 U13861 ( .A1(n10901), .A2(n10900), .ZN(n10952) );
  AOI22_X1 U13862 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12571), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U13863 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U13864 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10905) );
  INV_X1 U13865 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11470) );
  INV_X1 U13866 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n21017) );
  OAI22_X1 U13867 ( .A1(n12653), .A2(n11470), .B1(n12654), .B2(n21017), .ZN(
        n10903) );
  INV_X1 U13868 ( .A(n10903), .ZN(n10904) );
  NAND4_X1 U13869 ( .A1(n10907), .A2(n10906), .A3(n10905), .A4(n10904), .ZN(
        n10913) );
  AOI22_X1 U13870 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13871 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13872 ( .A1(n12572), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13873 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10908) );
  NAND4_X1 U13874 ( .A1(n10911), .A2(n10910), .A3(n10909), .A4(n10908), .ZN(
        n10912) );
  NOR2_X1 U13875 ( .A1(n10913), .A2(n10912), .ZN(n11494) );
  OR2_X1 U13876 ( .A1(n11494), .A2(n15614), .ZN(n10953) );
  INV_X1 U13877 ( .A(n10953), .ZN(n13014) );
  INV_X1 U13878 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11544) );
  INV_X1 U13879 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12538) );
  OAI22_X1 U13880 ( .A1(n11544), .A2(n12653), .B1(n12654), .B2(n12538), .ZN(
        n10916) );
  INV_X1 U13881 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10914) );
  INV_X1 U13882 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11541) );
  OAI22_X1 U13883 ( .A1(n10914), .A2(n12656), .B1(n15588), .B2(n11541), .ZN(
        n10915) );
  NOR2_X1 U13884 ( .A1(n10916), .A2(n10915), .ZN(n10931) );
  INV_X1 U13885 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10917) );
  INV_X1 U13886 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12536) );
  OAI22_X1 U13887 ( .A1(n10917), .A2(n11631), .B1(n11629), .B2(n12536), .ZN(
        n10924) );
  NAND2_X1 U13888 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10922) );
  NAND2_X1 U13889 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10921) );
  NAND2_X1 U13890 ( .A1(n10918), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10920) );
  NAND2_X1 U13891 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10919) );
  NAND4_X1 U13892 ( .A1(n10922), .A2(n10921), .A3(n10920), .A4(n10919), .ZN(
        n10923) );
  NOR2_X1 U13893 ( .A1(n10924), .A2(n10923), .ZN(n10930) );
  AOI22_X1 U13894 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12661), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10928) );
  NAND2_X1 U13895 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10927) );
  NAND2_X1 U13896 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10926) );
  AOI22_X1 U13897 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10925) );
  NAND3_X1 U13898 ( .A1(n10931), .A2(n10930), .A3(n10929), .ZN(n11505) );
  NAND2_X1 U13899 ( .A1(n13014), .A2(n11505), .ZN(n10956) );
  INV_X1 U13900 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11565) );
  INV_X1 U13901 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11561) );
  OAI22_X1 U13902 ( .A1(n11565), .A2(n12653), .B1(n12654), .B2(n11561), .ZN(
        n10934) );
  INV_X1 U13903 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11562) );
  INV_X1 U13904 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10932) );
  OAI22_X1 U13905 ( .A1(n11562), .A2(n15588), .B1(n11629), .B2(n10932), .ZN(
        n10933) );
  NOR2_X1 U13906 ( .A1(n10934), .A2(n10933), .ZN(n10950) );
  INV_X1 U13907 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10936) );
  INV_X1 U13908 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10935) );
  OAI22_X1 U13909 ( .A1(n10936), .A2(n12656), .B1(n11631), .B2(n10935), .ZN(
        n10943) );
  NAND2_X1 U13910 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10941) );
  NAND2_X1 U13911 ( .A1(n10918), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10940) );
  NAND2_X1 U13912 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10939) );
  NAND2_X1 U13913 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10938) );
  NAND4_X1 U13914 ( .A1(n10941), .A2(n10940), .A3(n10939), .A4(n10938), .ZN(
        n10942) );
  NOR2_X1 U13915 ( .A1(n10943), .A2(n10942), .ZN(n10949) );
  AOI22_X1 U13916 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12661), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10948) );
  NAND2_X1 U13917 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10947) );
  NAND2_X1 U13918 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10946) );
  AOI22_X1 U13919 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10945) );
  AND2_X1 U13920 ( .A1(n10953), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13013) );
  XNOR2_X1 U13921 ( .A(n11494), .B(n11505), .ZN(n10954) );
  NAND2_X1 U13922 ( .A1(n13013), .A2(n10954), .ZN(n10955) );
  XOR2_X1 U13923 ( .A(n10954), .B(n13013), .Z(n13006) );
  NAND2_X1 U13924 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13006), .ZN(
        n13005) );
  NAND2_X1 U13925 ( .A1(n10955), .A2(n13005), .ZN(n10957) );
  XNOR2_X1 U13926 ( .A(n9801), .B(n10957), .ZN(n14335) );
  XNOR2_X1 U13927 ( .A(n11515), .B(n10956), .ZN(n14334) );
  NAND2_X1 U13928 ( .A1(n14335), .A2(n14334), .ZN(n14333) );
  NAND2_X1 U13929 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10957), .ZN(
        n10958) );
  NAND2_X1 U13930 ( .A1(n14333), .A2(n10958), .ZN(n10959) );
  INV_X1 U13931 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21168) );
  XNOR2_X1 U13932 ( .A(n10959), .B(n21168), .ZN(n13548) );
  NAND2_X1 U13933 ( .A1(n13547), .A2(n13548), .ZN(n10961) );
  NAND2_X1 U13934 ( .A1(n10959), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10960) );
  INV_X1 U13935 ( .A(n10985), .ZN(n10981) );
  AOI22_X1 U13936 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11020), .B1(
        n10902), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U13937 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12569), .B1(
        n12570), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10973) );
  INV_X1 U13938 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10965) );
  INV_X1 U13939 ( .A(n12661), .ZN(n10964) );
  INV_X1 U13940 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10963) );
  OAI22_X1 U13941 ( .A1(n10965), .A2(n10964), .B1(n11015), .B2(n10963), .ZN(
        n10970) );
  INV_X1 U13942 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10967) );
  INV_X1 U13943 ( .A(n12660), .ZN(n10966) );
  INV_X1 U13944 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15634) );
  OAI22_X1 U13945 ( .A1(n10968), .A2(n10967), .B1(n10966), .B2(n15634), .ZN(
        n10969) );
  NOR2_X1 U13946 ( .A1(n10970), .A2(n10969), .ZN(n10972) );
  AOI22_X1 U13947 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12572), .B1(
        n12571), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10971) );
  NAND4_X1 U13948 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(
        n10980) );
  AOI22_X1 U13949 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12667), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U13950 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U13951 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10937), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10976) );
  NAND3_X1 U13952 ( .A1(n10978), .A2(n10977), .A3(n10976), .ZN(n10979) );
  INV_X1 U13953 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13623) );
  AOI22_X1 U13954 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19408), .B1(
        n10986), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U13955 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n15603), .B1(
        n10987), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U13956 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n10988), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U13957 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19316), .B1(
        n10990), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U13958 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n11004), .B1(
        n10995), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U13959 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19346), .B1(
        n13565), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U13960 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19436), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U13961 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19281), .B1(
        n10997), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10998) );
  INV_X1 U13962 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13624) );
  AOI22_X1 U13963 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11004), .B1(
        n10995), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U13964 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19346), .B1(
        n10996), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11007) );
  AOI22_X1 U13965 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10986), .B1(
        n10997), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U13966 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n15603), .B1(
        n10990), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11005) );
  NAND4_X1 U13967 ( .A1(n11008), .A2(n11007), .A3(n11006), .A4(n11005), .ZN(
        n11014) );
  AOI22_X1 U13968 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n13565), .B1(
        n19436), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11012) );
  AOI22_X1 U13969 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19281), .B1(
        n19408), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U13970 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10987), .B1(
        n10988), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U13971 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19316), .B1(
        n10989), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11009) );
  NAND4_X1 U13972 ( .A1(n11012), .A2(n11011), .A3(n11010), .A4(n11009), .ZN(
        n11013) );
  AOI22_X1 U13973 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10857), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U13974 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10975), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11018) );
  NAND2_X1 U13975 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11017) );
  NAND2_X1 U13976 ( .A1(n12570), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11016) );
  NAND4_X1 U13977 ( .A1(n11019), .A2(n11018), .A3(n11017), .A4(n11016), .ZN(
        n11026) );
  NAND2_X1 U13978 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11024) );
  NAND2_X1 U13979 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11023) );
  NAND2_X1 U13980 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11022) );
  NAND2_X1 U13981 ( .A1(n12572), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11021) );
  NAND4_X1 U13982 ( .A1(n11024), .A2(n11023), .A3(n11022), .A4(n11021), .ZN(
        n11025) );
  NOR2_X1 U13983 ( .A1(n11026), .A2(n11025), .ZN(n11031) );
  AOI22_X1 U13984 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n12667), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U13985 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n12660), .ZN(n11028) );
  AOI22_X1 U13986 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10937), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11027) );
  AND3_X1 U13987 ( .A1(n11029), .A2(n11028), .A3(n11027), .ZN(n11030) );
  NAND2_X1 U13988 ( .A1(n11535), .A2(n19903), .ZN(n11032) );
  NAND2_X1 U13989 ( .A1(n13620), .A2(n11035), .ZN(n11038) );
  NAND2_X1 U13990 ( .A1(n11036), .A2(n11039), .ZN(n11037) );
  NAND2_X1 U13991 ( .A1(n15531), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15532) );
  NAND2_X1 U13992 ( .A1(n11039), .A2(n11040), .ZN(n11042) );
  NAND2_X1 U13993 ( .A1(n11042), .A2(n11041), .ZN(n11043) );
  NAND2_X1 U13994 ( .A1(n15532), .A2(n11043), .ZN(n15274) );
  AOI22_X1 U13995 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10975), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U13996 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12661), .B1(
        n10857), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11046) );
  NAND2_X1 U13997 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11045) );
  NAND2_X1 U13998 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11044) );
  NAND2_X1 U13999 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11051) );
  NAND2_X1 U14000 ( .A1(n12570), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11050) );
  NAND2_X1 U14001 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11049) );
  NAND2_X1 U14002 ( .A1(n12668), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11048) );
  INV_X1 U14003 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11053) );
  INV_X1 U14004 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11052) );
  OAI22_X1 U14005 ( .A1(n11053), .A2(n12656), .B1(n11631), .B2(n11052), .ZN(
        n11054) );
  INV_X1 U14006 ( .A(n11054), .ZN(n11060) );
  NAND2_X1 U14007 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11058) );
  NAND2_X1 U14008 ( .A1(n10918), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11057) );
  NAND2_X1 U14009 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11056) );
  NAND2_X1 U14010 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11055) );
  NAND4_X1 U14011 ( .A1(n11062), .A2(n11061), .A3(n11060), .A4(n11059), .ZN(
        n11160) );
  NAND2_X1 U14012 ( .A1(n11063), .A2(n11539), .ZN(n11064) );
  XNOR2_X1 U14013 ( .A(n11065), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15273) );
  NAND2_X1 U14014 ( .A1(n15274), .A2(n15273), .ZN(n15275) );
  INV_X1 U14015 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15527) );
  NAND2_X1 U14016 ( .A1(n15275), .A2(n11066), .ZN(n16121) );
  NAND2_X1 U14017 ( .A1(n16121), .A2(n16120), .ZN(n16119) );
  INV_X1 U14018 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11488) );
  INV_X1 U14019 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15497) );
  INV_X1 U14020 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16109) );
  NOR2_X1 U14021 ( .A1(n15497), .A2(n16109), .ZN(n15496) );
  AND2_X1 U14022 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15496), .ZN(
        n16154) );
  AND2_X1 U14023 ( .A1(n16154), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11755) );
  INV_X1 U14024 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16089) );
  INV_X1 U14025 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16155) );
  NAND2_X1 U14026 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11757) );
  INV_X1 U14027 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15425) );
  INV_X1 U14028 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15404) );
  INV_X1 U14029 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n20968) );
  INV_X1 U14030 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15359) );
  INV_X1 U14031 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15332) );
  INV_X1 U14032 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11069) );
  INV_X1 U14033 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15284) );
  NAND2_X1 U14034 ( .A1(n15112), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11070) );
  NAND2_X1 U14035 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19883), .ZN(
        n11097) );
  OAI21_X1 U14036 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19883), .A(
        n11097), .ZN(n11399) );
  MUX2_X1 U14037 ( .A(n11494), .B(n11399), .S(n11084), .Z(n11117) );
  NAND2_X1 U14038 ( .A1(n19873), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11073) );
  NAND2_X1 U14039 ( .A1(n10795), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11072) );
  NAND2_X1 U14040 ( .A1(n11073), .A2(n11072), .ZN(n11398) );
  NAND2_X1 U14041 ( .A1(n11074), .A2(n11073), .ZN(n11077) );
  MUX2_X1 U14042 ( .A(n19864), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11076) );
  XNOR2_X1 U14043 ( .A(n11077), .B(n11076), .ZN(n11096) );
  INV_X1 U14044 ( .A(n11096), .ZN(n11396) );
  NAND2_X1 U14045 ( .A1(n11084), .A2(n11396), .ZN(n11394) );
  OAI21_X2 U14046 ( .B1(n11084), .B2(n11515), .A(n11394), .ZN(n11111) );
  INV_X1 U14047 ( .A(n11111), .ZN(n11075) );
  OAI21_X1 U14048 ( .B1(n11117), .B2(n11398), .A(n11075), .ZN(n11086) );
  NAND2_X1 U14049 ( .A1(n11077), .A2(n11076), .ZN(n11079) );
  NAND2_X1 U14050 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19864), .ZN(
        n11078) );
  XNOR2_X1 U14051 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11081) );
  XNOR2_X1 U14052 ( .A(n11082), .B(n11081), .ZN(n11093) );
  NOR2_X1 U14053 ( .A1(n10676), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11080) );
  AOI21_X1 U14054 ( .B1(n11082), .B2(n11081), .A(n11080), .ZN(n11088) );
  NOR2_X1 U14055 ( .A1(n16246), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11083) );
  NAND2_X1 U14056 ( .A1(n11088), .A2(n11083), .ZN(n11094) );
  MUX2_X1 U14057 ( .A(n11526), .B(n11094), .S(n11084), .Z(n11129) );
  NAND3_X1 U14058 ( .A1(n11086), .A2(n11085), .A3(n11129), .ZN(n11091) );
  NAND2_X1 U14059 ( .A1(n16246), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11087) );
  NAND2_X1 U14060 ( .A1(n11088), .A2(n11087), .ZN(n11090) );
  NAND2_X1 U14061 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16240), .ZN(
        n11089) );
  NAND2_X1 U14062 ( .A1(n11091), .A2(n11409), .ZN(n19887) );
  INV_X1 U14063 ( .A(n11092), .ZN(n16232) );
  AND2_X1 U14064 ( .A1(n19903), .A2(n16231), .ZN(n11441) );
  NAND2_X1 U14065 ( .A1(n16232), .A2(n11441), .ZN(n19885) );
  INV_X1 U14066 ( .A(n11093), .ZN(n11095) );
  NAND2_X1 U14067 ( .A1(n11095), .A2(n11094), .ZN(n11410) );
  NOR2_X1 U14068 ( .A1(n11096), .A2(n11410), .ZN(n11099) );
  INV_X1 U14069 ( .A(n11099), .ZN(n11101) );
  INV_X1 U14070 ( .A(n11097), .ZN(n11098) );
  XNOR2_X1 U14071 ( .A(n11398), .B(n11098), .ZN(n11400) );
  NAND2_X1 U14072 ( .A1(n11400), .A2(n11099), .ZN(n11100) );
  OAI21_X1 U14073 ( .B1(n11399), .B2(n11101), .A(n16226), .ZN(n11105) );
  NAND2_X1 U14074 ( .A1(n9799), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11102) );
  NAND2_X1 U14075 ( .A1(n11102), .A2(n16240), .ZN(n16233) );
  OR2_X1 U14076 ( .A1(n10918), .A2(n16233), .ZN(n11103) );
  INV_X1 U14077 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n15736) );
  NAND2_X1 U14078 ( .A1(n11103), .A2(n15736), .ZN(n19875) );
  INV_X1 U14079 ( .A(n19875), .ZN(n11104) );
  MUX2_X1 U14080 ( .A(n11105), .B(n11104), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n15734) );
  NAND2_X1 U14081 ( .A1(n16232), .A2(n15614), .ZN(n11106) );
  NAND2_X1 U14082 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n11393), .ZN(n19761) );
  INV_X1 U14083 ( .A(n19761), .ZN(n11107) );
  NAND2_X1 U14084 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11107), .ZN(n19134) );
  AND2_X1 U14085 ( .A1(n16231), .A2(n13032), .ZN(n11108) );
  NAND2_X1 U14086 ( .A1(n11463), .A2(n11108), .ZN(n12980) );
  INV_X1 U14087 ( .A(n12980), .ZN(n11292) );
  NAND2_X1 U14088 ( .A1(n11292), .A2(n19903), .ZN(n16145) );
  NAND2_X1 U14089 ( .A1(n9830), .A2(n19241), .ZN(n11431) );
  INV_X1 U14090 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13073) );
  MUX2_X2 U14091 ( .A(n13073), .B(n11111), .S(n11236), .Z(n11122) );
  NOR2_X1 U14092 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11112) );
  MUX2_X1 U14093 ( .A(n11112), .B(n11505), .S(n11236), .Z(n11121) );
  NAND2_X1 U14094 ( .A1(n11122), .A2(n11121), .ZN(n11113) );
  INV_X1 U14095 ( .A(n11133), .ZN(n11116) );
  NAND2_X1 U14096 ( .A1(n11114), .A2(n11113), .ZN(n11115) );
  NAND2_X1 U14097 ( .A1(n11116), .A2(n11115), .ZN(n13426) );
  INV_X1 U14098 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13044) );
  MUX2_X1 U14099 ( .A(n11117), .B(n13044), .S(n12817), .Z(n19071) );
  INV_X1 U14100 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13015) );
  INV_X1 U14101 ( .A(n11121), .ZN(n11119) );
  NAND3_X1 U14102 ( .A1(n12817), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n11118) );
  NAND2_X1 U14103 ( .A1(n11119), .A2(n11118), .ZN(n19052) );
  NOR2_X1 U14104 ( .A1(n10342), .A2(n19052), .ZN(n11120) );
  NAND2_X1 U14105 ( .A1(n10342), .A2(n19052), .ZN(n13003) );
  OAI21_X1 U14106 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11120), .A(
        n13003), .ZN(n14342) );
  XNOR2_X1 U14107 ( .A(n11122), .B(n11121), .ZN(n13504) );
  XNOR2_X1 U14108 ( .A(n13504), .B(n9801), .ZN(n14341) );
  OR2_X1 U14109 ( .A1(n14342), .A2(n14341), .ZN(n14356) );
  INV_X1 U14110 ( .A(n13504), .ZN(n11123) );
  NAND2_X1 U14111 ( .A1(n11123), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11124) );
  NAND2_X1 U14112 ( .A1(n14356), .A2(n11124), .ZN(n13545) );
  INV_X1 U14113 ( .A(n13545), .ZN(n11125) );
  NAND2_X1 U14114 ( .A1(n13543), .A2(n11125), .ZN(n11127) );
  NAND2_X1 U14115 ( .A1(n11127), .A2(n13544), .ZN(n13592) );
  INV_X1 U14116 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11128) );
  MUX2_X1 U14117 ( .A(n11129), .B(n11128), .S(n12817), .Z(n11132) );
  INV_X1 U14118 ( .A(n11132), .ZN(n11130) );
  XNOR2_X1 U14119 ( .A(n11133), .B(n11130), .ZN(n19031) );
  XNOR2_X1 U14120 ( .A(n19031), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13591) );
  NAND2_X1 U14121 ( .A1(n19031), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11131) );
  INV_X1 U14122 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n21112) );
  INV_X1 U14123 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11630) );
  INV_X1 U14124 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12612) );
  OAI22_X1 U14125 ( .A1(n12653), .A2(n11630), .B1(n12654), .B2(n12612), .ZN(
        n11136) );
  INV_X1 U14126 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11626) );
  INV_X1 U14127 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11134) );
  OAI22_X1 U14128 ( .A1(n15588), .A2(n11626), .B1(n12656), .B2(n11134), .ZN(
        n11135) );
  NOR2_X1 U14129 ( .A1(n11136), .A2(n11135), .ZN(n11140) );
  AOI22_X1 U14130 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U14131 ( .A1(n12661), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11138) );
  AOI22_X1 U14132 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10902), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11137) );
  NAND4_X1 U14133 ( .A1(n11140), .A2(n11139), .A3(n11138), .A4(n11137), .ZN(
        n11146) );
  AOI22_X1 U14134 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11144) );
  AOI22_X1 U14135 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11143) );
  NAND2_X1 U14136 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11142) );
  NAND2_X1 U14137 ( .A1(n12668), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11141) );
  NAND4_X1 U14138 ( .A1(n11144), .A2(n11143), .A3(n11142), .A4(n11141), .ZN(
        n11145) );
  MUX2_X1 U14139 ( .A(n21112), .B(n11532), .S(n11236), .Z(n11147) );
  OAI21_X1 U14140 ( .B1(n11148), .B2(n11147), .A(n11154), .ZN(n19020) );
  XNOR2_X1 U14141 ( .A(n11150), .B(n13624), .ZN(n13616) );
  NAND2_X1 U14142 ( .A1(n13615), .A2(n13616), .ZN(n11152) );
  NAND2_X1 U14143 ( .A1(n11150), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11151) );
  NAND2_X1 U14144 ( .A1(n11152), .A2(n11151), .ZN(n15544) );
  MUX2_X1 U14145 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n11535), .S(n11236), .Z(
        n11153) );
  AND2_X1 U14146 ( .A1(n11154), .A2(n11153), .ZN(n11155) );
  OR2_X1 U14147 ( .A1(n11155), .A2(n11166), .ZN(n19009) );
  INV_X1 U14148 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15540) );
  XNOR2_X1 U14149 ( .A(n11157), .B(n15540), .ZN(n15545) );
  NAND2_X1 U14150 ( .A1(n15544), .A2(n15545), .ZN(n11159) );
  NAND2_X1 U14151 ( .A1(n11157), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11158) );
  INV_X1 U14152 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13144) );
  MUX2_X1 U14153 ( .A(n13144), .B(n11160), .S(n11236), .Z(n11164) );
  OR2_X1 U14154 ( .A1(n11162), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11161) );
  NAND2_X2 U14155 ( .A1(n11257), .A2(n11161), .ZN(n11172) );
  AND3_X1 U14156 ( .A1(n11162), .A2(P2_EBX_REG_8__SCAN_IN), .A3(n12817), .ZN(
        n11163) );
  OR2_X1 U14157 ( .A1(n11172), .A2(n11163), .ZN(n18987) );
  NOR2_X1 U14158 ( .A1(n18987), .A2(n11539), .ZN(n11167) );
  AND2_X1 U14159 ( .A1(n11167), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16126) );
  INV_X1 U14160 ( .A(n11164), .ZN(n11165) );
  XNOR2_X1 U14161 ( .A(n11166), .B(n11165), .ZN(n19000) );
  AND2_X1 U14162 ( .A1(n19000), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16123) );
  INV_X1 U14163 ( .A(n11167), .ZN(n11168) );
  NAND2_X1 U14164 ( .A1(n11168), .A2(n11488), .ZN(n16125) );
  INV_X1 U14165 ( .A(n19000), .ZN(n11169) );
  NAND2_X1 U14166 ( .A1(n11169), .A2(n15527), .ZN(n16124) );
  AND2_X1 U14167 ( .A1(n16125), .A2(n16124), .ZN(n11170) );
  AND2_X1 U14168 ( .A1(n12817), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11171) );
  XNOR2_X1 U14169 ( .A(n11172), .B(n11171), .ZN(n18975) );
  AOI21_X1 U14170 ( .B1(n18975), .B2(n11289), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15259) );
  NAND2_X1 U14171 ( .A1(n12817), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11173) );
  INV_X1 U14172 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n20978) );
  MUX2_X1 U14173 ( .A(n11173), .B(P2_EBX_REG_10__SCAN_IN), .S(n11179), .Z(
        n11174) );
  NAND2_X1 U14174 ( .A1(n11174), .A2(n11257), .ZN(n11175) );
  OAI21_X1 U14175 ( .B1(n11175), .B2(n11539), .A(n16109), .ZN(n16113) );
  INV_X1 U14176 ( .A(n11175), .ZN(n18968) );
  AND2_X1 U14177 ( .A1(n11289), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11176) );
  NAND2_X1 U14178 ( .A1(n18968), .A2(n11176), .ZN(n16112) );
  AND2_X1 U14179 ( .A1(n11289), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11177) );
  NAND2_X1 U14180 ( .A1(n18975), .A2(n11177), .ZN(n15258) );
  AND2_X1 U14181 ( .A1(n16112), .A2(n15258), .ZN(n11178) );
  INV_X1 U14182 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13315) );
  NAND2_X1 U14183 ( .A1(n12817), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11180) );
  OR2_X1 U14184 ( .A1(n11181), .A2(n11180), .ZN(n11183) );
  INV_X1 U14185 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n18954) );
  INV_X1 U14186 ( .A(n11186), .ZN(n11182) );
  NAND2_X1 U14187 ( .A1(n11183), .A2(n11182), .ZN(n18955) );
  NOR2_X1 U14188 ( .A1(n18955), .A2(n11539), .ZN(n11184) );
  AND2_X1 U14189 ( .A1(n11184), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15493) );
  INV_X1 U14190 ( .A(n11184), .ZN(n11185) );
  NAND2_X1 U14191 ( .A1(n12817), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11187) );
  NAND2_X1 U14192 ( .A1(n10003), .A2(n11188), .ZN(n11189) );
  NAND2_X1 U14193 ( .A1(n11214), .A2(n11189), .ZN(n18947) );
  XNOR2_X1 U14194 ( .A(n11190), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15476) );
  INV_X1 U14195 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11193) );
  NOR2_X1 U14196 ( .A1(n11236), .A2(n11193), .ZN(n11213) );
  INV_X1 U14197 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11194) );
  INV_X1 U14198 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11195) );
  OR2_X2 U14199 ( .A1(n11205), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11206) );
  NAND2_X1 U14200 ( .A1(n12817), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11208) );
  AND2_X1 U14201 ( .A1(n12817), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11200) );
  AND2_X1 U14202 ( .A1(n12817), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11197) );
  INV_X1 U14203 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n15007) );
  NAND3_X1 U14204 ( .A1(n11237), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n12817), 
        .ZN(n11196) );
  OAI211_X1 U14205 ( .C1(n11237), .C2(P2_EBX_REG_21__SCAN_IN), .A(n11196), .B(
        n11257), .ZN(n12921) );
  OAI21_X1 U14206 ( .B1(n12921), .B2(n11539), .A(n20968), .ZN(n15185) );
  AND2_X1 U14207 ( .A1(n11202), .A2(n11197), .ZN(n11198) );
  NOR2_X1 U14208 ( .A1(n11218), .A2(n11198), .ZN(n18872) );
  NAND2_X1 U14209 ( .A1(n18872), .A2(n11289), .ZN(n11228) );
  NAND2_X1 U14210 ( .A1(n11228), .A2(n15404), .ZN(n15208) );
  NAND2_X1 U14211 ( .A1(n11199), .A2(n11200), .ZN(n11201) );
  NAND2_X1 U14212 ( .A1(n11202), .A2(n11201), .ZN(n11230) );
  OAI21_X1 U14213 ( .B1(n11230), .B2(n11539), .A(n15425), .ZN(n15221) );
  AND2_X2 U14214 ( .A1(n15208), .A2(n15221), .ZN(n15197) );
  AND2_X1 U14215 ( .A1(n12817), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11204) );
  INV_X1 U14216 ( .A(n11257), .ZN(n11203) );
  AOI21_X1 U14217 ( .B1(n11205), .B2(n11204), .A(n11203), .ZN(n11207) );
  AND2_X1 U14218 ( .A1(n11207), .A2(n11206), .ZN(n18905) );
  NAND2_X1 U14219 ( .A1(n18905), .A2(n11289), .ZN(n11222) );
  XNOR2_X1 U14220 ( .A(n11222), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15240) );
  OR2_X1 U14221 ( .A1(n11209), .A2(n11208), .ZN(n11210) );
  NAND2_X1 U14222 ( .A1(n11210), .A2(n11199), .ZN(n18896) );
  NOR2_X1 U14223 ( .A1(n18896), .A2(n11539), .ZN(n11220) );
  NOR2_X1 U14224 ( .A1(n11220), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15180) );
  AND2_X1 U14225 ( .A1(n12817), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11211) );
  XNOR2_X1 U14226 ( .A(n11212), .B(n11211), .ZN(n18914) );
  AOI21_X1 U14227 ( .B1(n18914), .B2(n11289), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15249) );
  XNOR2_X1 U14228 ( .A(n11216), .B(n9919), .ZN(n18924) );
  AOI21_X1 U14229 ( .B1(n18924), .B2(n11289), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15177) );
  NAND2_X1 U14230 ( .A1(n11214), .A2(n11213), .ZN(n11215) );
  AND2_X1 U14231 ( .A1(n11216), .A2(n11215), .ZN(n18935) );
  AOI21_X1 U14232 ( .B1(n18935), .B2(n11289), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16086) );
  NOR4_X1 U14233 ( .A1(n15180), .A2(n15249), .A3(n15177), .A4(n16086), .ZN(
        n11217) );
  NAND2_X1 U14234 ( .A1(n11289), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11219) );
  OR2_X1 U14235 ( .A1(n12921), .A2(n11219), .ZN(n15184) );
  INV_X1 U14236 ( .A(n11220), .ZN(n11221) );
  INV_X1 U14237 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11689) );
  NOR2_X1 U14238 ( .A1(n11221), .A2(n11689), .ZN(n15181) );
  INV_X1 U14239 ( .A(n11222), .ZN(n11223) );
  NAND2_X1 U14240 ( .A1(n11223), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15179) );
  AND2_X1 U14241 ( .A1(n11289), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11224) );
  NAND2_X1 U14242 ( .A1(n18914), .A2(n11224), .ZN(n15250) );
  AND2_X1 U14243 ( .A1(n11289), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11225) );
  NAND2_X1 U14244 ( .A1(n18924), .A2(n11225), .ZN(n16076) );
  AND2_X1 U14245 ( .A1(n11289), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11226) );
  NAND2_X1 U14246 ( .A1(n18935), .A2(n11226), .ZN(n16084) );
  NAND4_X1 U14247 ( .A1(n15179), .A2(n15250), .A3(n16076), .A4(n16084), .ZN(
        n11227) );
  NOR2_X1 U14248 ( .A1(n15181), .A2(n11227), .ZN(n11232) );
  INV_X1 U14249 ( .A(n11228), .ZN(n11229) );
  NAND2_X1 U14250 ( .A1(n11229), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15209) );
  INV_X1 U14251 ( .A(n11230), .ZN(n18881) );
  AND2_X1 U14252 ( .A1(n11289), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11231) );
  NAND2_X1 U14253 ( .A1(n18881), .A2(n11231), .ZN(n15220) );
  NAND4_X1 U14254 ( .A1(n15184), .A2(n11232), .A3(n15209), .A4(n15220), .ZN(
        n11234) );
  AND2_X1 U14255 ( .A1(n11289), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11233) );
  INV_X1 U14256 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11235) );
  NOR2_X1 U14257 ( .A1(n11236), .A2(n11235), .ZN(n11241) );
  INV_X1 U14258 ( .A(n11238), .ZN(n11240) );
  AOI21_X1 U14259 ( .B1(n11241), .B2(n11240), .A(n11245), .ZN(n15682) );
  AOI21_X1 U14260 ( .B1(n15682), .B2(n11289), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15169) );
  NAND3_X1 U14261 ( .A1(n15682), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n11289), .ZN(n15170) );
  NAND2_X1 U14262 ( .A1(n12817), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11244) );
  INV_X1 U14263 ( .A(n11244), .ZN(n11242) );
  NAND2_X1 U14264 ( .A1(n11243), .A2(n11242), .ZN(n11246) );
  NAND2_X1 U14265 ( .A1(n11246), .A2(n11254), .ZN(n12934) );
  OR2_X1 U14266 ( .A1(n12934), .A2(n11539), .ZN(n11247) );
  NAND2_X1 U14267 ( .A1(n15157), .A2(n15158), .ZN(n11248) );
  INV_X1 U14268 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15342) );
  NAND2_X1 U14269 ( .A1(n12817), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11249) );
  MUX2_X1 U14270 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n11249), .S(n11254), .Z(
        n11250) );
  NAND2_X1 U14271 ( .A1(n11250), .A2(n11257), .ZN(n16047) );
  NOR2_X1 U14272 ( .A1(n16047), .A2(n11539), .ZN(n15149) );
  INV_X1 U14273 ( .A(n15149), .ZN(n11251) );
  NAND2_X1 U14274 ( .A1(n12817), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11255) );
  MUX2_X1 U14275 ( .A(P2_EBX_REG_25__SCAN_IN), .B(n11255), .S(n9870), .Z(
        n11256) );
  NAND2_X1 U14276 ( .A1(n11256), .A2(n11257), .ZN(n16038) );
  NOR2_X1 U14277 ( .A1(n11273), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15138) );
  AND2_X1 U14278 ( .A1(n12817), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11258) );
  AOI21_X1 U14279 ( .B1(n11259), .B2(n11258), .A(n11285), .ZN(n16028) );
  INV_X1 U14280 ( .A(n16028), .ZN(n11260) );
  NOR2_X1 U14281 ( .A1(n11260), .A2(n11539), .ZN(n11261) );
  NAND3_X1 U14282 ( .A1(n16028), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n11289), .ZN(n11274) );
  OAI21_X1 U14283 ( .B1(n11261), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11274), .ZN(n15131) );
  NAND2_X1 U14284 ( .A1(n12817), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11262) );
  INV_X1 U14285 ( .A(n11262), .ZN(n11263) );
  NAND2_X1 U14286 ( .A1(n11263), .A2(n9855), .ZN(n11264) );
  NAND2_X1 U14287 ( .A1(n11267), .A2(n11264), .ZN(n12946) );
  INV_X1 U14288 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11265) );
  NOR2_X1 U14289 ( .A1(n11236), .A2(n11265), .ZN(n11266) );
  NAND2_X1 U14290 ( .A1(n11267), .A2(n11266), .ZN(n11268) );
  NAND2_X1 U14291 ( .A1(n11276), .A2(n11268), .ZN(n12962) );
  OAI21_X1 U14292 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n12439), .ZN(n11269) );
  NAND2_X1 U14293 ( .A1(n11270), .A2(n11269), .ZN(n11272) );
  INV_X1 U14294 ( .A(n12439), .ZN(n11271) );
  INV_X1 U14295 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15297) );
  NAND2_X1 U14296 ( .A1(n11273), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15139) );
  NAND2_X1 U14297 ( .A1(n15139), .A2(n11274), .ZN(n12434) );
  INV_X1 U14298 ( .A(n12434), .ZN(n11275) );
  NAND2_X1 U14299 ( .A1(n12817), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11277) );
  XNOR2_X1 U14300 ( .A(n11278), .B(n11277), .ZN(n11281) );
  OAI21_X1 U14301 ( .B1(n11281), .B2(n11539), .A(n15284), .ZN(n15105) );
  NAND2_X1 U14302 ( .A1(n12817), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11279) );
  AOI21_X1 U14303 ( .B1(n11280), .B2(n11289), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11774) );
  INV_X1 U14304 ( .A(n11280), .ZN(n12896) );
  INV_X1 U14305 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11386) );
  INV_X1 U14306 ( .A(n11281), .ZN(n16017) );
  NAND3_X1 U14307 ( .A1(n16017), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11289), .ZN(n15106) );
  NOR2_X1 U14308 ( .A1(n11283), .A2(n11282), .ZN(n11284) );
  INV_X1 U14309 ( .A(n11285), .ZN(n11288) );
  NOR2_X1 U14310 ( .A1(n11286), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11287) );
  MUX2_X1 U14311 ( .A(n11288), .B(n11287), .S(n12817), .Z(n16005) );
  NAND2_X1 U14312 ( .A1(n16005), .A2(n11289), .ZN(n11290) );
  XOR2_X1 U14313 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11290), .Z(
        n11291) );
  NAND2_X1 U14314 ( .A1(n11294), .A2(n11293), .ZN(n11299) );
  INV_X1 U14315 ( .A(n11295), .ZN(n11296) );
  OR2_X1 U14316 ( .A1(n11297), .A2(n11296), .ZN(n11298) );
  NAND2_X1 U14317 ( .A1(n11299), .A2(n11298), .ZN(n13159) );
  INV_X1 U14318 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U14319 ( .A1(n11387), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11302) );
  NAND2_X1 U14320 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11301) );
  OAI211_X1 U14321 ( .C1(n11303), .C2(n11380), .A(n11302), .B(n11301), .ZN(
        n11304) );
  AOI21_X1 U14322 ( .B1(n10820), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11304), .ZN(n13158) );
  INV_X1 U14323 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11308) );
  NAND2_X1 U14324 ( .A1(n11387), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11307) );
  NAND2_X1 U14325 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11306) );
  OAI211_X1 U14326 ( .C1(n11308), .C2(n11380), .A(n11307), .B(n11306), .ZN(
        n11309) );
  AOI21_X1 U14327 ( .B1(n10820), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11309), .ZN(n13076) );
  INV_X1 U14328 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n11312) );
  NAND2_X1 U14329 ( .A1(n11387), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11311) );
  NAND2_X1 U14330 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11310) );
  OAI211_X1 U14331 ( .C1(n11312), .C2(n11380), .A(n11311), .B(n11310), .ZN(
        n11313) );
  AOI21_X1 U14332 ( .B1(n10820), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11313), .ZN(n13128) );
  AOI22_X1 U14333 ( .A1(n11387), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11316) );
  NAND2_X1 U14334 ( .A1(n11314), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11315) );
  OAI211_X1 U14335 ( .C1(n11390), .C2(n15527), .A(n11316), .B(n11315), .ZN(
        n13141) );
  NAND2_X1 U14336 ( .A1(n13142), .A2(n13141), .ZN(n13200) );
  INV_X1 U14337 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n11491) );
  NAND2_X1 U14338 ( .A1(n11387), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11318) );
  NAND2_X1 U14339 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11317) );
  OAI211_X1 U14340 ( .C1(n11491), .C2(n11380), .A(n11318), .B(n11317), .ZN(
        n11319) );
  AOI21_X1 U14341 ( .B1(n10820), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11319), .ZN(n13199) );
  INV_X1 U14342 ( .A(n11390), .ZN(n11326) );
  INV_X1 U14343 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U14344 ( .A1(n11387), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11323) );
  NAND2_X1 U14345 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11322) );
  OAI211_X1 U14346 ( .C1(n11324), .C2(n11380), .A(n11323), .B(n11322), .ZN(
        n11325) );
  AOI21_X1 U14347 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11325), .ZN(n13286) );
  AOI22_X1 U14348 ( .A1(n11387), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11328) );
  NAND2_X1 U14349 ( .A1(n11314), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11327) );
  OAI211_X1 U14350 ( .C1(n11390), .C2(n16109), .A(n11328), .B(n11327), .ZN(
        n13313) );
  AOI22_X1 U14351 ( .A1(n11387), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11330) );
  NAND2_X1 U14352 ( .A1(n11314), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11329) );
  OAI211_X1 U14353 ( .C1(n11390), .C2(n15497), .A(n11330), .B(n11329), .ZN(
        n13414) );
  INV_X1 U14354 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11333) );
  NAND2_X1 U14355 ( .A1(n11387), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U14356 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11331) );
  OAI211_X1 U14357 ( .C1(n11333), .C2(n11380), .A(n11332), .B(n11331), .ZN(
        n11334) );
  AOI21_X1 U14358 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11334), .ZN(n13468) );
  INV_X1 U14359 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11337) );
  NAND2_X1 U14360 ( .A1(n11387), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11336) );
  NAND2_X1 U14361 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11335) );
  OAI211_X1 U14362 ( .C1(n11337), .C2(n11380), .A(n11336), .B(n11335), .ZN(
        n11338) );
  AOI21_X1 U14363 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11338), .ZN(n13474) );
  INV_X1 U14364 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11341) );
  NAND2_X1 U14365 ( .A1(n11387), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11340) );
  NAND2_X1 U14366 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11339) );
  OAI211_X1 U14367 ( .C1(n11341), .C2(n11380), .A(n11340), .B(n11339), .ZN(
        n11342) );
  AOI21_X1 U14368 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11342), .ZN(n13586) );
  INV_X1 U14369 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15466) );
  AOI22_X1 U14370 ( .A1(n11387), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11344) );
  NAND2_X1 U14371 ( .A1(n11314), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11343) );
  OAI211_X1 U14372 ( .C1(n11390), .C2(n15466), .A(n11344), .B(n11343), .ZN(
        n13605) );
  INV_X1 U14373 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15451) );
  NAND2_X1 U14374 ( .A1(n11387), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11346) );
  NAND2_X1 U14375 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11345) );
  OAI211_X1 U14376 ( .C1(n15451), .C2(n11380), .A(n11346), .B(n11345), .ZN(
        n11347) );
  AOI21_X1 U14377 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11347), .ZN(n15033) );
  INV_X1 U14378 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19808) );
  NAND2_X1 U14379 ( .A1(n11387), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11349) );
  NAND2_X1 U14380 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11348) );
  OAI211_X1 U14381 ( .C1(n19808), .C2(n11380), .A(n11349), .B(n11348), .ZN(
        n11350) );
  AOI21_X1 U14382 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11350), .ZN(n15024) );
  AOI22_X1 U14383 ( .A1(n11387), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11352) );
  NAND2_X1 U14384 ( .A1(n11314), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11351) );
  OAI211_X1 U14385 ( .C1(n11390), .C2(n15425), .A(n11352), .B(n11351), .ZN(
        n15015) );
  AOI22_X1 U14386 ( .A1(n11387), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11354) );
  NAND2_X1 U14387 ( .A1(n11314), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11353) );
  OAI211_X1 U14388 ( .C1(n11390), .C2(n15404), .A(n11354), .B(n11353), .ZN(
        n15008) );
  NAND2_X1 U14389 ( .A1(n15017), .A2(n15008), .ZN(n14998) );
  INV_X1 U14390 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15201) );
  NAND2_X1 U14391 ( .A1(n11387), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11356) );
  NAND2_X1 U14392 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11355) );
  OAI211_X1 U14393 ( .C1(n15201), .C2(n11380), .A(n11356), .B(n11355), .ZN(
        n11357) );
  AOI21_X1 U14394 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11357), .ZN(n15001) );
  INV_X1 U14395 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19814) );
  NAND2_X1 U14396 ( .A1(n11387), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11359) );
  NAND2_X1 U14397 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11358) );
  OAI211_X1 U14398 ( .C1(n19814), .C2(n11380), .A(n11359), .B(n11358), .ZN(
        n11360) );
  AOI21_X1 U14399 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11360), .ZN(n12922) );
  INV_X1 U14400 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15372) );
  AOI22_X1 U14401 ( .A1(n11387), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11362) );
  NAND2_X1 U14402 ( .A1(n11314), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11361) );
  OAI211_X1 U14403 ( .C1(n11390), .C2(n15372), .A(n11362), .B(n11361), .ZN(
        n14989) );
  INV_X1 U14404 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19818) );
  NAND2_X1 U14405 ( .A1(n11387), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11364) );
  NAND2_X1 U14406 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11363) );
  OAI211_X1 U14407 ( .C1(n19818), .C2(n11380), .A(n11364), .B(n11363), .ZN(
        n11365) );
  AOI21_X1 U14408 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11365), .ZN(n12935) );
  INV_X1 U14409 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19820) );
  NAND2_X1 U14410 ( .A1(n11387), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11367) );
  NAND2_X1 U14411 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11366) );
  OAI211_X1 U14412 ( .C1(n19820), .C2(n11380), .A(n11367), .B(n11366), .ZN(
        n11368) );
  AOI21_X1 U14413 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11368), .ZN(n14978) );
  INV_X1 U14414 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19822) );
  NAND2_X1 U14415 ( .A1(n11387), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11370) );
  NAND2_X1 U14416 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11369) );
  OAI211_X1 U14417 ( .C1(n19822), .C2(n11380), .A(n11370), .B(n11369), .ZN(
        n11371) );
  AOI21_X1 U14418 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11371), .ZN(n14965) );
  INV_X1 U14419 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14420 ( .A1(n11387), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11373) );
  NAND2_X1 U14421 ( .A1(n11314), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11372) );
  OAI211_X1 U14422 ( .C1(n11390), .C2(n11374), .A(n11373), .B(n11372), .ZN(
        n14955) );
  NAND2_X1 U14423 ( .A1(n14966), .A2(n14955), .ZN(n12948) );
  INV_X1 U14424 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19827) );
  NAND2_X1 U14425 ( .A1(n11387), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11376) );
  NAND2_X1 U14426 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11375) );
  OAI211_X1 U14427 ( .C1(n19827), .C2(n11380), .A(n11376), .B(n11375), .ZN(
        n11377) );
  AOI21_X1 U14428 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11377), .ZN(n12949) );
  INV_X1 U14429 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19828) );
  NAND2_X1 U14430 ( .A1(n11387), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11379) );
  NAND2_X1 U14431 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11378) );
  OAI211_X1 U14432 ( .C1(n19828), .C2(n11380), .A(n11379), .B(n11378), .ZN(
        n11381) );
  AOI21_X1 U14433 ( .B1(n11326), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11381), .ZN(n12442) );
  AOI22_X1 U14434 ( .A1(n11387), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11383) );
  NAND2_X1 U14435 ( .A1(n11314), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11382) );
  OAI211_X1 U14436 ( .C1(n11390), .C2(n15284), .A(n11383), .B(n11382), .ZN(
        n12834) );
  AOI22_X1 U14437 ( .A1(n11387), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11385) );
  NAND2_X1 U14438 ( .A1(n11314), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11384) );
  OAI211_X1 U14439 ( .C1(n11390), .C2(n11386), .A(n11385), .B(n11384), .ZN(
        n11432) );
  INV_X1 U14440 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12849) );
  AOI22_X1 U14441 ( .A1(n11387), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11389) );
  NAND2_X1 U14442 ( .A1(n11314), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11388) );
  OAI211_X1 U14443 ( .C1(n11390), .C2(n12849), .A(n11389), .B(n11388), .ZN(
        n11391) );
  INV_X1 U14444 ( .A(n11391), .ZN(n11392) );
  INV_X1 U14445 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n11393) );
  NAND2_X1 U14446 ( .A1(n19654), .A2(n11393), .ZN(n19900) );
  INV_X1 U14447 ( .A(n11394), .ZN(n11408) );
  NAND2_X1 U14448 ( .A1(n16231), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19142) );
  AOI21_X1 U14449 ( .B1(n19142), .B2(n15614), .A(n11396), .ZN(n11407) );
  NAND2_X1 U14450 ( .A1(n11395), .A2(n11396), .ZN(n11404) );
  OAI21_X1 U14451 ( .B1(n11399), .B2(n11398), .A(n11397), .ZN(n11403) );
  INV_X1 U14452 ( .A(n11399), .ZN(n11401) );
  OAI211_X1 U14453 ( .C1(n15614), .C2(n11401), .A(n11443), .B(n11400), .ZN(
        n11402) );
  NAND3_X1 U14454 ( .A1(n11404), .A2(n11403), .A3(n11402), .ZN(n11406) );
  INV_X1 U14455 ( .A(n11410), .ZN(n11405) );
  OAI211_X1 U14456 ( .C1(n11408), .C2(n11407), .A(n11406), .B(n11405), .ZN(
        n11412) );
  AOI21_X1 U14457 ( .B1(n11397), .B2(n11410), .A(n11415), .ZN(n11411) );
  NAND2_X1 U14458 ( .A1(n11412), .A2(n11411), .ZN(n11413) );
  MUX2_X1 U14459 ( .A(n11413), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19904), .Z(n11435) );
  INV_X1 U14460 ( .A(n19142), .ZN(n11414) );
  NAND2_X1 U14461 ( .A1(n11415), .A2(n11414), .ZN(n11416) );
  NAND2_X1 U14462 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19140) );
  NAND2_X1 U14463 ( .A1(n11393), .A2(n19469), .ZN(n15592) );
  NAND2_X1 U14464 ( .A1(n15596), .A2(n15592), .ZN(n19874) );
  NAND2_X1 U14465 ( .A1(n19874), .A2(n19904), .ZN(n11417) );
  NAND2_X1 U14466 ( .A1(n19904), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12504) );
  NAND2_X1 U14467 ( .A1(n19902), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11418) );
  NAND2_X1 U14468 ( .A1(n12504), .A2(n11418), .ZN(n13018) );
  NAND2_X1 U14469 ( .A1(n12859), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12856) );
  INV_X1 U14470 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16106) );
  INV_X1 U14471 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15234) );
  INV_X1 U14472 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15214) );
  AND2_X1 U14473 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12869) );
  AND2_X1 U14474 ( .A1(n12869), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11421) );
  INV_X1 U14475 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15145) );
  INV_X1 U14476 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15122) );
  INV_X1 U14477 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12878) );
  OR2_X1 U14478 ( .A1(n15122), .A2(n12878), .ZN(n11422) );
  AND2_X1 U14479 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11423) );
  NAND2_X1 U14480 ( .A1(n12840), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11425) );
  INV_X1 U14481 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11424) );
  NOR2_X1 U14482 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n15592), .ZN(n12972) );
  AND2_X1 U14483 ( .A1(n12972), .A2(n19904), .ZN(n16202) );
  NAND2_X1 U14484 ( .A1(n19236), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11790) );
  NAND2_X1 U14485 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11426) );
  OAI211_X1 U14486 ( .C1(n19247), .C2(n12850), .A(n11790), .B(n11426), .ZN(
        n11427) );
  INV_X1 U14487 ( .A(n11427), .ZN(n11428) );
  NAND2_X1 U14488 ( .A1(n10353), .A2(n11428), .ZN(n11429) );
  AOI21_X1 U14489 ( .B1(n11782), .B2(n19242), .A(n11429), .ZN(n11430) );
  NAND2_X1 U14490 ( .A1(n11431), .A2(n11430), .ZN(P2_U2983) );
  NAND2_X1 U14491 ( .A1(n12826), .A2(n15614), .ZN(n19138) );
  INV_X1 U14492 ( .A(n19138), .ZN(n11434) );
  NOR2_X1 U14493 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19778) );
  AOI211_X1 U14494 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19778), .ZN(n19906) );
  NAND2_X1 U14495 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19901) );
  NAND2_X1 U14496 ( .A1(n19906), .A2(n19901), .ZN(n12886) );
  INV_X1 U14497 ( .A(n12886), .ZN(n12978) );
  NAND2_X1 U14498 ( .A1(n11434), .A2(n12978), .ZN(n13030) );
  AOI21_X1 U14499 ( .B1(n11435), .B2(n11443), .A(n13457), .ZN(n11436) );
  NAND2_X1 U14500 ( .A1(n19138), .A2(n11436), .ZN(n11460) );
  OAI21_X1 U14501 ( .B1(n12804), .B2(n13457), .A(n13572), .ZN(n11439) );
  NAND2_X1 U14502 ( .A1(n19135), .A2(n11439), .ZN(n11450) );
  NAND2_X1 U14503 ( .A1(n11442), .A2(n11441), .ZN(n11729) );
  INV_X1 U14504 ( .A(n11734), .ZN(n11447) );
  NAND2_X1 U14505 ( .A1(n19903), .A2(n11732), .ZN(n11725) );
  NAND2_X1 U14506 ( .A1(n11725), .A2(n11443), .ZN(n11444) );
  NAND2_X1 U14507 ( .A1(n11445), .A2(n13572), .ZN(n11446) );
  INV_X1 U14508 ( .A(n16226), .ZN(n11452) );
  NOR2_X1 U14509 ( .A1(n12886), .A2(n11452), .ZN(n11453) );
  NAND2_X1 U14510 ( .A1(n11451), .A2(n11453), .ZN(n11454) );
  NAND2_X1 U14511 ( .A1(n11727), .A2(n11454), .ZN(n13023) );
  MUX2_X1 U14512 ( .A(n11455), .B(n13572), .S(n19903), .Z(n11457) );
  NAND2_X1 U14513 ( .A1(n16226), .A2(n19901), .ZN(n11456) );
  NOR2_X1 U14514 ( .A1(n11457), .A2(n11456), .ZN(n11458) );
  NOR2_X1 U14515 ( .A1(n13023), .A2(n11458), .ZN(n11459) );
  AND2_X1 U14516 ( .A1(n11460), .A2(n11459), .ZN(n11461) );
  OAI21_X1 U14517 ( .B1(n13030), .B2(n13572), .A(n11461), .ZN(n11462) );
  OAI21_X2 U14518 ( .B1(n11463), .B2(n11462), .A(n13032), .ZN(n11779) );
  NAND2_X1 U14519 ( .A1(n11464), .A2(n19903), .ZN(n11465) );
  AND2_X1 U14520 ( .A1(n10786), .A2(n11465), .ZN(n11466) );
  NOR2_X1 U14521 ( .A1(n12817), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11468) );
  INV_X1 U14522 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11469) );
  INV_X1 U14523 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n19543) );
  OAI22_X1 U14524 ( .A1(n12653), .A2(n11469), .B1(n12654), .B2(n19543), .ZN(
        n11472) );
  OAI22_X1 U14525 ( .A1(n11631), .A2(n11470), .B1(n15588), .B2(n21017), .ZN(
        n11471) );
  NOR2_X1 U14526 ( .A1(n11472), .A2(n11471), .ZN(n11486) );
  INV_X1 U14527 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15612) );
  INV_X1 U14528 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11473) );
  OAI22_X1 U14529 ( .A1(n11629), .A2(n15612), .B1(n12656), .B2(n11473), .ZN(
        n11479) );
  NAND2_X1 U14530 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11477) );
  NAND2_X1 U14531 ( .A1(n10918), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11476) );
  NAND2_X1 U14532 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11475) );
  NAND2_X1 U14533 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11474) );
  NAND4_X1 U14534 ( .A1(n11477), .A2(n11476), .A3(n11475), .A4(n11474), .ZN(
        n11478) );
  NOR2_X1 U14535 ( .A1(n11479), .A2(n11478), .ZN(n11485) );
  AOI22_X1 U14536 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14537 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11482) );
  NAND2_X1 U14538 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11481) );
  NAND2_X1 U14539 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11480) );
  AND4_X1 U14540 ( .A1(n11483), .A2(n11482), .A3(n11481), .A4(n11480), .ZN(
        n11484) );
  NAND3_X1 U14541 ( .A1(n11486), .A2(n11485), .A3(n11484), .ZN(n13203) );
  INV_X1 U14542 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n11489) );
  AND2_X1 U14543 ( .A1(n15614), .A2(n19469), .ZN(n11528) );
  INV_X1 U14544 ( .A(n11713), .ZN(n11700) );
  OAI22_X1 U14545 ( .A1(n11701), .A2(n11489), .B1(n11700), .B2(n11488), .ZN(
        n11493) );
  AND3_X4 U14546 ( .A1(n11490), .A2(n19903), .A3(n12817), .ZN(n11784) );
  NOR2_X1 U14547 ( .A1(n11702), .A2(n11491), .ZN(n11492) );
  AOI211_X1 U14548 ( .C1(n11495), .C2(n13203), .A(n11493), .B(n11492), .ZN(
        n16191) );
  INV_X1 U14549 ( .A(n11494), .ZN(n11496) );
  NAND2_X1 U14550 ( .A1(n12804), .A2(n11528), .ZN(n11513) );
  AND2_X1 U14551 ( .A1(n11497), .A2(n11513), .ZN(n11498) );
  NAND2_X1 U14552 ( .A1(n11784), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11502) );
  INV_X1 U14553 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n11501) );
  NAND2_X1 U14554 ( .A1(n15614), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11500) );
  NAND2_X1 U14555 ( .A1(n11502), .A2(n9875), .ZN(n13038) );
  AOI22_X1 U14556 ( .A1(n11487), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11528), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11504) );
  NAND2_X1 U14557 ( .A1(n11784), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11503) );
  NAND2_X1 U14558 ( .A1(n11504), .A2(n11503), .ZN(n11510) );
  INV_X1 U14559 ( .A(n11505), .ZN(n11508) );
  MUX2_X1 U14560 ( .A(n11506), .B(n19873), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11507) );
  OAI21_X1 U14561 ( .B1(n11508), .B2(n11681), .A(n11507), .ZN(n13080) );
  NOR2_X1 U14562 ( .A1(n13081), .A2(n13080), .ZN(n11512) );
  NOR2_X1 U14563 ( .A1(n11509), .A2(n11510), .ZN(n11511) );
  NOR2_X2 U14564 ( .A1(n11512), .A2(n11511), .ZN(n11519) );
  NAND2_X1 U14565 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11514) );
  OAI211_X1 U14566 ( .C1(n11681), .C2(n11515), .A(n11514), .B(n11513), .ZN(
        n11518) );
  XNOR2_X1 U14567 ( .A(n11519), .B(n11518), .ZN(n13266) );
  INV_X2 U14568 ( .A(n11701), .ZN(n11716) );
  AOI22_X1 U14569 ( .A1(n11716), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11713), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11517) );
  NAND2_X1 U14570 ( .A1(n11784), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11516) );
  NAND2_X1 U14571 ( .A1(n11517), .A2(n11516), .ZN(n13265) );
  NOR2_X1 U14572 ( .A1(n11519), .A2(n11518), .ZN(n11520) );
  OR2_X1 U14573 ( .A1(n11681), .A2(n11521), .ZN(n11525) );
  AOI22_X1 U14574 ( .A1(n11713), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11524) );
  NAND2_X1 U14575 ( .A1(n11784), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11523) );
  NAND2_X1 U14576 ( .A1(n11716), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11522) );
  NAND4_X1 U14577 ( .A1(n11525), .A2(n11524), .A3(n11523), .A4(n11522), .ZN(
        n13422) );
  INV_X1 U14578 ( .A(n11526), .ZN(n11527) );
  OR2_X1 U14579 ( .A1(n11681), .A2(n11527), .ZN(n11531) );
  AOI22_X1 U14580 ( .A1(n11716), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11713), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11530) );
  NAND2_X1 U14581 ( .A1(n11784), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14582 ( .A1(n11495), .A2(n11532), .B1(P2_REIP_REG_5__SCAN_IN), 
        .B2(n11784), .ZN(n11534) );
  AOI22_X1 U14583 ( .A1(n11716), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11713), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U14584 ( .A1(n11534), .A2(n11533), .ZN(n13629) );
  NAND2_X1 U14585 ( .A1(n13630), .A2(n13629), .ZN(n13628) );
  OR2_X1 U14586 ( .A1(n11681), .A2(n11535), .ZN(n15534) );
  NAND2_X1 U14587 ( .A1(n13628), .A2(n15534), .ZN(n11538) );
  AOI22_X1 U14588 ( .A1(n11716), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11713), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11537) );
  NAND2_X1 U14589 ( .A1(n11784), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11536) );
  NAND2_X1 U14590 ( .A1(n11537), .A2(n11536), .ZN(n15533) );
  NAND2_X1 U14591 ( .A1(n11538), .A2(n15533), .ZN(n15537) );
  INV_X1 U14592 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19188) );
  INV_X1 U14593 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19794) );
  OAI222_X1 U14594 ( .A1(n11700), .A2(n15527), .B1(n11701), .B2(n19188), .C1(
        n11702), .C2(n19794), .ZN(n15521) );
  INV_X1 U14595 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11540) );
  INV_X1 U14596 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12539) );
  OAI22_X1 U14597 ( .A1(n11540), .A2(n12653), .B1(n12654), .B2(n12539), .ZN(
        n11543) );
  OAI22_X1 U14598 ( .A1(n11541), .A2(n12656), .B1(n15588), .B2(n12538), .ZN(
        n11542) );
  NOR2_X1 U14599 ( .A1(n11543), .A2(n11542), .ZN(n11556) );
  INV_X1 U14600 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15618) );
  OAI22_X1 U14601 ( .A1(n15618), .A2(n11629), .B1(n11631), .B2(n11544), .ZN(
        n11550) );
  NAND2_X1 U14602 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11548) );
  NAND2_X1 U14603 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11547) );
  NAND2_X1 U14604 ( .A1(n10918), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11546) );
  NAND2_X1 U14605 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11545) );
  NAND4_X1 U14606 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n11549) );
  NOR2_X1 U14607 ( .A1(n11550), .A2(n11549), .ZN(n11555) );
  AOI22_X1 U14608 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12661), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11554) );
  NAND2_X1 U14609 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11553) );
  NAND2_X1 U14610 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11552) );
  AOI22_X1 U14611 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14612 ( .A1(n11716), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11713), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11558) );
  NAND2_X1 U14613 ( .A1(n11784), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11557) );
  OAI211_X1 U14614 ( .C1(n11681), .C2(n13284), .A(n11558), .B(n11557), .ZN(
        n15509) );
  INV_X1 U14615 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11560) );
  INV_X1 U14616 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11559) );
  OAI22_X1 U14617 ( .A1(n11560), .A2(n12653), .B1(n12654), .B2(n11559), .ZN(
        n11564) );
  OAI22_X1 U14618 ( .A1(n11562), .A2(n12656), .B1(n15588), .B2(n11561), .ZN(
        n11563) );
  NOR2_X1 U14619 ( .A1(n11564), .A2(n11563), .ZN(n11578) );
  INV_X1 U14620 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15623) );
  OAI22_X1 U14621 ( .A1(n15623), .A2(n11629), .B1(n11631), .B2(n11565), .ZN(
        n11571) );
  NAND2_X1 U14622 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11569) );
  NAND2_X1 U14623 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11568) );
  NAND2_X1 U14624 ( .A1(n10918), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11567) );
  NAND2_X1 U14625 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11566) );
  NAND4_X1 U14626 ( .A1(n11569), .A2(n11568), .A3(n11567), .A4(n11566), .ZN(
        n11570) );
  NOR2_X1 U14627 ( .A1(n11571), .A2(n11570), .ZN(n11577) );
  AOI22_X1 U14628 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12661), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11575) );
  NAND2_X1 U14629 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11574) );
  NAND2_X1 U14630 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11573) );
  AOI22_X1 U14631 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11572) );
  AND4_X1 U14632 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11576) );
  NAND3_X1 U14633 ( .A1(n11578), .A2(n11577), .A3(n11576), .ZN(n13312) );
  INV_X1 U14634 ( .A(n13312), .ZN(n13407) );
  NOR2_X1 U14635 ( .A1(n11681), .A2(n13407), .ZN(n11581) );
  INV_X1 U14636 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n11579) );
  OAI22_X1 U14637 ( .A1(n11701), .A2(n11579), .B1(n11700), .B2(n16109), .ZN(
        n11580) );
  AOI211_X1 U14638 ( .C1(n11784), .C2(P2_REIP_REG_10__SCAN_IN), .A(n11581), 
        .B(n11580), .ZN(n16175) );
  INV_X1 U14639 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11583) );
  INV_X1 U14640 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11582) );
  OAI22_X1 U14641 ( .A1(n11583), .A2(n12653), .B1(n12654), .B2(n11582), .ZN(
        n11587) );
  INV_X1 U14642 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11585) );
  INV_X1 U14643 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11584) );
  OAI22_X1 U14644 ( .A1(n11585), .A2(n12656), .B1(n15588), .B2(n11584), .ZN(
        n11586) );
  NOR2_X1 U14645 ( .A1(n11587), .A2(n11586), .ZN(n11601) );
  INV_X1 U14646 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15629) );
  INV_X1 U14647 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11588) );
  OAI22_X1 U14648 ( .A1(n15629), .A2(n11629), .B1(n11631), .B2(n11588), .ZN(
        n11594) );
  NAND2_X1 U14649 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11592) );
  NAND2_X1 U14650 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11591) );
  NAND2_X1 U14651 ( .A1(n10918), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11590) );
  NAND2_X1 U14652 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11589) );
  NAND4_X1 U14653 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n11589), .ZN(
        n11593) );
  NOR2_X1 U14654 ( .A1(n11594), .A2(n11593), .ZN(n11600) );
  AOI22_X1 U14655 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12661), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11598) );
  NAND2_X1 U14656 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11597) );
  NAND2_X1 U14657 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11596) );
  AOI22_X1 U14658 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11595) );
  AND4_X1 U14659 ( .A1(n11598), .A2(n11597), .A3(n11596), .A4(n11595), .ZN(
        n11599) );
  NAND3_X1 U14660 ( .A1(n11601), .A2(n11600), .A3(n11599), .ZN(n13411) );
  AOI22_X1 U14661 ( .A1(n11495), .A2(n13411), .B1(n11784), .B2(
        P2_REIP_REG_11__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14662 ( .A1(n11716), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11602) );
  NAND2_X1 U14663 ( .A1(n11603), .A2(n11602), .ZN(n15501) );
  INV_X1 U14664 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11604) );
  OAI22_X1 U14665 ( .A1(n15634), .A2(n11629), .B1(n11631), .B2(n11604), .ZN(
        n11610) );
  NAND2_X1 U14666 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11608) );
  NAND2_X1 U14667 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11607) );
  NAND2_X1 U14668 ( .A1(n10918), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11606) );
  NAND2_X1 U14669 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11605) );
  NAND4_X1 U14670 ( .A1(n11608), .A2(n11607), .A3(n11606), .A4(n11605), .ZN(
        n11609) );
  NOR2_X1 U14671 ( .A1(n11610), .A2(n11609), .ZN(n11620) );
  AOI22_X1 U14672 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10944), .B1(
        n10857), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14673 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10975), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11613) );
  NAND2_X1 U14674 ( .A1(n12570), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11612) );
  NAND2_X1 U14675 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11611) );
  AND4_X1 U14676 ( .A1(n11614), .A2(n11613), .A3(n11612), .A4(n11611), .ZN(
        n11619) );
  AOI22_X1 U14677 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12569), .B1(
        n10902), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11618) );
  INV_X1 U14678 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11615) );
  INV_X1 U14679 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12590) );
  OAI22_X1 U14680 ( .A1(n11615), .A2(n12656), .B1(n15588), .B2(n12590), .ZN(
        n11616) );
  INV_X1 U14681 ( .A(n11616), .ZN(n11617) );
  NAND4_X1 U14682 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n13471) );
  INV_X1 U14683 ( .A(n13471), .ZN(n11621) );
  OR2_X1 U14684 ( .A1(n11681), .A2(n11621), .ZN(n11624) );
  AOI22_X1 U14685 ( .A1(n11716), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11623) );
  NAND2_X1 U14686 ( .A1(n11784), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11622) );
  INV_X1 U14687 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11625) );
  INV_X1 U14688 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12613) );
  OAI22_X1 U14689 ( .A1(n12653), .A2(n11625), .B1(n12654), .B2(n12613), .ZN(
        n11628) );
  OAI22_X1 U14690 ( .A1(n15588), .A2(n12612), .B1(n12656), .B2(n11626), .ZN(
        n11627) );
  NOR2_X1 U14691 ( .A1(n11628), .A2(n11627), .ZN(n11644) );
  INV_X1 U14692 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15639) );
  OAI22_X1 U14693 ( .A1(n11631), .A2(n11630), .B1(n11629), .B2(n15639), .ZN(
        n11637) );
  NAND2_X1 U14694 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11635) );
  NAND2_X1 U14695 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11634) );
  NAND2_X1 U14696 ( .A1(n10918), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11633) );
  NAND2_X1 U14697 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11632) );
  NAND4_X1 U14698 ( .A1(n11635), .A2(n11634), .A3(n11633), .A4(n11632), .ZN(
        n11636) );
  NOR2_X1 U14699 ( .A1(n11637), .A2(n11636), .ZN(n11643) );
  AOI22_X1 U14700 ( .A1(n12661), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11641) );
  NAND2_X1 U14701 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11640) );
  NAND2_X1 U14702 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11639) );
  AOI22_X1 U14703 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11638) );
  AND4_X1 U14704 ( .A1(n11641), .A2(n11640), .A3(n11639), .A4(n11638), .ZN(
        n11642) );
  NAND3_X1 U14705 ( .A1(n11644), .A2(n11643), .A3(n11642), .ZN(n13479) );
  AOI22_X1 U14706 ( .A1(n11495), .A2(n13479), .B1(n11784), .B2(
        P2_REIP_REG_13__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14707 ( .A1(n11716), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11645) );
  NAND2_X1 U14708 ( .A1(n11646), .A2(n11645), .ZN(n16166) );
  NAND2_X1 U14709 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11650) );
  NAND2_X1 U14710 ( .A1(n12570), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11649) );
  NAND2_X1 U14711 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11648) );
  NAND2_X1 U14712 ( .A1(n12572), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11647) );
  NAND4_X1 U14713 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(
        n11656) );
  AOI22_X1 U14714 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12661), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U14715 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11653) );
  NAND2_X1 U14716 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11652) );
  AOI22_X1 U14717 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11651) );
  NAND4_X1 U14718 ( .A1(n11654), .A2(n11653), .A3(n11652), .A4(n11651), .ZN(
        n11655) );
  OR2_X1 U14719 ( .A1(n11656), .A2(n11655), .ZN(n11662) );
  AOI22_X1 U14720 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10937), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14721 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11659) );
  NAND2_X1 U14722 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11658) );
  NAND2_X1 U14723 ( .A1(n12668), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11657) );
  NAND4_X1 U14724 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n11661) );
  NOR2_X1 U14725 ( .A1(n11662), .A2(n11661), .ZN(n13609) );
  AOI22_X1 U14726 ( .A1(n11716), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11664) );
  NAND2_X1 U14727 ( .A1(n11784), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11663) );
  OAI211_X1 U14728 ( .C1(n11681), .C2(n13609), .A(n11664), .B(n11663), .ZN(
        n15462) );
  INV_X1 U14729 ( .A(n15462), .ZN(n11685) );
  NAND2_X1 U14730 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11668) );
  NAND2_X1 U14731 ( .A1(n12570), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11667) );
  NAND2_X1 U14732 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11666) );
  NAND2_X1 U14733 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11665) );
  NAND4_X1 U14734 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(
        n11674) );
  AOI22_X1 U14735 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12661), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11672) );
  NAND2_X1 U14736 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11671) );
  NAND2_X1 U14737 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11670) );
  AOI22_X1 U14738 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11669) );
  NAND4_X1 U14739 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11673) );
  OR2_X1 U14740 ( .A1(n11674), .A2(n11673), .ZN(n11680) );
  AOI22_X1 U14741 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10937), .B1(
        n12666), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14742 ( .A1(n10918), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11677) );
  NAND2_X1 U14743 ( .A1(n12572), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11676) );
  NAND2_X1 U14744 ( .A1(n12668), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11675) );
  NAND4_X1 U14745 ( .A1(n11678), .A2(n11677), .A3(n11676), .A4(n11675), .ZN(
        n11679) );
  NOR2_X1 U14746 ( .A1(n11680), .A2(n11679), .ZN(n13587) );
  OR2_X1 U14747 ( .A1(n11681), .A2(n13587), .ZN(n11684) );
  AOI22_X1 U14748 ( .A1(n11716), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11683) );
  NAND2_X1 U14749 ( .A1(n11784), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11682) );
  NOR2_X4 U14750 ( .A1(n16164), .A2(n11686), .ZN(n15460) );
  AOI22_X1 U14751 ( .A1(n11716), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11688) );
  NAND2_X1 U14752 ( .A1(n11784), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11687) );
  NAND2_X1 U14753 ( .A1(n11688), .A2(n11687), .ZN(n15448) );
  INV_X1 U14754 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19169) );
  OAI222_X1 U14755 ( .A1(n11702), .A2(n19808), .B1(n11701), .B2(n19169), .C1(
        n11689), .C2(n11700), .ZN(n13759) );
  AOI22_X1 U14756 ( .A1(n11716), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11691) );
  NAND2_X1 U14757 ( .A1(n11784), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11690) );
  AND2_X1 U14758 ( .A1(n11691), .A2(n11690), .ZN(n15416) );
  AOI22_X1 U14759 ( .A1(n11716), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11693) );
  NAND2_X1 U14760 ( .A1(n11784), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11692) );
  AND2_X1 U14761 ( .A1(n11693), .A2(n11692), .ZN(n15097) );
  AOI22_X1 U14762 ( .A1(n11716), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11695) );
  NAND2_X1 U14763 ( .A1(n11784), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11694) );
  NAND2_X1 U14764 ( .A1(n11695), .A2(n11694), .ZN(n15392) );
  AOI22_X1 U14765 ( .A1(n11716), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11697) );
  NAND2_X1 U14766 ( .A1(n11784), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11696) );
  AND2_X1 U14767 ( .A1(n11697), .A2(n11696), .ZN(n12925) );
  AOI22_X1 U14768 ( .A1(n11716), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11699) );
  NAND2_X1 U14769 ( .A1(n11784), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11698) );
  AND2_X1 U14770 ( .A1(n11699), .A2(n11698), .ZN(n15369) );
  INV_X1 U14771 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19157) );
  OAI222_X1 U14772 ( .A1(n11702), .A2(n19818), .B1(n11701), .B2(n19157), .C1(
        n15359), .C2(n11700), .ZN(n12938) );
  AOI22_X1 U14773 ( .A1(n11716), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11704) );
  NAND2_X1 U14774 ( .A1(n11784), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11703) );
  AND2_X1 U14775 ( .A1(n11704), .A2(n11703), .ZN(n15080) );
  AOI22_X1 U14776 ( .A1(n11716), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11706) );
  NAND2_X1 U14777 ( .A1(n11784), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11705) );
  AND2_X1 U14778 ( .A1(n11706), .A2(n11705), .ZN(n15067) );
  AOI22_X1 U14779 ( .A1(n11716), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11708) );
  NAND2_X1 U14780 ( .A1(n11784), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11707) );
  AND2_X1 U14781 ( .A1(n11708), .A2(n11707), .ZN(n15060) );
  AOI22_X1 U14782 ( .A1(n11716), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11710) );
  NAND2_X1 U14783 ( .A1(n11784), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11709) );
  NAND2_X1 U14784 ( .A1(n11710), .A2(n11709), .ZN(n12953) );
  AOI22_X1 U14785 ( .A1(n11716), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11712) );
  NAND2_X1 U14786 ( .A1(n11784), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11711) );
  AND2_X1 U14787 ( .A1(n11712), .A2(n11711), .ZN(n12964) );
  AOI22_X1 U14788 ( .A1(n11716), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11715) );
  NAND2_X1 U14789 ( .A1(n11784), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11714) );
  AND2_X1 U14790 ( .A1(n11715), .A2(n11714), .ZN(n12805) );
  AOI22_X1 U14791 ( .A1(n11716), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11713), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11718) );
  NAND2_X1 U14792 ( .A1(n11784), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11717) );
  NAND2_X1 U14793 ( .A1(n11718), .A2(n11717), .ZN(n11719) );
  INV_X1 U14794 ( .A(n14325), .ZN(n12900) );
  NAND2_X1 U14795 ( .A1(n10796), .A2(n19135), .ZN(n16224) );
  NAND2_X1 U14796 ( .A1(n16224), .A2(n15614), .ZN(n11723) );
  NAND2_X1 U14797 ( .A1(n15559), .A2(n11722), .ZN(n16227) );
  AND2_X1 U14798 ( .A1(n11723), .A2(n16227), .ZN(n11724) );
  INV_X1 U14799 ( .A(n11725), .ZN(n11726) );
  NAND2_X1 U14800 ( .A1(n11727), .A2(n11726), .ZN(n13530) );
  NAND2_X1 U14801 ( .A1(n11728), .A2(n15614), .ZN(n15560) );
  NAND2_X1 U14802 ( .A1(n15560), .A2(n11729), .ZN(n11730) );
  NAND2_X1 U14803 ( .A1(n11730), .A2(n15625), .ZN(n11745) );
  INV_X1 U14804 ( .A(n11731), .ZN(n12976) );
  OAI21_X1 U14805 ( .B1(n11734), .B2(n11732), .A(n12976), .ZN(n11737) );
  NAND3_X1 U14806 ( .A1(n11735), .A2(n11734), .A3(n11733), .ZN(n11736) );
  AND2_X1 U14807 ( .A1(n11737), .A2(n11736), .ZN(n11742) );
  NAND2_X1 U14808 ( .A1(n11739), .A2(n11738), .ZN(n12800) );
  NAND2_X1 U14809 ( .A1(n11740), .A2(n16231), .ZN(n11741) );
  AND4_X1 U14810 ( .A1(n11743), .A2(n11742), .A3(n12800), .A4(n11741), .ZN(
        n11744) );
  NAND2_X1 U14811 ( .A1(n11745), .A2(n11744), .ZN(n15576) );
  NOR2_X1 U14812 ( .A1(n15576), .A2(n11746), .ZN(n11747) );
  NAND2_X1 U14813 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11748) );
  OR2_X1 U14814 ( .A1(n15342), .A2(n11748), .ZN(n11769) );
  INV_X1 U14815 ( .A(n11769), .ZN(n11749) );
  OR2_X1 U14816 ( .A1(n15481), .A2(n11749), .ZN(n11760) );
  NOR2_X1 U14817 ( .A1(n15359), .A2(n15372), .ZN(n15354) );
  INV_X1 U14818 ( .A(n15481), .ZN(n15551) );
  NOR2_X1 U14819 ( .A1(n13624), .A2(n13623), .ZN(n13622) );
  OR2_X1 U14820 ( .A1(n15481), .A2(n13622), .ZN(n11752) );
  AND2_X1 U14821 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14338) );
  NOR2_X1 U14822 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14338), .ZN(
        n11764) );
  INV_X1 U14823 ( .A(n11764), .ZN(n11750) );
  NOR2_X1 U14824 ( .A1(n15437), .A2(n11750), .ZN(n14337) );
  NOR2_X1 U14825 ( .A1(n15443), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14340) );
  OR2_X1 U14826 ( .A1(n15443), .A2(n14338), .ZN(n11751) );
  INV_X2 U14827 ( .A(n16202), .ZN(n19034) );
  NAND2_X1 U14828 ( .A1(n11779), .A2(n19034), .ZN(n15552) );
  NAND2_X1 U14829 ( .A1(n11751), .A2(n15552), .ZN(n14343) );
  NOR3_X1 U14830 ( .A1(n14337), .A2(n14340), .A3(n14343), .ZN(n13549) );
  OAI21_X1 U14831 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15481), .A(
        n13549), .ZN(n13627) );
  INV_X1 U14832 ( .A(n13627), .ZN(n13596) );
  NAND2_X1 U14833 ( .A1(n11752), .A2(n13596), .ZN(n15541) );
  NOR2_X1 U14834 ( .A1(n15481), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11753) );
  NOR2_X1 U14835 ( .A1(n15541), .A2(n11753), .ZN(n16189) );
  NAND2_X1 U14836 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16203) );
  NAND2_X1 U14837 ( .A1(n15551), .A2(n16203), .ZN(n11754) );
  AND2_X1 U14838 ( .A1(n11755), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11766) );
  AND2_X1 U14839 ( .A1(n11766), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11756) );
  NAND2_X1 U14840 ( .A1(n15513), .A2(n11756), .ZN(n15441) );
  INV_X1 U14841 ( .A(n11757), .ZN(n15433) );
  NAND2_X1 U14842 ( .A1(n15433), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15424) );
  NOR2_X1 U14843 ( .A1(n15441), .A2(n15424), .ZN(n15421) );
  NAND2_X1 U14844 ( .A1(n15421), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15408) );
  NAND2_X1 U14845 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11768) );
  OAI21_X1 U14846 ( .B1(n15408), .B2(n11768), .A(n15440), .ZN(n15383) );
  INV_X1 U14847 ( .A(n15383), .ZN(n11758) );
  AOI21_X1 U14848 ( .B1(n20968), .B2(n15551), .A(n11758), .ZN(n15373) );
  OAI21_X1 U14849 ( .B1(n15354), .B2(n15481), .A(n15373), .ZN(n15322) );
  INV_X1 U14850 ( .A(n15322), .ZN(n11759) );
  NAND2_X1 U14851 ( .A1(n11760), .A2(n11759), .ZN(n15311) );
  NAND2_X1 U14852 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15282) );
  NOR2_X1 U14853 ( .A1(n15282), .A2(n15284), .ZN(n11788) );
  OAI21_X1 U14854 ( .B1(n15481), .B2(n11788), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11761) );
  NOR2_X1 U14855 ( .A1(n15311), .A2(n11761), .ZN(n11792) );
  INV_X1 U14856 ( .A(n15443), .ZN(n11762) );
  NAND3_X1 U14857 ( .A1(n11762), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        n14338), .ZN(n11763) );
  OAI21_X1 U14858 ( .B1(n11764), .B2(n15437), .A(n11763), .ZN(n13551) );
  NAND2_X1 U14859 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13551), .ZN(
        n13621) );
  INV_X1 U14860 ( .A(n13622), .ZN(n11765) );
  NOR2_X1 U14861 ( .A1(n13621), .A2(n11765), .ZN(n15539) );
  NAND2_X1 U14862 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15539), .ZN(
        n15519) );
  NAND2_X1 U14863 ( .A1(n16153), .A2(n11766), .ZN(n16163) );
  NOR2_X1 U14864 ( .A1(n15424), .A2(n15425), .ZN(n11767) );
  NAND2_X1 U14865 ( .A1(n15467), .A2(n11767), .ZN(n15410) );
  NOR2_X1 U14866 ( .A1(n15410), .A2(n11768), .ZN(n15385) );
  NAND2_X1 U14867 ( .A1(n15353), .A2(n15354), .ZN(n15341) );
  AOI21_X1 U14868 ( .B1(n11788), .B2(n15283), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11770) );
  NAND2_X1 U14869 ( .A1(n19236), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12842) );
  XNOR2_X1 U14870 ( .A(n15112), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12839) );
  NAND2_X1 U14871 ( .A1(n11773), .A2(n15106), .ZN(n11778) );
  INV_X1 U14872 ( .A(n11774), .ZN(n11776) );
  NAND2_X1 U14873 ( .A1(n11776), .A2(n11775), .ZN(n11777) );
  NAND2_X1 U14874 ( .A1(n16232), .A2(n11397), .ZN(n19891) );
  NAND3_X1 U14875 ( .A1(n10341), .A2(n11781), .A3(n11780), .ZN(P2_U3016) );
  NAND2_X1 U14876 ( .A1(n9830), .A2(n16183), .ZN(n11798) );
  NAND2_X1 U14877 ( .A1(n11782), .A2(n16196), .ZN(n11797) );
  AOI222_X1 U14878 ( .A1(n11784), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11716), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11713), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11785) );
  INV_X1 U14879 ( .A(n11785), .ZN(n11786) );
  NAND2_X1 U14880 ( .A1(n15440), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11791) );
  NAND4_X1 U14881 ( .A1(n11788), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12849), .A4(n15283), .ZN(n11789) );
  OAI211_X1 U14882 ( .C1(n11792), .C2(n11791), .A(n11790), .B(n11789), .ZN(
        n11793) );
  OAI21_X1 U14883 ( .B1(n11783), .B2(n16194), .A(n11794), .ZN(n11795) );
  INV_X1 U14884 ( .A(n11795), .ZN(n11796) );
  NAND3_X1 U14885 ( .A1(n11798), .A2(n11797), .A3(n11796), .ZN(P2_U3015) );
  XNOR2_X1 U14886 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11810) );
  NAND2_X1 U14887 ( .A1(n20581), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U14888 ( .A1(n11810), .A2(n11809), .ZN(n11800) );
  NAND2_X1 U14889 ( .A1(n20660), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11799) );
  NAND2_X1 U14890 ( .A1(n11800), .A2(n11799), .ZN(n11812) );
  XNOR2_X1 U14891 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11811) );
  NAND2_X1 U14892 ( .A1(n11812), .A2(n11811), .ZN(n11802) );
  NAND2_X1 U14893 ( .A1(n20420), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11801) );
  NAND2_X1 U14894 ( .A1(n11802), .A2(n11801), .ZN(n11814) );
  MUX2_X1 U14895 ( .A(n20618), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11813) );
  NAND2_X1 U14896 ( .A1(n11814), .A2(n11813), .ZN(n11804) );
  NAND2_X1 U14897 ( .A1(n20618), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11803) );
  NAND2_X1 U14898 ( .A1(n11804), .A2(n11803), .ZN(n11808) );
  NOR2_X1 U14899 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15995), .ZN(
        n11805) );
  XNOR2_X1 U14900 ( .A(n11810), .B(n11809), .ZN(n11950) );
  XNOR2_X1 U14901 ( .A(n11812), .B(n11811), .ZN(n11960) );
  XNOR2_X1 U14902 ( .A(n11814), .B(n11813), .ZN(n11965) );
  NOR4_X1 U14903 ( .A1(n11969), .A2(n11950), .A3(n11960), .A4(n11965), .ZN(
        n11815) );
  NOR2_X1 U14904 ( .A1(n11939), .A2(n11815), .ZN(n13061) );
  NAND2_X1 U14905 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20828) );
  NAND2_X1 U14906 ( .A1(n13061), .A2(n20828), .ZN(n13112) );
  NAND2_X1 U14907 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11819) );
  NAND2_X1 U14908 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11818) );
  NAND2_X1 U14909 ( .A1(n11877), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11817) );
  NOR2_X4 U14910 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11832) );
  AND2_X4 U14911 ( .A1(n11832), .A2(n11820), .ZN(n12288) );
  NAND2_X1 U14912 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11816) );
  NAND2_X1 U14913 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11824) );
  NAND2_X1 U14914 ( .A1(n12308), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11823) );
  AND2_X4 U14915 ( .A1(n11831), .A2(n11832), .ZN(n12307) );
  NAND2_X1 U14916 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11822) );
  AND2_X4 U14917 ( .A1(n11820), .A2(n14937), .ZN(n12282) );
  NAND2_X1 U14918 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11821) );
  AND2_X4 U14919 ( .A1(n11831), .A2(n11825), .ZN(n12203) );
  NAND2_X1 U14920 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11830) );
  NAND2_X1 U14921 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11829) );
  AND2_X4 U14922 ( .A1(n11826), .A2(n14937), .ZN(n12315) );
  NAND2_X1 U14923 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11828) );
  NAND2_X1 U14924 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11827) );
  NAND2_X1 U14925 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11836) );
  NAND2_X1 U14926 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11835) );
  NAND2_X1 U14928 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11834) );
  NAND2_X1 U14929 ( .A1(n12309), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11833) );
  INV_X1 U14930 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n11841) );
  XNOR2_X1 U14931 ( .A(n11841), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n12140) );
  NAND2_X1 U14932 ( .A1(n12140), .A2(n20735), .ZN(n15731) );
  AND2_X1 U14933 ( .A1(n12026), .A2(n15731), .ZN(n11842) );
  OR2_X1 U14934 ( .A1(n13112), .A2(n11842), .ZN(n11981) );
  AOI22_X1 U14935 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14936 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U14937 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14938 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U14939 ( .A1(n11877), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14940 ( .A1(n12308), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U14941 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14942 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14943 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14944 ( .A1(n12308), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U14945 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U14946 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11851) );
  NAND4_X1 U14947 ( .A1(n11854), .A2(n11853), .A3(n11852), .A4(n11851), .ZN(
        n11860) );
  AOI22_X1 U14948 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11877), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U14949 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U14950 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U14951 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11855) );
  NAND4_X1 U14952 ( .A1(n11858), .A2(n11857), .A3(n11856), .A4(n11855), .ZN(
        n11859) );
  AOI22_X1 U14953 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14954 ( .A1(n12308), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U14955 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U14956 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11861) );
  NAND4_X1 U14957 ( .A1(n11864), .A2(n11863), .A3(n11862), .A4(n11861), .ZN(
        n11872) );
  AOI22_X1 U14958 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11865), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14959 ( .A1(n11877), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14960 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U14961 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11867) );
  NAND4_X1 U14962 ( .A1(n11870), .A2(n11869), .A3(n11868), .A4(n11867), .ZN(
        n11871) );
  AOI22_X1 U14963 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U14964 ( .A1(n12308), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U14965 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14966 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11873) );
  NAND4_X1 U14967 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n11883) );
  AOI22_X1 U14968 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U14969 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U14970 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11877), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U14971 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11878) );
  NAND4_X1 U14972 ( .A1(n11881), .A2(n11880), .A3(n11879), .A4(n11878), .ZN(
        n11882) );
  OR2_X2 U14973 ( .A1(n11883), .A2(n11882), .ZN(n12256) );
  NAND2_X1 U14974 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11887) );
  NAND2_X1 U14975 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11886) );
  NAND2_X1 U14976 ( .A1(n11877), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11885) );
  NAND2_X1 U14977 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11884) );
  NAND2_X1 U14978 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11891) );
  NAND2_X1 U14979 ( .A1(n12308), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11890) );
  NAND2_X1 U14980 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11889) );
  NAND2_X1 U14981 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11888) );
  NAND2_X1 U14982 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11895) );
  NAND2_X1 U14983 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11894) );
  NAND2_X1 U14984 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11893) );
  NAND2_X1 U14985 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11892) );
  NAND2_X1 U14986 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11899) );
  NAND2_X1 U14987 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11898) );
  NAND2_X1 U14988 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11897) );
  NAND2_X1 U14989 ( .A1(n12309), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11896) );
  AOI22_X1 U14990 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11877), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U14991 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U14992 ( .A1(n12308), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U14993 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14994 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U14995 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U14996 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U14997 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11911) );
  NAND3_X2 U14998 ( .A1(n10356), .A2(n11914), .A3(n11913), .ZN(n11982) );
  NAND2_X1 U14999 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11920) );
  NAND2_X1 U15000 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11919) );
  NAND2_X1 U15001 ( .A1(n11877), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11918) );
  NAND2_X1 U15002 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11917) );
  NAND2_X1 U15003 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11924) );
  NAND2_X1 U15004 ( .A1(n12308), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11923) );
  NAND2_X1 U15005 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11922) );
  NAND2_X1 U15006 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11921) );
  NAND2_X1 U15007 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11928) );
  NAND2_X1 U15008 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11927) );
  NAND2_X1 U15009 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11926) );
  NAND2_X1 U15010 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11925) );
  NAND2_X1 U15011 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11932) );
  NAND2_X1 U15012 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11931) );
  NAND2_X1 U15013 ( .A1(n11865), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11930) );
  NAND2_X1 U15014 ( .A1(n12309), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11929) );
  AOI21_X1 U15015 ( .B1(n13118), .B2(n20828), .A(n20152), .ZN(n11938) );
  INV_X1 U15016 ( .A(n15731), .ZN(n15718) );
  NOR2_X1 U15017 ( .A1(n20821), .A2(n15718), .ZN(n11937) );
  OAI21_X1 U15018 ( .B1(n11938), .B2(n11937), .A(n13171), .ZN(n11979) );
  NAND2_X1 U15019 ( .A1(n12256), .A2(n12026), .ZN(n12391) );
  NAND2_X1 U15020 ( .A1(n11966), .A2(n11939), .ZN(n11978) );
  NAND2_X1 U15021 ( .A1(n11939), .A2(n12377), .ZN(n11976) );
  INV_X1 U15022 ( .A(n11940), .ZN(n12217) );
  NOR2_X1 U15023 ( .A1(n12217), .A2(n12426), .ZN(n11942) );
  OAI21_X1 U15024 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20581), .A(
        n11941), .ZN(n11943) );
  AOI21_X1 U15025 ( .B1(n20199), .B2(n13669), .A(n12026), .ZN(n11958) );
  NOR3_X1 U15026 ( .A1(n11942), .A2(n11943), .A3(n11958), .ZN(n11946) );
  INV_X1 U15027 ( .A(n11943), .ZN(n11944) );
  AOI21_X1 U15028 ( .B1(n11944), .B2(n12377), .A(n11966), .ZN(n11945) );
  INV_X1 U15029 ( .A(n11951), .ZN(n11955) );
  NAND2_X1 U15030 ( .A1(n20199), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11948) );
  OAI21_X1 U15031 ( .B1(n11956), .B2(n20169), .A(n11948), .ZN(n11947) );
  AOI21_X1 U15032 ( .B1(n12365), .B2(n11950), .A(n11947), .ZN(n11952) );
  INV_X1 U15033 ( .A(n11952), .ZN(n11954) );
  AND2_X1 U15034 ( .A1(n11948), .A2(n12026), .ZN(n11949) );
  NAND2_X1 U15035 ( .A1(n11956), .A2(n11949), .ZN(n11968) );
  AOI22_X1 U15036 ( .A1(n11952), .A2(n11951), .B1(n11950), .B2(n11968), .ZN(
        n11953) );
  AOI21_X1 U15037 ( .B1(n11955), .B2(n11954), .A(n11953), .ZN(n11962) );
  NOR2_X1 U15038 ( .A1(n11956), .A2(n11960), .ZN(n11957) );
  AOI211_X1 U15039 ( .C1(n12365), .C2(n11960), .A(n11958), .B(n11957), .ZN(
        n11961) );
  NAND2_X1 U15040 ( .A1(n11958), .A2(n12377), .ZN(n11959) );
  OAI22_X1 U15041 ( .A1(n11962), .A2(n11961), .B1(n11960), .B2(n11959), .ZN(
        n11964) );
  NAND2_X1 U15042 ( .A1(n12380), .A2(n11965), .ZN(n11963) );
  AOI22_X1 U15043 ( .A1(n11966), .A2(n11965), .B1(n11964), .B2(n11963), .ZN(
        n11973) );
  INV_X1 U15044 ( .A(n11969), .ZN(n11967) );
  NOR2_X1 U15045 ( .A1(n12365), .A2(n11967), .ZN(n11972) );
  INV_X1 U15046 ( .A(n11968), .ZN(n11970) );
  NAND3_X1 U15047 ( .A1(n12365), .A2(n11970), .A3(n11969), .ZN(n11971) );
  OAI21_X1 U15048 ( .B1(n11973), .B2(n11972), .A(n11971), .ZN(n11974) );
  AOI21_X1 U15049 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20824), .A(
        n11974), .ZN(n11975) );
  NAND2_X1 U15050 ( .A1(n11976), .A2(n11975), .ZN(n11977) );
  NAND2_X1 U15051 ( .A1(n11979), .A2(n13293), .ZN(n11980) );
  MUX2_X1 U15052 ( .A(n11981), .B(n11980), .S(n20177), .Z(n12001) );
  NAND2_X1 U15053 ( .A1(n20199), .A2(n13191), .ZN(n11983) );
  OR2_X1 U15054 ( .A1(n11989), .A2(n12120), .ZN(n11985) );
  NAND2_X1 U15055 ( .A1(n14933), .A2(n20152), .ZN(n11987) );
  NAND3_X1 U15056 ( .A1(n11988), .A2(n12257), .A3(n11987), .ZN(n12427) );
  INV_X1 U15057 ( .A(n12427), .ZN(n11991) );
  NAND2_X1 U15058 ( .A1(n11988), .A2(n20192), .ZN(n12019) );
  OR2_X1 U15059 ( .A1(n11989), .A2(n20169), .ZN(n12022) );
  AND2_X1 U15060 ( .A1(n12022), .A2(n13669), .ZN(n11990) );
  NAND2_X1 U15061 ( .A1(n12019), .A2(n11990), .ZN(n12010) );
  NAND2_X1 U15062 ( .A1(n11991), .A2(n12010), .ZN(n11999) );
  NAND2_X1 U15063 ( .A1(n13171), .A2(n11993), .ZN(n11995) );
  NAND3_X1 U15064 ( .A1(n13191), .A2(n20177), .A3(n12256), .ZN(n11994) );
  AND2_X2 U15065 ( .A1(n11997), .A2(n11996), .ZN(n12009) );
  NOR2_X1 U15066 ( .A1(n12426), .A2(n13669), .ZN(n11998) );
  INV_X1 U15067 ( .A(n12142), .ZN(n13060) );
  NAND2_X1 U15068 ( .A1(n11999), .A2(n13060), .ZN(n13115) );
  OR2_X1 U15069 ( .A1(n13293), .A2(n12022), .ZN(n12000) );
  NAND3_X1 U15070 ( .A1(n12001), .A2(n13115), .A3(n12000), .ZN(n12002) );
  INV_X1 U15071 ( .A(n13192), .ZN(n13097) );
  NAND2_X1 U15072 ( .A1(n11988), .A2(n13097), .ZN(n12007) );
  NAND2_X1 U15073 ( .A1(n13056), .A2(n14364), .ZN(n12005) );
  NAND2_X1 U15074 ( .A1(n20152), .A2(n12026), .ZN(n13113) );
  INV_X1 U15075 ( .A(n13113), .ZN(n13661) );
  NAND2_X1 U15076 ( .A1(n13661), .A2(n12426), .ZN(n12004) );
  NAND2_X1 U15077 ( .A1(n12005), .A2(n12004), .ZN(n12006) );
  AOI21_X1 U15078 ( .B1(n12007), .B2(n12026), .A(n12006), .ZN(n12012) );
  NAND2_X1 U15079 ( .A1(n12426), .A2(n12003), .ZN(n12008) );
  NAND2_X1 U15080 ( .A1(n12163), .A2(n13684), .ZN(n12011) );
  NAND2_X1 U15081 ( .A1(n13192), .A2(n11984), .ZN(n12159) );
  MUX2_X1 U15082 ( .A(n12017), .B(n20177), .S(n13669), .Z(n12013) );
  NAND3_X1 U15083 ( .A1(n13100), .A2(n12159), .A3(n12013), .ZN(n12014) );
  NAND2_X1 U15084 ( .A1(n12425), .A2(n12014), .ZN(n14870) );
  NAND2_X1 U15085 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20128) );
  NAND2_X1 U15086 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20106) );
  INV_X1 U15087 ( .A(n20106), .ZN(n12015) );
  NAND2_X1 U15088 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12015), .ZN(
        n14894) );
  NOR2_X1 U15089 ( .A1(n20128), .A2(n14894), .ZN(n14896) );
  INV_X1 U15090 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14737) );
  INV_X1 U15091 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15951) );
  NAND3_X1 U15092 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15939) );
  NOR3_X1 U15093 ( .A1(n12061), .A2(n15951), .A3(n15939), .ZN(n14895) );
  NAND2_X1 U15094 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14895), .ZN(
        n14898) );
  NOR2_X1 U15095 ( .A1(n14737), .A2(n14898), .ZN(n14871) );
  NAND2_X1 U15096 ( .A1(n14896), .A2(n14871), .ZN(n14869) );
  NOR2_X1 U15097 ( .A1(n14870), .A2(n14869), .ZN(n12024) );
  NAND2_X1 U15098 ( .A1(n12003), .A2(n13669), .ZN(n12016) );
  NAND2_X1 U15099 ( .A1(n12163), .A2(n20152), .ZN(n12021) );
  AND2_X1 U15100 ( .A1(n13097), .A2(n13113), .ZN(n12020) );
  NAND4_X1 U15101 ( .A1(n12154), .A2(n12166), .A3(n12021), .A4(n12020), .ZN(
        n12145) );
  NOR2_X1 U15102 ( .A1(n12145), .A2(n12022), .ZN(n13109) );
  NAND2_X1 U15103 ( .A1(n12425), .A2(n13109), .ZN(n20132) );
  INV_X1 U15104 ( .A(n20132), .ZN(n14899) );
  INV_X1 U15105 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20129) );
  INV_X1 U15106 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20122) );
  INV_X1 U15107 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21116) );
  OAI21_X1 U15108 ( .B1(n20129), .B2(n20122), .A(n21116), .ZN(n20127) );
  INV_X1 U15109 ( .A(n20127), .ZN(n15923) );
  NOR2_X1 U15110 ( .A1(n15923), .A2(n14894), .ZN(n15931) );
  NAND2_X1 U15111 ( .A1(n14871), .A2(n15931), .ZN(n12125) );
  INV_X1 U15112 ( .A(n12125), .ZN(n12023) );
  AOI22_X1 U15113 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n12024), .B1(
        n14899), .B2(n12023), .ZN(n14865) );
  INV_X1 U15114 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12404) );
  NOR2_X1 U15115 ( .A1(n14865), .A2(n12404), .ZN(n14847) );
  NOR2_X1 U15116 ( .A1(n12404), .A2(n14869), .ZN(n14867) );
  AND2_X1 U15117 ( .A1(n12142), .A2(n12026), .ZN(n15691) );
  NAND2_X1 U15118 ( .A1(n12425), .A2(n15691), .ZN(n14868) );
  INV_X1 U15119 ( .A(n14868), .ZN(n14846) );
  NOR2_X1 U15120 ( .A1(n14846), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14915) );
  OAI221_X1 U15121 ( .B1(n14847), .B2(n14867), .C1(n14847), .C2(n14892), .A(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15891) );
  NAND2_X1 U15122 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15893) );
  NOR2_X1 U15123 ( .A1(n15891), .A2(n15893), .ZN(n14874) );
  NAND2_X1 U15124 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n14874), .ZN(
        n15890) );
  INV_X1 U15125 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15828) );
  AND2_X1 U15126 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12130) );
  NAND2_X1 U15127 ( .A1(n15881), .A2(n12130), .ZN(n14841) );
  NAND2_X1 U15128 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12133) );
  AND2_X1 U15129 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14797) );
  NAND2_X1 U15130 ( .A1(n14797), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14624) );
  INV_X1 U15131 ( .A(n14624), .ZN(n14799) );
  NAND2_X1 U15132 ( .A1(n14799), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12025) );
  NOR2_X1 U15133 ( .A1(n14796), .A2(n12025), .ZN(n14793) );
  NAND2_X1 U15134 ( .A1(n14793), .A2(n10349), .ZN(n14770) );
  INV_X1 U15135 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12027) );
  NAND2_X1 U15136 ( .A1(n12105), .A2(n12027), .ZN(n12031) );
  NAND2_X1 U15137 ( .A1(n12112), .A2(n20122), .ZN(n12029) );
  OAI211_X1 U15138 ( .C1(n14360), .C2(P1_EBX_REG_1__SCAN_IN), .A(n12029), .B(
        n12099), .ZN(n12030) );
  NAND2_X1 U15139 ( .A1(n12031), .A2(n12030), .ZN(n12035) );
  NAND2_X1 U15140 ( .A1(n12112), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12034) );
  INV_X1 U15141 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12032) );
  NAND2_X1 U15142 ( .A1(n12099), .A2(n12032), .ZN(n12033) );
  NAND2_X1 U15143 ( .A1(n12034), .A2(n12033), .ZN(n13189) );
  INV_X1 U15144 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12036) );
  NAND2_X1 U15145 ( .A1(n12105), .A2(n12036), .ZN(n12039) );
  NAND2_X1 U15146 ( .A1(n12112), .A2(n21116), .ZN(n12037) );
  OAI211_X1 U15147 ( .C1(n14360), .C2(P1_EBX_REG_2__SCAN_IN), .A(n12037), .B(
        n12099), .ZN(n12038) );
  NAND2_X1 U15148 ( .A1(n12039), .A2(n12038), .ZN(n13243) );
  OR2_X1 U15149 ( .A1(n14364), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12041) );
  MUX2_X1 U15150 ( .A(n12109), .B(n12099), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12040) );
  AND2_X1 U15151 ( .A1(n12041), .A2(n12040), .ZN(n13404) );
  INV_X1 U15152 ( .A(n12112), .ZN(n12084) );
  MUX2_X1 U15153 ( .A(n12105), .B(n12084), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12043) );
  INV_X1 U15154 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20109) );
  OR2_X1 U15155 ( .A1(n12112), .A2(n13291), .ZN(n12069) );
  OAI21_X1 U15156 ( .B1(n13291), .B2(n20109), .A(n12069), .ZN(n12042) );
  NOR2_X1 U15157 ( .A1(n12043), .A2(n12042), .ZN(n13493) );
  OR2_X1 U15158 ( .A1(n12109), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n12048) );
  NAND2_X1 U15159 ( .A1(n12099), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12046) );
  OAI211_X1 U15160 ( .C1(n14360), .C2(P1_EBX_REG_5__SCAN_IN), .A(n12112), .B(
        n12046), .ZN(n12047) );
  NAND2_X1 U15161 ( .A1(n12048), .A2(n12047), .ZN(n15980) );
  MUX2_X1 U15162 ( .A(n12117), .B(n12112), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12051) );
  NAND2_X1 U15163 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14360), .ZN(
        n12049) );
  AND2_X1 U15164 ( .A1(n12069), .A2(n12049), .ZN(n12050) );
  NAND2_X1 U15165 ( .A1(n12051), .A2(n12050), .ZN(n15965) );
  OR2_X1 U15166 ( .A1(n12109), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n12054) );
  NAND2_X1 U15167 ( .A1(n12099), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12052) );
  OAI211_X1 U15168 ( .C1(n14360), .C2(P1_EBX_REG_7__SCAN_IN), .A(n12112), .B(
        n12052), .ZN(n12053) );
  AND2_X1 U15169 ( .A1(n12054), .A2(n12053), .ZN(n15964) );
  MUX2_X1 U15170 ( .A(n12117), .B(n12112), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12057) );
  NAND2_X1 U15171 ( .A1(n14360), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12055) );
  AND2_X1 U15172 ( .A1(n12069), .A2(n12055), .ZN(n12056) );
  NAND2_X1 U15173 ( .A1(n12057), .A2(n12056), .ZN(n13708) );
  OR2_X1 U15174 ( .A1(n12109), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n12060) );
  NAND2_X1 U15175 ( .A1(n12099), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12058) );
  OAI211_X1 U15176 ( .C1(n14360), .C2(P1_EBX_REG_9__SCAN_IN), .A(n12112), .B(
        n12058), .ZN(n12059) );
  NAND2_X1 U15177 ( .A1(n12060), .A2(n12059), .ZN(n15942) );
  INV_X1 U15178 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13787) );
  NAND2_X1 U15179 ( .A1(n12105), .A2(n13787), .ZN(n12064) );
  INV_X1 U15180 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12061) );
  NAND2_X1 U15181 ( .A1(n12112), .A2(n12061), .ZN(n12062) );
  OAI211_X1 U15182 ( .C1(n14360), .C2(P1_EBX_REG_10__SCAN_IN), .A(n12062), .B(
        n12099), .ZN(n12063) );
  OR2_X1 U15183 ( .A1(n14364), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12067) );
  MUX2_X1 U15184 ( .A(n12109), .B(n12099), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12066) );
  AND2_X1 U15185 ( .A1(n12067), .A2(n12066), .ZN(n13830) );
  MUX2_X1 U15186 ( .A(n12117), .B(n12112), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12071) );
  NAND2_X1 U15187 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14360), .ZN(
        n12068) );
  AND2_X1 U15188 ( .A1(n12069), .A2(n12068), .ZN(n12070) );
  NAND2_X1 U15189 ( .A1(n12071), .A2(n12070), .ZN(n13919) );
  INV_X1 U15190 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n12072) );
  MUX2_X1 U15191 ( .A(n14382), .B(n12109), .S(n12072), .Z(n12073) );
  OAI21_X1 U15192 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14364), .A(
        n12073), .ZN(n13871) );
  INV_X1 U15193 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n13906) );
  NAND2_X1 U15194 ( .A1(n12105), .A2(n13906), .ZN(n12076) );
  INV_X1 U15195 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15903) );
  NAND2_X1 U15196 ( .A1(n12112), .A2(n15903), .ZN(n12074) );
  OAI211_X1 U15197 ( .C1(n14360), .C2(P1_EBX_REG_14__SCAN_IN), .A(n12074), .B(
        n12099), .ZN(n12075) );
  INV_X1 U15198 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15800) );
  MUX2_X1 U15199 ( .A(n12099), .B(n12109), .S(n15800), .Z(n12078) );
  OR2_X1 U15200 ( .A1(n14364), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12077) );
  AND2_X1 U15201 ( .A1(n12078), .A2(n12077), .ZN(n14883) );
  INV_X1 U15202 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n13965) );
  NAND2_X1 U15203 ( .A1(n12105), .A2(n13965), .ZN(n12081) );
  INV_X1 U15204 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14860) );
  NAND2_X1 U15205 ( .A1(n12112), .A2(n14860), .ZN(n12079) );
  OAI211_X1 U15206 ( .C1(n14360), .C2(P1_EBX_REG_16__SCAN_IN), .A(n12079), .B(
        n14382), .ZN(n12080) );
  NAND2_X1 U15207 ( .A1(n12081), .A2(n12080), .ZN(n13963) );
  NAND2_X1 U15208 ( .A1(n14885), .A2(n13963), .ZN(n14525) );
  MUX2_X1 U15209 ( .A(n12109), .B(n12099), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12083) );
  OR2_X1 U15210 ( .A1(n14364), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12082) );
  NAND2_X1 U15211 ( .A1(n12083), .A2(n12082), .ZN(n14526) );
  MUX2_X1 U15212 ( .A(n12105), .B(n12084), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12086) );
  AND2_X1 U15213 ( .A1(n14360), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12085) );
  NOR2_X1 U15214 ( .A1(n12086), .A2(n12085), .ZN(n14518) );
  MUX2_X1 U15215 ( .A(n12109), .B(n12099), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12088) );
  OR2_X1 U15216 ( .A1(n14364), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12087) );
  NAND2_X1 U15217 ( .A1(n12088), .A2(n12087), .ZN(n14512) );
  MUX2_X1 U15218 ( .A(n12117), .B(n12112), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12090) );
  NAND2_X1 U15219 ( .A1(n14360), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12089) );
  NAND2_X1 U15220 ( .A1(n12090), .A2(n12089), .ZN(n14505) );
  MUX2_X1 U15221 ( .A(n12109), .B(n12099), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12092) );
  OR2_X1 U15222 ( .A1(n14364), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12091) );
  NAND2_X1 U15223 ( .A1(n12092), .A2(n12091), .ZN(n14499) );
  INV_X1 U15224 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n12093) );
  NAND2_X1 U15225 ( .A1(n12105), .A2(n12093), .ZN(n12096) );
  INV_X1 U15226 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14833) );
  NAND2_X1 U15227 ( .A1(n12112), .A2(n14833), .ZN(n12094) );
  OAI211_X1 U15228 ( .C1(n12028), .C2(P1_EBX_REG_22__SCAN_IN), .A(n12094), .B(
        n12099), .ZN(n12095) );
  AND2_X1 U15229 ( .A1(n12096), .A2(n12095), .ZN(n14493) );
  MUX2_X1 U15230 ( .A(n12109), .B(n12099), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12098) );
  OR2_X1 U15231 ( .A1(n14364), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12097) );
  AND2_X1 U15232 ( .A1(n12098), .A2(n12097), .ZN(n14459) );
  INV_X1 U15233 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14489) );
  NAND2_X1 U15234 ( .A1(n12105), .A2(n14489), .ZN(n12102) );
  INV_X1 U15235 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14819) );
  NAND2_X1 U15236 ( .A1(n12112), .A2(n14819), .ZN(n12100) );
  OAI211_X1 U15237 ( .C1(n14360), .C2(P1_EBX_REG_24__SCAN_IN), .A(n12100), .B(
        n12099), .ZN(n12101) );
  NAND2_X1 U15238 ( .A1(n12102), .A2(n12101), .ZN(n14454) );
  MUX2_X1 U15239 ( .A(n12109), .B(n12099), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12104) );
  OR2_X1 U15240 ( .A1(n14364), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12103) );
  NAND2_X1 U15241 ( .A1(n12104), .A2(n12103), .ZN(n14433) );
  INV_X1 U15242 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14485) );
  NAND2_X1 U15243 ( .A1(n12105), .A2(n14485), .ZN(n12108) );
  INV_X1 U15244 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14798) );
  NAND2_X1 U15245 ( .A1(n12112), .A2(n14798), .ZN(n12106) );
  OAI211_X1 U15246 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n14360), .A(n12106), .B(
        n12099), .ZN(n12107) );
  AND2_X1 U15247 ( .A1(n12108), .A2(n12107), .ZN(n14417) );
  MUX2_X1 U15248 ( .A(n12109), .B(n12099), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12111) );
  OR2_X1 U15249 ( .A1(n14364), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12110) );
  AND2_X1 U15250 ( .A1(n12111), .A2(n12110), .ZN(n14405) );
  INV_X1 U15251 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U15252 ( .A1(n12112), .A2(n14782), .ZN(n12113) );
  OAI211_X1 U15253 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n14360), .A(n12113), .B(
        n12099), .ZN(n12114) );
  OAI21_X1 U15254 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(n12117), .A(n12114), .ZN(
        n14226) );
  OR2_X1 U15255 ( .A1(n14364), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12116) );
  OR2_X1 U15256 ( .A1(n12028), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12115) );
  NAND2_X1 U15257 ( .A1(n12116), .A2(n12115), .ZN(n14380) );
  INV_X1 U15258 ( .A(n14382), .ZN(n13053) );
  OAI22_X1 U15259 ( .A1(n14380), .A2(n13053), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12117), .ZN(n12118) );
  NOR2_X1 U15260 ( .A1(n14379), .A2(n12118), .ZN(n12119) );
  NAND3_X1 U15261 ( .A1(n13192), .A2(n13684), .A3(n20199), .ZN(n13093) );
  NAND2_X1 U15262 ( .A1(n12141), .A2(n20169), .ZN(n15721) );
  OAI21_X1 U15263 ( .B1(n12429), .B2(n12120), .A(n15721), .ZN(n12121) );
  NOR2_X1 U15264 ( .A1(n14870), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12123) );
  NAND2_X1 U15265 ( .A1(n15992), .A2(n20824), .ZN(n13182) );
  OR2_X2 U15266 ( .A1(n13182), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20135) );
  NOR2_X1 U15267 ( .A1(n12425), .A2(n12122), .ZN(n14910) );
  INV_X1 U15268 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15892) );
  INV_X1 U15269 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14863) );
  NOR4_X1 U15270 ( .A1(n15903), .A2(n15892), .A3(n14860), .A4(n14863), .ZN(
        n14873) );
  AND2_X1 U15271 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14873), .ZN(
        n12126) );
  AND2_X1 U15272 ( .A1(n14867), .A2(n12126), .ZN(n12124) );
  NOR2_X1 U15273 ( .A1(n15930), .A2(n12124), .ZN(n12129) );
  NOR2_X1 U15274 ( .A1(n12404), .A2(n12125), .ZN(n15902) );
  AND2_X1 U15275 ( .A1(n15902), .A2(n12126), .ZN(n12127) );
  NOR2_X1 U15276 ( .A1(n20132), .A2(n12127), .ZN(n12128) );
  OR3_X1 U15277 ( .A1(n20120), .A2(n12129), .A3(n12128), .ZN(n15880) );
  INV_X1 U15278 ( .A(n12130), .ZN(n12132) );
  INV_X1 U15279 ( .A(n20120), .ZN(n12131) );
  NAND2_X1 U15280 ( .A1(n12131), .A2(n15952), .ZN(n15932) );
  OAI21_X1 U15281 ( .B1(n15880), .B2(n12132), .A(n15932), .ZN(n14840) );
  NAND2_X1 U15282 ( .A1(n15932), .A2(n12133), .ZN(n12134) );
  AND2_X1 U15283 ( .A1(n14840), .A2(n12134), .ZN(n14825) );
  OR2_X1 U15284 ( .A1(n15952), .A2(n14797), .ZN(n12135) );
  NAND2_X1 U15285 ( .A1(n14809), .A2(n15952), .ZN(n14761) );
  NAND3_X1 U15286 ( .A1(n14809), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12136) );
  NAND2_X1 U15287 ( .A1(n14761), .A2(n12136), .ZN(n14788) );
  OR2_X1 U15288 ( .A1(n15952), .A2(n10349), .ZN(n12137) );
  NAND2_X1 U15289 ( .A1(n14788), .A2(n12137), .ZN(n14760) );
  INV_X1 U15290 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20792) );
  NOR2_X1 U15291 ( .A1(n20135), .A2(n20792), .ZN(n14615) );
  AOI21_X1 U15292 ( .B1(n14760), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14615), .ZN(n12138) );
  OAI21_X1 U15293 ( .B1(n14482), .B2(n15936), .A(n12138), .ZN(n12139) );
  INV_X1 U15294 ( .A(n12139), .ZN(n12433) );
  NAND2_X1 U15295 ( .A1(n12141), .A2(n12140), .ZN(n12143) );
  NAND2_X1 U15296 ( .A1(n13118), .A2(n13291), .ZN(n13247) );
  NAND4_X1 U15297 ( .A1(n12143), .A2(n12428), .A3(n13247), .A4(n12429), .ZN(
        n12144) );
  NAND2_X1 U15298 ( .A1(n12145), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12146) );
  NAND2_X1 U15299 ( .A1(n12170), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12149) );
  NAND2_X1 U15300 ( .A1(n20660), .A2(n20581), .ZN(n20545) );
  NAND2_X1 U15301 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20656) );
  NAND2_X1 U15302 ( .A1(n20545), .A2(n20656), .ZN(n20619) );
  OR2_X1 U15303 ( .A1(n15726), .A2(n20660), .ZN(n12167) );
  OAI21_X1 U15304 ( .B1(n20619), .B2(n13182), .A(n12167), .ZN(n12147) );
  INV_X1 U15305 ( .A(n12147), .ZN(n12148) );
  NAND2_X1 U15306 ( .A1(n12149), .A2(n12148), .ZN(n12151) );
  NAND2_X1 U15307 ( .A1(n12170), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12153) );
  MUX2_X1 U15308 ( .A(n15726), .B(n13182), .S(n20581), .Z(n12152) );
  INV_X1 U15309 ( .A(n12154), .ZN(n12161) );
  INV_X1 U15310 ( .A(n12155), .ZN(n12156) );
  NAND2_X1 U15311 ( .A1(n12156), .A2(n12397), .ZN(n12158) );
  INV_X1 U15312 ( .A(n15992), .ZN(n20807) );
  NOR2_X1 U15313 ( .A1(n20807), .A2(n20824), .ZN(n12157) );
  NAND4_X1 U15314 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n13113), .ZN(
        n12160) );
  INV_X1 U15315 ( .A(n13684), .ZN(n13250) );
  NAND3_X1 U15316 ( .A1(n13250), .A2(n11989), .A3(n12250), .ZN(n12162) );
  NAND2_X1 U15317 ( .A1(n12163), .A2(n12162), .ZN(n12164) );
  NAND2_X2 U15318 ( .A1(n20277), .A2(n12239), .ZN(n12242) );
  INV_X1 U15319 ( .A(n12150), .ZN(n12169) );
  NAND2_X1 U15320 ( .A1(n12167), .A2(n9984), .ZN(n12168) );
  NAND2_X1 U15321 ( .A1(n12169), .A2(n12168), .ZN(n12175) );
  NAND2_X1 U15322 ( .A1(n12242), .A2(n12175), .ZN(n12173) );
  NOR2_X1 U15323 ( .A1(n15726), .A2(n20420), .ZN(n12171) );
  INV_X1 U15324 ( .A(n13182), .ZN(n12278) );
  XNOR2_X1 U15325 ( .A(n20656), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20161) );
  NAND2_X1 U15326 ( .A1(n12278), .A2(n20161), .ZN(n12174) );
  NAND2_X1 U15327 ( .A1(n12176), .A2(n12174), .ZN(n12172) );
  NAND2_X2 U15328 ( .A1(n12173), .A2(n12172), .ZN(n13335) );
  NAND4_X1 U15329 ( .A1(n12242), .A2(n12176), .A3(n12175), .A4(n12174), .ZN(
        n12177) );
  AOI22_X1 U15330 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15331 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15332 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15333 ( .A1(n14199), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12178) );
  NAND4_X1 U15334 ( .A1(n12181), .A2(n12180), .A3(n12179), .A4(n12178), .ZN(
        n12187) );
  BUF_X1 U15335 ( .A(n12314), .Z(n12287) );
  AOI22_X1 U15336 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U15337 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15338 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15339 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12182) );
  NAND4_X1 U15340 ( .A1(n12185), .A2(n12184), .A3(n12183), .A4(n12182), .ZN(
        n12186) );
  INV_X1 U15341 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n21161) );
  OAI22_X1 U15342 ( .A1(n12380), .A2(n21161), .B1(n12297), .B2(n12222), .ZN(
        n12188) );
  INV_X1 U15343 ( .A(n12190), .ZN(n12191) );
  AOI22_X1 U15344 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15345 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15346 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15347 ( .A1(n14199), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12193) );
  NAND4_X1 U15348 ( .A1(n12196), .A2(n12195), .A3(n12194), .A4(n12193), .ZN(
        n12202) );
  AOI22_X1 U15349 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U15350 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15351 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15352 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12197) );
  NAND4_X1 U15353 ( .A1(n12200), .A2(n12199), .A3(n12198), .A4(n12197), .ZN(
        n12201) );
  NAND2_X1 U15354 ( .A1(n20192), .A2(n12396), .ZN(n12219) );
  NOR2_X1 U15355 ( .A1(n12243), .A2(n12396), .ZN(n12235) );
  AOI22_X1 U15356 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15357 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15358 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15359 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12204) );
  NAND4_X1 U15360 ( .A1(n12207), .A2(n12206), .A3(n12205), .A4(n12204), .ZN(
        n12213) );
  AOI22_X1 U15361 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15362 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15363 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15364 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12208) );
  NAND4_X1 U15365 ( .A1(n12211), .A2(n12210), .A3(n12209), .A4(n12208), .ZN(
        n12212) );
  MUX2_X1 U15366 ( .A(n12220), .B(n12235), .S(n12265), .Z(n12214) );
  INV_X1 U15367 ( .A(n12214), .ZN(n12215) );
  INV_X1 U15368 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n21141) );
  OAI21_X1 U15369 ( .B1(n12265), .B2(n20824), .A(n12217), .ZN(n12218) );
  OAI211_X1 U15370 ( .C1(n12380), .C2(n21141), .A(n12219), .B(n12218), .ZN(
        n12262) );
  NAND2_X1 U15371 ( .A1(n12263), .A2(n12262), .ZN(n12221) );
  INV_X1 U15372 ( .A(n12220), .ZN(n12392) );
  NAND2_X1 U15373 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12238) );
  INV_X1 U15374 ( .A(n12222), .ZN(n12234) );
  BUF_X1 U15375 ( .A(n12306), .Z(n12223) );
  AOI22_X1 U15376 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15377 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12281), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15378 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15379 ( .A1(n14199), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12224) );
  NAND4_X1 U15380 ( .A1(n12227), .A2(n12226), .A3(n12225), .A4(n12224), .ZN(
        n12233) );
  AOI22_X1 U15381 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15382 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15383 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15384 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12228) );
  NAND4_X1 U15385 ( .A1(n12231), .A2(n12230), .A3(n12229), .A4(n12228), .ZN(
        n12232) );
  NAND2_X1 U15386 ( .A1(n12234), .A2(n12255), .ZN(n12237) );
  INV_X1 U15387 ( .A(n12235), .ZN(n12236) );
  INV_X1 U15388 ( .A(n20277), .ZN(n12241) );
  INV_X1 U15389 ( .A(n12239), .ZN(n12240) );
  INV_X1 U15390 ( .A(n12243), .ZN(n12244) );
  NAND2_X1 U15391 ( .A1(n13207), .A2(n13208), .ZN(n12249) );
  INV_X1 U15392 ( .A(n12245), .ZN(n12246) );
  INV_X1 U15393 ( .A(n12391), .ZN(n12382) );
  NAND2_X1 U15394 ( .A1(n12255), .A2(n12265), .ZN(n12298) );
  XNOR2_X1 U15395 ( .A(n12298), .B(n12297), .ZN(n12252) );
  NAND2_X1 U15396 ( .A1(n20152), .A2(n12250), .ZN(n12264) );
  INV_X1 U15397 ( .A(n12264), .ZN(n12251) );
  AOI21_X1 U15398 ( .B1(n12252), .B2(n12397), .A(n12251), .ZN(n12253) );
  NAND2_X1 U15399 ( .A1(n12254), .A2(n12253), .ZN(n13277) );
  XNOR2_X1 U15400 ( .A(n12255), .B(n12265), .ZN(n12258) );
  OAI211_X1 U15401 ( .C1(n12258), .C2(n20821), .A(n12257), .B(n12256), .ZN(
        n12259) );
  INV_X1 U15402 ( .A(n12259), .ZN(n12260) );
  OAI21_X1 U15403 ( .B1(n20821), .B2(n12265), .A(n12264), .ZN(n12266) );
  INV_X1 U15404 ( .A(n12266), .ZN(n12267) );
  INV_X1 U15405 ( .A(n12268), .ZN(n12269) );
  NAND2_X1 U15406 ( .A1(n9806), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12272) );
  INV_X1 U15407 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20118) );
  INV_X1 U15408 ( .A(n12273), .ZN(n12274) );
  NAND2_X1 U15409 ( .A1(n12170), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12280) );
  INV_X1 U15410 ( .A(n20656), .ZN(n15694) );
  INV_X1 U15411 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20618) );
  NAND2_X1 U15412 ( .A1(n20618), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20363) );
  INV_X1 U15413 ( .A(n20363), .ZN(n12275) );
  NAND2_X1 U15414 ( .A1(n15694), .A2(n12275), .ZN(n20391) );
  OAI21_X1 U15415 ( .B1(n20656), .B2(n20420), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12276) );
  NAND2_X1 U15416 ( .A1(n20391), .A2(n12276), .ZN(n20422) );
  INV_X1 U15417 ( .A(n15726), .ZN(n12277) );
  AOI22_X1 U15418 ( .A1(n20422), .A2(n12278), .B1(n12277), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12279) );
  XNOR2_X2 U15419 ( .A(n13335), .B(n20309), .ZN(n20421) );
  AOI22_X1 U15420 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15421 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15422 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15423 ( .A1(n14199), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12283) );
  NAND4_X1 U15424 ( .A1(n12286), .A2(n12285), .A3(n12284), .A4(n12283), .ZN(
        n12294) );
  AOI22_X1 U15425 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15426 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15427 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15428 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12289) );
  NAND4_X1 U15429 ( .A1(n12292), .A2(n12291), .A3(n12290), .A4(n12289), .ZN(
        n12293) );
  AOI22_X1 U15430 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12377), .B2(n12346), .ZN(n12295) );
  NAND2_X1 U15431 ( .A1(n20146), .A2(n12382), .ZN(n12302) );
  NAND2_X1 U15432 ( .A1(n12298), .A2(n12297), .ZN(n12348) );
  INV_X1 U15433 ( .A(n12346), .ZN(n12299) );
  XNOR2_X1 U15434 ( .A(n12348), .B(n12299), .ZN(n12300) );
  NAND2_X1 U15435 ( .A1(n12300), .A2(n12397), .ZN(n12301) );
  NAND2_X1 U15436 ( .A1(n12302), .A2(n12301), .ZN(n13462) );
  NAND2_X1 U15437 ( .A1(n12303), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12304) );
  NAND2_X2 U15438 ( .A1(n13461), .A2(n12304), .ZN(n12329) );
  INV_X1 U15439 ( .A(n12332), .ZN(n12324) );
  INV_X1 U15440 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U15441 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14015), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15442 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12307), .B1(
        n12281), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15443 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11906), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15444 ( .A1(n14199), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12310) );
  NAND4_X1 U15445 ( .A1(n12313), .A2(n12312), .A3(n12311), .A4(n12310), .ZN(
        n12321) );
  AOI22_X1 U15446 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U15447 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U15448 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15449 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12316) );
  NAND4_X1 U15450 ( .A1(n12319), .A2(n12318), .A3(n12317), .A4(n12316), .ZN(
        n12320) );
  NAND2_X1 U15451 ( .A1(n12377), .A2(n12345), .ZN(n12322) );
  XNOR2_X1 U15452 ( .A(n12324), .B(n12331), .ZN(n13490) );
  NAND2_X1 U15453 ( .A1(n13490), .A2(n12382), .ZN(n12328) );
  NAND2_X1 U15454 ( .A1(n12348), .A2(n12346), .ZN(n12325) );
  XNOR2_X1 U15455 ( .A(n12325), .B(n12345), .ZN(n12326) );
  NAND2_X1 U15456 ( .A1(n12326), .A2(n12397), .ZN(n12327) );
  NAND2_X1 U15457 ( .A1(n12328), .A2(n12327), .ZN(n20092) );
  NAND2_X1 U15458 ( .A1(n12329), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12330) );
  INV_X1 U15459 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U15460 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15461 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15462 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15463 ( .A1(n14199), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12333) );
  NAND4_X1 U15464 ( .A1(n12336), .A2(n12335), .A3(n12334), .A4(n12333), .ZN(
        n12342) );
  AOI22_X1 U15465 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15466 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15467 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15468 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12337) );
  NAND4_X1 U15469 ( .A1(n12340), .A2(n12339), .A3(n12338), .A4(n12337), .ZN(
        n12341) );
  NAND2_X1 U15470 ( .A1(n12377), .A2(n12368), .ZN(n12343) );
  OAI21_X1 U15471 ( .B1(n12380), .B2(n12344), .A(n12343), .ZN(n12354) );
  XNOR2_X1 U15472 ( .A(n12353), .B(n12354), .ZN(n13519) );
  NAND2_X1 U15473 ( .A1(n13519), .A2(n12382), .ZN(n12351) );
  AND2_X1 U15474 ( .A1(n12346), .A2(n12345), .ZN(n12347) );
  NAND2_X1 U15475 ( .A1(n12348), .A2(n12347), .ZN(n12370) );
  XNOR2_X1 U15476 ( .A(n12370), .B(n12368), .ZN(n12349) );
  NAND2_X1 U15477 ( .A1(n12349), .A2(n12397), .ZN(n12350) );
  NAND2_X1 U15478 ( .A1(n12351), .A2(n12350), .ZN(n12352) );
  INV_X1 U15479 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15988) );
  XNOR2_X1 U15480 ( .A(n12352), .B(n15988), .ZN(n15872) );
  AOI22_X1 U15481 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15482 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15483 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15484 ( .A1(n14199), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12355) );
  NAND4_X1 U15485 ( .A1(n12358), .A2(n12357), .A3(n12356), .A4(n12355), .ZN(
        n12364) );
  AOI22_X1 U15486 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15487 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15488 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15489 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12359) );
  NAND4_X1 U15490 ( .A1(n12362), .A2(n12361), .A3(n12360), .A4(n12359), .ZN(
        n12363) );
  AOI22_X1 U15491 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12377), .B2(n12384), .ZN(n12366) );
  NAND2_X1 U15492 ( .A1(n12367), .A2(n12366), .ZN(n13642) );
  NAND3_X1 U15493 ( .A1(n12394), .A2(n13642), .A3(n12382), .ZN(n12373) );
  INV_X1 U15494 ( .A(n12368), .ZN(n12369) );
  OR2_X1 U15495 ( .A1(n12370), .A2(n12369), .ZN(n12383) );
  XNOR2_X1 U15496 ( .A(n12383), .B(n12384), .ZN(n12371) );
  NAND2_X1 U15497 ( .A1(n12371), .A2(n12397), .ZN(n12372) );
  INV_X1 U15498 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15961) );
  NAND2_X1 U15499 ( .A1(n15867), .A2(n15961), .ZN(n12374) );
  INV_X1 U15500 ( .A(n15867), .ZN(n12375) );
  NAND2_X1 U15501 ( .A1(n12375), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12376) );
  INV_X1 U15502 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12379) );
  NAND2_X1 U15503 ( .A1(n12377), .A2(n12396), .ZN(n12378) );
  OAI21_X1 U15504 ( .B1(n12380), .B2(n12379), .A(n12378), .ZN(n12381) );
  NAND2_X1 U15505 ( .A1(n13649), .A2(n12382), .ZN(n12388) );
  INV_X1 U15506 ( .A(n12383), .ZN(n12385) );
  NAND2_X1 U15507 ( .A1(n12385), .A2(n12384), .ZN(n12395) );
  XNOR2_X1 U15508 ( .A(n12395), .B(n12396), .ZN(n12386) );
  NAND2_X1 U15509 ( .A1(n12386), .A2(n12397), .ZN(n12387) );
  NAND2_X1 U15510 ( .A1(n12388), .A2(n12387), .ZN(n12389) );
  OR2_X1 U15511 ( .A1(n12389), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15862) );
  NAND2_X1 U15512 ( .A1(n15860), .A2(n15862), .ZN(n12390) );
  NAND2_X1 U15513 ( .A1(n12389), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15861) );
  NOR2_X1 U15514 ( .A1(n12392), .A2(n12391), .ZN(n12393) );
  INV_X4 U15515 ( .A(n10332), .ZN(n15852) );
  INV_X1 U15516 ( .A(n12395), .ZN(n12398) );
  NAND3_X1 U15517 ( .A1(n12398), .A2(n12397), .A3(n12396), .ZN(n12399) );
  INV_X1 U15518 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12400) );
  NAND2_X1 U15519 ( .A1(n13800), .A2(n12400), .ZN(n12401) );
  INV_X1 U15520 ( .A(n13800), .ZN(n12402) );
  NAND2_X1 U15521 ( .A1(n12402), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12403) );
  NAND2_X1 U15522 ( .A1(n10332), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14724) );
  NAND2_X1 U15523 ( .A1(n15852), .A2(n12404), .ZN(n12405) );
  NAND2_X1 U15524 ( .A1(n14724), .A2(n12405), .ZN(n14739) );
  AND2_X1 U15525 ( .A1(n15852), .A2(n14737), .ZN(n14738) );
  NAND2_X1 U15526 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12406) );
  NAND2_X1 U15527 ( .A1(n15852), .A2(n12406), .ZN(n14733) );
  NAND2_X1 U15528 ( .A1(n15852), .A2(n15903), .ZN(n12407) );
  AND2_X1 U15529 ( .A1(n14733), .A2(n12407), .ZN(n12408) );
  NAND2_X1 U15530 ( .A1(n14723), .A2(n12408), .ZN(n14707) );
  NAND2_X1 U15531 ( .A1(n10332), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12409) );
  NAND2_X1 U15532 ( .A1(n14724), .A2(n12409), .ZN(n12412) );
  NOR2_X1 U15533 ( .A1(n15852), .A2(n15892), .ZN(n14711) );
  NOR2_X1 U15534 ( .A1(n12412), .A2(n14711), .ZN(n14856) );
  XNOR2_X1 U15535 ( .A(n15852), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14713) );
  NAND2_X1 U15536 ( .A1(n15852), .A2(n15892), .ZN(n14878) );
  NAND2_X1 U15537 ( .A1(n14713), .A2(n14878), .ZN(n12410) );
  NAND2_X1 U15538 ( .A1(n14857), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12411) );
  INV_X1 U15539 ( .A(n12412), .ZN(n12414) );
  NOR2_X1 U15540 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14734) );
  NAND2_X1 U15541 ( .A1(n14734), .A2(n14737), .ZN(n12413) );
  NAND2_X1 U15542 ( .A1(n10332), .A2(n12413), .ZN(n14722) );
  NAND2_X1 U15543 ( .A1(n12414), .A2(n14722), .ZN(n14708) );
  OAI21_X2 U15544 ( .B1(n14685), .B2(n12417), .A(n10332), .ZN(n14677) );
  XNOR2_X1 U15545 ( .A(n15852), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14700) );
  INV_X1 U15546 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21133) );
  NOR2_X1 U15547 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14653) );
  INV_X1 U15548 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14808) );
  NOR2_X1 U15549 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12420) );
  NAND2_X1 U15550 ( .A1(n12421), .A2(n12420), .ZN(n14292) );
  NAND2_X1 U15551 ( .A1(n12422), .A2(n14292), .ZN(n14297) );
  AND2_X1 U15552 ( .A1(n15852), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14605) );
  INV_X1 U15553 ( .A(n14605), .ZN(n12423) );
  INV_X1 U15554 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14757) );
  NAND2_X1 U15555 ( .A1(n10332), .A2(n14757), .ZN(n14293) );
  AND2_X1 U15556 ( .A1(n12423), .A2(n14293), .ZN(n12424) );
  XNOR2_X1 U15557 ( .A(n14297), .B(n12424), .ZN(n14621) );
  INV_X1 U15558 ( .A(n12425), .ZN(n12432) );
  NOR2_X1 U15559 ( .A1(n12427), .A2(n12426), .ZN(n15707) );
  NOR2_X1 U15560 ( .A1(n12427), .A2(n13250), .ZN(n13110) );
  OR2_X1 U15561 ( .A1(n15707), .A2(n13110), .ZN(n13057) );
  OAI211_X1 U15562 ( .C1(n20192), .C2(n12429), .A(n12428), .B(n13247), .ZN(
        n12430) );
  NOR2_X1 U15563 ( .A1(n13057), .A2(n12430), .ZN(n12431) );
  OAI211_X1 U15564 ( .C1(n14770), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12433), .B(n10348), .ZN(P1_U3002) );
  XNOR2_X1 U15565 ( .A(n12436), .B(n12438), .ZN(n15116) );
  INV_X1 U15566 ( .A(n12436), .ZN(n12437) );
  XNOR2_X1 U15567 ( .A(n12439), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12440) );
  XNOR2_X1 U15568 ( .A(n12441), .B(n12440), .ZN(n15307) );
  INV_X1 U15569 ( .A(n19242), .ZN(n12452) );
  INV_X1 U15570 ( .A(n12835), .ZN(n12444) );
  NAND2_X1 U15571 ( .A1(n12951), .A2(n12442), .ZN(n12443) );
  INV_X1 U15572 ( .A(n15296), .ZN(n12450) );
  INV_X1 U15573 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12448) );
  AND2_X1 U15574 ( .A1(n12445), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12882) );
  NOR2_X1 U15575 ( .A1(n12445), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12446) );
  NOR2_X1 U15576 ( .A1(n12882), .A2(n12446), .ZN(n12961) );
  NAND2_X1 U15577 ( .A1(n16143), .A2(n12961), .ZN(n12447) );
  NAND2_X1 U15578 ( .A1(n19236), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15300) );
  OAI211_X1 U15579 ( .C1(n16150), .C2(n12448), .A(n12447), .B(n15300), .ZN(
        n12449) );
  NOR4_X1 U15580 ( .A1(n18813), .A2(n18199), .A3(n18608), .A4(n12453), .ZN(
        n12465) );
  INV_X1 U15581 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18684) );
  NOR2_X2 U15582 ( .A1(n16410), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18754) );
  NOR2_X1 U15583 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16415) );
  INV_X1 U15584 ( .A(n16415), .ZN(n18683) );
  NAND3_X1 U15585 ( .A1(n18684), .A2(n18757), .A3(n18683), .ZN(n18811) );
  NAND2_X1 U15586 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18814) );
  INV_X1 U15587 ( .A(n18814), .ZN(n18693) );
  AOI21_X1 U15588 ( .B1(n18811), .B2(n12454), .A(n18693), .ZN(n16416) );
  AND3_X1 U15589 ( .A1(n12456), .A2(n12455), .A3(n16416), .ZN(n12464) );
  AOI21_X1 U15590 ( .B1(n18190), .B2(n12457), .A(n13975), .ZN(n12463) );
  INV_X1 U15591 ( .A(n12458), .ZN(n12461) );
  OAI211_X1 U15592 ( .C1(n12462), .C2(n12461), .A(n12460), .B(n12459), .ZN(
        n13974) );
  NOR4_X1 U15593 ( .A1(n12465), .A2(n12464), .A3(n12463), .A4(n13974), .ZN(
        n12466) );
  NOR3_X4 U15594 ( .A1(n12467), .A2(n18142), .A3(n17327), .ZN(n18078) );
  NAND2_X1 U15595 ( .A1(n18134), .A2(n18076), .ZN(n18110) );
  INV_X1 U15596 ( .A(n18110), .ZN(n18145) );
  NOR3_X1 U15597 ( .A1(n18085), .A2(n18091), .A3(n18070), .ZN(n12469) );
  NAND2_X1 U15598 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18108) );
  NAND3_X1 U15599 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17964) );
  NOR2_X1 U15600 ( .A1(n18108), .A2(n17964), .ZN(n18073) );
  NAND2_X1 U15601 ( .A1(n12469), .A2(n18073), .ZN(n17972) );
  NOR2_X1 U15602 ( .A1(n21150), .A2(n17972), .ZN(n18035) );
  INV_X1 U15603 ( .A(n18035), .ZN(n18058) );
  NOR2_X1 U15604 ( .A1(n17967), .A2(n18058), .ZN(n17934) );
  INV_X1 U15605 ( .A(n17934), .ZN(n17975) );
  NOR2_X1 U15606 ( .A1(n17853), .A2(n17975), .ZN(n17924) );
  INV_X1 U15607 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17862) );
  NOR2_X1 U15608 ( .A1(n17851), .A2(n17862), .ZN(n16314) );
  NAND2_X1 U15609 ( .A1(n17924), .A2(n16314), .ZN(n12472) );
  AOI21_X1 U15610 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18106) );
  NOR2_X1 U15611 ( .A1(n18106), .A2(n17964), .ZN(n18071) );
  NAND2_X1 U15612 ( .A1(n12469), .A2(n18071), .ZN(n17973) );
  NOR3_X1 U15613 ( .A1(n17620), .A2(n17967), .A3(n17973), .ZN(n17956) );
  NAND2_X1 U15614 ( .A1(n16312), .A2(n17956), .ZN(n17900) );
  NOR2_X1 U15615 ( .A1(n17882), .A2(n17900), .ZN(n17852) );
  NAND2_X1 U15616 ( .A1(n12470), .A2(n17852), .ZN(n12477) );
  NOR2_X1 U15617 ( .A1(n17967), .A2(n17972), .ZN(n17957) );
  NAND2_X1 U15618 ( .A1(n12471), .A2(n17957), .ZN(n12476) );
  AOI222_X1 U15619 ( .A1(n18637), .A2(n12472), .B1(n12477), .B2(n18635), .C1(
        n12476), .C2(n18623), .ZN(n15672) );
  OAI21_X1 U15620 ( .B1(n15672), .B2(n18142), .A(n18109), .ZN(n12473) );
  AOI21_X1 U15621 ( .B1(n18145), .B2(n12474), .A(n12473), .ZN(n16300) );
  NOR2_X1 U15622 ( .A1(n16282), .A2(n16317), .ZN(n12475) );
  NAND2_X1 U15623 ( .A1(n18609), .A2(n18134), .ZN(n18154) );
  NAND2_X1 U15624 ( .A1(n18066), .A2(n18150), .ZN(n18156) );
  INV_X1 U15625 ( .A(n16277), .ZN(n16296) );
  AOI22_X1 U15626 ( .A1(n12475), .A2(n18141), .B1(n18139), .B2(n16296), .ZN(
        n15673) );
  AOI21_X1 U15627 ( .B1(n16300), .B2(n15673), .A(n16265), .ZN(n12483) );
  AOI21_X1 U15628 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18637), .A(
        n18623), .ZN(n18125) );
  OAI22_X1 U15629 ( .A1(n18612), .A2(n12477), .B1(n12476), .B2(n18125), .ZN(
        n16303) );
  NAND2_X1 U15630 ( .A1(n18609), .A2(n17327), .ZN(n18015) );
  OAI22_X1 U15631 ( .A1(n18611), .A2(n17858), .B1(n17855), .B2(n18015), .ZN(
        n12478) );
  OAI21_X1 U15632 ( .B1(n16303), .B2(n12478), .A(n18150), .ZN(n15675) );
  OAI21_X1 U15633 ( .B1(n10754), .B2(n19904), .A(n19469), .ZN(n12507) );
  NOR2_X1 U15634 ( .A1(n15596), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12486) );
  AOI21_X1 U15635 ( .B1(n12507), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12486), .ZN(n12487) );
  AND2_X1 U15636 ( .A1(n12758), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12495) );
  NAND2_X1 U15637 ( .A1(n12489), .A2(n12505), .ZN(n12493) );
  NAND2_X1 U15638 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19312) );
  NOR2_X1 U15639 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19466) );
  INV_X1 U15640 ( .A(n19466), .ZN(n12490) );
  NAND2_X1 U15641 ( .A1(n19312), .A2(n12490), .ZN(n19407) );
  OR2_X1 U15642 ( .A1(n19407), .A2(n15596), .ZN(n19539) );
  INV_X1 U15643 ( .A(n19539), .ZN(n12491) );
  AOI21_X1 U15644 ( .B1(n12507), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12491), .ZN(n12492) );
  INV_X1 U15645 ( .A(n12494), .ZN(n12497) );
  INV_X1 U15646 ( .A(n12495), .ZN(n12496) );
  NAND2_X1 U15647 ( .A1(n12497), .A2(n12496), .ZN(n12498) );
  NAND2_X1 U15648 ( .A1(n19312), .A2(n19864), .ZN(n12500) );
  NOR2_X1 U15649 ( .A1(n19864), .A2(n19873), .ZN(n19699) );
  NAND2_X1 U15650 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19699), .ZN(
        n15598) );
  NAND2_X1 U15651 ( .A1(n12500), .A2(n15598), .ZN(n19343) );
  NOR2_X1 U15652 ( .A1(n19343), .A2(n15596), .ZN(n12501) );
  AOI21_X1 U15653 ( .B1(n12507), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12501), .ZN(n12502) );
  NAND2_X1 U15654 ( .A1(n12758), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12511) );
  NAND2_X1 U15655 ( .A1(n13072), .A2(n13071), .ZN(n13136) );
  INV_X1 U15656 ( .A(n12504), .ZN(n12505) );
  INV_X1 U15657 ( .A(n19312), .ZN(n16212) );
  NOR2_X1 U15658 ( .A1(n19864), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19402) );
  NAND2_X1 U15659 ( .A1(n16212), .A2(n19402), .ZN(n19471) );
  NAND2_X1 U15660 ( .A1(n15598), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12506) );
  AOI21_X1 U15661 ( .B1(n19471), .B2(n12506), .A(n15596), .ZN(n19582) );
  AOI21_X1 U15662 ( .B1(n12507), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19582), .ZN(n12508) );
  NAND2_X1 U15663 ( .A1(n13134), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12513) );
  INV_X1 U15664 ( .A(n12511), .ZN(n12512) );
  AND3_X1 U15665 ( .A1(n10754), .A2(n15614), .A3(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12514) );
  AND2_X1 U15666 ( .A1(n12758), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13133) );
  AND2_X1 U15667 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12515) );
  INV_X1 U15668 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15654) );
  AND2_X2 U15669 ( .A1(n13204), .A2(n13203), .ZN(n13285) );
  AND2_X1 U15670 ( .A1(n13479), .A2(n13471), .ZN(n12517) );
  NOR2_X2 U15671 ( .A1(n13588), .A2(n13609), .ZN(n13610) );
  NAND2_X1 U15672 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12522) );
  NAND2_X1 U15673 ( .A1(n12570), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12521) );
  NAND2_X1 U15674 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12520) );
  NAND2_X1 U15675 ( .A1(n12572), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12519) );
  NAND4_X1 U15676 ( .A1(n12522), .A2(n12521), .A3(n12520), .A4(n12519), .ZN(
        n12528) );
  AOI22_X1 U15677 ( .A1(n12661), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12526) );
  NAND2_X1 U15678 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12525) );
  NAND2_X1 U15679 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12524) );
  AOI22_X1 U15680 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12523) );
  NAND4_X1 U15681 ( .A1(n12526), .A2(n12525), .A3(n12524), .A4(n12523), .ZN(
        n12527) );
  OR2_X1 U15682 ( .A1(n12528), .A2(n12527), .ZN(n12534) );
  AOI22_X1 U15683 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U15684 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12531) );
  NAND2_X1 U15685 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12530) );
  NAND2_X1 U15686 ( .A1(n12668), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12529) );
  NAND4_X1 U15687 ( .A1(n12532), .A2(n12531), .A3(n12530), .A4(n12529), .ZN(
        n12533) );
  NOR2_X1 U15688 ( .A1(n12534), .A2(n12533), .ZN(n15028) );
  INV_X1 U15689 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12537) );
  OAI22_X1 U15690 ( .A1(n12537), .A2(n12654), .B1(n12653), .B2(n12536), .ZN(
        n12541) );
  OAI22_X1 U15691 ( .A1(n12539), .A2(n15588), .B1(n12656), .B2(n12538), .ZN(
        n12540) );
  NOR2_X1 U15692 ( .A1(n12541), .A2(n12540), .ZN(n12545) );
  AOI22_X1 U15693 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12544) );
  AOI22_X1 U15694 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12661), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15695 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11020), .B1(
        n10902), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12542) );
  NAND4_X1 U15696 ( .A1(n12545), .A2(n12544), .A3(n12543), .A4(n12542), .ZN(
        n12551) );
  AOI22_X1 U15697 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10937), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15698 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12548) );
  NAND2_X1 U15699 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12547) );
  NAND2_X1 U15700 ( .A1(n12668), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12546) );
  NAND4_X1 U15701 ( .A1(n12549), .A2(n12548), .A3(n12547), .A4(n12546), .ZN(
        n12550) );
  OR2_X1 U15702 ( .A1(n12551), .A2(n12550), .ZN(n13758) );
  NAND2_X1 U15703 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12555) );
  NAND2_X1 U15704 ( .A1(n12570), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12554) );
  NAND2_X1 U15705 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12553) );
  NAND2_X1 U15706 ( .A1(n12572), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12552) );
  NAND4_X1 U15707 ( .A1(n12555), .A2(n12554), .A3(n12553), .A4(n12552), .ZN(
        n12561) );
  AOI22_X1 U15708 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12661), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12559) );
  NAND2_X1 U15709 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12558) );
  NAND2_X1 U15710 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12557) );
  AOI22_X1 U15711 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12556) );
  NAND4_X1 U15712 ( .A1(n12559), .A2(n12558), .A3(n12557), .A4(n12556), .ZN(
        n12560) );
  OR2_X1 U15713 ( .A1(n12561), .A2(n12560), .ZN(n12567) );
  AOI22_X1 U15714 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10937), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U15715 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12564) );
  NAND2_X1 U15716 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12563) );
  NAND2_X1 U15717 ( .A1(n12668), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12562) );
  NAND4_X1 U15718 ( .A1(n12565), .A2(n12564), .A3(n12563), .A4(n12562), .ZN(
        n12566) );
  NOR2_X1 U15719 ( .A1(n12567), .A2(n12566), .ZN(n15020) );
  NAND2_X1 U15720 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12576) );
  NAND2_X1 U15721 ( .A1(n12570), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12575) );
  NAND2_X1 U15722 ( .A1(n12571), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12574) );
  NAND2_X1 U15723 ( .A1(n12572), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12573) );
  NAND4_X1 U15724 ( .A1(n12576), .A2(n12575), .A3(n12574), .A4(n12573), .ZN(
        n12582) );
  AOI22_X1 U15725 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12661), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12580) );
  NAND2_X1 U15726 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12579) );
  NAND2_X1 U15727 ( .A1(n10902), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12578) );
  INV_X1 U15728 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n19294) );
  AOI22_X1 U15729 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12577) );
  NAND4_X1 U15730 ( .A1(n12580), .A2(n12579), .A3(n12578), .A4(n12577), .ZN(
        n12581) );
  OR2_X1 U15731 ( .A1(n12582), .A2(n12581), .ZN(n12588) );
  AOI22_X1 U15732 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10937), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15733 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U15734 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12584) );
  NAND2_X1 U15735 ( .A1(n12668), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12583) );
  NAND4_X1 U15736 ( .A1(n12586), .A2(n12585), .A3(n12584), .A4(n12583), .ZN(
        n12587) );
  NOR2_X1 U15737 ( .A1(n12588), .A2(n12587), .ZN(n15011) );
  NOR2_X2 U15738 ( .A1(n15010), .A2(n15011), .ZN(n15002) );
  INV_X1 U15739 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13460) );
  INV_X1 U15740 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12589) );
  OAI22_X1 U15741 ( .A1(n13460), .A2(n12654), .B1(n12653), .B2(n12589), .ZN(
        n12593) );
  INV_X1 U15742 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12591) );
  OAI22_X1 U15743 ( .A1(n12591), .A2(n15588), .B1(n12656), .B2(n12590), .ZN(
        n12592) );
  NOR2_X1 U15744 ( .A1(n12593), .A2(n12592), .ZN(n12597) );
  AOI22_X1 U15745 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15746 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12661), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15747 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11020), .B1(
        n10902), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12594) );
  NAND4_X1 U15748 ( .A1(n12597), .A2(n12596), .A3(n12595), .A4(n12594), .ZN(
        n12603) );
  AOI22_X1 U15749 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10937), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12601) );
  AOI22_X1 U15750 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12600) );
  NAND2_X1 U15751 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12599) );
  NAND2_X1 U15752 ( .A1(n12668), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12598) );
  NAND4_X1 U15753 ( .A1(n12601), .A2(n12600), .A3(n12599), .A4(n12598), .ZN(
        n12602) );
  OR2_X1 U15754 ( .A1(n12603), .A2(n12602), .ZN(n15003) );
  AOI22_X1 U15755 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10902), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U15756 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U15757 ( .A1(n12661), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12604) );
  NAND3_X1 U15758 ( .A1(n12606), .A2(n12605), .A3(n12604), .ZN(n12617) );
  AOI22_X1 U15759 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12668), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U15760 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U15761 ( .A1(n10937), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12607) );
  NAND3_X1 U15762 ( .A1(n12609), .A2(n12608), .A3(n12607), .ZN(n12616) );
  INV_X1 U15763 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12611) );
  INV_X1 U15764 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12610) );
  OAI22_X1 U15765 ( .A1(n12653), .A2(n12611), .B1(n12654), .B2(n12610), .ZN(
        n12615) );
  OAI22_X1 U15766 ( .A1(n15588), .A2(n12613), .B1(n12656), .B2(n12612), .ZN(
        n12614) );
  NOR4_X1 U15767 ( .A1(n12617), .A2(n12616), .A3(n12615), .A4(n12614), .ZN(
        n14995) );
  AOI22_X1 U15768 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11020), .B1(
        n10902), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U15769 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U15770 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10944), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12618) );
  NAND3_X1 U15771 ( .A1(n12620), .A2(n12619), .A3(n12618), .ZN(n12627) );
  INV_X1 U15772 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12622) );
  INV_X1 U15773 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12621) );
  OAI22_X1 U15774 ( .A1(n12622), .A2(n12654), .B1(n12653), .B2(n12621), .ZN(
        n12626) );
  INV_X1 U15775 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12624) );
  INV_X1 U15776 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12623) );
  OAI22_X1 U15777 ( .A1(n12624), .A2(n15588), .B1(n12656), .B2(n12623), .ZN(
        n12625) );
  NOR3_X1 U15778 ( .A1(n12627), .A2(n12626), .A3(n12625), .ZN(n12631) );
  AOI22_X1 U15779 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12668), .B1(
        n12667), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U15780 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15781 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10937), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12628) );
  NAND4_X1 U15782 ( .A1(n12631), .A2(n12630), .A3(n12629), .A4(n12628), .ZN(
        n14988) );
  AOI22_X1 U15783 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12643) );
  AOI22_X1 U15784 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12780), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12642) );
  AND2_X1 U15785 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12634) );
  OR2_X1 U15786 ( .A1(n12634), .A2(n12633), .ZN(n14313) );
  INV_X1 U15787 ( .A(n14313), .ZN(n12783) );
  NAND2_X1 U15788 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12638) );
  NAND2_X1 U15789 ( .A1(n10878), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12637) );
  AND3_X1 U15790 ( .A1(n12783), .A2(n12638), .A3(n12637), .ZN(n12641) );
  AOI22_X1 U15791 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12640) );
  NAND4_X1 U15792 ( .A1(n12643), .A2(n12642), .A3(n12641), .A4(n12640), .ZN(
        n12651) );
  AOI22_X1 U15793 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U15794 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12780), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U15795 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12647) );
  NAND2_X1 U15796 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12645) );
  NAND2_X1 U15797 ( .A1(n10878), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12644) );
  AND3_X1 U15798 ( .A1(n12645), .A2(n12644), .A3(n14313), .ZN(n12646) );
  NAND4_X1 U15799 ( .A1(n12649), .A2(n12648), .A3(n12647), .A4(n12646), .ZN(
        n12650) );
  AND2_X1 U15800 ( .A1(n12651), .A2(n12650), .ZN(n12698) );
  AND2_X1 U15801 ( .A1(n15614), .A2(n12698), .ZN(n12675) );
  INV_X1 U15802 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12655) );
  INV_X1 U15803 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12652) );
  OAI22_X1 U15804 ( .A1(n12655), .A2(n12654), .B1(n12653), .B2(n12652), .ZN(
        n12659) );
  INV_X1 U15805 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12657) );
  INV_X1 U15806 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14309) );
  OAI22_X1 U15807 ( .A1(n12657), .A2(n12656), .B1(n15588), .B2(n14309), .ZN(
        n12658) );
  NOR2_X1 U15808 ( .A1(n12659), .A2(n12658), .ZN(n12665) );
  AOI22_X1 U15809 ( .A1(n10857), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U15810 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10944), .B1(
        n12661), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U15811 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11020), .B1(
        n10902), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12662) );
  NAND4_X1 U15812 ( .A1(n12665), .A2(n12664), .A3(n12663), .A4(n12662), .ZN(
        n12674) );
  AOI22_X1 U15813 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10937), .B1(
        n10918), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U15814 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12671) );
  NAND2_X1 U15815 ( .A1(n12667), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12670) );
  NAND2_X1 U15816 ( .A1(n12668), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12669) );
  NAND4_X1 U15817 ( .A1(n12672), .A2(n12671), .A3(n12670), .A4(n12669), .ZN(
        n12673) );
  OR2_X1 U15818 ( .A1(n12674), .A2(n12673), .ZN(n12693) );
  INV_X1 U15819 ( .A(n12698), .ZN(n12676) );
  NOR2_X1 U15820 ( .A1(n15614), .A2(n12676), .ZN(n14982) );
  NAND2_X1 U15821 ( .A1(n10225), .A2(n10333), .ZN(n12678) );
  NAND2_X1 U15822 ( .A1(n14981), .A2(n12678), .ZN(n14971) );
  AOI22_X1 U15823 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U15824 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10878), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12683) );
  NAND2_X1 U15825 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12680) );
  NAND2_X1 U15826 ( .A1(n12780), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12679) );
  AND3_X1 U15827 ( .A1(n12783), .A2(n12680), .A3(n12679), .ZN(n12682) );
  AOI22_X1 U15828 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12681) );
  NAND4_X1 U15829 ( .A1(n12684), .A2(n12683), .A3(n12682), .A4(n12681), .ZN(
        n12692) );
  AOI22_X1 U15830 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12690) );
  AOI22_X1 U15831 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10878), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U15832 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12688) );
  NAND2_X1 U15833 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12686) );
  NAND2_X1 U15834 ( .A1(n12780), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12685) );
  AND3_X1 U15835 ( .A1(n12686), .A2(n14313), .A3(n12685), .ZN(n12687) );
  NAND4_X1 U15836 ( .A1(n12690), .A2(n12689), .A3(n12688), .A4(n12687), .ZN(
        n12691) );
  AND2_X1 U15837 ( .A1(n12692), .A2(n12691), .ZN(n12694) );
  INV_X1 U15838 ( .A(n12694), .ZN(n12697) );
  AND2_X1 U15839 ( .A1(n12693), .A2(n12698), .ZN(n12695) );
  INV_X1 U15840 ( .A(n12695), .ZN(n12696) );
  AND2_X1 U15841 ( .A1(n12695), .A2(n12694), .ZN(n12714) );
  INV_X1 U15842 ( .A(n12758), .ZN(n13164) );
  AOI211_X1 U15843 ( .C1(n12697), .C2(n12696), .A(n12714), .B(n13164), .ZN(
        n14972) );
  NAND2_X1 U15844 ( .A1(n14971), .A2(n14972), .ZN(n14970) );
  NOR2_X1 U15845 ( .A1(n15614), .A2(n12697), .ZN(n14974) );
  NAND2_X1 U15846 ( .A1(n10333), .A2(n10350), .ZN(n12699) );
  NAND2_X1 U15847 ( .A1(n14970), .A2(n12699), .ZN(n12717) );
  AOI22_X1 U15848 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15849 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10878), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12704) );
  NAND2_X1 U15850 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12701) );
  NAND2_X1 U15851 ( .A1(n12780), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12700) );
  AND3_X1 U15852 ( .A1(n12783), .A2(n12701), .A3(n12700), .ZN(n12703) );
  AOI22_X1 U15853 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12702) );
  NAND4_X1 U15854 ( .A1(n12705), .A2(n12704), .A3(n12703), .A4(n12702), .ZN(
        n12713) );
  AOI22_X1 U15855 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15856 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10878), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12710) );
  AOI22_X1 U15857 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12709) );
  NAND2_X1 U15858 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12707) );
  NAND2_X1 U15859 ( .A1(n12780), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12706) );
  AND3_X1 U15860 ( .A1(n12707), .A2(n14313), .A3(n12706), .ZN(n12708) );
  NAND4_X1 U15861 ( .A1(n12711), .A2(n12710), .A3(n12709), .A4(n12708), .ZN(
        n12712) );
  AND2_X1 U15862 ( .A1(n12713), .A2(n12712), .ZN(n12715) );
  NAND2_X1 U15863 ( .A1(n12714), .A2(n12715), .ZN(n12736) );
  OAI211_X1 U15864 ( .C1(n12714), .C2(n12715), .A(n12758), .B(n12736), .ZN(
        n12718) );
  INV_X1 U15865 ( .A(n12715), .ZN(n12716) );
  NOR2_X1 U15866 ( .A1(n15614), .A2(n12716), .ZN(n14964) );
  INV_X1 U15867 ( .A(n12717), .ZN(n12719) );
  INV_X1 U15868 ( .A(n12736), .ZN(n12737) );
  AOI22_X1 U15869 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U15870 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10878), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12725) );
  NAND2_X1 U15871 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12722) );
  NAND2_X1 U15872 ( .A1(n12780), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12721) );
  AND3_X1 U15873 ( .A1(n12783), .A2(n12722), .A3(n12721), .ZN(n12724) );
  AOI22_X1 U15874 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12723) );
  NAND4_X1 U15875 ( .A1(n12726), .A2(n12725), .A3(n12724), .A4(n12723), .ZN(
        n12734) );
  AOI22_X1 U15876 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U15877 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10878), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12731) );
  AOI22_X1 U15878 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12730) );
  NAND2_X1 U15879 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12728) );
  NAND2_X1 U15880 ( .A1(n12780), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12727) );
  AND3_X1 U15881 ( .A1(n12728), .A2(n14313), .A3(n12727), .ZN(n12729) );
  NAND4_X1 U15882 ( .A1(n12732), .A2(n12731), .A3(n12730), .A4(n12729), .ZN(
        n12733) );
  NAND2_X1 U15883 ( .A1(n12734), .A2(n12733), .ZN(n12735) );
  INV_X1 U15884 ( .A(n12735), .ZN(n12739) );
  OR2_X1 U15885 ( .A1(n12736), .A2(n12735), .ZN(n12743) );
  OAI211_X1 U15886 ( .C1(n12737), .C2(n12739), .A(n12758), .B(n12743), .ZN(
        n12741) );
  INV_X1 U15887 ( .A(n12741), .ZN(n12738) );
  NAND2_X1 U15888 ( .A1(n19903), .A2(n12739), .ZN(n14958) );
  NOR2_X2 U15889 ( .A1(n14959), .A2(n14958), .ZN(n14957) );
  INV_X1 U15890 ( .A(n12743), .ZN(n12759) );
  AOI22_X1 U15891 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U15892 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10878), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12748) );
  NAND2_X1 U15893 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12745) );
  NAND2_X1 U15894 ( .A1(n12780), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12744) );
  AND3_X1 U15895 ( .A1(n12783), .A2(n12745), .A3(n12744), .ZN(n12747) );
  AOI22_X1 U15896 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12746) );
  NAND4_X1 U15897 ( .A1(n12749), .A2(n12748), .A3(n12747), .A4(n12746), .ZN(
        n12757) );
  AOI22_X1 U15898 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15899 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10878), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U15900 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12753) );
  NAND2_X1 U15901 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12751) );
  NAND2_X1 U15902 ( .A1(n12780), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12750) );
  AND3_X1 U15903 ( .A1(n12751), .A2(n14313), .A3(n12750), .ZN(n12752) );
  NAND4_X1 U15904 ( .A1(n12755), .A2(n12754), .A3(n12753), .A4(n12752), .ZN(
        n12756) );
  AND2_X1 U15905 ( .A1(n12757), .A2(n12756), .ZN(n12761) );
  NAND2_X1 U15906 ( .A1(n12759), .A2(n12761), .ZN(n14944) );
  OAI211_X1 U15907 ( .C1(n12759), .C2(n12761), .A(n12758), .B(n14944), .ZN(
        n12760) );
  INV_X1 U15908 ( .A(n12761), .ZN(n12762) );
  NOR2_X1 U15909 ( .A1(n15614), .A2(n12762), .ZN(n14951) );
  INV_X1 U15910 ( .A(n12763), .ZN(n14945) );
  AOI22_X1 U15911 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U15912 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10878), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12768) );
  NAND2_X1 U15913 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12765) );
  NAND2_X1 U15914 ( .A1(n12780), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12764) );
  AND3_X1 U15915 ( .A1(n12783), .A2(n12765), .A3(n12764), .ZN(n12767) );
  AOI22_X1 U15916 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12766) );
  NAND4_X1 U15917 ( .A1(n12769), .A2(n12768), .A3(n12767), .A4(n12766), .ZN(
        n12777) );
  AOI22_X1 U15918 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12775) );
  AOI22_X1 U15919 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10878), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U15920 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12773) );
  NAND2_X1 U15921 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12771) );
  NAND2_X1 U15922 ( .A1(n12780), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12770) );
  AND3_X1 U15923 ( .A1(n12771), .A2(n14313), .A3(n12770), .ZN(n12772) );
  NAND4_X1 U15924 ( .A1(n12775), .A2(n12774), .A3(n12773), .A4(n12772), .ZN(
        n12776) );
  NAND2_X1 U15925 ( .A1(n12777), .A2(n12776), .ZN(n14947) );
  INV_X1 U15926 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n21029) );
  INV_X1 U15927 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12778) );
  OAI22_X1 U15928 ( .A1(n21029), .A2(n10869), .B1(n10853), .B2(n12778), .ZN(
        n12779) );
  INV_X1 U15929 ( .A(n12779), .ZN(n12787) );
  AOI22_X1 U15930 ( .A1(n14310), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12780), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12786) );
  NAND2_X1 U15931 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12782) );
  NAND2_X1 U15932 ( .A1(n10878), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12781) );
  AND3_X1 U15933 ( .A1(n12783), .A2(n12782), .A3(n12781), .ZN(n12785) );
  AOI22_X1 U15934 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12784) );
  NAND4_X1 U15935 ( .A1(n12787), .A2(n12786), .A3(n12785), .A4(n12784), .ZN(
        n12795) );
  AOI22_X1 U15936 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12793) );
  AOI22_X1 U15937 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12780), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U15938 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12791) );
  NAND2_X1 U15939 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12789) );
  NAND2_X1 U15940 ( .A1(n10878), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12788) );
  AND3_X1 U15941 ( .A1(n12789), .A2(n12788), .A3(n14313), .ZN(n12790) );
  NAND4_X1 U15942 ( .A1(n12793), .A2(n12792), .A3(n12791), .A4(n12790), .ZN(
        n12794) );
  NAND2_X1 U15943 ( .A1(n12795), .A2(n12794), .ZN(n12797) );
  OR3_X1 U15944 ( .A1(n14944), .A2(n19903), .A3(n14947), .ZN(n12796) );
  NOR2_X1 U15945 ( .A1(n12796), .A2(n12797), .ZN(n14303) );
  AOI21_X1 U15946 ( .B1(n12797), .B2(n12796), .A(n14303), .ZN(n12798) );
  NOR2_X1 U15947 ( .A1(n12799), .A2(n12798), .ZN(n12831) );
  INV_X1 U15948 ( .A(n13530), .ZN(n16229) );
  NAND2_X1 U15949 ( .A1(n16229), .A2(n12826), .ZN(n13027) );
  NAND2_X1 U15950 ( .A1(n13027), .A2(n12800), .ZN(n12801) );
  NAND2_X1 U15951 ( .A1(n12801), .A2(n13032), .ZN(n12803) );
  AND2_X1 U15952 ( .A1(n11731), .A2(n19901), .ZN(n13024) );
  NAND2_X1 U15953 ( .A1(n19895), .A2(n13024), .ZN(n12802) );
  NAND2_X1 U15954 ( .A1(n19121), .A2(n12804), .ZN(n19093) );
  NAND2_X1 U15955 ( .A1(n19121), .A2(n12830), .ZN(n19092) );
  AND2_X1 U15956 ( .A1(n19121), .A2(n9882), .ZN(n13035) );
  NOR4_X1 U15957 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12810) );
  NOR4_X1 U15958 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12809) );
  NOR4_X1 U15959 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12808) );
  NOR4_X1 U15960 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12807) );
  NAND4_X1 U15961 ( .A1(n12810), .A2(n12809), .A3(n12808), .A4(n12807), .ZN(
        n12815) );
  NOR4_X1 U15962 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12813) );
  NOR4_X1 U15963 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12812) );
  NOR4_X1 U15964 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n12811) );
  INV_X1 U15965 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19790) );
  NAND4_X1 U15966 ( .A1(n12813), .A2(n12812), .A3(n12811), .A4(n19790), .ZN(
        n12814) );
  OAI21_X1 U15967 ( .B1(n12815), .B2(n12814), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12816) );
  INV_X1 U15968 ( .A(n19088), .ZN(n15082) );
  INV_X1 U15969 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14535) );
  OR2_X1 U15970 ( .A1(n19100), .A2(n14535), .ZN(n12819) );
  NAND2_X1 U15971 ( .A1(n19100), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12818) );
  AND2_X1 U15972 ( .A1(n12819), .A2(n12818), .ZN(n19230) );
  INV_X1 U15973 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19145) );
  OAI22_X1 U15974 ( .A1(n15082), .A2(n19230), .B1(n19121), .B2(n19145), .ZN(
        n12822) );
  INV_X1 U15975 ( .A(n19090), .ZN(n15054) );
  INV_X1 U15976 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n12820) );
  NOR2_X1 U15977 ( .A1(n15054), .A2(n12820), .ZN(n12821) );
  AOI211_X1 U15978 ( .C1(BUF1_REG_29__SCAN_IN), .C2(n19089), .A(n12822), .B(
        n12821), .ZN(n12823) );
  INV_X1 U15979 ( .A(n12824), .ZN(n12825) );
  INV_X1 U15980 ( .A(n12826), .ZN(n16230) );
  INV_X1 U15981 ( .A(n16227), .ZN(n12827) );
  NAND2_X1 U15982 ( .A1(n16230), .A2(n12827), .ZN(n13026) );
  NAND2_X1 U15983 ( .A1(n13026), .A2(n12828), .ZN(n12829) );
  INV_X2 U15984 ( .A(n15036), .ZN(n14984) );
  INV_X1 U15985 ( .A(n12832), .ZN(n12833) );
  OAI21_X1 U15986 ( .B1(n12835), .B2(n12834), .A(n12833), .ZN(n16024) );
  NAND2_X1 U15987 ( .A1(n14984), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12836) );
  OR2_X1 U15988 ( .A1(n12839), .A2(n16145), .ZN(n12848) );
  NOR2_X1 U15989 ( .A1(n14329), .A2(n16130), .ZN(n12844) );
  XNOR2_X1 U15990 ( .A(n12840), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16012) );
  NAND2_X1 U15991 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12841) );
  OAI211_X1 U15992 ( .C1(n19247), .C2(n16012), .A(n12842), .B(n12841), .ZN(
        n12843) );
  NAND3_X1 U15993 ( .A1(n12848), .A2(n12847), .A3(n12846), .ZN(P2_U2984) );
  INV_X1 U15994 ( .A(n12870), .ZN(n12868) );
  OAI21_X1 U15995 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12851), .A(
        n12868), .ZN(n15203) );
  INV_X1 U15996 ( .A(n15203), .ZN(n18859) );
  AOI21_X1 U15997 ( .B1(n21083), .B2(n12852), .A(n12853), .ZN(n18920) );
  AOI21_X1 U15998 ( .B1(n10216), .B2(n9903), .A(n12854), .ZN(n18941) );
  NOR2_X1 U15999 ( .A1(n12855), .A2(n16106), .ZN(n12864) );
  AOI21_X1 U16000 ( .B1(n16106), .B2(n12855), .A(n12864), .ZN(n18960) );
  AOI21_X1 U16001 ( .B1(n15264), .B2(n12856), .A(n12857), .ZN(n18981) );
  AOI21_X1 U16002 ( .B1(n15276), .B2(n12858), .A(n12859), .ZN(n18997) );
  AOI21_X1 U16003 ( .B1(n19019), .B2(n12860), .A(n12861), .ZN(n19026) );
  INV_X1 U16004 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13576) );
  NOR2_X1 U16005 ( .A1(n13576), .A2(n12862), .ZN(n12863) );
  AOI21_X1 U16006 ( .B1(n13576), .B2(n12862), .A(n12863), .ZN(n13578) );
  OAI22_X1 U16007 ( .A1(n19904), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19084) );
  INV_X1 U16008 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19057) );
  OAI22_X1 U16009 ( .A1(n19904), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19057), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13537) );
  AND2_X1 U16010 ( .A1(n19084), .A2(n13537), .ZN(n13498) );
  OAI21_X1 U16011 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12862), .ZN(n14352) );
  NAND2_X1 U16012 ( .A1(n13498), .A2(n14352), .ZN(n13420) );
  NOR2_X1 U16013 ( .A1(n13578), .A2(n13420), .ZN(n19040) );
  OAI21_X1 U16014 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12863), .A(
        n12860), .ZN(n19246) );
  NAND2_X1 U16015 ( .A1(n19040), .A2(n19246), .ZN(n19023) );
  NOR2_X1 U16016 ( .A1(n19026), .A2(n19023), .ZN(n19012) );
  OAI21_X1 U16017 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12861), .A(
        n12858), .ZN(n19013) );
  NAND2_X1 U16018 ( .A1(n19012), .A2(n19013), .ZN(n18996) );
  NOR2_X1 U16019 ( .A1(n18997), .A2(n18996), .ZN(n18989) );
  OAI21_X1 U16020 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12859), .A(
        n12856), .ZN(n18990) );
  NAND2_X1 U16021 ( .A1(n18989), .A2(n18990), .ZN(n18979) );
  NOR2_X1 U16022 ( .A1(n18981), .A2(n18979), .ZN(n18965) );
  OAI21_X1 U16023 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12857), .A(
        n12855), .ZN(n18967) );
  NAND2_X1 U16024 ( .A1(n18965), .A2(n18967), .ZN(n18958) );
  NOR2_X1 U16025 ( .A1(n18960), .A2(n18958), .ZN(n18944) );
  OAI21_X1 U16026 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12864), .A(
        n9903), .ZN(n18945) );
  NAND2_X1 U16027 ( .A1(n18944), .A2(n18945), .ZN(n18934) );
  NOR2_X1 U16028 ( .A1(n18941), .A2(n18934), .ZN(n18933) );
  OAI21_X1 U16029 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12854), .A(
        n12852), .ZN(n18927) );
  NAND2_X1 U16030 ( .A1(n18933), .A2(n18927), .ZN(n18919) );
  NOR2_X1 U16031 ( .A1(n18920), .A2(n18919), .ZN(n18918) );
  OAI21_X1 U16032 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12853), .A(
        n9840), .ZN(n12865) );
  INV_X1 U16033 ( .A(n12865), .ZN(n18904) );
  NOR2_X1 U16034 ( .A1(n18903), .A2(n18904), .ZN(n18902) );
  NOR2_X1 U16035 ( .A1(n19041), .A2(n18902), .ZN(n18891) );
  AOI21_X1 U16036 ( .B1(n9840), .B2(n15234), .A(n12866), .ZN(n18892) );
  NOR2_X1 U16037 ( .A1(n18891), .A2(n18892), .ZN(n18890) );
  OAI21_X1 U16038 ( .B1(n12866), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n12867), .ZN(n15227) );
  INV_X1 U16039 ( .A(n15227), .ZN(n18880) );
  AOI21_X1 U16040 ( .B1(n15214), .B2(n12867), .A(n12851), .ZN(n18869) );
  NOR2_X1 U16041 ( .A1(n18867), .A2(n19041), .ZN(n18857) );
  NOR2_X1 U16042 ( .A1(n18859), .A2(n18857), .ZN(n18858) );
  NOR2_X1 U16043 ( .A1(n19041), .A2(n18858), .ZN(n12918) );
  INV_X1 U16044 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15189) );
  AND2_X1 U16045 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12870), .ZN(
        n12871) );
  AOI21_X1 U16046 ( .B1(n12868), .B2(n15189), .A(n12871), .ZN(n15191) );
  NOR2_X1 U16047 ( .A1(n12918), .A2(n15191), .ZN(n12919) );
  NOR2_X1 U16048 ( .A1(n19041), .A2(n12919), .ZN(n15679) );
  NAND2_X1 U16049 ( .A1(n12870), .A2(n12869), .ZN(n12873) );
  OAI21_X1 U16050 ( .B1(n12871), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n12873), .ZN(n15168) );
  INV_X1 U16051 ( .A(n15168), .ZN(n15681) );
  INV_X1 U16052 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15160) );
  AOI21_X1 U16053 ( .B1(n15160), .B2(n12873), .A(n12872), .ZN(n15163) );
  OR2_X1 U16054 ( .A1(n12872), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12875) );
  NAND2_X1 U16055 ( .A1(n12874), .A2(n12875), .ZN(n15154) );
  INV_X1 U16056 ( .A(n15154), .ZN(n16053) );
  NOR2_X1 U16057 ( .A1(n16051), .A2(n16053), .ZN(n16052) );
  INV_X1 U16058 ( .A(n12876), .ZN(n12877) );
  AOI21_X1 U16059 ( .B1(n15145), .B2(n12874), .A(n12877), .ZN(n16037) );
  OR2_X1 U16060 ( .A1(n12876), .A2(n12878), .ZN(n12880) );
  NAND2_X1 U16061 ( .A1(n12876), .A2(n12878), .ZN(n12879) );
  NAND2_X1 U16062 ( .A1(n12880), .A2(n12879), .ZN(n15134) );
  INV_X1 U16063 ( .A(n15134), .ZN(n16027) );
  NOR2_X1 U16064 ( .A1(n19041), .A2(n16026), .ZN(n12945) );
  AND2_X1 U16065 ( .A1(n12880), .A2(n15122), .ZN(n12881) );
  NOR2_X1 U16066 ( .A1(n12445), .A2(n12881), .ZN(n15120) );
  NOR2_X1 U16067 ( .A1(n12945), .A2(n15120), .ZN(n12944) );
  NOR2_X1 U16068 ( .A1(n12882), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12883) );
  OR2_X1 U16069 ( .A1(n12840), .A2(n12883), .ZN(n15110) );
  INV_X1 U16070 ( .A(n15110), .ZN(n16016) );
  NOR2_X1 U16071 ( .A1(n19041), .A2(n16011), .ZN(n12884) );
  XNOR2_X1 U16072 ( .A(n12884), .B(n16012), .ZN(n12885) );
  NAND4_X1 U16073 ( .A1(n19654), .A2(n19904), .A3(n19902), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19061) );
  INV_X1 U16074 ( .A(n19061), .ZN(n19764) );
  NAND2_X1 U16075 ( .A1(n12885), .A2(n19764), .ZN(n12902) );
  NOR2_X1 U16076 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n12886), .ZN(n16249) );
  AND2_X1 U16077 ( .A1(n15614), .A2(n19901), .ZN(n12887) );
  INV_X1 U16078 ( .A(n16249), .ZN(n16006) );
  NAND2_X1 U16079 ( .A1(n19231), .A2(n16006), .ZN(n12890) );
  NAND2_X1 U16080 ( .A1(n19902), .A2(n19901), .ZN(n12888) );
  AND2_X1 U16081 ( .A1(n12973), .A2(n12888), .ZN(n12892) );
  INV_X1 U16082 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n20980) );
  NAND2_X1 U16083 ( .A1(n12892), .A2(n20980), .ZN(n12889) );
  AND2_X1 U16084 ( .A1(n15614), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12891) );
  NAND2_X1 U16085 ( .A1(n12892), .A2(n12891), .ZN(n19070) );
  NAND2_X1 U16086 ( .A1(n19061), .A2(n19034), .ZN(n12893) );
  NAND2_X1 U16087 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19654), .ZN(n19762) );
  NOR3_X1 U16088 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19469), .A3(n19762), 
        .ZN(n16247) );
  OR2_X1 U16089 ( .A1(n12893), .A2(n16247), .ZN(n12894) );
  NAND2_X1 U16090 ( .A1(n19069), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19035) );
  AOI22_X1 U16091 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19080), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19049), .ZN(n12895) );
  OAI21_X1 U16092 ( .B1(n12896), .B2(n19070), .A(n12895), .ZN(n12897) );
  AOI21_X1 U16093 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19063), .A(n12897), .ZN(
        n12898) );
  NAND2_X1 U16094 ( .A1(n12902), .A2(n12901), .ZN(P2_U2825) );
  NOR4_X1 U16095 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n12906) );
  NOR4_X1 U16096 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12905) );
  NOR4_X1 U16097 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n12904) );
  NOR4_X1 U16098 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_11__SCAN_IN), .A3(P1_ADDRESS_REG_10__SCAN_IN), .A4(
        P1_ADDRESS_REG_9__SCAN_IN), .ZN(n12903) );
  AND4_X1 U16099 ( .A1(n12906), .A2(n12905), .A3(n12904), .A4(n12903), .ZN(
        n12911) );
  NOR4_X1 U16100 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12909) );
  NOR4_X1 U16101 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12908) );
  NOR4_X1 U16102 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_3__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12907) );
  INV_X1 U16103 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20745) );
  AND4_X1 U16104 ( .A1(n12909), .A2(n12908), .A3(n12907), .A4(n20745), .ZN(
        n12910) );
  NAND2_X1 U16105 ( .A1(n12911), .A2(n12910), .ZN(n12912) );
  INV_X1 U16106 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21065) );
  NOR3_X1 U16107 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21065), .ZN(n12914) );
  NOR4_X1 U16108 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12913) );
  NAND4_X1 U16109 ( .A1(n20145), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n12914), .A4(
        n12913), .ZN(U214) );
  NOR2_X1 U16110 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12916) );
  NOR4_X1 U16111 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12915) );
  NAND4_X1 U16112 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12916), .A4(n12915), .ZN(n12917) );
  NOR2_X1 U16113 ( .A1(n19100), .A2(n12917), .ZN(n16332) );
  NAND2_X1 U16114 ( .A1(n16332), .A2(U214), .ZN(U212) );
  NOR2_X1 U16115 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12917), .ZN(n16390)
         );
  AOI211_X1 U16116 ( .C1(n15191), .C2(n12918), .A(n12919), .B(n19061), .ZN(
        n12932) );
  OAI22_X1 U16117 ( .A1(n15189), .A2(n19035), .B1(n19814), .B2(n19069), .ZN(
        n12931) );
  INV_X1 U16118 ( .A(n19063), .ZN(n19008) );
  INV_X1 U16119 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12920) );
  OAI22_X1 U16120 ( .A1(n12921), .A2(n19070), .B1(n19008), .B2(n12920), .ZN(
        n12930) );
  AND2_X1 U16121 ( .A1(n14999), .A2(n12922), .ZN(n12923) );
  OR2_X1 U16122 ( .A1(n12923), .A2(n14990), .ZN(n15387) );
  INV_X1 U16123 ( .A(n15387), .ZN(n12927) );
  NAND2_X1 U16124 ( .A1(n12924), .A2(n12925), .ZN(n12926) );
  AND2_X1 U16125 ( .A1(n15368), .A2(n12926), .ZN(n15380) );
  AOI22_X1 U16126 ( .A1(n12927), .A2(n19062), .B1(n15380), .B2(n19064), .ZN(
        n12928) );
  INV_X1 U16127 ( .A(n12928), .ZN(n12929) );
  OR4_X1 U16128 ( .A1(n12932), .A2(n12931), .A3(n12930), .A4(n12929), .ZN(
        P2_U2834) );
  AOI211_X1 U16129 ( .C1(n15163), .C2(n12933), .A(n10189), .B(n19061), .ZN(
        n12943) );
  OAI22_X1 U16130 ( .A1(n12934), .A2(n19070), .B1(n19818), .B2(n19069), .ZN(
        n12942) );
  INV_X1 U16131 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n14985) );
  OAI22_X1 U16132 ( .A1(n19008), .A2(n14985), .B1(n15160), .B2(n19035), .ZN(
        n12941) );
  INV_X1 U16133 ( .A(n12935), .ZN(n12936) );
  OAI21_X1 U16134 ( .B1(n9899), .B2(n12936), .A(n14977), .ZN(n15352) );
  OR2_X1 U16135 ( .A1(n15367), .A2(n12938), .ZN(n12939) );
  NAND2_X1 U16136 ( .A1(n12937), .A2(n12939), .ZN(n15355) );
  OAI22_X1 U16137 ( .A1(n15352), .A2(n19047), .B1(n15355), .B2(n19053), .ZN(
        n12940) );
  OR4_X1 U16138 ( .A1(n12943), .A2(n12942), .A3(n12941), .A4(n12940), .ZN(
        P2_U2832) );
  AOI211_X1 U16139 ( .C1(n15120), .C2(n12945), .A(n12944), .B(n19061), .ZN(
        n12958) );
  OAI22_X1 U16140 ( .A1(n12946), .A2(n19070), .B1(n19827), .B2(n19069), .ZN(
        n12957) );
  AOI22_X1 U16141 ( .A1(n19063), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19080), .ZN(n12947) );
  INV_X1 U16142 ( .A(n12947), .ZN(n12956) );
  NAND2_X1 U16143 ( .A1(n12948), .A2(n12949), .ZN(n12950) );
  NAND2_X1 U16144 ( .A1(n12951), .A2(n12950), .ZN(n15119) );
  OR2_X1 U16145 ( .A1(n15062), .A2(n12953), .ZN(n12954) );
  NAND2_X1 U16146 ( .A1(n12952), .A2(n12954), .ZN(n15314) );
  OAI22_X1 U16147 ( .A1(n15119), .A2(n19047), .B1(n15314), .B2(n19053), .ZN(
        n12955) );
  OR4_X1 U16148 ( .A1(n12958), .A2(n12957), .A3(n12956), .A4(n12955), .ZN(
        P2_U2828) );
  AOI211_X1 U16149 ( .C1(n12961), .C2(n12959), .A(n12960), .B(n19061), .ZN(
        n12969) );
  OAI22_X1 U16150 ( .A1(n12962), .A2(n19070), .B1(n19035), .B2(n12448), .ZN(
        n12968) );
  AOI22_X1 U16151 ( .A1(n19063), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19049), .ZN(n12963) );
  INV_X1 U16152 ( .A(n12963), .ZN(n12967) );
  NAND2_X1 U16153 ( .A1(n12952), .A2(n12964), .ZN(n12965) );
  NAND2_X1 U16154 ( .A1(n9883), .A2(n12965), .ZN(n15301) );
  OAI22_X1 U16155 ( .A1(n15296), .A2(n19047), .B1(n15301), .B2(n19053), .ZN(
        n12966) );
  OR4_X1 U16156 ( .A1(n12969), .A2(n12968), .A3(n12967), .A4(n12966), .ZN(
        P2_U2827) );
  INV_X1 U16157 ( .A(n12970), .ZN(n12971) );
  OR2_X1 U16158 ( .A1(n19135), .A2(n12971), .ZN(n13510) );
  INV_X1 U16159 ( .A(n13510), .ZN(n19077) );
  INV_X1 U16160 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12975) );
  INV_X1 U16161 ( .A(n12972), .ZN(n18832) );
  INV_X1 U16162 ( .A(n12973), .ZN(n12974) );
  OAI211_X1 U16163 ( .C1(n19077), .C2(n12975), .A(n18832), .B(n12974), .ZN(
        P2_U2814) );
  NOR2_X1 U16164 ( .A1(n19895), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n12977)
         );
  AOI22_X1 U16165 ( .A1(n12977), .A2(n18832), .B1(n12976), .B2(n19895), .ZN(
        P2_U3612) );
  INV_X1 U16166 ( .A(n13025), .ZN(n12979) );
  NOR3_X1 U16167 ( .A1(n12979), .A2(n13024), .A3(n12978), .ZN(n16235) );
  NOR2_X1 U16168 ( .A1(n16235), .A2(n19134), .ZN(n19892) );
  OAI21_X1 U16169 ( .B1(n19892), .B2(n15736), .A(n12980), .ZN(P2_U2819) );
  INV_X1 U16170 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n12981) );
  OR2_X1 U16171 ( .A1(n19205), .A2(n19231), .ZN(n12998) );
  INV_X1 U16172 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n21118) );
  INV_X1 U16173 ( .A(n19205), .ZN(n19234) );
  OAI22_X1 U16174 ( .A1(n19100), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19101), .ZN(n19220) );
  OAI222_X1 U16175 ( .A1(n12981), .A2(n12998), .B1(n19136), .B2(n21118), .C1(
        n19234), .C2(n19220), .ZN(P2_U2958) );
  INV_X1 U16176 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19194) );
  NAND2_X1 U16177 ( .A1(n19232), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n12982) );
  INV_X1 U16178 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16363) );
  INV_X1 U16179 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18189) );
  AOI22_X1 U16180 ( .A1(n19101), .A2(n16363), .B1(n18189), .B2(n19100), .ZN(
        n16066) );
  NAND2_X1 U16181 ( .A1(n19205), .A2(n16066), .ZN(n12994) );
  OAI211_X1 U16182 ( .C1(n19194), .C2(n19136), .A(n12982), .B(n12994), .ZN(
        P2_U2971) );
  INV_X1 U16183 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19198) );
  NAND2_X1 U16184 ( .A1(n19232), .A2(P2_LWORD_REG_2__SCAN_IN), .ZN(n12983) );
  INV_X1 U16185 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16366) );
  INV_X1 U16186 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18180) );
  AOI22_X1 U16187 ( .A1(n19101), .A2(n16366), .B1(n18180), .B2(n19100), .ZN(
        n16071) );
  NAND2_X1 U16188 ( .A1(n19205), .A2(n16071), .ZN(n12990) );
  OAI211_X1 U16189 ( .C1(n19198), .C2(n19136), .A(n12983), .B(n12990), .ZN(
        P2_U2969) );
  INV_X1 U16190 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19151) );
  NAND2_X1 U16191 ( .A1(n19232), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12986) );
  NAND2_X1 U16192 ( .A1(n19100), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12985) );
  INV_X1 U16193 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16354) );
  OR2_X1 U16194 ( .A1(n19100), .A2(n16354), .ZN(n12984) );
  NAND2_X1 U16195 ( .A1(n12985), .A2(n12984), .ZN(n19111) );
  NAND2_X1 U16196 ( .A1(n19205), .A2(n19111), .ZN(n12996) );
  OAI211_X1 U16197 ( .C1(n19151), .C2(n19136), .A(n12986), .B(n12996), .ZN(
        P2_U2962) );
  INV_X1 U16198 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12988) );
  NAND2_X1 U16199 ( .A1(n19232), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12987) );
  MUX2_X1 U16200 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n19100), .Z(n19104) );
  NAND2_X1 U16201 ( .A1(n19205), .A2(n19104), .ZN(n12992) );
  OAI211_X1 U16202 ( .C1(n12988), .C2(n19136), .A(n12987), .B(n12992), .ZN(
        P2_U2966) );
  INV_X1 U16203 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19155) );
  NAND2_X1 U16204 ( .A1(n19232), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12989) );
  MUX2_X1 U16205 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n19100), .Z(n19116) );
  NAND2_X1 U16206 ( .A1(n19205), .A2(n19116), .ZN(n12999) );
  OAI211_X1 U16207 ( .C1(n19155), .C2(n19136), .A(n12989), .B(n12999), .ZN(
        P2_U2960) );
  INV_X1 U16208 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19166) );
  NAND2_X1 U16209 ( .A1(n19232), .A2(P2_UWORD_REG_2__SCAN_IN), .ZN(n12991) );
  OAI211_X1 U16210 ( .C1(n19166), .C2(n19136), .A(n12991), .B(n12990), .ZN(
        P2_U2954) );
  INV_X1 U16211 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19176) );
  NAND2_X1 U16212 ( .A1(n19232), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12993) );
  OAI211_X1 U16213 ( .C1(n19176), .C2(n19136), .A(n12993), .B(n12992), .ZN(
        P2_U2981) );
  INV_X1 U16214 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19162) );
  NAND2_X1 U16215 ( .A1(n19232), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n12995) );
  OAI211_X1 U16216 ( .C1(n19162), .C2(n19136), .A(n12995), .B(n12994), .ZN(
        P2_U2956) );
  NAND2_X1 U16217 ( .A1(n19232), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12997) );
  OAI211_X1 U16218 ( .C1(n11579), .C2(n19136), .A(n12997), .B(n12996), .ZN(
        P2_U2977) );
  INV_X2 U16219 ( .A(n12998), .ZN(n19232) );
  NAND2_X1 U16220 ( .A1(n19232), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13000) );
  OAI211_X1 U16221 ( .C1(n11489), .C2(n19136), .A(n13000), .B(n12999), .ZN(
        P2_U2975) );
  AOI22_X1 U16222 ( .A1(n19101), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19100), .ZN(n19214) );
  INV_X1 U16223 ( .A(n19214), .ZN(n13761) );
  AOI222_X1 U16224 ( .A1(P2_EAX_REG_17__SCAN_IN), .A2(n19231), .B1(n19205), 
        .B2(n13761), .C1(n19232), .C2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13001) );
  INV_X1 U16225 ( .A(n13001), .ZN(P2_U2953) );
  AOI22_X1 U16226 ( .A1(n19101), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19100), .ZN(n19216) );
  INV_X1 U16227 ( .A(n19216), .ZN(n15099) );
  AOI222_X1 U16228 ( .A1(P2_EAX_REG_19__SCAN_IN), .A2(n19231), .B1(n15099), 
        .B2(n19205), .C1(n19232), .C2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13002) );
  INV_X1 U16229 ( .A(n13002), .ZN(P2_U2955) );
  OAI21_X1 U16230 ( .B1(n10342), .B2(n19052), .A(n13003), .ZN(n13004) );
  XOR2_X1 U16231 ( .A(n13004), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n13082) );
  NOR2_X1 U16232 ( .A1(n16150), .A2(n19057), .ZN(n13008) );
  OAI21_X1 U16233 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13006), .A(
        n13005), .ZN(n13087) );
  NAND2_X1 U16234 ( .A1(n19236), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13085) );
  OAI21_X1 U16235 ( .B1(n16145), .B2(n13087), .A(n13085), .ZN(n13007) );
  AOI211_X1 U16236 ( .C1(n16143), .C2(n19057), .A(n13008), .B(n13007), .ZN(
        n13010) );
  NAND2_X1 U16237 ( .A1(n12489), .A2(n9787), .ZN(n13009) );
  OAI211_X1 U16238 ( .C1(n13082), .C2(n12452), .A(n13010), .B(n13009), .ZN(
        P2_U3013) );
  AOI22_X1 U16239 ( .A1(n19101), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19100), .ZN(n19218) );
  INV_X1 U16240 ( .A(n19218), .ZN(n19124) );
  AOI222_X1 U16241 ( .A1(P2_EAX_REG_21__SCAN_IN), .A2(n19231), .B1(n19205), 
        .B2(n19124), .C1(P2_UWORD_REG_5__SCAN_IN), .C2(n19232), .ZN(n13011) );
  INV_X1 U16242 ( .A(n13011), .ZN(P2_U2957) );
  INV_X1 U16243 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16359) );
  INV_X1 U16244 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18203) );
  OAI22_X1 U16245 ( .A1(n19100), .A2(n16359), .B1(n18203), .B2(n19101), .ZN(
        n15645) );
  AOI222_X1 U16246 ( .A1(P2_EAX_REG_23__SCAN_IN), .A2(n19231), .B1(n19205), 
        .B2(n15645), .C1(P2_UWORD_REG_7__SCAN_IN), .C2(n19232), .ZN(n13012) );
  INV_X1 U16247 ( .A(n13012), .ZN(P2_U2959) );
  AOI21_X1 U16248 ( .B1(n13015), .B2(n13014), .A(n13013), .ZN(n15553) );
  NAND2_X1 U16249 ( .A1(n19071), .A2(n13015), .ZN(n13016) );
  NAND2_X1 U16250 ( .A1(n10342), .A2(n13016), .ZN(n15549) );
  NAND2_X1 U16251 ( .A1(n19236), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n15556) );
  OAI21_X1 U16252 ( .B1(n12452), .B2(n15549), .A(n15556), .ZN(n13017) );
  AOI21_X1 U16253 ( .B1(n19241), .B2(n15553), .A(n13017), .ZN(n13020) );
  OAI21_X1 U16254 ( .B1(n19237), .B2(n13018), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13019) );
  OAI211_X1 U16255 ( .C1(n16130), .C2(n9968), .A(n13020), .B(n13019), .ZN(
        P2_U3014) );
  AND2_X1 U16256 ( .A1(n12142), .A2(n13061), .ZN(n13066) );
  NAND2_X1 U16257 ( .A1(n13066), .A2(n13294), .ZN(n13052) );
  INV_X1 U16258 ( .A(n13052), .ZN(n13022) );
  INV_X1 U16259 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20833) );
  NOR2_X2 U16260 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20671) );
  AND2_X1 U16261 ( .A1(n20671), .A2(n15722), .ZN(n13051) );
  INV_X1 U16262 ( .A(n13051), .ZN(n13021) );
  OAI211_X1 U16263 ( .C1(n13022), .C2(n20833), .A(n13348), .B(n13021), .ZN(
        P1_U2801) );
  AOI21_X1 U16264 ( .B1(n13025), .B2(n13024), .A(n13023), .ZN(n13028) );
  AND3_X1 U16265 ( .A1(n13028), .A2(n13027), .A3(n13026), .ZN(n13029) );
  OAI21_X1 U16266 ( .B1(n13030), .B2(n19135), .A(n13029), .ZN(n16239) );
  NOR2_X1 U16267 ( .A1(n19904), .A2(n19140), .ZN(n16259) );
  INV_X1 U16268 ( .A(n16259), .ZN(n15735) );
  OAI22_X1 U16269 ( .A1(n15735), .A2(n15736), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n19469), .ZN(n13031) );
  AOI21_X1 U16270 ( .B1(n16239), .B2(n13032), .A(n13031), .ZN(n15594) );
  INV_X1 U16271 ( .A(n15594), .ZN(n13034) );
  NOR2_X1 U16272 ( .A1(n10771), .A2(n10313), .ZN(n16234) );
  INV_X1 U16273 ( .A(n15592), .ZN(n13540) );
  NAND4_X1 U16274 ( .A1(n13034), .A2(n16234), .A3(n16233), .A4(n13540), .ZN(
        n13033) );
  OAI21_X1 U16275 ( .B1(n16240), .B2(n13034), .A(n13033), .ZN(P2_U3595) );
  INV_X1 U16276 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16373) );
  INV_X1 U16277 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18167) );
  AOI22_X1 U16278 ( .A1(n19101), .A2(n16373), .B1(n18167), .B2(n19100), .ZN(
        n19204) );
  INV_X1 U16279 ( .A(n19204), .ZN(n13043) );
  NAND2_X1 U16280 ( .A1(n15614), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13036) );
  AND4_X1 U16281 ( .A1(n10754), .A2(n13036), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19469), .ZN(n13037) );
  NOR2_X1 U16282 ( .A1(n13039), .A2(n13038), .ZN(n13040) );
  NOR2_X1 U16283 ( .A1(n11509), .A2(n13040), .ZN(n19065) );
  NAND2_X1 U16284 ( .A1(n19078), .A2(n19065), .ZN(n13153) );
  OAI211_X1 U16285 ( .C1(n19078), .C2(n19065), .A(n13153), .B(n19127), .ZN(
        n13042) );
  AOI22_X1 U16286 ( .A1(n19099), .A2(n19065), .B1(n19125), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13041) );
  OAI211_X1 U16287 ( .C1(n19120), .C2(n13043), .A(n13042), .B(n13041), .ZN(
        P2_U2919) );
  MUX2_X1 U16288 ( .A(n9968), .B(n13044), .S(n14984), .Z(n13045) );
  OAI21_X1 U16289 ( .B1(n19878), .B2(n15038), .A(n13045), .ZN(P2_U2887) );
  INV_X1 U16290 ( .A(n13046), .ZN(n13048) );
  INV_X1 U16291 ( .A(n12489), .ZN(n13090) );
  NOR2_X1 U16292 ( .A1(n13090), .A2(n14984), .ZN(n13049) );
  AOI21_X1 U16293 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n14984), .A(n13049), .ZN(
        n13050) );
  OAI21_X1 U16294 ( .B1(n19868), .B2(n15038), .A(n13050), .ZN(P2_U2886) );
  NOR2_X1 U16295 ( .A1(n13051), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13055)
         );
  OAI21_X1 U16296 ( .B1(n13684), .B2(n13053), .A(n20826), .ZN(n13054) );
  OAI21_X1 U16297 ( .B1(n13055), .B2(n20826), .A(n13054), .ZN(P1_U3487) );
  NOR2_X1 U16298 ( .A1(n13056), .A2(n20152), .ZN(n13058) );
  AOI21_X1 U16299 ( .B1(n13059), .B2(n13058), .A(n13057), .ZN(n13062) );
  OAI22_X1 U16300 ( .A1(n13062), .A2(n13293), .B1(n13061), .B2(n13060), .ZN(
        n13065) );
  INV_X1 U16301 ( .A(n13109), .ZN(n13063) );
  INV_X1 U16302 ( .A(n13293), .ZN(n13108) );
  NOR2_X1 U16303 ( .A1(n13063), .A2(n13108), .ZN(n13064) );
  OAI21_X1 U16304 ( .B1(n13065), .B2(n13064), .A(n11986), .ZN(n15710) );
  OAI22_X1 U16305 ( .A1(n13066), .A2(n12141), .B1(n13684), .B2(n13293), .ZN(
        n19917) );
  NAND2_X1 U16306 ( .A1(n14360), .A2(n15731), .ZN(n13116) );
  OR2_X1 U16307 ( .A1(n13116), .A2(n13684), .ZN(n20820) );
  AND2_X1 U16308 ( .A1(n20820), .A2(n20828), .ZN(n13067) );
  NOR2_X1 U16309 ( .A1(n19917), .A2(n13067), .ZN(n15708) );
  INV_X1 U16310 ( .A(n13294), .ZN(n19916) );
  OR2_X1 U16311 ( .A1(n15708), .A2(n19916), .ZN(n13070) );
  INV_X1 U16312 ( .A(n13070), .ZN(n19924) );
  INV_X1 U16313 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13068) );
  OR2_X1 U16314 ( .A1(n19924), .A2(n13068), .ZN(n13069) );
  OAI21_X1 U16315 ( .B1(n15710), .B2(n13070), .A(n13069), .ZN(P1_U3484) );
  MUX2_X1 U16316 ( .A(n13073), .B(n14359), .S(n15036), .Z(n13074) );
  OAI21_X1 U16317 ( .B1(n19860), .B2(n15038), .A(n13074), .ZN(P2_U2885) );
  XNOR2_X1 U16318 ( .A(n13075), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13079) );
  NAND2_X1 U16319 ( .A1(n13161), .A2(n13076), .ZN(n13077) );
  AND2_X1 U16320 ( .A1(n13129), .A2(n13077), .ZN(n19027) );
  INV_X1 U16321 ( .A(n19027), .ZN(n13631) );
  MUX2_X1 U16322 ( .A(n13631), .B(n21112), .S(n14984), .Z(n13078) );
  OAI21_X1 U16323 ( .B1(n13079), .B2(n15038), .A(n13078), .ZN(P2_U2882) );
  XNOR2_X1 U16324 ( .A(n13081), .B(n13080), .ZN(n19871) );
  INV_X1 U16325 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20994) );
  AOI211_X1 U16326 ( .C1(n13015), .C2(n20994), .A(n15481), .B(n14338), .ZN(
        n13084) );
  OAI22_X1 U16327 ( .A1(n20994), .A2(n15552), .B1(n16187), .B2(n13082), .ZN(
        n13083) );
  NOR2_X1 U16328 ( .A1(n13084), .A2(n13083), .ZN(n13086) );
  OAI211_X1 U16329 ( .C1(n16199), .C2(n13087), .A(n13086), .B(n13085), .ZN(
        n13088) );
  AOI21_X1 U16330 ( .B1(n16192), .B2(n19871), .A(n13088), .ZN(n13089) );
  OAI21_X1 U16331 ( .B1(n13090), .B2(n16194), .A(n13089), .ZN(P2_U3045) );
  INV_X1 U16332 ( .A(n13092), .ZN(n13094) );
  NAND2_X1 U16333 ( .A1(n13094), .A2(n13093), .ZN(n13098) );
  NOR2_X1 U16334 ( .A1(n13098), .A2(n13118), .ZN(n13095) );
  AND2_X1 U16335 ( .A1(n12428), .A2(n13095), .ZN(n13096) );
  NAND2_X1 U16336 ( .A1(n13100), .A2(n13096), .ZN(n14936) );
  INV_X1 U16337 ( .A(n14936), .ZN(n13148) );
  OR2_X1 U16338 ( .A1(n13109), .A2(n13110), .ZN(n13327) );
  XNOR2_X1 U16339 ( .A(n14937), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13104) );
  NOR2_X1 U16340 ( .A1(n13098), .A2(n13097), .ZN(n13099) );
  NAND2_X1 U16341 ( .A1(n13100), .A2(n13099), .ZN(n13325) );
  INV_X1 U16342 ( .A(n15691), .ZN(n14932) );
  XNOR2_X1 U16343 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13101) );
  OAI22_X1 U16344 ( .A1(n13325), .A2(n13104), .B1(n14932), .B2(n13101), .ZN(
        n13102) );
  AOI21_X1 U16345 ( .B1(n13327), .B2(n13104), .A(n13102), .ZN(n13103) );
  OAI21_X1 U16346 ( .B1(n13091), .B2(n13148), .A(n13103), .ZN(n13331) );
  INV_X1 U16347 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14762) );
  OAI22_X1 U16348 ( .A1(n14762), .A2(n20122), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14940) );
  INV_X1 U16349 ( .A(n14940), .ZN(n13107) );
  NOR2_X1 U16350 ( .A1(n15722), .A2(n20129), .ZN(n14939) );
  INV_X1 U16351 ( .A(n20805), .ZN(n13106) );
  INV_X1 U16352 ( .A(n13104), .ZN(n13105) );
  AOI222_X1 U16353 ( .A1(n13331), .A2(n15992), .B1(n13107), .B2(n14939), .C1(
        n13106), .C2(n13105), .ZN(n13124) );
  NAND2_X1 U16354 ( .A1(n13109), .A2(n13108), .ZN(n13195) );
  NAND2_X1 U16355 ( .A1(n13110), .A2(n13293), .ZN(n13111) );
  OAI21_X1 U16356 ( .B1(n12428), .B2(n13112), .A(n13111), .ZN(n13253) );
  INV_X1 U16357 ( .A(n13253), .ZN(n13122) );
  OR2_X1 U16358 ( .A1(n13113), .A2(n12003), .ZN(n13114) );
  AND2_X1 U16359 ( .A1(n13115), .A2(n13114), .ZN(n13120) );
  AND2_X1 U16360 ( .A1(n13116), .A2(n20828), .ZN(n13117) );
  OAI211_X1 U16361 ( .C1(n15691), .C2(n13118), .A(n13117), .B(n13293), .ZN(
        n13119) );
  AND2_X1 U16362 ( .A1(n13120), .A2(n13119), .ZN(n13121) );
  NAND3_X1 U16363 ( .A1(n13195), .A2(n13122), .A3(n13121), .ZN(n13337) );
  INV_X1 U16364 ( .A(n13337), .ZN(n15692) );
  INV_X2 U16365 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n13230) );
  NOR2_X1 U16366 ( .A1(n13230), .A2(n15722), .ZN(n16002) );
  NAND2_X1 U16367 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16002), .ZN(n16003) );
  INV_X1 U16368 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19923) );
  OAI22_X1 U16369 ( .A1(n15692), .A2(n19916), .B1(n16003), .B2(n19923), .ZN(
        n15990) );
  INV_X1 U16370 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20551) );
  NOR2_X1 U16371 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20551), .ZN(n20151) );
  OR2_X1 U16372 ( .A1(n15990), .A2(n20151), .ZN(n20809) );
  INV_X1 U16373 ( .A(n20809), .ZN(n13151) );
  NAND2_X1 U16374 ( .A1(n13151), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13123) );
  OAI21_X1 U16375 ( .B1(n13124), .B2(n13151), .A(n13123), .ZN(P1_U3472) );
  INV_X1 U16376 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19007) );
  INV_X1 U16377 ( .A(n13075), .ZN(n13125) );
  NOR2_X1 U16378 ( .A1(n13125), .A2(n15639), .ZN(n13127) );
  OAI211_X1 U16379 ( .C1(n13127), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15021), .B(n13126), .ZN(n13132) );
  AND2_X1 U16380 ( .A1(n13129), .A2(n13128), .ZN(n13130) );
  NOR2_X1 U16381 ( .A1(n13142), .A2(n13130), .ZN(n19015) );
  NAND2_X1 U16382 ( .A1(n19015), .A2(n15036), .ZN(n13131) );
  OAI211_X1 U16383 ( .C1(n15036), .C2(n19007), .A(n13132), .B(n13131), .ZN(
        P2_U2881) );
  NAND2_X1 U16384 ( .A1(n13134), .A2(n13133), .ZN(n13163) );
  INV_X1 U16385 ( .A(n13138), .ZN(n15578) );
  NOR2_X1 U16386 ( .A1(n15578), .A2(n14984), .ZN(n13139) );
  AOI21_X1 U16387 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n14984), .A(n13139), .ZN(
        n13140) );
  OAI21_X1 U16388 ( .B1(n19846), .B2(n15038), .A(n13140), .ZN(P2_U2884) );
  XOR2_X1 U16389 ( .A(n13126), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13146)
         );
  OR2_X1 U16390 ( .A1(n13142), .A2(n13141), .ZN(n13143) );
  NAND2_X1 U16391 ( .A1(n13200), .A2(n13143), .ZN(n19002) );
  MUX2_X1 U16392 ( .A(n19002), .B(n13144), .S(n14984), .Z(n13145) );
  OAI21_X1 U16393 ( .B1(n13146), .B2(n15038), .A(n13145), .ZN(P2_U2880) );
  AOI21_X1 U16394 ( .B1(n15691), .B2(n15992), .A(n13151), .ZN(n13152) );
  INV_X1 U16395 ( .A(n13147), .ZN(n13343) );
  OAI22_X1 U16396 ( .A1(n13343), .A2(n13148), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14933), .ZN(n15690) );
  OAI22_X1 U16397 ( .A1(n15722), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20805), .ZN(n13149) );
  AOI21_X1 U16398 ( .B1(n15690), .B2(n15992), .A(n13149), .ZN(n13150) );
  OAI22_X1 U16399 ( .A1(n13152), .A2(n10159), .B1(n13151), .B2(n13150), .ZN(
        P1_U3474) );
  INV_X1 U16400 ( .A(n19871), .ZN(n19054) );
  NOR2_X1 U16401 ( .A1(n19342), .A2(n19871), .ZN(n13269) );
  AOI21_X1 U16402 ( .B1(n19871), .B2(n19342), .A(n13269), .ZN(n13154) );
  NAND2_X1 U16403 ( .A1(n13154), .A2(n13153), .ZN(n13271) );
  OAI21_X1 U16404 ( .B1(n13154), .B2(n13153), .A(n13271), .ZN(n13155) );
  NAND2_X1 U16405 ( .A1(n13155), .A2(n19127), .ZN(n13157) );
  AOI22_X1 U16406 ( .A1(n19123), .A2(n13761), .B1(n19125), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13156) );
  OAI211_X1 U16407 ( .C1(n19054), .C2(n19092), .A(n13157), .B(n13156), .ZN(
        P2_U2918) );
  NAND2_X1 U16408 ( .A1(n13159), .A2(n13158), .ZN(n13160) );
  NAND2_X1 U16409 ( .A1(n13161), .A2(n13160), .ZN(n19048) );
  NAND2_X1 U16410 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15640), .ZN(
        n13162) );
  OAI211_X1 U16411 ( .C1(n13164), .C2(n15634), .A(n13163), .B(n13162), .ZN(
        n13165) );
  AOI21_X1 U16412 ( .B1(n13167), .B2(n13166), .A(n13165), .ZN(n13168) );
  NOR2_X1 U16413 ( .A1(n13168), .A2(n13075), .ZN(n19128) );
  NAND2_X1 U16414 ( .A1(n19128), .A2(n15021), .ZN(n13170) );
  NAND2_X1 U16415 ( .A1(n14984), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n13169) );
  OAI211_X1 U16416 ( .C1(n19048), .C2(n14984), .A(n13170), .B(n13169), .ZN(
        P2_U2883) );
  NOR2_X2 U16417 ( .A1(n13191), .A2(n13230), .ZN(n13951) );
  INV_X1 U16418 ( .A(n13171), .ZN(n14220) );
  NAND2_X1 U16419 ( .A1(n14220), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13487) );
  NAND2_X1 U16420 ( .A1(n14287), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n13173) );
  NAND2_X1 U16421 ( .A1(n13230), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13172) );
  OAI211_X1 U16422 ( .C1(n13487), .C2(n10159), .A(n13173), .B(n13172), .ZN(
        n13174) );
  AOI21_X1 U16423 ( .B1(n13147), .B2(n13951), .A(n13174), .ZN(n13216) );
  NAND2_X1 U16424 ( .A1(n13175), .A2(n11984), .ZN(n13176) );
  NAND2_X1 U16425 ( .A1(n13176), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13178) );
  OR2_X1 U16426 ( .A1(n13178), .A2(n13216), .ZN(n13219) );
  INV_X1 U16427 ( .A(n13219), .ZN(n13177) );
  AOI21_X1 U16428 ( .B1(n13216), .B2(n13178), .A(n13177), .ZN(n13197) );
  NAND3_X1 U16429 ( .A1(n20824), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15997) );
  INV_X1 U16430 ( .A(n15997), .ZN(n13179) );
  AND2_X2 U16431 ( .A1(n13179), .A2(n20671), .ZN(n20096) );
  OAI21_X1 U16432 ( .B1(n13181), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13180), .ZN(n13263) );
  NAND2_X1 U16433 ( .A1(n12122), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13257) );
  INV_X1 U16434 ( .A(n20671), .ZN(n20669) );
  NAND2_X1 U16435 ( .A1(n20669), .A2(n13182), .ZN(n20827) );
  AND2_X1 U16436 ( .A1(n20827), .A2(n20824), .ZN(n13183) );
  NAND2_X1 U16437 ( .A1(n20824), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13185) );
  INV_X1 U16438 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20622) );
  NAND2_X1 U16439 ( .A1(n20622), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13184) );
  NAND2_X1 U16440 ( .A1(n13185), .A2(n13184), .ZN(n13223) );
  OAI21_X1 U16441 ( .B1(n20090), .B2(n13223), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13186) );
  OAI211_X1 U16442 ( .C1(n13263), .C2(n19922), .A(n13257), .B(n13186), .ZN(
        n13187) );
  AOI21_X1 U16443 ( .B1(n13197), .B2(n20096), .A(n13187), .ZN(n13188) );
  INV_X1 U16444 ( .A(n13188), .ZN(P1_U2999) );
  OR2_X1 U16445 ( .A1(n14364), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13190) );
  AND2_X1 U16446 ( .A1(n13190), .A2(n13189), .ZN(n13673) );
  INV_X1 U16447 ( .A(n13673), .ZN(n13198) );
  NAND4_X1 U16448 ( .A1(n13193), .A2(n20214), .A3(n13192), .A4(n13191), .ZN(
        n13251) );
  OR2_X1 U16449 ( .A1(n13251), .A2(n14360), .ZN(n13194) );
  NAND2_X1 U16450 ( .A1(n13195), .A2(n13194), .ZN(n13196) );
  INV_X1 U16451 ( .A(n13197), .ZN(n13686) );
  OAI222_X1 U16452 ( .A1(n13198), .A2(n20015), .B1(n12032), .B2(n20029), .C1(
        n13686), .C2(n14529), .ZN(P1_U2872) );
  NAND2_X1 U16453 ( .A1(n13200), .A2(n13199), .ZN(n13201) );
  NAND2_X1 U16454 ( .A1(n13287), .A2(n13201), .ZN(n18995) );
  OAI211_X1 U16455 ( .C1(n13204), .C2(n13203), .A(n13202), .B(n15021), .ZN(
        n13206) );
  NAND2_X1 U16456 ( .A1(n14984), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13205) );
  OAI211_X1 U16457 ( .C1(n18995), .C2(n14984), .A(n13206), .B(n13205), .ZN(
        P2_U2879) );
  NAND2_X1 U16458 ( .A1(n14919), .A2(n13951), .ZN(n13215) );
  NAND2_X1 U16459 ( .A1(n14287), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n13212) );
  NAND2_X1 U16460 ( .A1(n13230), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13211) );
  OAI211_X1 U16461 ( .C1(n13487), .C2(n9984), .A(n13212), .B(n13211), .ZN(
        n13213) );
  INV_X1 U16462 ( .A(n13213), .ZN(n13214) );
  NAND2_X1 U16463 ( .A1(n13215), .A2(n13214), .ZN(n13221) );
  INV_X1 U16464 ( .A(n13216), .ZN(n13217) );
  OR2_X1 U16465 ( .A1(n13217), .A2(n10352), .ZN(n13218) );
  NAND2_X1 U16466 ( .A1(n13219), .A2(n13218), .ZN(n13220) );
  NAND2_X1 U16467 ( .A1(n13221), .A2(n13220), .ZN(n13238) );
  OAI21_X1 U16468 ( .B1(n13221), .B2(n13220), .A(n13238), .ZN(n13732) );
  INV_X1 U16469 ( .A(n20096), .ZN(n14748) );
  INV_X1 U16470 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13222) );
  NOR2_X1 U16471 ( .A1(n20135), .A2(n13222), .ZN(n14913) );
  NOR2_X1 U16472 ( .A1(n20101), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13224) );
  AOI211_X1 U16473 ( .C1(n20090), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14913), .B(n13224), .ZN(n13228) );
  OR2_X1 U16474 ( .A1(n13225), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14908) );
  NAND3_X1 U16475 ( .A1(n14908), .A2(n9815), .A3(n20097), .ZN(n13227) );
  OAI211_X1 U16476 ( .C1(n13732), .C2(n14748), .A(n13228), .B(n13227), .ZN(
        P1_U2998) );
  NAND2_X1 U16477 ( .A1(n13229), .A2(n13951), .ZN(n13236) );
  XNOR2_X1 U16478 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20003) );
  NAND2_X1 U16479 ( .A1(n13230), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13514) );
  AOI21_X1 U16480 ( .B1(n14282), .B2(n20003), .A(n14286), .ZN(n13232) );
  NAND2_X1 U16481 ( .A1(n14287), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n13231) );
  OAI211_X1 U16482 ( .C1(n13487), .C2(n13233), .A(n13232), .B(n13231), .ZN(
        n13234) );
  INV_X1 U16483 ( .A(n13234), .ZN(n13235) );
  NAND2_X1 U16484 ( .A1(n13236), .A2(n13235), .ZN(n13237) );
  NAND2_X1 U16485 ( .A1(n14286), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13388) );
  NAND2_X1 U16486 ( .A1(n13237), .A2(n13388), .ZN(n13241) );
  NAND2_X1 U16487 ( .A1(n13241), .A2(n13238), .ZN(n13242) );
  NAND2_X1 U16488 ( .A1(n13389), .A2(n13242), .ZN(n20005) );
  NOR2_X1 U16489 ( .A1(n13244), .A2(n13243), .ZN(n13245) );
  OR2_X1 U16490 ( .A1(n13405), .A2(n13245), .ZN(n20011) );
  INV_X1 U16491 ( .A(n20011), .ZN(n20125) );
  AOI22_X1 U16492 ( .A1(n20024), .A2(n20125), .B1(n14527), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13246) );
  OAI21_X1 U16493 ( .B1(n20005), .B2(n14529), .A(n13246), .ZN(P1_U2870) );
  INV_X1 U16494 ( .A(n13247), .ZN(n13248) );
  NAND3_X1 U16495 ( .A1(n13248), .A2(n13293), .A3(n20828), .ZN(n13249) );
  OAI21_X1 U16496 ( .B1(n13251), .B2(n13250), .A(n13249), .ZN(n13252) );
  NAND2_X1 U16497 ( .A1(n11989), .A2(n11986), .ZN(n13255) );
  NAND2_X2 U16498 ( .A1(n14600), .A2(n13255), .ZN(n14603) );
  INV_X1 U16499 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20059) );
  MUX2_X1 U16500 ( .A(DATAI_0_), .B(BUF1_REG_0__SCAN_IN), .S(n20145), .Z(
        n20159) );
  INV_X1 U16501 ( .A(n20159), .ZN(n13256) );
  OAI222_X1 U16502 ( .A1(n14603), .A2(n13686), .B1(n14600), .B2(n20059), .C1(
        n14602), .C2(n13256), .ZN(P1_U2904) );
  INV_X1 U16503 ( .A(n13257), .ZN(n13260) );
  INV_X1 U16504 ( .A(n14870), .ZN(n13258) );
  NOR2_X1 U16505 ( .A1(n13258), .A2(n14899), .ZN(n13259) );
  NOR2_X1 U16506 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13259), .ZN(
        n14909) );
  AOI211_X1 U16507 ( .C1(n20126), .C2(n13673), .A(n13260), .B(n14909), .ZN(
        n13262) );
  OAI21_X1 U16508 ( .B1(n14910), .B2(n14846), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13261) );
  OAI211_X1 U16509 ( .C1(n13263), .C2(n15935), .A(n13262), .B(n13261), .ZN(
        P1_U3031) );
  INV_X1 U16510 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20053) );
  MUX2_X1 U16511 ( .A(DATAI_2_), .B(BUF1_REG_2__SCAN_IN), .S(n20145), .Z(
        n20178) );
  INV_X1 U16512 ( .A(n20178), .ZN(n13264) );
  OAI222_X1 U16513 ( .A1(n14603), .A2(n20005), .B1(n14600), .B2(n20053), .C1(
        n14602), .C2(n13264), .ZN(P1_U2902) );
  NAND2_X1 U16514 ( .A1(n13266), .A2(n13265), .ZN(n13268) );
  AND2_X1 U16515 ( .A1(n13268), .A2(n10122), .ZN(n13505) );
  INV_X1 U16516 ( .A(n19860), .ZN(n13539) );
  INV_X1 U16517 ( .A(n13505), .ZN(n19862) );
  NOR2_X1 U16518 ( .A1(n13539), .A2(n19862), .ZN(n13442) );
  AOI21_X1 U16519 ( .B1(n13539), .B2(n19862), .A(n13442), .ZN(n13273) );
  INV_X1 U16520 ( .A(n13269), .ZN(n13270) );
  NAND2_X1 U16521 ( .A1(n13271), .A2(n13270), .ZN(n13272) );
  NAND2_X1 U16522 ( .A1(n13273), .A2(n13272), .ZN(n13444) );
  OAI21_X1 U16523 ( .B1(n13273), .B2(n13272), .A(n13444), .ZN(n13274) );
  NAND2_X1 U16524 ( .A1(n13274), .A2(n19127), .ZN(n13276) );
  AOI22_X1 U16525 ( .A1(n19123), .A2(n16071), .B1(n19125), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13275) );
  OAI211_X1 U16526 ( .C1(n13505), .C2(n19092), .A(n13276), .B(n13275), .ZN(
        P2_U2917) );
  OR2_X1 U16527 ( .A1(n13278), .A2(n13277), .ZN(n20124) );
  NAND3_X1 U16528 ( .A1(n20124), .A2(n9813), .A3(n20097), .ZN(n13283) );
  INV_X1 U16529 ( .A(n20003), .ZN(n13281) );
  INV_X1 U16530 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20993) );
  INV_X1 U16531 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n19999) );
  OAI22_X1 U16532 ( .A1(n14742), .A2(n20993), .B1(n20135), .B2(n19999), .ZN(
        n13280) );
  AOI21_X1 U16533 ( .B1(n13281), .B2(n15847), .A(n13280), .ZN(n13282) );
  OAI211_X1 U16534 ( .C1(n20005), .C2(n14748), .A(n13283), .B(n13282), .ZN(
        P1_U2997) );
  OAI211_X1 U16535 ( .C1(n13285), .C2(n12516), .A(n15021), .B(n13408), .ZN(
        n13290) );
  AND2_X1 U16536 ( .A1(n13287), .A2(n13286), .ZN(n13288) );
  OR2_X1 U16537 ( .A1(n13288), .A2(n9918), .ZN(n15265) );
  INV_X1 U16538 ( .A(n15265), .ZN(n18982) );
  NAND2_X1 U16539 ( .A1(n18982), .A2(n15036), .ZN(n13289) );
  OAI211_X1 U16540 ( .C1(n15036), .C2(n20978), .A(n13290), .B(n13289), .ZN(
        P2_U2878) );
  XNOR2_X1 U16541 ( .A(n13726), .B(n13291), .ZN(n14914) );
  AOI22_X1 U16542 ( .A1(n20024), .A2(n14914), .B1(n14527), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13292) );
  OAI21_X1 U16543 ( .B1(n13732), .B2(n14529), .A(n13292), .ZN(P1_U2871) );
  INV_X1 U16544 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13298) );
  NAND3_X1 U16545 ( .A1(n15691), .A2(n13294), .A3(n13293), .ZN(n13295) );
  NAND2_X1 U16546 ( .A1(n16002), .A2(n20824), .ZN(n20046) );
  INV_X1 U16547 ( .A(n20046), .ZN(n20051) );
  AOI22_X1 U16548 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13297) );
  OAI21_X1 U16549 ( .B1(n13298), .B2(n20030), .A(n13297), .ZN(P1_U2910) );
  INV_X1 U16550 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13300) );
  AOI22_X1 U16551 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13299) );
  OAI21_X1 U16552 ( .B1(n13300), .B2(n20030), .A(n13299), .ZN(P1_U2915) );
  INV_X1 U16553 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13302) );
  AOI22_X1 U16554 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13301) );
  OAI21_X1 U16555 ( .B1(n13302), .B2(n20030), .A(n13301), .ZN(P1_U2917) );
  INV_X1 U16556 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U16557 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13303) );
  OAI21_X1 U16558 ( .B1(n13304), .B2(n20030), .A(n13303), .ZN(P1_U2920) );
  INV_X1 U16559 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13306) );
  AOI22_X1 U16560 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13305) );
  OAI21_X1 U16561 ( .B1(n13306), .B2(n20030), .A(n13305), .ZN(P1_U2918) );
  INV_X1 U16562 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13308) );
  AOI22_X1 U16563 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13307) );
  OAI21_X1 U16564 ( .B1(n13308), .B2(n20030), .A(n13307), .ZN(P1_U2909) );
  INV_X1 U16565 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13310) );
  AOI22_X1 U16566 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13309) );
  OAI21_X1 U16567 ( .B1(n13310), .B2(n20030), .A(n13309), .ZN(P1_U2916) );
  INV_X1 U16568 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n21052) );
  AOI22_X1 U16569 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13311) );
  OAI21_X1 U16570 ( .B1(n21052), .B2(n20030), .A(n13311), .ZN(P1_U2919) );
  XOR2_X1 U16571 ( .A(n13408), .B(n13312), .Z(n13317) );
  NOR2_X1 U16572 ( .A1(n9918), .A2(n13313), .ZN(n13314) );
  OR2_X1 U16573 ( .A1(n13415), .A2(n13314), .ZN(n18970) );
  MUX2_X1 U16574 ( .A(n18970), .B(n13315), .S(n14984), .Z(n13316) );
  OAI21_X1 U16575 ( .B1(n13317), .B2(n15038), .A(n13316), .ZN(P2_U2877) );
  INV_X1 U16576 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n16341) );
  INV_X1 U16577 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n21134) );
  INV_X1 U16578 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n20997) );
  OAI222_X1 U16579 ( .A1(n20045), .A2(n16341), .B1(n20030), .B2(n21134), .C1(
        n20046), .C2(n20997), .ZN(P1_U2914) );
  NAND2_X1 U16580 ( .A1(n20421), .A2(n14936), .ZN(n13330) );
  MUX2_X1 U16581 ( .A(n11826), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14937), .Z(n13319) );
  NOR2_X1 U16582 ( .A1(n13319), .A2(n13318), .ZN(n13328) );
  AOI21_X1 U16583 ( .B1(n14937), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13397), .ZN(n13320) );
  NOR2_X1 U16584 ( .A1(n12282), .A2(n13320), .ZN(n20806) );
  NAND2_X1 U16585 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13321) );
  INV_X1 U16586 ( .A(n13321), .ZN(n13322) );
  MUX2_X1 U16587 ( .A(n13322), .B(n13321), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13323) );
  NAND2_X1 U16588 ( .A1(n15691), .A2(n13323), .ZN(n13324) );
  OAI21_X1 U16589 ( .B1(n13325), .B2(n20806), .A(n13324), .ZN(n13326) );
  AOI21_X1 U16590 ( .B1(n13328), .B2(n13327), .A(n13326), .ZN(n13329) );
  NAND2_X1 U16591 ( .A1(n13330), .A2(n13329), .ZN(n20804) );
  MUX2_X1 U16592 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20804), .S(
        n13337), .Z(n15702) );
  NOR2_X1 U16593 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15722), .ZN(n13338) );
  AOI22_X1 U16594 ( .A1(n15702), .A2(n15722), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13338), .ZN(n13333) );
  MUX2_X1 U16595 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13331), .S(
        n13337), .Z(n15698) );
  AOI22_X1 U16596 ( .A1(n13338), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15698), .B2(n15722), .ZN(n13332) );
  NOR2_X1 U16597 ( .A1(n13333), .A2(n13332), .ZN(n15714) );
  INV_X1 U16598 ( .A(n11832), .ZN(n13334) );
  NAND2_X1 U16599 ( .A1(n15714), .A2(n13334), .ZN(n13342) );
  INV_X1 U16600 ( .A(n20309), .ZN(n20542) );
  OR2_X1 U16601 ( .A1(n13335), .A2(n20542), .ZN(n13336) );
  XNOR2_X1 U16602 ( .A(n13336), .B(n15995), .ZN(n19991) );
  OAI21_X1 U16603 ( .B1(n19991), .B2(n12428), .A(n13337), .ZN(n13340) );
  AOI21_X1 U16604 ( .B1(n15692), .B2(n15995), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13339) );
  AOI22_X1 U16605 ( .A1(n13340), .A2(n13339), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13338), .ZN(n15712) );
  AND3_X1 U16606 ( .A1(n13342), .A2(n15712), .A3(n19923), .ZN(n13341) );
  NAND2_X1 U16607 ( .A1(n13230), .A2(n15722), .ZN(n20823) );
  INV_X1 U16608 ( .A(n20823), .ZN(n13662) );
  OAI21_X1 U16609 ( .B1(n13341), .B2(n16003), .A(n20315), .ZN(n20142) );
  NAND3_X1 U16610 ( .A1(n13342), .A2(n15712), .A3(n16002), .ZN(n15723) );
  INV_X1 U16611 ( .A(n15723), .ZN(n13345) );
  NAND2_X1 U16612 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20551), .ZN(n14928) );
  INV_X1 U16613 ( .A(n14928), .ZN(n14922) );
  OAI22_X1 U16614 ( .A1(n13175), .A2(n20669), .B1(n13343), .B2(n14922), .ZN(
        n13344) );
  OAI21_X1 U16615 ( .B1(n13345), .B2(n13344), .A(n20142), .ZN(n13346) );
  OAI21_X1 U16616 ( .B1(n20142), .B2(n20581), .A(n13346), .ZN(P1_U3478) );
  INV_X1 U16617 ( .A(n20828), .ZN(n15730) );
  AND2_X1 U16618 ( .A1(n20821), .A2(n15730), .ZN(n13347) );
  OR2_X2 U16619 ( .A1(n13348), .A2(n13347), .ZN(n20086) );
  AOI22_X1 U16620 ( .A1(n20087), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20086), .ZN(n13349) );
  NOR2_X2 U16621 ( .A1(n20086), .A2(n20169), .ZN(n20074) );
  MUX2_X1 U16622 ( .A(DATAI_3_), .B(BUF1_REG_3__SCAN_IN), .S(n20145), .Z(
        n20186) );
  NAND2_X1 U16623 ( .A1(n20074), .A2(n20186), .ZN(n13376) );
  NAND2_X1 U16624 ( .A1(n13349), .A2(n13376), .ZN(P1_U2955) );
  AOI22_X1 U16625 ( .A1(n20087), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20086), .ZN(n13350) );
  MUX2_X1 U16626 ( .A(DATAI_7_), .B(BUF1_REG_7__SCAN_IN), .S(n20145), .Z(
        n20217) );
  NAND2_X1 U16627 ( .A1(n20074), .A2(n20217), .ZN(n13361) );
  NAND2_X1 U16628 ( .A1(n13350), .A2(n13361), .ZN(P1_U2959) );
  INV_X2 U16629 ( .A(n13385), .ZN(n20087) );
  AOI22_X1 U16630 ( .A1(n20087), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20086), .ZN(n13351) );
  MUX2_X1 U16631 ( .A(DATAI_5_), .B(BUF1_REG_5__SCAN_IN), .S(n20145), .Z(
        n20200) );
  NAND2_X1 U16632 ( .A1(n20074), .A2(n20200), .ZN(n13374) );
  NAND2_X1 U16633 ( .A1(n13351), .A2(n13374), .ZN(P1_U2942) );
  AOI22_X1 U16634 ( .A1(n20087), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20086), .ZN(n13354) );
  INV_X1 U16635 ( .A(n20145), .ZN(n20144) );
  INV_X1 U16636 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16357) );
  NOR2_X1 U16637 ( .A1(n20144), .A2(n16357), .ZN(n13352) );
  AOI21_X1 U16638 ( .B1(DATAI_8_), .B2(n20144), .A(n13352), .ZN(n14554) );
  INV_X1 U16639 ( .A(n14554), .ZN(n13353) );
  NAND2_X1 U16640 ( .A1(n20074), .A2(n13353), .ZN(n13359) );
  NAND2_X1 U16641 ( .A1(n13354), .A2(n13359), .ZN(P1_U2960) );
  AOI22_X1 U16642 ( .A1(n20087), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20086), .ZN(n13355) );
  NAND2_X1 U16643 ( .A1(n20074), .A2(n20159), .ZN(n13372) );
  NAND2_X1 U16644 ( .A1(n13355), .A2(n13372), .ZN(P1_U2937) );
  AOI22_X1 U16645 ( .A1(n20087), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20086), .ZN(n13356) );
  MUX2_X1 U16646 ( .A(DATAI_1_), .B(BUF1_REG_1__SCAN_IN), .S(n20145), .Z(
        n20170) );
  NAND2_X1 U16647 ( .A1(n20074), .A2(n20170), .ZN(n13370) );
  NAND2_X1 U16648 ( .A1(n13356), .A2(n13370), .ZN(P1_U2938) );
  AOI22_X1 U16649 ( .A1(n20087), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20086), .ZN(n13357) );
  MUX2_X1 U16650 ( .A(DATAI_4_), .B(BUF1_REG_4__SCAN_IN), .S(n20145), .Z(
        n20193) );
  NAND2_X1 U16651 ( .A1(n20074), .A2(n20193), .ZN(n13366) );
  NAND2_X1 U16652 ( .A1(n13357), .A2(n13366), .ZN(P1_U2941) );
  AOI22_X1 U16653 ( .A1(n20087), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20086), .ZN(n13358) );
  MUX2_X1 U16654 ( .A(DATAI_6_), .B(BUF1_REG_6__SCAN_IN), .S(n20145), .Z(
        n20206) );
  NAND2_X1 U16655 ( .A1(n20074), .A2(n20206), .ZN(n13363) );
  NAND2_X1 U16656 ( .A1(n13358), .A2(n13363), .ZN(P1_U2958) );
  AOI22_X1 U16657 ( .A1(n20087), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20086), .ZN(n13360) );
  NAND2_X1 U16658 ( .A1(n13360), .A2(n13359), .ZN(P1_U2945) );
  AOI22_X1 U16659 ( .A1(n20087), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20086), .ZN(n13362) );
  NAND2_X1 U16660 ( .A1(n13362), .A2(n13361), .ZN(P1_U2944) );
  AOI22_X1 U16661 ( .A1(n20087), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20086), .ZN(n13364) );
  NAND2_X1 U16662 ( .A1(n13364), .A2(n13363), .ZN(P1_U2943) );
  AOI22_X1 U16663 ( .A1(n20087), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20086), .ZN(n13365) );
  NAND2_X1 U16664 ( .A1(n20074), .A2(n20178), .ZN(n13368) );
  NAND2_X1 U16665 ( .A1(n13365), .A2(n13368), .ZN(P1_U2939) );
  AOI22_X1 U16666 ( .A1(n20087), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20086), .ZN(n13367) );
  NAND2_X1 U16667 ( .A1(n13367), .A2(n13366), .ZN(P1_U2956) );
  AOI22_X1 U16668 ( .A1(n20087), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20086), .ZN(n13369) );
  NAND2_X1 U16669 ( .A1(n13369), .A2(n13368), .ZN(P1_U2954) );
  AOI22_X1 U16670 ( .A1(n20087), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20086), .ZN(n13371) );
  NAND2_X1 U16671 ( .A1(n13371), .A2(n13370), .ZN(P1_U2953) );
  AOI22_X1 U16672 ( .A1(n20087), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20086), .ZN(n13373) );
  NAND2_X1 U16673 ( .A1(n13373), .A2(n13372), .ZN(P1_U2952) );
  AOI22_X1 U16674 ( .A1(n20087), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20086), .ZN(n13375) );
  NAND2_X1 U16675 ( .A1(n13375), .A2(n13374), .ZN(P1_U2957) );
  AOI22_X1 U16676 ( .A1(n20087), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20086), .ZN(n13377) );
  NAND2_X1 U16677 ( .A1(n13377), .A2(n13376), .ZN(P1_U2940) );
  INV_X1 U16678 ( .A(P1_UWORD_REG_9__SCAN_IN), .ZN(n21113) );
  MUX2_X1 U16679 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n20145), .Z(
        n14548) );
  NAND2_X1 U16680 ( .A1(n20074), .A2(n14548), .ZN(n20076) );
  NAND2_X1 U16681 ( .A1(n20087), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n13378) );
  OAI211_X1 U16682 ( .C1(n13381), .C2(n21113), .A(n20076), .B(n13378), .ZN(
        P1_U2946) );
  INV_X1 U16683 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13384) );
  INV_X1 U16684 ( .A(n20074), .ZN(n13383) );
  INV_X1 U16685 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13379) );
  NOR2_X1 U16686 ( .A1(n20144), .A2(n13379), .ZN(n13380) );
  AOI21_X1 U16687 ( .B1(DATAI_15_), .B2(n20144), .A(n13380), .ZN(n14598) );
  INV_X1 U16688 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13382) );
  OAI222_X1 U16689 ( .A1(n13385), .A2(n13384), .B1(n13383), .B2(n14598), .C1(
        n13382), .C2(n13381), .ZN(P1_U2967) );
  INV_X1 U16690 ( .A(P1_UWORD_REG_14__SCAN_IN), .ZN(n13387) );
  INV_X1 U16691 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14530) );
  INV_X1 U16692 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13386) );
  OAI222_X1 U16693 ( .A1(n13387), .A2(n20046), .B1(n20030), .B2(n14530), .C1(
        n13386), .C2(n20045), .ZN(P1_U2906) );
  NAND2_X1 U16694 ( .A1(n20146), .A2(n13951), .ZN(n13400) );
  INV_X1 U16695 ( .A(n13391), .ZN(n13390) );
  INV_X1 U16696 ( .A(n13484), .ZN(n13394) );
  INV_X1 U16697 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13392) );
  NAND2_X1 U16698 ( .A1(n13392), .A2(n13391), .ZN(n13393) );
  NAND2_X1 U16699 ( .A1(n13394), .A2(n13393), .ZN(n13710) );
  AOI22_X1 U16700 ( .A1(n13710), .A2(n14282), .B1(n14286), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13396) );
  NAND2_X1 U16701 ( .A1(n14287), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n13395) );
  OAI211_X1 U16702 ( .C1(n13487), .C2(n13397), .A(n13396), .B(n13395), .ZN(
        n13398) );
  INV_X1 U16703 ( .A(n13398), .ZN(n13399) );
  NAND2_X1 U16704 ( .A1(n13400), .A2(n13399), .ZN(n13401) );
  OAI21_X1 U16705 ( .B1(n13402), .B2(n13401), .A(n13520), .ZN(n13717) );
  INV_X1 U16706 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20050) );
  INV_X1 U16707 ( .A(n20186), .ZN(n13403) );
  OAI222_X1 U16708 ( .A1(n14603), .A2(n13717), .B1(n14600), .B2(n20050), .C1(
        n14602), .C2(n13403), .ZN(P1_U2901) );
  OAI21_X1 U16709 ( .B1(n13405), .B2(n13404), .A(n13494), .ZN(n20110) );
  INV_X1 U16710 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13406) );
  OAI222_X1 U16711 ( .A1(n20110), .A2(n20015), .B1(n13406), .B2(n20029), .C1(
        n13717), .C2(n14529), .ZN(P1_U2869) );
  NOR2_X1 U16712 ( .A1(n13408), .A2(n13407), .ZN(n13412) );
  INV_X1 U16713 ( .A(n13409), .ZN(n13410) );
  OAI211_X1 U16714 ( .C1(n13412), .C2(n13411), .A(n13410), .B(n15021), .ZN(
        n13418) );
  OAI21_X1 U16715 ( .B1(n13415), .B2(n13414), .A(n13413), .ZN(n13416) );
  INV_X1 U16716 ( .A(n13416), .ZN(n18961) );
  NAND2_X1 U16717 ( .A1(n18961), .A2(n15036), .ZN(n13417) );
  OAI211_X1 U16718 ( .C1(n15036), .C2(n18954), .A(n13418), .B(n13417), .ZN(
        P2_U2876) );
  NAND2_X1 U16719 ( .A1(n9925), .A2(n13420), .ZN(n13421) );
  XNOR2_X1 U16720 ( .A(n13578), .B(n13421), .ZN(n13432) );
  OR2_X1 U16721 ( .A1(n13423), .A2(n13422), .ZN(n13425) );
  NAND2_X1 U16722 ( .A1(n13425), .A2(n13424), .ZN(n19850) );
  INV_X1 U16723 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19789) );
  INV_X1 U16724 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n20955) );
  OAI22_X1 U16725 ( .A1(n19008), .A2(n20955), .B1(n13576), .B2(n19035), .ZN(
        n13428) );
  NOR2_X1 U16726 ( .A1(n13426), .A2(n19070), .ZN(n13427) );
  AOI211_X1 U16727 ( .C1(n19049), .C2(P2_REIP_REG_3__SCAN_IN), .A(n13428), .B(
        n13427), .ZN(n13430) );
  NAND2_X1 U16728 ( .A1(n13138), .A2(n19062), .ZN(n13429) );
  OAI211_X1 U16729 ( .C1(n19850), .C2(n19053), .A(n13430), .B(n13429), .ZN(
        n13431) );
  AOI21_X1 U16730 ( .B1(n13432), .B2(n19764), .A(n13431), .ZN(n13433) );
  OAI21_X1 U16731 ( .B1(n19846), .B2(n13510), .A(n13433), .ZN(P2_U2852) );
  INV_X1 U16732 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U16733 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13434) );
  OAI21_X1 U16734 ( .B1(n13435), .B2(n20030), .A(n13434), .ZN(P1_U2908) );
  INV_X1 U16735 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13437) );
  AOI22_X1 U16736 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13436) );
  OAI21_X1 U16737 ( .B1(n13437), .B2(n20030), .A(n13436), .ZN(P1_U2907) );
  AOI22_X1 U16738 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13438) );
  OAI21_X1 U16739 ( .B1(n14553), .B2(n20030), .A(n13438), .ZN(P1_U2912) );
  INV_X1 U16740 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13440) );
  AOI22_X1 U16741 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13439) );
  OAI21_X1 U16742 ( .B1(n13440), .B2(n20030), .A(n13439), .ZN(P1_U2913) );
  INV_X1 U16743 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20055) );
  INV_X1 U16744 ( .A(n20170), .ZN(n13441) );
  OAI222_X1 U16745 ( .A1(n14603), .A2(n13732), .B1(n14600), .B2(n20055), .C1(
        n14602), .C2(n13441), .ZN(P1_U2903) );
  XOR2_X1 U16746 ( .A(n19850), .B(n19846), .Z(n13446) );
  INV_X1 U16747 ( .A(n13442), .ZN(n13443) );
  NAND2_X1 U16748 ( .A1(n13444), .A2(n13443), .ZN(n13445) );
  NAND2_X1 U16749 ( .A1(n13445), .A2(n13446), .ZN(n13561) );
  OAI21_X1 U16750 ( .B1(n13446), .B2(n13445), .A(n13561), .ZN(n13447) );
  NAND2_X1 U16751 ( .A1(n13447), .A2(n19127), .ZN(n13449) );
  AOI22_X1 U16752 ( .A1(n19123), .A2(n15099), .B1(n19125), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n13448) );
  OAI211_X1 U16753 ( .C1(n19850), .C2(n19092), .A(n13449), .B(n13448), .ZN(
        P2_U2916) );
  OR2_X1 U16754 ( .A1(n19846), .A2(n19902), .ZN(n19706) );
  NAND2_X1 U16755 ( .A1(n19864), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19540) );
  OAI22_X1 U16756 ( .A1(n19706), .A2(n19847), .B1(n19873), .B2(n19540), .ZN(
        n13453) );
  NAND2_X1 U16757 ( .A1(n10986), .A2(n19469), .ZN(n13451) );
  INV_X1 U16758 ( .A(n19540), .ZN(n19497) );
  NAND2_X1 U16759 ( .A1(n16212), .A2(n19497), .ZN(n13454) );
  AND2_X1 U16760 ( .A1(n13454), .A2(n15596), .ZN(n13450) );
  AOI21_X1 U16761 ( .B1(n13451), .B2(n13450), .A(n19536), .ZN(n13452) );
  NAND2_X1 U16762 ( .A1(n13453), .A2(n13452), .ZN(n19573) );
  INV_X1 U16763 ( .A(n19573), .ZN(n19581) );
  NOR2_X2 U16764 ( .A1(n19650), .A2(n19847), .ZN(n19578) );
  INV_X1 U16765 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20191) );
  INV_X1 U16766 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n17222) );
  OAI22_X2 U16767 ( .A1(n20191), .A2(n15651), .B1(n17222), .B2(n15650), .ZN(
        n19734) );
  NOR2_X2 U16768 ( .A1(n19620), .A2(n19847), .ZN(n19609) );
  INV_X1 U16769 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20189) );
  INV_X1 U16770 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18188) );
  OAI22_X2 U16771 ( .A1(n20189), .A2(n15651), .B1(n18188), .B2(n15650), .ZN(
        n19678) );
  AOI22_X1 U16772 ( .A1(n19578), .A2(n19734), .B1(n19609), .B2(n19678), .ZN(
        n13459) );
  NAND2_X1 U16773 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19497), .ZN(
        n13456) );
  INV_X1 U16774 ( .A(n13454), .ZN(n19576) );
  OAI21_X1 U16775 ( .B1(n10986), .B2(n19576), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13455) );
  OAI21_X1 U16776 ( .B1(n13456), .B2(n15596), .A(n13455), .ZN(n19577) );
  NAND2_X1 U16777 ( .A1(n16066), .A2(n19707), .ZN(n19681) );
  INV_X1 U16778 ( .A(n19681), .ZN(n19733) );
  NOR2_X2 U16779 ( .A1(n13457), .A2(n15608), .ZN(n19732) );
  AOI22_X1 U16780 ( .A1(n19577), .A2(n19733), .B1(n19732), .B2(n19576), .ZN(
        n13458) );
  OAI211_X1 U16781 ( .C1(n19581), .C2(n13460), .A(n13459), .B(n13458), .ZN(
        P2_U3140) );
  OAI21_X1 U16782 ( .B1(n13463), .B2(n13462), .A(n13461), .ZN(n20113) );
  INV_X1 U16783 ( .A(n13717), .ZN(n13466) );
  AOI22_X1 U16784 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13464) );
  OAI21_X1 U16785 ( .B1(n20101), .B2(n13710), .A(n13464), .ZN(n13465) );
  AOI21_X1 U16786 ( .B1(n13466), .B2(n20096), .A(n13465), .ZN(n13467) );
  OAI21_X1 U16787 ( .B1(n20113), .B2(n19922), .A(n13467), .ZN(P1_U2996) );
  NAND2_X1 U16788 ( .A1(n13413), .A2(n13468), .ZN(n13469) );
  AND2_X1 U16789 ( .A1(n13475), .A2(n13469), .ZN(n18950) );
  INV_X1 U16790 ( .A(n18950), .ZN(n15488) );
  AND2_X1 U16791 ( .A1(n13409), .A2(n13471), .ZN(n13480) );
  INV_X1 U16792 ( .A(n13480), .ZN(n13470) );
  OAI211_X1 U16793 ( .C1(n13409), .C2(n13471), .A(n13470), .B(n15021), .ZN(
        n13473) );
  NAND2_X1 U16794 ( .A1(n14984), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13472) );
  OAI211_X1 U16795 ( .C1(n15488), .C2(n14984), .A(n13473), .B(n13472), .ZN(
        P2_U2875) );
  NAND2_X1 U16796 ( .A1(n13475), .A2(n13474), .ZN(n13476) );
  AND2_X1 U16797 ( .A1(n13585), .A2(n13476), .ZN(n18940) );
  INV_X1 U16798 ( .A(n18940), .ZN(n13483) );
  INV_X1 U16799 ( .A(n13477), .ZN(n13478) );
  OAI211_X1 U16800 ( .C1(n13480), .C2(n13479), .A(n13478), .B(n15021), .ZN(
        n13482) );
  NAND2_X1 U16801 ( .A1(n14984), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13481) );
  OAI211_X1 U16802 ( .C1(n13483), .C2(n14984), .A(n13482), .B(n13481), .ZN(
        P2_U2874) );
  INV_X1 U16803 ( .A(n20193), .ZN(n13492) );
  OAI21_X1 U16804 ( .B1(n13484), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13511), .ZN(n20100) );
  NAND2_X1 U16805 ( .A1(n13230), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13486) );
  NAND2_X1 U16806 ( .A1(n14287), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n13485) );
  OAI211_X1 U16807 ( .C1(n13487), .C2(n15995), .A(n13486), .B(n13485), .ZN(
        n13488) );
  MUX2_X1 U16808 ( .A(n20100), .B(n13488), .S(n10352), .Z(n13489) );
  INV_X1 U16809 ( .A(n13521), .ZN(n13491) );
  XNOR2_X1 U16810 ( .A(n13520), .B(n13491), .ZN(n20095) );
  INV_X1 U16811 ( .A(n20095), .ZN(n13496) );
  INV_X1 U16812 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20048) );
  OAI222_X1 U16813 ( .A1(n14602), .A2(n13492), .B1(n14603), .B2(n13496), .C1(
        n20048), .C2(n14600), .ZN(P1_U2900) );
  NAND2_X1 U16814 ( .A1(n13494), .A2(n13493), .ZN(n13495) );
  AND2_X1 U16815 ( .A1(n15981), .A2(n13495), .ZN(n20105) );
  INV_X1 U16816 ( .A(n20105), .ZN(n13497) );
  INV_X1 U16817 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n19983) );
  OAI222_X1 U16818 ( .A1(n20015), .A2(n13497), .B1(n19983), .B2(n20029), .C1(
        n14529), .C2(n13496), .ZN(P1_U2868) );
  INV_X1 U16819 ( .A(n14352), .ZN(n13500) );
  NOR2_X1 U16820 ( .A1(n19041), .A2(n13498), .ZN(n13536) );
  INV_X1 U16821 ( .A(n13536), .ZN(n13499) );
  AOI221_X1 U16822 ( .B1(n13500), .B2(n13536), .C1(n14352), .C2(n13499), .A(
        n19061), .ZN(n13501) );
  INV_X1 U16823 ( .A(n13501), .ZN(n13509) );
  NAND2_X1 U16824 ( .A1(n19063), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n13503) );
  AOI22_X1 U16825 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19080), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19049), .ZN(n13502) );
  OAI211_X1 U16826 ( .C1(n19070), .C2(n13504), .A(n13503), .B(n13502), .ZN(
        n13507) );
  NOR2_X1 U16827 ( .A1(n13505), .A2(n19053), .ZN(n13506) );
  AOI211_X1 U16828 ( .C1(n19062), .C2(n9956), .A(n13507), .B(n13506), .ZN(
        n13508) );
  OAI211_X1 U16829 ( .C1(n19860), .C2(n13510), .A(n13509), .B(n13508), .ZN(
        P2_U2853) );
  INV_X1 U16830 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13517) );
  AND2_X1 U16831 ( .A1(n13511), .A2(n13513), .ZN(n13512) );
  OR2_X1 U16832 ( .A1(n13512), .A2(n13637), .ZN(n19978) );
  NOR2_X1 U16833 ( .A1(n13514), .A2(n13513), .ZN(n13515) );
  AOI21_X1 U16834 ( .B1(n19978), .B2(n14282), .A(n13515), .ZN(n13516) );
  OAI21_X1 U16835 ( .B1(n13654), .B2(n13517), .A(n13516), .ZN(n13518) );
  OAI21_X1 U16836 ( .B1(n13520), .B2(n13521), .A(n13522), .ZN(n13525) );
  AND2_X1 U16837 ( .A1(n13525), .A2(n13644), .ZN(n20026) );
  INV_X1 U16838 ( .A(n20026), .ZN(n13527) );
  INV_X1 U16839 ( .A(n20200), .ZN(n13526) );
  OAI222_X1 U16840 ( .A1(n14603), .A2(n13527), .B1(n14600), .B2(n13517), .C1(
        n14602), .C2(n13526), .ZN(P1_U2899) );
  INV_X1 U16841 ( .A(n15567), .ZN(n13528) );
  NAND2_X1 U16842 ( .A1(n13528), .A2(n16211), .ZN(n15584) );
  NAND2_X1 U16843 ( .A1(n13529), .A2(n15584), .ZN(n13535) );
  NAND2_X1 U16844 ( .A1(n9956), .A2(n15576), .ZN(n13534) );
  NAND2_X1 U16845 ( .A1(n13530), .A2(n16227), .ZN(n15585) );
  NOR2_X1 U16846 ( .A1(n13531), .A2(n9799), .ZN(n13532) );
  AOI22_X1 U16847 ( .A1(n15585), .A2(n13535), .B1(n13532), .B2(n11464), .ZN(
        n13533) );
  OAI211_X1 U16848 ( .C1(n15582), .C2(n13535), .A(n13534), .B(n13533), .ZN(
        n16210) );
  OAI21_X1 U16849 ( .B1(n19084), .B2(n13537), .A(n13536), .ZN(n19060) );
  OAI21_X1 U16850 ( .B1(n9925), .B2(n20994), .A(n19060), .ZN(n15573) );
  INV_X1 U16851 ( .A(n19084), .ZN(n13538) );
  AOI22_X1 U16852 ( .A1(n19041), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n13538), .B2(n9925), .ZN(n15564) );
  NOR2_X1 U16853 ( .A1(n15564), .A2(n11393), .ZN(n15572) );
  AOI222_X1 U16854 ( .A1(n16210), .A2(n13540), .B1(n15573), .B2(n15572), .C1(
        n13539), .C2(n16252), .ZN(n13542) );
  NAND2_X1 U16855 ( .A1(n15594), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13541) );
  OAI21_X1 U16856 ( .B1(n13542), .B2(n15594), .A(n13541), .ZN(P2_U3599) );
  NAND2_X1 U16857 ( .A1(n13544), .A2(n13543), .ZN(n13546) );
  XNOR2_X1 U16858 ( .A(n13546), .B(n13545), .ZN(n13583) );
  XNOR2_X1 U16859 ( .A(n13547), .B(n13548), .ZN(n13580) );
  INV_X1 U16860 ( .A(n13549), .ZN(n13552) );
  NOR2_X1 U16861 ( .A1(n19789), .A2(n19034), .ZN(n13550) );
  AOI221_X1 U16862 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13552), .C1(
        n21168), .C2(n13551), .A(n13550), .ZN(n13555) );
  OAI22_X1 U16863 ( .A1(n19850), .A2(n16177), .B1(n15578), .B2(n16194), .ZN(
        n13553) );
  INV_X1 U16864 ( .A(n13553), .ZN(n13554) );
  OAI211_X1 U16865 ( .C1(n13580), .C2(n16199), .A(n13555), .B(n13554), .ZN(
        n13556) );
  AOI21_X1 U16866 ( .B1(n13583), .B2(n16196), .A(n13556), .ZN(n13557) );
  INV_X1 U16867 ( .A(n13557), .ZN(P2_U3043) );
  NAND2_X1 U16868 ( .A1(n19846), .A2(n19850), .ZN(n13560) );
  INV_X1 U16869 ( .A(n13424), .ZN(n13558) );
  XNOR2_X1 U16870 ( .A(n13559), .B(n13558), .ZN(n19032) );
  AOI21_X1 U16871 ( .B1(n13561), .B2(n13560), .A(n19032), .ZN(n19126) );
  XOR2_X1 U16872 ( .A(n19128), .B(n19126), .Z(n13564) );
  AOI22_X1 U16873 ( .A1(n19099), .A2(n19032), .B1(n19125), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13563) );
  NAND2_X1 U16874 ( .A1(n19123), .A2(n16066), .ZN(n13562) );
  OAI211_X1 U16875 ( .C1(n13564), .C2(n19093), .A(n13563), .B(n13562), .ZN(
        P2_U2915) );
  NAND2_X1 U16876 ( .A1(n19846), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19434) );
  NOR2_X1 U16877 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16209) );
  NAND2_X1 U16878 ( .A1(n19873), .A2(n16209), .ZN(n13569) );
  OAI21_X1 U16879 ( .B1(n19434), .B2(n19502), .A(n13569), .ZN(n13568) );
  NOR2_X1 U16880 ( .A1(n19883), .A2(n13569), .ZN(n19270) );
  OAI211_X1 U16881 ( .C1(n19270), .C2(n19469), .A(n19707), .B(n13571), .ZN(
        n13566) );
  INV_X1 U16882 ( .A(n13566), .ZN(n13567) );
  NAND2_X1 U16883 ( .A1(n13568), .A2(n13567), .ZN(n19272) );
  INV_X1 U16884 ( .A(n19272), .ZN(n19255) );
  INV_X1 U16885 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13575) );
  INV_X1 U16886 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20176) );
  INV_X1 U16887 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n17232) );
  OAI22_X2 U16888 ( .A1(n20176), .A2(n15651), .B1(n17232), .B2(n15650), .ZN(
        n19722) );
  NOR2_X2 U16889 ( .A1(n19502), .A2(n19441), .ZN(n19305) );
  INV_X1 U16890 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20173) );
  INV_X1 U16891 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18179) );
  OAI22_X2 U16892 ( .A1(n20173), .A2(n15651), .B1(n18179), .B2(n15650), .ZN(
        n19670) );
  AOI22_X1 U16893 ( .A1(n19265), .A2(n19722), .B1(n19305), .B2(n19670), .ZN(
        n13574) );
  INV_X1 U16894 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19654) );
  OAI21_X1 U16895 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n13569), .A(n19654), 
        .ZN(n13570) );
  AND2_X1 U16896 ( .A1(n13571), .A2(n13570), .ZN(n19271) );
  NAND2_X1 U16897 ( .A1(n16071), .A2(n19707), .ZN(n19673) );
  NOR2_X2 U16898 ( .A1(n13572), .A2(n15608), .ZN(n19720) );
  AOI22_X1 U16899 ( .A1(n19271), .A2(n19721), .B1(n19720), .B2(n19270), .ZN(
        n13573) );
  OAI211_X1 U16900 ( .C1(n19255), .C2(n13575), .A(n13574), .B(n13573), .ZN(
        P2_U3058) );
  OAI22_X1 U16901 ( .A1(n16150), .A2(n13576), .B1(n19789), .B2(n19034), .ZN(
        n13577) );
  AOI21_X1 U16902 ( .B1(n16143), .B2(n13578), .A(n13577), .ZN(n13579) );
  OAI21_X1 U16903 ( .B1(n15578), .B2(n16130), .A(n13579), .ZN(n13582) );
  NOR2_X1 U16904 ( .A1(n13580), .A2(n16145), .ZN(n13581) );
  AOI211_X1 U16905 ( .C1(n13583), .C2(n19242), .A(n13582), .B(n13581), .ZN(
        n13584) );
  INV_X1 U16906 ( .A(n13584), .ZN(P2_U3011) );
  AOI21_X1 U16907 ( .B1(n13586), .B2(n13585), .A(n13606), .ZN(n16158) );
  INV_X1 U16908 ( .A(n16158), .ZN(n18932) );
  OAI211_X1 U16909 ( .C1(n13477), .C2(n12518), .A(n15021), .B(n13608), .ZN(
        n13590) );
  NAND2_X1 U16910 ( .A1(n14984), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13589) );
  OAI211_X1 U16911 ( .C1(n18932), .C2(n14984), .A(n13590), .B(n13589), .ZN(
        P2_U2873) );
  XOR2_X1 U16912 ( .A(n13592), .B(n13591), .Z(n19243) );
  INV_X1 U16913 ( .A(n19243), .ZN(n13603) );
  NAND2_X1 U16914 ( .A1(n13594), .A2(n13593), .ZN(n13595) );
  XNOR2_X1 U16915 ( .A(n13595), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19240) );
  NOR2_X1 U16916 ( .A1(n11303), .A2(n19034), .ZN(n13598) );
  NOR2_X1 U16917 ( .A1(n13623), .A2(n13596), .ZN(n13597) );
  AOI211_X1 U16918 ( .C1(n16192), .C2(n19032), .A(n13598), .B(n13597), .ZN(
        n13600) );
  INV_X1 U16919 ( .A(n19048), .ZN(n19238) );
  NAND2_X1 U16920 ( .A1(n19238), .A2(n16182), .ZN(n13599) );
  OAI211_X1 U16921 ( .C1(n13621), .C2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13600), .B(n13599), .ZN(n13601) );
  AOI21_X1 U16922 ( .B1(n19240), .B2(n16183), .A(n13601), .ZN(n13602) );
  OAI21_X1 U16923 ( .B1(n13603), .B2(n16187), .A(n13602), .ZN(P2_U3042) );
  OR2_X1 U16924 ( .A1(n13606), .A2(n13605), .ZN(n13607) );
  NAND2_X1 U16925 ( .A1(n13604), .A2(n13607), .ZN(n18917) );
  INV_X1 U16926 ( .A(n13608), .ZN(n13612) );
  INV_X1 U16927 ( .A(n13609), .ZN(n13611) );
  INV_X1 U16928 ( .A(n13610), .ZN(n15029) );
  OAI211_X1 U16929 ( .C1(n13612), .C2(n13611), .A(n15021), .B(n15029), .ZN(
        n13614) );
  NAND2_X1 U16930 ( .A1(n14984), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n13613) );
  OAI211_X1 U16931 ( .C1(n18917), .C2(n14984), .A(n13614), .B(n13613), .ZN(
        P2_U2872) );
  XNOR2_X1 U16932 ( .A(n13615), .B(n13616), .ZN(n16146) );
  OAI21_X1 U16933 ( .B1(n13620), .B2(n13618), .A(n13617), .ZN(n13619) );
  OAI21_X1 U16934 ( .B1(n11039), .B2(n13620), .A(n13619), .ZN(n16144) );
  NOR2_X1 U16935 ( .A1(n11308), .A2(n19034), .ZN(n13626) );
  AOI211_X1 U16936 ( .C1(n13624), .C2(n13623), .A(n13622), .B(n13621), .ZN(
        n13625) );
  AOI211_X1 U16937 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n13627), .A(
        n13626), .B(n13625), .ZN(n13634) );
  OAI21_X1 U16938 ( .B1(n13630), .B2(n13629), .A(n13628), .ZN(n19132) );
  OAI22_X1 U16939 ( .A1(n19132), .A2(n16177), .B1(n16194), .B2(n13631), .ZN(
        n13632) );
  INV_X1 U16940 ( .A(n13632), .ZN(n13633) );
  OAI211_X1 U16941 ( .C1(n16144), .C2(n16199), .A(n13634), .B(n13633), .ZN(
        n13635) );
  INV_X1 U16942 ( .A(n13635), .ZN(n13636) );
  OAI21_X1 U16943 ( .B1(n16146), .B2(n16187), .A(n13636), .ZN(P2_U3041) );
  INV_X1 U16944 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13640) );
  NOR2_X1 U16945 ( .A1(n13637), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13638) );
  OR2_X1 U16946 ( .A1(n13650), .A2(n13638), .ZN(n19970) );
  AOI22_X1 U16947 ( .A1(n19970), .A2(n14282), .B1(n14286), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13639) );
  OAI21_X1 U16948 ( .B1(n13654), .B2(n13640), .A(n13639), .ZN(n13641) );
  AND2_X1 U16949 ( .A1(n13644), .A2(n13643), .ZN(n13645) );
  NOR2_X1 U16950 ( .A1(n13656), .A2(n13645), .ZN(n19966) );
  INV_X1 U16951 ( .A(n19966), .ZN(n13648) );
  XNOR2_X1 U16952 ( .A(n15983), .B(n15965), .ZN(n19964) );
  AOI22_X1 U16953 ( .A1(n19964), .A2(n20024), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14527), .ZN(n13646) );
  OAI21_X1 U16954 ( .B1(n13648), .B2(n14529), .A(n13646), .ZN(P1_U2866) );
  INV_X1 U16955 ( .A(n20206), .ZN(n13647) );
  OAI222_X1 U16956 ( .A1(n14603), .A2(n13648), .B1(n14600), .B2(n13640), .C1(
        n14602), .C2(n13647), .ZN(P1_U2898) );
  INV_X1 U16957 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13658) );
  OR2_X1 U16958 ( .A1(n13650), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13651) );
  NAND2_X1 U16959 ( .A1(n13651), .A2(n13700), .ZN(n19960) );
  AOI22_X1 U16960 ( .A1(n19960), .A2(n14282), .B1(n14286), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13652) );
  NAND2_X1 U16961 ( .A1(n13656), .A2(n13655), .ZN(n13705) );
  OR2_X1 U16962 ( .A1(n13656), .A2(n13655), .ZN(n13657) );
  AND2_X1 U16963 ( .A1(n13705), .A2(n13657), .ZN(n20020) );
  INV_X1 U16964 ( .A(n20020), .ZN(n13660) );
  INV_X1 U16965 ( .A(n20217), .ZN(n13659) );
  OAI222_X1 U16966 ( .A1(n14603), .A2(n13660), .B1(n14602), .B2(n13659), .C1(
        n13658), .C2(n14600), .ZN(P1_U2897) );
  NAND2_X1 U16967 ( .A1(n20826), .A2(n13661), .ZN(n19990) );
  INV_X1 U16968 ( .A(n19990), .ZN(n20008) );
  OAI221_X1 U16969 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20551), .C1(n20824), 
        .C2(P1_STATE2_REG_3__SCAN_IN), .A(n13662), .ZN(n13665) );
  NOR2_X1 U16970 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15722), .ZN(n13663) );
  NAND2_X1 U16971 ( .A1(n14282), .A2(n13663), .ZN(n13664) );
  NAND2_X1 U16972 ( .A1(n13665), .A2(n13664), .ZN(n13666) );
  AND2_X1 U16973 ( .A1(n20828), .A2(n20622), .ZN(n15717) );
  OAI21_X1 U16974 ( .B1(n12026), .B2(n15718), .A(n15717), .ZN(n13668) );
  NOR2_X1 U16975 ( .A1(n13668), .A2(n20152), .ZN(n13667) );
  NAND2_X1 U16976 ( .A1(n19951), .A2(n19940), .ZN(n19972) );
  INV_X1 U16977 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n21140) );
  INV_X1 U16978 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14480) );
  OR2_X1 U16979 ( .A1(n14360), .A2(n14480), .ZN(n13671) );
  AND3_X1 U16980 ( .A1(n13671), .A2(n13669), .A3(n13668), .ZN(n13670) );
  NAND2_X1 U16981 ( .A1(n20826), .A2(n13670), .ZN(n19984) );
  NOR2_X1 U16982 ( .A1(n13671), .A2(n15717), .ZN(n13672) );
  AOI22_X1 U16983 ( .A1(P1_EBX_REG_0__SCAN_IN), .A2(n19996), .B1(n19988), .B2(
        n13673), .ZN(n13682) );
  INV_X1 U16984 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15784) );
  INV_X1 U16985 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14117) );
  INV_X1 U16986 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14434) );
  INV_X1 U16987 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14179) );
  INV_X1 U16988 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14629) );
  INV_X1 U16989 ( .A(n14281), .ZN(n13677) );
  NAND2_X1 U16990 ( .A1(n13677), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13678) );
  INV_X1 U16991 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14371) );
  NAND2_X1 U16992 ( .A1(n19986), .A2(n20002), .ZN(n13680) );
  NAND2_X1 U16993 ( .A1(n13680), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13681) );
  OAI211_X1 U16994 ( .C1(n15816), .C2(n21140), .A(n13682), .B(n13681), .ZN(
        n13688) );
  NOR2_X1 U16995 ( .A1(n14300), .A2(n15722), .ZN(n13683) );
  NAND2_X1 U16996 ( .A1(n20826), .A2(n13684), .ZN(n13685) );
  NAND2_X1 U16997 ( .A1(n19947), .A2(n13685), .ZN(n19982) );
  NOR2_X1 U16998 ( .A1(n13686), .A2(n20004), .ZN(n13687) );
  AOI211_X1 U16999 ( .C1(n20008), .C2(n13147), .A(n13688), .B(n13687), .ZN(
        n13689) );
  INV_X1 U17000 ( .A(n13689), .ZN(P1_U2840) );
  AOI22_X1 U17001 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13693) );
  AOI22_X1 U17002 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13692) );
  AOI22_X1 U17003 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13691) );
  AOI22_X1 U17004 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13690) );
  NAND4_X1 U17005 ( .A1(n13693), .A2(n13692), .A3(n13691), .A4(n13690), .ZN(
        n13699) );
  AOI22_X1 U17006 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U17007 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13696) );
  AOI22_X1 U17008 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13695) );
  AOI22_X1 U17009 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13694) );
  NAND4_X1 U17010 ( .A1(n13697), .A2(n13696), .A3(n13695), .A4(n13694), .ZN(
        n13698) );
  OAI21_X1 U17011 ( .B1(n13699), .B2(n13698), .A(n13951), .ZN(n13704) );
  NAND2_X1 U17012 ( .A1(n14287), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n13703) );
  INV_X1 U17013 ( .A(n13700), .ZN(n13701) );
  XNOR2_X1 U17014 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n13701), .ZN(
        n13803) );
  AOI22_X1 U17015 ( .A1(n14282), .A2(n13803), .B1(n14286), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13702) );
  NOR2_X2 U17016 ( .A1(n13705), .A2(n13707), .ZN(n13752) );
  AOI21_X1 U17017 ( .B1(n13707), .B2(n13705), .A(n13706), .ZN(n13805) );
  INV_X1 U17018 ( .A(n13805), .ZN(n13724) );
  INV_X1 U17019 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13709) );
  OAI21_X1 U17020 ( .B1(n15967), .B2(n13708), .A(n15943), .ZN(n15957) );
  OAI222_X1 U17021 ( .A1(n13724), .A2(n14529), .B1(n20029), .B2(n13709), .C1(
        n15957), .C2(n20015), .ZN(P1_U2864) );
  INV_X1 U17022 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20999) );
  OAI222_X1 U17023 ( .A1(n14603), .A2(n13724), .B1(n14600), .B2(n20999), .C1(
        n14602), .C2(n14554), .ZN(P1_U2896) );
  NOR2_X1 U17024 ( .A1(n19940), .A2(n13222), .ZN(n20000) );
  NAND2_X1 U17025 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n19981) );
  OAI211_X1 U17026 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(P1_REIP_REG_2__SCAN_IN), 
        .A(n20000), .B(n19981), .ZN(n13716) );
  INV_X1 U17027 ( .A(n13710), .ZN(n13711) );
  OAI21_X1 U17028 ( .B1(n19940), .B2(P1_REIP_REG_1__SCAN_IN), .A(n19951), .ZN(
        n19997) );
  AOI22_X1 U17029 ( .A1(n13711), .A2(n15809), .B1(n19997), .B2(
        P1_REIP_REG_3__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U17030 ( .A1(n19998), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n19996), .B2(P1_EBX_REG_3__SCAN_IN), .ZN(n13712) );
  OAI211_X1 U17031 ( .C1(n20012), .C2(n20110), .A(n13713), .B(n13712), .ZN(
        n13714) );
  AOI21_X1 U17032 ( .B1(n20421), .B2(n20008), .A(n13714), .ZN(n13715) );
  OAI211_X1 U17033 ( .C1(n13717), .C2(n20004), .A(n13716), .B(n13715), .ZN(
        P1_U2837) );
  INV_X1 U17034 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20982) );
  INV_X1 U17035 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20747) );
  NOR3_X1 U17036 ( .A1(n13222), .A2(n20747), .A3(n19981), .ZN(n19952) );
  NAND4_X1 U17037 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19952), .A3(
        P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n19939) );
  NOR2_X1 U17038 ( .A1(n20982), .A2(n19939), .ZN(n14230) );
  NAND2_X1 U17039 ( .A1(n14230), .A2(n19951), .ZN(n13870) );
  INV_X1 U17040 ( .A(n13870), .ZN(n15739) );
  NOR2_X1 U17041 ( .A1(n15816), .A2(n15739), .ZN(n19945) );
  OAI21_X1 U17042 ( .B1(n19940), .B2(n19939), .A(n20982), .ZN(n13722) );
  OAI21_X1 U17043 ( .B1(n19984), .B2(n13709), .A(n20135), .ZN(n13719) );
  NOR2_X1 U17044 ( .A1(n20002), .A2(n13803), .ZN(n13718) );
  AOI211_X1 U17045 ( .C1(n19998), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n13719), .B(n13718), .ZN(n13720) );
  OAI21_X1 U17046 ( .B1(n15957), .B2(n20012), .A(n13720), .ZN(n13721) );
  AOI21_X1 U17047 ( .B1(n19945), .B2(n13722), .A(n13721), .ZN(n13723) );
  OAI21_X1 U17048 ( .B1(n13724), .B2(n19947), .A(n13723), .ZN(P1_U2832) );
  INV_X1 U17049 ( .A(n13725), .ZN(n20625) );
  MUX2_X1 U17050 ( .A(n15809), .B(n19998), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13730) );
  INV_X1 U17051 ( .A(n19940), .ZN(n15741) );
  AOI22_X1 U17052 ( .A1(n15741), .A2(n13222), .B1(n19996), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13728) );
  NAND2_X1 U17053 ( .A1(n19988), .A2(n13726), .ZN(n13727) );
  OAI211_X1 U17054 ( .C1(n13222), .C2(n19951), .A(n13728), .B(n13727), .ZN(
        n13729) );
  AOI211_X1 U17055 ( .C1(n20625), .C2(n20008), .A(n13730), .B(n13729), .ZN(
        n13731) );
  OAI21_X1 U17056 ( .B1(n13732), .B2(n20004), .A(n13731), .ZN(P1_U2839) );
  XOR2_X1 U17057 ( .A(n19942), .B(n13733), .Z(n13827) );
  INV_X1 U17058 ( .A(n13827), .ZN(n19946) );
  AOI22_X1 U17059 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13738) );
  AOI22_X1 U17060 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13737) );
  AOI22_X1 U17061 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13736) );
  AOI22_X1 U17062 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13735) );
  NAND4_X1 U17063 ( .A1(n13738), .A2(n13737), .A3(n13736), .A4(n13735), .ZN(
        n13744) );
  AOI22_X1 U17064 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13742) );
  AOI22_X1 U17065 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13741) );
  AOI22_X1 U17066 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13740) );
  AOI22_X1 U17067 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13739) );
  NAND4_X1 U17068 ( .A1(n13742), .A2(n13741), .A3(n13740), .A4(n13739), .ZN(
        n13743) );
  OAI21_X1 U17069 ( .B1(n13744), .B2(n13743), .A(n13951), .ZN(n13747) );
  NAND2_X1 U17070 ( .A1(n14287), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13746) );
  NAND2_X1 U17071 ( .A1(n14286), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13745) );
  NAND3_X1 U17072 ( .A1(n13747), .A2(n13746), .A3(n13745), .ZN(n13748) );
  AOI21_X1 U17073 ( .B1(n19946), .B2(n14282), .A(n13748), .ZN(n13750) );
  AND2_X1 U17074 ( .A1(n13749), .A2(n13750), .ZN(n13753) );
  OR2_X1 U17075 ( .A1(n13753), .A2(n13782), .ZN(n20016) );
  INV_X1 U17076 ( .A(n14602), .ZN(n13754) );
  AOI22_X1 U17077 ( .A1(n13754), .A2(n14548), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14587), .ZN(n13755) );
  OAI21_X1 U17078 ( .B1(n20016), .B2(n14603), .A(n13755), .ZN(P1_U2895) );
  OAI21_X1 U17079 ( .B1(n13756), .B2(n13758), .A(n13757), .ZN(n15027) );
  OR2_X1 U17080 ( .A1(n15450), .A2(n13759), .ZN(n13760) );
  NAND2_X1 U17081 ( .A1(n15417), .A2(n13760), .ZN(n18901) );
  AOI22_X1 U17082 ( .A1(n19089), .A2(BUF1_REG_17__SCAN_IN), .B1(n19090), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U17083 ( .A1(n19088), .A2(n13761), .B1(n19125), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n13762) );
  OAI211_X1 U17084 ( .C1(n19092), .C2(n18901), .A(n13763), .B(n13762), .ZN(
        n13764) );
  INV_X1 U17085 ( .A(n13764), .ZN(n13765) );
  OAI21_X1 U17086 ( .B1(n15027), .B2(n19093), .A(n13765), .ZN(P2_U2902) );
  AOI22_X1 U17087 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13769) );
  AOI22_X1 U17088 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11906), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13768) );
  AOI22_X1 U17089 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13767) );
  AOI22_X1 U17090 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13766) );
  NAND4_X1 U17091 ( .A1(n13769), .A2(n13768), .A3(n13767), .A4(n13766), .ZN(
        n13775) );
  AOI22_X1 U17092 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13773) );
  AOI22_X1 U17093 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13772) );
  AOI22_X1 U17094 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13771) );
  AOI22_X1 U17095 ( .A1(n14199), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13770) );
  NAND4_X1 U17096 ( .A1(n13773), .A2(n13772), .A3(n13771), .A4(n13770), .ZN(
        n13774) );
  NOR2_X1 U17097 ( .A1(n13775), .A2(n13774), .ZN(n13780) );
  INV_X1 U17098 ( .A(n13951), .ZN(n13779) );
  XNOR2_X1 U17099 ( .A(n13776), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14752) );
  NAND2_X1 U17100 ( .A1(n14752), .A2(n14282), .ZN(n13778) );
  AOI22_X1 U17101 ( .A1(n14287), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n14286), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13777) );
  OAI211_X1 U17102 ( .C1(n13780), .C2(n13779), .A(n13778), .B(n13777), .ZN(
        n13781) );
  INV_X1 U17103 ( .A(n13781), .ZN(n13783) );
  AOI21_X1 U17104 ( .B1(n13783), .B2(n9803), .A(n13867), .ZN(n14754) );
  AND2_X1 U17105 ( .A1(n15945), .A2(n13785), .ZN(n13786) );
  OR2_X1 U17106 ( .A1(n13786), .A2(n9868), .ZN(n15937) );
  OAI22_X1 U17107 ( .A1(n15937), .A2(n20015), .B1(n13787), .B2(n20029), .ZN(
        n13788) );
  AOI21_X1 U17108 ( .B1(n14754), .B2(n20025), .A(n13788), .ZN(n13789) );
  INV_X1 U17109 ( .A(n13789), .ZN(P1_U2862) );
  INV_X1 U17110 ( .A(n14754), .ZN(n13798) );
  INV_X1 U17111 ( .A(n14752), .ZN(n13792) );
  AOI22_X1 U17112 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19998), .B1(
        n19996), .B2(P1_EBX_REG_10__SCAN_IN), .ZN(n13790) );
  OAI211_X1 U17113 ( .C1(n15937), .C2(n20012), .A(n13790), .B(n20135), .ZN(
        n13791) );
  AOI21_X1 U17114 ( .B1(n15809), .B2(n13792), .A(n13791), .ZN(n13795) );
  INV_X1 U17115 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20755) );
  NOR4_X1 U17116 ( .A1(n19940), .A2(n20982), .A3(n19939), .A4(n20755), .ZN(
        n13793) );
  NAND2_X1 U17117 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n13793), .ZN(n15817) );
  OAI211_X1 U17118 ( .C1(n13793), .C2(P1_REIP_REG_10__SCAN_IN), .A(n15817), 
        .B(n19972), .ZN(n13794) );
  OAI211_X1 U17119 ( .C1(n13798), .C2(n19947), .A(n13795), .B(n13794), .ZN(
        P1_U2830) );
  NOR2_X1 U17120 ( .A1(n20144), .A2(n16354), .ZN(n13796) );
  AOI21_X1 U17121 ( .B1(DATAI_10_), .B2(n20144), .A(n13796), .ZN(n20060) );
  INV_X1 U17122 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13797) );
  OAI222_X1 U17123 ( .A1(n14603), .A2(n13798), .B1(n14602), .B2(n20060), .C1(
        n13797), .C2(n14600), .ZN(P1_U2894) );
  XNOR2_X1 U17124 ( .A(n13800), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13801) );
  XNOR2_X1 U17125 ( .A(n9816), .B(n13801), .ZN(n15958) );
  AOI22_X1 U17126 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13802) );
  OAI21_X1 U17127 ( .B1(n20101), .B2(n13803), .A(n13802), .ZN(n13804) );
  AOI21_X1 U17128 ( .B1(n13805), .B2(n20096), .A(n13804), .ZN(n13806) );
  OAI21_X1 U17129 ( .B1(n15958), .B2(n19922), .A(n13806), .ZN(P1_U2991) );
  NAND2_X1 U17130 ( .A1(n14287), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n13809) );
  OAI21_X1 U17131 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13807), .A(
        n13835), .ZN(n15859) );
  AOI22_X1 U17132 ( .A1(n14282), .A2(n15859), .B1(n14286), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13808) );
  NAND2_X1 U17133 ( .A1(n13809), .A2(n13808), .ZN(n13810) );
  OAI21_X1 U17134 ( .B1(n13867), .B2(n13810), .A(n13865), .ZN(n13834) );
  AOI22_X1 U17135 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12203), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13814) );
  AOI22_X1 U17136 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12281), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13813) );
  AOI22_X1 U17137 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13812) );
  AOI22_X1 U17138 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13811) );
  NAND4_X1 U17139 ( .A1(n13814), .A2(n13813), .A3(n13812), .A4(n13811), .ZN(
        n13820) );
  AOI22_X1 U17140 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11906), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13818) );
  AOI22_X1 U17141 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13817) );
  AOI22_X1 U17142 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13816) );
  AOI22_X1 U17143 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13815) );
  NAND4_X1 U17144 ( .A1(n13818), .A2(n13817), .A3(n13816), .A4(n13815), .ZN(
        n13819) );
  OR2_X1 U17145 ( .A1(n13820), .A2(n13819), .ZN(n13821) );
  AND2_X1 U17146 ( .A1(n13951), .A2(n13821), .ZN(n13866) );
  XNOR2_X1 U17147 ( .A(n13834), .B(n13866), .ZN(n15856) );
  INV_X1 U17148 ( .A(n15856), .ZN(n13832) );
  INV_X1 U17149 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13823) );
  INV_X1 U17150 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n15048) );
  NOR2_X1 U17151 ( .A1(n20144), .A2(n15048), .ZN(n13822) );
  AOI21_X1 U17152 ( .B1(DATAI_11_), .B2(n20144), .A(n13822), .ZN(n20063) );
  OAI222_X1 U17153 ( .A1(n13832), .A2(n14603), .B1(n13823), .B2(n14600), .C1(
        n14602), .C2(n20063), .ZN(P1_U2893) );
  MUX2_X1 U17154 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n15951), .S(
        n15852), .Z(n13824) );
  XNOR2_X1 U17155 ( .A(n13825), .B(n13824), .ZN(n15947) );
  NAND2_X1 U17156 ( .A1(n15947), .A2(n20097), .ZN(n13829) );
  OAI22_X1 U17157 ( .A1(n14742), .A2(n19942), .B1(n20135), .B2(n20755), .ZN(
        n13826) );
  AOI21_X1 U17158 ( .B1(n15847), .B2(n13827), .A(n13826), .ZN(n13828) );
  OAI211_X1 U17159 ( .C1(n14748), .C2(n20016), .A(n13829), .B(n13828), .ZN(
        P1_U2990) );
  NOR2_X1 U17160 ( .A1(n9868), .A2(n13830), .ZN(n13831) );
  OR2_X1 U17161 ( .A1(n13918), .A2(n13831), .ZN(n15920) );
  INV_X1 U17162 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15818) );
  OAI222_X1 U17163 ( .A1(n15920), .A2(n20015), .B1(n15818), .B2(n20029), .C1(
        n13832), .C2(n14529), .ZN(P1_U2861) );
  INV_X1 U17164 ( .A(n13866), .ZN(n13833) );
  OAI21_X1 U17165 ( .B1(n13834), .B2(n13833), .A(n13865), .ZN(n13913) );
  XOR2_X1 U17166 ( .A(n13836), .B(n13835), .Z(n15846) );
  AOI22_X1 U17167 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n11906), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13840) );
  AOI22_X1 U17168 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12307), .B1(
        n12281), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13839) );
  AOI22_X1 U17169 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14053), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13838) );
  AOI22_X1 U17170 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13837) );
  NAND4_X1 U17171 ( .A1(n13840), .A2(n13839), .A3(n13838), .A4(n13837), .ZN(
        n13846) );
  AOI22_X1 U17172 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17173 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14015), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13843) );
  AOI22_X1 U17174 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13842) );
  AOI22_X1 U17175 ( .A1(n14186), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13841) );
  NAND4_X1 U17176 ( .A1(n13844), .A2(n13843), .A3(n13842), .A4(n13841), .ZN(
        n13845) );
  OAI21_X1 U17177 ( .B1(n13846), .B2(n13845), .A(n13951), .ZN(n13849) );
  NAND2_X1 U17178 ( .A1(n14287), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n13848) );
  NAND2_X1 U17179 ( .A1(n14286), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13847) );
  AND3_X1 U17180 ( .A1(n13849), .A2(n13848), .A3(n13847), .ZN(n13850) );
  OAI21_X1 U17181 ( .B1(n15846), .B2(n10352), .A(n13850), .ZN(n13914) );
  AND2_X1 U17182 ( .A1(n13913), .A2(n13914), .ZN(n13915) );
  XOR2_X1 U17183 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n13851), .Z(
        n14744) );
  AOI22_X1 U17184 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12203), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13855) );
  AOI22_X1 U17185 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11906), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13854) );
  AOI22_X1 U17186 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13853) );
  AOI22_X1 U17187 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13852) );
  NAND4_X1 U17188 ( .A1(n13855), .A2(n13854), .A3(n13853), .A4(n13852), .ZN(
        n13861) );
  AOI22_X1 U17189 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13859) );
  AOI22_X1 U17190 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13858) );
  AOI22_X1 U17191 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13857) );
  AOI22_X1 U17192 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13856) );
  NAND4_X1 U17193 ( .A1(n13859), .A2(n13858), .A3(n13857), .A4(n13856), .ZN(
        n13860) );
  OR2_X1 U17194 ( .A1(n13861), .A2(n13860), .ZN(n13862) );
  AOI22_X1 U17195 ( .A1(n13951), .A2(n13862), .B1(n14286), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13864) );
  NAND2_X1 U17196 ( .A1(n14287), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n13863) );
  OAI211_X1 U17197 ( .C1(n14744), .C2(n10352), .A(n13864), .B(n13863), .ZN(
        n13869) );
  OAI21_X1 U17198 ( .B1(n13915), .B2(n13869), .A(n13894), .ZN(n14747) );
  INV_X1 U17199 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20758) );
  INV_X1 U17200 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20760) );
  NOR3_X1 U17201 ( .A1(n20758), .A2(n20760), .A3(n15817), .ZN(n15765) );
  INV_X1 U17202 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20763) );
  NAND4_X1 U17203 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .A4(P1_REIP_REG_12__SCAN_IN), .ZN(n14229) );
  OAI21_X1 U17204 ( .B1(n14229), .B2(n13870), .A(n19972), .ZN(n15775) );
  INV_X1 U17205 ( .A(n15775), .ZN(n15810) );
  NAND2_X1 U17206 ( .A1(n13872), .A2(n13871), .ZN(n13873) );
  NAND2_X1 U17207 ( .A1(n13898), .A2(n13873), .ZN(n15919) );
  AOI21_X1 U17208 ( .B1(n19998), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n12122), .ZN(n13875) );
  AOI22_X1 U17209 ( .A1(n15809), .A2(n14744), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n19996), .ZN(n13874) );
  OAI211_X1 U17210 ( .C1(n20012), .C2(n15919), .A(n13875), .B(n13874), .ZN(
        n13876) );
  AOI221_X1 U17211 ( .B1(n15765), .B2(n20763), .C1(n15810), .C2(
        P1_REIP_REG_13__SCAN_IN), .A(n13876), .ZN(n13877) );
  OAI21_X1 U17212 ( .B1(n14747), .B2(n19947), .A(n13877), .ZN(P1_U2827) );
  XNOR2_X1 U17213 ( .A(n13878), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14729) );
  AOI22_X1 U17214 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11906), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13882) );
  AOI22_X1 U17215 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13881) );
  AOI22_X1 U17216 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13880) );
  AOI22_X1 U17217 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13879) );
  NAND4_X1 U17218 ( .A1(n13882), .A2(n13881), .A3(n13880), .A4(n13879), .ZN(
        n13888) );
  AOI22_X1 U17219 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13886) );
  AOI22_X1 U17220 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13885) );
  AOI22_X1 U17221 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13884) );
  AOI22_X1 U17222 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13883) );
  NAND4_X1 U17223 ( .A1(n13886), .A2(n13885), .A3(n13884), .A4(n13883), .ZN(
        n13887) );
  OAI21_X1 U17224 ( .B1(n13888), .B2(n13887), .A(n13951), .ZN(n13891) );
  NAND2_X1 U17225 ( .A1(n14287), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n13890) );
  NAND2_X1 U17226 ( .A1(n14286), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13889) );
  NAND3_X1 U17227 ( .A1(n13891), .A2(n13890), .A3(n13889), .ZN(n13892) );
  AOI21_X1 U17228 ( .B1(n14729), .B2(n14282), .A(n13892), .ZN(n13895) );
  AOI21_X1 U17229 ( .B1(n13895), .B2(n13894), .A(n13960), .ZN(n14731) );
  INV_X1 U17230 ( .A(n14731), .ZN(n13912) );
  AOI21_X1 U17231 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15765), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n13896) );
  INV_X1 U17232 ( .A(n13896), .ZN(n13904) );
  INV_X1 U17233 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20765) );
  NOR2_X1 U17234 ( .A1(n20765), .A2(n20763), .ZN(n14472) );
  OAI21_X1 U17235 ( .B1(n15816), .B2(n14472), .A(n15775), .ZN(n15799) );
  AND2_X1 U17236 ( .A1(n13898), .A2(n13897), .ZN(n13899) );
  OR2_X1 U17237 ( .A1(n13899), .A2(n9917), .ZN(n15910) );
  OAI21_X1 U17238 ( .B1(n13906), .B2(n19984), .A(n20135), .ZN(n13901) );
  NOR2_X1 U17239 ( .A1(n20002), .A2(n14729), .ZN(n13900) );
  AOI211_X1 U17240 ( .C1(n19998), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n13901), .B(n13900), .ZN(n13902) );
  OAI21_X1 U17241 ( .B1(n15910), .B2(n20012), .A(n13902), .ZN(n13903) );
  AOI21_X1 U17242 ( .B1(n13904), .B2(n15799), .A(n13903), .ZN(n13905) );
  OAI21_X1 U17243 ( .B1(n13912), .B2(n19947), .A(n13905), .ZN(P1_U2826) );
  OAI22_X1 U17244 ( .A1(n15910), .A2(n20015), .B1(n13906), .B2(n20029), .ZN(
        n13907) );
  AOI21_X1 U17245 ( .B1(n14731), .B2(n20025), .A(n13907), .ZN(n13908) );
  INV_X1 U17246 ( .A(n13908), .ZN(P1_U2858) );
  INV_X1 U17247 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n13911) );
  INV_X1 U17248 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13909) );
  NOR2_X1 U17249 ( .A1(n20144), .A2(n13909), .ZN(n13910) );
  AOI21_X1 U17250 ( .B1(DATAI_14_), .B2(n20144), .A(n13910), .ZN(n20072) );
  OAI222_X1 U17251 ( .A1(n13912), .A2(n14603), .B1(n13911), .B2(n14600), .C1(
        n14602), .C2(n20072), .ZN(P1_U2890) );
  INV_X1 U17252 ( .A(n13913), .ZN(n13917) );
  INV_X1 U17253 ( .A(n13914), .ZN(n13916) );
  AOI21_X1 U17254 ( .B1(n13917), .B2(n13916), .A(n13915), .ZN(n15845) );
  INV_X1 U17255 ( .A(n15845), .ZN(n13923) );
  XOR2_X1 U17256 ( .A(n13919), .B(n13918), .Z(n15808) );
  AOI22_X1 U17257 ( .A1(n15808), .A2(n20024), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14527), .ZN(n13920) );
  OAI21_X1 U17258 ( .B1(n13923), .B2(n14529), .A(n13920), .ZN(P1_U2860) );
  INV_X1 U17259 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n13922) );
  INV_X1 U17260 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n15039) );
  NOR2_X1 U17261 ( .A1(n20144), .A2(n15039), .ZN(n13921) );
  AOI21_X1 U17262 ( .B1(DATAI_12_), .B2(n20144), .A(n13921), .ZN(n20066) );
  OAI222_X1 U17263 ( .A1(n13923), .A2(n14603), .B1(n13922), .B2(n14600), .C1(
        n14602), .C2(n20066), .ZN(P1_U2892) );
  INV_X1 U17264 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14716) );
  XNOR2_X1 U17265 ( .A(n13924), .B(n14716), .ZN(n14718) );
  NAND2_X1 U17266 ( .A1(n14718), .A2(n14282), .ZN(n13941) );
  AOI22_X1 U17267 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13928) );
  AOI22_X1 U17268 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14149), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13927) );
  AOI22_X1 U17269 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12281), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13926) );
  AOI22_X1 U17270 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13925) );
  NAND4_X1 U17271 ( .A1(n13928), .A2(n13927), .A3(n13926), .A4(n13925), .ZN(
        n13937) );
  NAND2_X1 U17272 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13930) );
  NAND2_X1 U17273 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13929) );
  AND3_X1 U17274 ( .A1(n13930), .A2(n13929), .A3(n10352), .ZN(n13934) );
  AOI22_X1 U17275 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13933) );
  AOI22_X1 U17276 ( .A1(n14186), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13932) );
  AOI22_X1 U17277 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13931) );
  NAND4_X1 U17278 ( .A1(n13934), .A2(n13933), .A3(n13932), .A4(n13931), .ZN(
        n13936) );
  INV_X1 U17279 ( .A(n14933), .ZN(n13935) );
  NAND2_X1 U17280 ( .A1(n14260), .A2(n10352), .ZN(n14084) );
  OAI21_X1 U17281 ( .B1(n13937), .B2(n13936), .A(n14084), .ZN(n13939) );
  AOI22_X1 U17282 ( .A1(n14287), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13230), .ZN(n13938) );
  NAND2_X1 U17283 ( .A1(n13939), .A2(n13938), .ZN(n13940) );
  NAND2_X1 U17284 ( .A1(n13941), .A2(n13940), .ZN(n13962) );
  XOR2_X1 U17285 ( .A(n15803), .B(n13942), .Z(n15840) );
  INV_X1 U17286 ( .A(n15840), .ZN(n13958) );
  AOI22_X1 U17287 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12203), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13946) );
  AOI22_X1 U17288 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13945) );
  AOI22_X1 U17289 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12281), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13944) );
  AOI22_X1 U17290 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13943) );
  NAND4_X1 U17291 ( .A1(n13946), .A2(n13945), .A3(n13944), .A4(n13943), .ZN(
        n13953) );
  AOI22_X1 U17292 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13950) );
  AOI22_X1 U17293 ( .A1(n14186), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13949) );
  AOI22_X1 U17294 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13948) );
  AOI22_X1 U17295 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13947) );
  NAND4_X1 U17296 ( .A1(n13950), .A2(n13949), .A3(n13948), .A4(n13947), .ZN(
        n13952) );
  OAI21_X1 U17297 ( .B1(n13953), .B2(n13952), .A(n13951), .ZN(n13956) );
  NAND2_X1 U17298 ( .A1(n14287), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13955) );
  NAND2_X1 U17299 ( .A1(n14286), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13954) );
  NAND3_X1 U17300 ( .A1(n13956), .A2(n13955), .A3(n13954), .ZN(n13957) );
  AOI21_X1 U17301 ( .B1(n13958), .B2(n14282), .A(n13957), .ZN(n14597) );
  AOI21_X1 U17302 ( .B1(n13962), .B2(n13961), .A(n13997), .ZN(n14471) );
  OR2_X1 U17303 ( .A1(n14885), .A2(n13963), .ZN(n13964) );
  NAND2_X1 U17304 ( .A1(n14525), .A2(n13964), .ZN(n15899) );
  OAI22_X1 U17305 ( .A1(n15899), .A2(n20015), .B1(n13965), .B2(n20029), .ZN(
        n13966) );
  AOI21_X1 U17306 ( .B1(n14471), .B2(n20025), .A(n13966), .ZN(n13967) );
  INV_X1 U17307 ( .A(n13967), .ZN(P1_U2856) );
  INV_X1 U17308 ( .A(n13968), .ZN(n13970) );
  OAI21_X1 U17309 ( .B1(n13971), .B2(n18775), .A(n18617), .ZN(n13981) );
  NAND2_X1 U17310 ( .A1(n16434), .A2(n13981), .ZN(n18615) );
  NOR2_X1 U17311 ( .A1(n18824), .A2(n18615), .ZN(n13980) );
  NOR2_X1 U17312 ( .A1(n18693), .A2(n18607), .ZN(n13977) );
  INV_X1 U17313 ( .A(n13972), .ZN(n13973) );
  NAND2_X1 U17314 ( .A1(n18813), .A2(n17417), .ZN(n18665) );
  AOI21_X1 U17315 ( .B1(n13977), .B2(n17358), .A(n13974), .ZN(n13978) );
  NAND2_X1 U17316 ( .A1(n13976), .A2(n18613), .ZN(n15656) );
  OAI221_X1 U17317 ( .B1(n16434), .B2(n17417), .C1(n16434), .C2(n16819), .A(
        n13977), .ZN(n15659) );
  NAND3_X1 U17318 ( .A1(n13978), .A2(n15656), .A3(n15659), .ZN(n18636) );
  INV_X1 U17319 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16419) );
  NAND2_X1 U17320 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18809), .ZN(n18680) );
  NOR2_X1 U17321 ( .A1(n16419), .A2(n18680), .ZN(n13979) );
  NOR2_X1 U17322 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18515), .ZN(n18171) );
  AOI211_X2 U17323 ( .C1(n18663), .C2(n18636), .A(n13979), .B(n18171), .ZN(
        n18797) );
  MUX2_X1 U17324 ( .A(n13980), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18797), .Z(P3_U3284) );
  NOR2_X1 U17325 ( .A1(n17144), .A2(n13981), .ZN(n18158) );
  OAI221_X1 U17326 ( .B1(n18680), .B2(n18158), .C1(n18680), .C2(n16419), .A(
        n18251), .ZN(n18165) );
  INV_X1 U17327 ( .A(n18165), .ZN(n18161) );
  NOR2_X1 U17328 ( .A1(n18808), .A2(n17803), .ZN(n15667) );
  AOI21_X1 U17329 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15667), .ZN(n15668) );
  NOR2_X1 U17330 ( .A1(n18161), .A2(n15668), .ZN(n13983) );
  INV_X1 U17331 ( .A(n18512), .ZN(n18168) );
  INV_X1 U17332 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18412) );
  NAND2_X1 U17333 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18412), .ZN(n18210) );
  NAND2_X1 U17334 ( .A1(n18210), .A2(n18165), .ZN(n15666) );
  OR2_X1 U17335 ( .A1(n18168), .A2(n15666), .ZN(n13982) );
  MUX2_X1 U17336 ( .A(n13983), .B(n13982), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  XOR2_X1 U17337 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n13984), .Z(
        n15835) );
  AOI22_X1 U17338 ( .A1(n14287), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n14286), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13996) );
  AOI22_X1 U17339 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12203), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13988) );
  AOI22_X1 U17340 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13987) );
  AOI22_X1 U17341 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13986) );
  AOI22_X1 U17342 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13985) );
  NAND4_X1 U17343 ( .A1(n13988), .A2(n13987), .A3(n13986), .A4(n13985), .ZN(
        n13994) );
  AOI22_X1 U17344 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13992) );
  AOI22_X1 U17345 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13991) );
  AOI22_X1 U17346 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13990) );
  AOI22_X1 U17347 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13989) );
  NAND4_X1 U17348 ( .A1(n13992), .A2(n13991), .A3(n13990), .A4(n13989), .ZN(
        n13993) );
  OAI21_X1 U17349 ( .B1(n13994), .B2(n13993), .A(n14277), .ZN(n13995) );
  OAI211_X1 U17350 ( .C1(n15835), .C2(n10352), .A(n13996), .B(n13995), .ZN(
        n14522) );
  XNOR2_X1 U17351 ( .A(n13998), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15788) );
  NAND2_X1 U17352 ( .A1(n15788), .A2(n14282), .ZN(n14014) );
  AOI22_X1 U17353 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14002) );
  AOI22_X1 U17354 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11906), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14001) );
  AOI22_X1 U17355 ( .A1(n14186), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14000) );
  AOI22_X1 U17356 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13999) );
  NAND4_X1 U17357 ( .A1(n14002), .A2(n14001), .A3(n14000), .A4(n13999), .ZN(
        n14010) );
  AOI22_X1 U17358 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14008) );
  AOI22_X1 U17359 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14015), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14007) );
  NAND2_X1 U17360 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n14004) );
  NAND2_X1 U17361 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14003) );
  AND3_X1 U17362 ( .A1(n14004), .A2(n14003), .A3(n10352), .ZN(n14006) );
  AOI22_X1 U17363 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14005) );
  NAND4_X1 U17364 ( .A1(n14008), .A2(n14007), .A3(n14006), .A4(n14005), .ZN(
        n14009) );
  OAI21_X1 U17365 ( .B1(n14010), .B2(n14009), .A(n14084), .ZN(n14012) );
  AOI22_X1 U17366 ( .A1(n14287), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n13230), .ZN(n14011) );
  NAND2_X1 U17367 ( .A1(n14012), .A2(n14011), .ZN(n14013) );
  NAND2_X1 U17368 ( .A1(n14014), .A2(n14013), .ZN(n14517) );
  AOI22_X1 U17369 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14015), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14019) );
  AOI22_X1 U17370 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12281), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14018) );
  AOI22_X1 U17371 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14017) );
  AOI22_X1 U17372 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14016) );
  NAND4_X1 U17373 ( .A1(n14019), .A2(n14018), .A3(n14017), .A4(n14016), .ZN(
        n14025) );
  AOI22_X1 U17374 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14023) );
  AOI22_X1 U17375 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14022) );
  AOI22_X1 U17376 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14021) );
  AOI22_X1 U17377 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14020) );
  NAND4_X1 U17378 ( .A1(n14023), .A2(n14022), .A3(n14021), .A4(n14020), .ZN(
        n14024) );
  NOR2_X1 U17379 ( .A1(n14025), .A2(n14024), .ZN(n14029) );
  NAND2_X1 U17380 ( .A1(n13230), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14026) );
  NAND2_X1 U17381 ( .A1(n10352), .A2(n14026), .ZN(n14027) );
  AOI21_X1 U17382 ( .B1(n14287), .B2(P1_EAX_REG_19__SCAN_IN), .A(n14027), .ZN(
        n14028) );
  OAI21_X1 U17383 ( .B1(n14260), .B2(n14029), .A(n14028), .ZN(n14036) );
  INV_X1 U17384 ( .A(n14050), .ZN(n14034) );
  INV_X1 U17385 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14032) );
  INV_X1 U17386 ( .A(n14030), .ZN(n14031) );
  NAND2_X1 U17387 ( .A1(n14032), .A2(n14031), .ZN(n14033) );
  NAND2_X1 U17388 ( .A1(n14034), .A2(n14033), .ZN(n15834) );
  NAND2_X1 U17389 ( .A1(n14036), .A2(n14035), .ZN(n14510) );
  AOI22_X1 U17390 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14053), .B1(
        n12314), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14040) );
  AOI22_X1 U17391 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11906), .B1(
        n14149), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14039) );
  AOI22_X1 U17392 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14038) );
  AOI22_X1 U17393 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14037) );
  NAND4_X1 U17394 ( .A1(n14040), .A2(n14039), .A3(n14038), .A4(n14037), .ZN(
        n14046) );
  AOI22_X1 U17395 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12203), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14044) );
  AOI22_X1 U17396 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12281), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14043) );
  AOI22_X1 U17397 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14042) );
  AOI22_X1 U17398 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12282), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14041) );
  NAND4_X1 U17399 ( .A1(n14044), .A2(n14043), .A3(n14042), .A4(n14041), .ZN(
        n14045) );
  NOR2_X1 U17400 ( .A1(n14046), .A2(n14045), .ZN(n14049) );
  INV_X1 U17401 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15773) );
  AOI21_X1 U17402 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15773), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14047) );
  AOI21_X1 U17403 ( .B1(n14287), .B2(P1_EAX_REG_20__SCAN_IN), .A(n14047), .ZN(
        n14048) );
  OAI21_X1 U17404 ( .B1(n14260), .B2(n14049), .A(n14048), .ZN(n14052) );
  XNOR2_X1 U17405 ( .A(n14050), .B(n15773), .ZN(n15763) );
  NAND2_X1 U17406 ( .A1(n15763), .A2(n14282), .ZN(n14051) );
  AOI22_X1 U17407 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14057) );
  AOI22_X1 U17408 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14056) );
  AOI22_X1 U17409 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14055) );
  AOI22_X1 U17410 ( .A1(n12282), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14054) );
  NAND4_X1 U17411 ( .A1(n14057), .A2(n14056), .A3(n14055), .A4(n14054), .ZN(
        n14063) );
  AOI22_X1 U17412 ( .A1(n14149), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11906), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14061) );
  AOI22_X1 U17413 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14060) );
  AOI22_X1 U17414 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14059) );
  AOI22_X1 U17415 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14058) );
  NAND4_X1 U17416 ( .A1(n14061), .A2(n14060), .A3(n14059), .A4(n14058), .ZN(
        n14062) );
  NOR2_X1 U17417 ( .A1(n14063), .A2(n14062), .ZN(n14067) );
  NAND2_X1 U17418 ( .A1(n13230), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14064) );
  NAND2_X1 U17419 ( .A1(n10352), .A2(n14064), .ZN(n14065) );
  AOI21_X1 U17420 ( .B1(n14287), .B2(P1_EAX_REG_21__SCAN_IN), .A(n14065), .ZN(
        n14066) );
  OAI21_X1 U17421 ( .B1(n14260), .B2(n14067), .A(n14066), .ZN(n14073) );
  INV_X1 U17422 ( .A(n14068), .ZN(n14070) );
  INV_X1 U17423 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14069) );
  NAND2_X1 U17424 ( .A1(n14070), .A2(n14069), .ZN(n14071) );
  NAND2_X1 U17425 ( .A1(n14089), .A2(n14071), .ZN(n15762) );
  AOI22_X1 U17426 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14077) );
  AOI22_X1 U17427 ( .A1(n14186), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14076) );
  AOI22_X1 U17428 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14075) );
  AOI22_X1 U17429 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14074) );
  NAND4_X1 U17430 ( .A1(n14077), .A2(n14076), .A3(n14075), .A4(n14074), .ZN(
        n14086) );
  AOI22_X1 U17431 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12314), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U17432 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14015), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14082) );
  NAND2_X1 U17433 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n14079) );
  NAND2_X1 U17434 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14078) );
  AND3_X1 U17435 ( .A1(n14079), .A2(n14078), .A3(n10352), .ZN(n14081) );
  AOI22_X1 U17436 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14080) );
  NAND4_X1 U17437 ( .A1(n14083), .A2(n14082), .A3(n14081), .A4(n14080), .ZN(
        n14085) );
  OAI21_X1 U17438 ( .B1(n14086), .B2(n14085), .A(n14084), .ZN(n14088) );
  AOI22_X1 U17439 ( .A1(n14287), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n13230), .ZN(n14087) );
  NAND2_X1 U17440 ( .A1(n14088), .A2(n14087), .ZN(n14091) );
  XNOR2_X1 U17441 ( .A(n14089), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15742) );
  NAND2_X1 U17442 ( .A1(n15742), .A2(n14282), .ZN(n14090) );
  NAND2_X1 U17443 ( .A1(n14091), .A2(n14090), .ZN(n14492) );
  AOI22_X1 U17444 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14096) );
  AOI22_X1 U17445 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14095) );
  AOI22_X1 U17446 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14094) );
  AOI22_X1 U17447 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14093) );
  NAND4_X1 U17448 ( .A1(n14096), .A2(n14095), .A3(n14094), .A4(n14093), .ZN(
        n14102) );
  AOI22_X1 U17449 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14100) );
  AOI22_X1 U17450 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14099) );
  AOI22_X1 U17451 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14098) );
  AOI22_X1 U17452 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14097) );
  NAND4_X1 U17453 ( .A1(n14100), .A2(n14099), .A3(n14098), .A4(n14097), .ZN(
        n14101) );
  NOR2_X1 U17454 ( .A1(n14102), .A2(n14101), .ZN(n14123) );
  AOI22_X1 U17455 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12287), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14106) );
  AOI22_X1 U17456 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14105) );
  AOI22_X1 U17457 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U17458 ( .A1(n14199), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14103) );
  NAND4_X1 U17459 ( .A1(n14106), .A2(n14105), .A3(n14104), .A4(n14103), .ZN(
        n14112) );
  AOI22_X1 U17460 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14110) );
  AOI22_X1 U17461 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14109) );
  AOI22_X1 U17462 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14108) );
  AOI22_X1 U17463 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14107) );
  NAND4_X1 U17464 ( .A1(n14110), .A2(n14109), .A3(n14108), .A4(n14107), .ZN(
        n14111) );
  NOR2_X1 U17465 ( .A1(n14112), .A2(n14111), .ZN(n14122) );
  XNOR2_X1 U17466 ( .A(n14123), .B(n14122), .ZN(n14116) );
  NAND2_X1 U17467 ( .A1(n13230), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14113) );
  NAND2_X1 U17468 ( .A1(n10352), .A2(n14113), .ZN(n14114) );
  AOI21_X1 U17469 ( .B1(n14287), .B2(P1_EAX_REG_23__SCAN_IN), .A(n14114), .ZN(
        n14115) );
  OAI21_X1 U17470 ( .B1(n14260), .B2(n14116), .A(n14115), .ZN(n14121) );
  NAND2_X1 U17471 ( .A1(n14118), .A2(n14117), .ZN(n14119) );
  NAND2_X1 U17472 ( .A1(n14138), .A2(n14119), .ZN(n14673) );
  NAND2_X1 U17473 ( .A1(n14121), .A2(n14120), .ZN(n14463) );
  NOR2_X1 U17474 ( .A1(n14123), .A2(n14122), .ZN(n14157) );
  AOI22_X1 U17475 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14127) );
  AOI22_X1 U17476 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14126) );
  AOI22_X1 U17477 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14125) );
  AOI22_X1 U17478 ( .A1(n14199), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14124) );
  NAND4_X1 U17479 ( .A1(n14127), .A2(n14126), .A3(n14125), .A4(n14124), .ZN(
        n14133) );
  AOI22_X1 U17480 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14131) );
  AOI22_X1 U17481 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14130) );
  AOI22_X1 U17482 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14129) );
  AOI22_X1 U17483 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14128) );
  NAND4_X1 U17484 ( .A1(n14131), .A2(n14130), .A3(n14129), .A4(n14128), .ZN(
        n14132) );
  OR2_X1 U17485 ( .A1(n14133), .A2(n14132), .ZN(n14156) );
  INV_X1 U17486 ( .A(n14156), .ZN(n14134) );
  XNOR2_X1 U17487 ( .A(n14157), .B(n14134), .ZN(n14135) );
  NAND2_X1 U17488 ( .A1(n14135), .A2(n14277), .ZN(n14141) );
  NAND2_X1 U17489 ( .A1(n13230), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14136) );
  NAND2_X1 U17490 ( .A1(n10352), .A2(n14136), .ZN(n14137) );
  AOI21_X1 U17491 ( .B1(n14287), .B2(P1_EAX_REG_24__SCAN_IN), .A(n14137), .ZN(
        n14140) );
  XNOR2_X1 U17492 ( .A(n14138), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14665) );
  AOI21_X1 U17493 ( .B1(n14141), .B2(n14140), .A(n14139), .ZN(n14443) );
  INV_X1 U17494 ( .A(n14142), .ZN(n14144) );
  OAI21_X1 U17495 ( .B1(n14144), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14143), .ZN(n14657) );
  AOI22_X1 U17496 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14148) );
  AOI22_X1 U17497 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14147) );
  AOI22_X1 U17498 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14146) );
  AOI22_X1 U17499 ( .A1(n14186), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14145) );
  NAND4_X1 U17500 ( .A1(n14148), .A2(n14147), .A3(n14146), .A4(n14145), .ZN(
        n14155) );
  AOI22_X1 U17501 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14153) );
  AOI22_X1 U17502 ( .A1(n12287), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14149), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14152) );
  AOI22_X1 U17503 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14151) );
  AOI22_X1 U17504 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14150) );
  NAND4_X1 U17505 ( .A1(n14153), .A2(n14152), .A3(n14151), .A4(n14150), .ZN(
        n14154) );
  NOR2_X1 U17506 ( .A1(n14155), .A2(n14154), .ZN(n14173) );
  NAND2_X1 U17507 ( .A1(n14157), .A2(n14156), .ZN(n14172) );
  XNOR2_X1 U17508 ( .A(n14173), .B(n14172), .ZN(n14160) );
  AOI21_X1 U17509 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n13230), .A(
        n14282), .ZN(n14159) );
  NAND2_X1 U17510 ( .A1(n14287), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n14158) );
  OAI211_X1 U17511 ( .C1(n14160), .C2(n14260), .A(n14159), .B(n14158), .ZN(
        n14161) );
  AOI22_X1 U17512 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14165) );
  AOI22_X1 U17513 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14164) );
  AOI22_X1 U17514 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14163) );
  AOI22_X1 U17515 ( .A1(n14199), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14162) );
  NAND4_X1 U17516 ( .A1(n14165), .A2(n14164), .A3(n14163), .A4(n14162), .ZN(
        n14171) );
  AOI22_X1 U17517 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14169) );
  AOI22_X1 U17518 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14168) );
  AOI22_X1 U17519 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14167) );
  AOI22_X1 U17520 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14166) );
  NAND4_X1 U17521 ( .A1(n14169), .A2(n14168), .A3(n14167), .A4(n14166), .ZN(
        n14170) );
  OR2_X1 U17522 ( .A1(n14171), .A2(n14170), .ZN(n14193) );
  NOR2_X1 U17523 ( .A1(n14173), .A2(n14172), .ZN(n14194) );
  XOR2_X1 U17524 ( .A(n14193), .B(n14194), .Z(n14174) );
  NAND2_X1 U17525 ( .A1(n14174), .A2(n14277), .ZN(n14178) );
  INV_X1 U17526 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14647) );
  NOR2_X1 U17527 ( .A1(n14647), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14175) );
  AOI211_X1 U17528 ( .C1(n14287), .C2(P1_EAX_REG_26__SCAN_IN), .A(n14282), .B(
        n14175), .ZN(n14177) );
  XOR2_X1 U17529 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B(n14176), .Z(
        n14651) );
  AOI22_X1 U17530 ( .A1(n14178), .A2(n14177), .B1(n14282), .B2(n14651), .ZN(
        n14416) );
  NAND2_X1 U17531 ( .A1(n14180), .A2(n14179), .ZN(n14181) );
  NAND2_X1 U17532 ( .A1(n14214), .A2(n14181), .ZN(n14640) );
  AOI22_X1 U17533 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14185) );
  AOI22_X1 U17534 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12281), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14184) );
  AOI22_X1 U17535 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14183) );
  AOI22_X1 U17536 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14182) );
  NAND4_X1 U17537 ( .A1(n14185), .A2(n14184), .A3(n14183), .A4(n14182), .ZN(
        n14192) );
  AOI22_X1 U17538 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11906), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14190) );
  AOI22_X1 U17539 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14189) );
  AOI22_X1 U17540 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14188) );
  AOI22_X1 U17541 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12306), .B1(
        n14186), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14187) );
  NAND4_X1 U17542 ( .A1(n14190), .A2(n14189), .A3(n14188), .A4(n14187), .ZN(
        n14191) );
  NOR2_X1 U17543 ( .A1(n14192), .A2(n14191), .ZN(n14211) );
  NAND2_X1 U17544 ( .A1(n14194), .A2(n14193), .ZN(n14210) );
  XNOR2_X1 U17545 ( .A(n14211), .B(n14210), .ZN(n14197) );
  AOI21_X1 U17546 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n13230), .A(
        n14282), .ZN(n14196) );
  NAND2_X1 U17547 ( .A1(n14287), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n14195) );
  OAI211_X1 U17548 ( .C1(n14197), .C2(n14260), .A(n14196), .B(n14195), .ZN(
        n14198) );
  AOI22_X1 U17549 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14203) );
  AOI22_X1 U17550 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14202) );
  AOI22_X1 U17551 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14201) );
  AOI22_X1 U17552 ( .A1(n14199), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14200) );
  NAND4_X1 U17553 ( .A1(n14203), .A2(n14202), .A3(n14201), .A4(n14200), .ZN(
        n14209) );
  AOI22_X1 U17554 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14207) );
  AOI22_X1 U17555 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14206) );
  AOI22_X1 U17556 ( .A1(n9820), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14205) );
  AOI22_X1 U17557 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14204) );
  NAND4_X1 U17558 ( .A1(n14207), .A2(n14206), .A3(n14205), .A4(n14204), .ZN(
        n14208) );
  OR2_X1 U17559 ( .A1(n14209), .A2(n14208), .ZN(n14246) );
  NOR2_X1 U17560 ( .A1(n14211), .A2(n14210), .ZN(n14247) );
  XOR2_X1 U17561 ( .A(n14246), .B(n14247), .Z(n14212) );
  NAND2_X1 U17562 ( .A1(n14212), .A2(n14277), .ZN(n14217) );
  NOR2_X1 U17563 ( .A1(n14629), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14213) );
  AOI211_X1 U17564 ( .C1(n14287), .C2(P1_EAX_REG_28__SCAN_IN), .A(n14282), .B(
        n14213), .ZN(n14216) );
  INV_X1 U17565 ( .A(n14214), .ZN(n14215) );
  XOR2_X1 U17566 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n14215), .Z(
        n14633) );
  AOI22_X1 U17567 ( .A1(n14217), .A2(n14216), .B1(n14282), .B2(n14633), .ZN(
        n14219) );
  OAI21_X2 U17568 ( .B1(n14218), .B2(n14219), .A(n14394), .ZN(n14630) );
  NAND2_X1 U17569 ( .A1(n14600), .A2(n14220), .ZN(n14223) );
  INV_X1 U17570 ( .A(n14223), .ZN(n14221) );
  NAND3_X1 U17571 ( .A1(n14600), .A2(n20199), .A3(n11986), .ZN(n14555) );
  OAI22_X1 U17572 ( .A1(n14555), .A2(n20066), .B1(n14600), .B2(n13435), .ZN(
        n14222) );
  AOI21_X1 U17573 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14557), .A(n14222), .ZN(
        n14225) );
  NOR2_X2 U17574 ( .A1(n14223), .A2(n20145), .ZN(n14593) );
  NAND2_X1 U17575 ( .A1(n14593), .A2(DATAI_28_), .ZN(n14224) );
  OAI211_X1 U17576 ( .C1(n14630), .C2(n14603), .A(n14225), .B(n14224), .ZN(
        P1_U2876) );
  NOR2_X1 U17577 ( .A1(n14404), .A2(n14226), .ZN(n14227) );
  NOR2_X1 U17578 ( .A1(n14379), .A2(n14227), .ZN(n14779) );
  AOI22_X1 U17579 ( .A1(n14779), .A2(n20024), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n14527), .ZN(n14228) );
  OAI21_X1 U17580 ( .B1(n14630), .B2(n14529), .A(n14228), .ZN(P1_U2844) );
  INV_X1 U17581 ( .A(n14633), .ZN(n14239) );
  INV_X1 U17582 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20948) );
  INV_X1 U17583 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20776) );
  NAND4_X1 U17584 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .A4(n14472), .ZN(n15764) );
  NAND2_X1 U17585 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15774) );
  NOR4_X1 U17586 ( .A1(n20776), .A2(n14229), .A3(n15764), .A4(n15774), .ZN(
        n15740) );
  NAND2_X1 U17587 ( .A1(n14230), .A2(n15740), .ZN(n15752) );
  NOR2_X1 U17588 ( .A1(n20948), .A2(n15752), .ZN(n14464) );
  NAND3_X1 U17589 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(n14464), .ZN(n14232) );
  OR2_X1 U17590 ( .A1(n19940), .A2(n14232), .ZN(n14451) );
  NAND3_X1 U17591 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(P1_REIP_REG_24__SCAN_IN), .ZN(n14231) );
  INV_X1 U17592 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20789) );
  NOR2_X1 U17593 ( .A1(n14409), .A2(n20789), .ZN(n14236) );
  INV_X1 U17594 ( .A(n14232), .ZN(n14233) );
  NAND2_X1 U17595 ( .A1(n19951), .A2(n14233), .ZN(n14447) );
  INV_X1 U17596 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20783) );
  NOR2_X1 U17597 ( .A1(n14447), .A2(n20783), .ZN(n14438) );
  AND2_X1 U17598 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14369) );
  INV_X1 U17599 ( .A(n14369), .ZN(n14234) );
  NAND2_X1 U17600 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14387) );
  NOR2_X1 U17601 ( .A1(n14234), .A2(n14387), .ZN(n14235) );
  AOI21_X1 U17602 ( .B1(n14438), .B2(n14235), .A(n15816), .ZN(n14401) );
  OAI21_X1 U17603 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14236), .A(n14401), 
        .ZN(n14238) );
  AOI22_X1 U17604 ( .A1(n19998), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n19996), .B2(P1_EBX_REG_28__SCAN_IN), .ZN(n14237) );
  OAI211_X1 U17605 ( .C1(n20002), .C2(n14239), .A(n14238), .B(n14237), .ZN(
        n14240) );
  AOI21_X1 U17606 ( .B1(n14779), .B2(n19988), .A(n14240), .ZN(n14241) );
  OAI21_X1 U17607 ( .B1(n14630), .B2(n19947), .A(n14241), .ZN(P1_U2812) );
  INV_X1 U17608 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20213) );
  INV_X1 U17609 ( .A(n14242), .ZN(n14244) );
  INV_X1 U17610 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14243) );
  NAND2_X1 U17611 ( .A1(n14244), .A2(n14243), .ZN(n14245) );
  NAND2_X1 U17612 ( .A1(n14281), .A2(n14245), .ZN(n14617) );
  NAND2_X1 U17613 ( .A1(n14247), .A2(n14246), .ZN(n14263) );
  AOI22_X1 U17614 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14251) );
  AOI22_X1 U17615 ( .A1(n12307), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14250) );
  AOI22_X1 U17616 ( .A1(n12288), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14249) );
  AOI22_X1 U17617 ( .A1(n14053), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14248) );
  NAND4_X1 U17618 ( .A1(n14251), .A2(n14250), .A3(n14249), .A4(n14248), .ZN(
        n14257) );
  AOI22_X1 U17619 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12203), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14255) );
  AOI22_X1 U17620 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11906), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14254) );
  AOI22_X1 U17621 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14253) );
  AOI22_X1 U17622 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14252) );
  NAND4_X1 U17623 ( .A1(n14255), .A2(n14254), .A3(n14253), .A4(n14252), .ZN(
        n14256) );
  NOR2_X1 U17624 ( .A1(n14257), .A2(n14256), .ZN(n14264) );
  XNOR2_X1 U17625 ( .A(n14263), .B(n14264), .ZN(n14261) );
  AOI21_X1 U17626 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n13230), .A(
        n14282), .ZN(n14259) );
  NAND2_X1 U17627 ( .A1(n14287), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n14258) );
  OAI211_X1 U17628 ( .C1(n14261), .C2(n14260), .A(n14259), .B(n14258), .ZN(
        n14262) );
  OAI21_X1 U17629 ( .B1(n10352), .B2(n14617), .A(n14262), .ZN(n14396) );
  NOR2_X1 U17630 ( .A1(n14264), .A2(n14263), .ZN(n14276) );
  AOI22_X1 U17631 ( .A1(n12281), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12307), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14268) );
  AOI22_X1 U17632 ( .A1(n14015), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12282), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14267) );
  AOI22_X1 U17633 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14266) );
  AOI22_X1 U17634 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14265) );
  NAND4_X1 U17635 ( .A1(n14268), .A2(n14267), .A3(n14266), .A4(n14265), .ZN(
        n14274) );
  AOI22_X1 U17636 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14053), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14272) );
  AOI22_X1 U17637 ( .A1(n12203), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12288), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14271) );
  AOI22_X1 U17638 ( .A1(n9791), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14270) );
  AOI22_X1 U17639 ( .A1(n11906), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12309), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14269) );
  NAND4_X1 U17640 ( .A1(n14272), .A2(n14271), .A3(n14270), .A4(n14269), .ZN(
        n14273) );
  NOR2_X1 U17641 ( .A1(n14274), .A2(n14273), .ZN(n14275) );
  XNOR2_X1 U17642 ( .A(n14276), .B(n14275), .ZN(n14278) );
  NAND2_X1 U17643 ( .A1(n14278), .A2(n14277), .ZN(n14285) );
  INV_X1 U17644 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14279) );
  AOI21_X1 U17645 ( .B1(n14279), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14280) );
  AOI21_X1 U17646 ( .B1(n14287), .B2(P1_EAX_REG_30__SCAN_IN), .A(n14280), .ZN(
        n14284) );
  XNOR2_X1 U17647 ( .A(n14281), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14386) );
  AOI21_X1 U17648 ( .B1(n14285), .B2(n14284), .A(n14283), .ZN(n14378) );
  AOI22_X1 U17649 ( .A1(n14287), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n14286), .ZN(n14288) );
  INV_X1 U17650 ( .A(n14288), .ZN(n14289) );
  NAND3_X1 U17651 ( .A1(n14367), .A2(n20214), .A3(n14600), .ZN(n14291) );
  AOI22_X1 U17652 ( .A1(n14593), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14587), .ZN(n14290) );
  OAI211_X1 U17653 ( .C1(n14591), .C2(n20213), .A(n14291), .B(n14290), .ZN(
        P1_U2873) );
  INV_X1 U17654 ( .A(n14292), .ZN(n14295) );
  INV_X1 U17655 ( .A(n14293), .ZN(n14294) );
  NAND2_X1 U17656 ( .A1(n14295), .A2(n14294), .ZN(n14608) );
  NAND2_X1 U17657 ( .A1(n14605), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14296) );
  OAI22_X2 U17658 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n14608), .B1(
        n14297), .B2(n14296), .ZN(n14298) );
  XNOR2_X1 U17659 ( .A(n14298), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14769) );
  INV_X1 U17660 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20794) );
  NOR2_X1 U17661 ( .A1(n20135), .A2(n20794), .ZN(n14765) );
  AOI21_X1 U17662 ( .B1(n20090), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14765), .ZN(n14299) );
  OAI21_X1 U17663 ( .B1(n20101), .B2(n14300), .A(n14299), .ZN(n14301) );
  OAI21_X1 U17664 ( .B1(n14769), .B2(n19922), .A(n14302), .ZN(P1_U2968) );
  AOI22_X1 U17665 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14306) );
  AOI22_X1 U17666 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12780), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14305) );
  NAND2_X1 U17667 ( .A1(n14306), .A2(n14305), .ZN(n14320) );
  AOI21_X1 U17668 ( .B1(n10878), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n14313), .ZN(n14308) );
  AOI22_X1 U17669 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14307) );
  OAI211_X1 U17670 ( .C1(n12635), .C2(n14309), .A(n14308), .B(n14307), .ZN(
        n14319) );
  AOI22_X1 U17671 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14310), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14312) );
  AOI22_X1 U17672 ( .A1(n10868), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10878), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14311) );
  NAND2_X1 U17673 ( .A1(n14312), .A2(n14311), .ZN(n14318) );
  AOI22_X1 U17674 ( .A1(n10867), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10880), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14316) );
  NAND2_X1 U17675 ( .A1(n12780), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n14315) );
  NAND2_X1 U17676 ( .A1(n10865), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14314) );
  NAND4_X1 U17677 ( .A1(n14316), .A2(n14315), .A3(n14314), .A4(n14313), .ZN(
        n14317) );
  OAI22_X1 U17678 ( .A1(n14320), .A2(n14319), .B1(n14318), .B2(n14317), .ZN(
        n14321) );
  XNOR2_X1 U17679 ( .A(n14322), .B(n14321), .ZN(n14332) );
  INV_X1 U17680 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n14324) );
  AOI22_X1 U17681 ( .A1(n19088), .A2(n19104), .B1(n19125), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14323) );
  OAI21_X1 U17682 ( .B1(n15054), .B2(n14324), .A(n14323), .ZN(n14327) );
  NOR2_X1 U17683 ( .A1(n14325), .A2(n19092), .ZN(n14326) );
  AOI211_X1 U17684 ( .C1(n19089), .C2(BUF1_REG_30__SCAN_IN), .A(n14327), .B(
        n14326), .ZN(n14328) );
  OAI21_X1 U17685 ( .B1(n14332), .B2(n19093), .A(n14328), .ZN(P2_U2889) );
  NOR2_X1 U17686 ( .A1(n14329), .A2(n14984), .ZN(n14330) );
  AOI21_X1 U17687 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n14984), .A(n14330), .ZN(
        n14331) );
  OAI21_X1 U17688 ( .B1(n14332), .B2(n15038), .A(n14331), .ZN(P2_U2857) );
  OAI21_X1 U17689 ( .B1(n14335), .B2(n14334), .A(n14333), .ZN(n14351) );
  NAND2_X1 U17690 ( .A1(n19236), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14350) );
  OAI21_X1 U17691 ( .B1(n14351), .B2(n16199), .A(n14350), .ZN(n14336) );
  NOR2_X1 U17692 ( .A1(n14337), .A2(n14336), .ZN(n14347) );
  NOR2_X1 U17693 ( .A1(n15437), .A2(n9801), .ZN(n14339) );
  OAI21_X1 U17694 ( .B1(n14340), .B2(n14339), .A(n14338), .ZN(n14346) );
  NAND2_X1 U17695 ( .A1(n14342), .A2(n14341), .ZN(n14355) );
  NAND3_X1 U17696 ( .A1(n14356), .A2(n16196), .A3(n14355), .ZN(n14345) );
  NAND2_X1 U17697 ( .A1(n14343), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14344) );
  NAND4_X1 U17698 ( .A1(n14347), .A2(n14346), .A3(n14345), .A4(n14344), .ZN(
        n14348) );
  AOI21_X1 U17699 ( .B1(n19862), .B2(n16192), .A(n14348), .ZN(n14349) );
  OAI21_X1 U17700 ( .B1(n14359), .B2(n16194), .A(n14349), .ZN(P2_U3044) );
  OAI21_X1 U17701 ( .B1(n14351), .B2(n16145), .A(n14350), .ZN(n14354) );
  NOR2_X1 U17702 ( .A1(n19247), .A2(n14352), .ZN(n14353) );
  AOI211_X1 U17703 ( .C1(n19237), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14354), .B(n14353), .ZN(n14358) );
  NAND3_X1 U17704 ( .A1(n14356), .A2(n19242), .A3(n14355), .ZN(n14357) );
  OAI211_X1 U17705 ( .C1(n16130), .C2(n14359), .A(n14358), .B(n14357), .ZN(
        P2_U3012) );
  AND2_X1 U17706 ( .A1(n14360), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14361) );
  AOI21_X1 U17707 ( .B1(n14364), .B2(P1_EBX_REG_30__SCAN_IN), .A(n14361), .ZN(
        n14384) );
  AOI22_X1 U17708 ( .A1(n14364), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n12028), .ZN(n14365) );
  XNOR2_X1 U17709 ( .A(n14366), .B(n14365), .ZN(n14756) );
  NAND2_X1 U17710 ( .A1(n14367), .A2(n19965), .ZN(n14377) );
  NAND2_X1 U17711 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14368) );
  NOR2_X1 U17712 ( .A1(n14387), .A2(n14368), .ZN(n14372) );
  NAND2_X1 U17713 ( .A1(n14438), .A2(n14369), .ZN(n14370) );
  NAND2_X1 U17714 ( .A1(n14370), .A2(n19972), .ZN(n14408) );
  OAI21_X1 U17715 ( .B1(n15816), .B2(n14372), .A(n14408), .ZN(n14388) );
  OAI22_X1 U17716 ( .A1(n19986), .A2(n14371), .B1(n14480), .B2(n19984), .ZN(
        n14375) );
  INV_X1 U17717 ( .A(n14372), .ZN(n14373) );
  NOR3_X1 U17718 ( .A1(n14409), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14373), 
        .ZN(n14374) );
  AOI211_X1 U17719 ( .C1(n14388), .C2(P1_REIP_REG_31__SCAN_IN), .A(n14375), 
        .B(n14374), .ZN(n14376) );
  OAI211_X1 U17720 ( .C1(n14756), .C2(n20012), .A(n14377), .B(n14376), .ZN(
        P1_U2809) );
  XOR2_X1 U17721 ( .A(n14378), .B(n14395), .Z(n14613) );
  INV_X1 U17722 ( .A(n14613), .ZN(n14534) );
  INV_X1 U17723 ( .A(n14379), .ZN(n14381) );
  OAI22_X1 U17724 ( .A1(n14383), .A2(n14382), .B1(n14381), .B2(n14380), .ZN(
        n14385) );
  XNOR2_X1 U17725 ( .A(n14385), .B(n14384), .ZN(n14776) );
  INV_X1 U17726 ( .A(n14386), .ZN(n14611) );
  OR2_X1 U17727 ( .A1(n14409), .A2(n14387), .ZN(n14397) );
  NOR2_X1 U17728 ( .A1(n14397), .A2(n20792), .ZN(n14389) );
  OAI21_X1 U17729 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14389), .A(n14388), 
        .ZN(n14391) );
  AOI22_X1 U17730 ( .A1(n19998), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n19996), .ZN(n14390) );
  OAI211_X1 U17731 ( .C1(n14611), .C2(n20002), .A(n14391), .B(n14390), .ZN(
        n14392) );
  AOI21_X1 U17732 ( .B1(n14776), .B2(n19988), .A(n14392), .ZN(n14393) );
  OAI21_X1 U17733 ( .B1(n14534), .B2(n19947), .A(n14393), .ZN(P1_U2810) );
  AOI21_X1 U17734 ( .B1(n14396), .B2(n14394), .A(n14395), .ZN(n14619) );
  NAND2_X1 U17735 ( .A1(n14619), .A2(n19965), .ZN(n14403) );
  NOR2_X1 U17736 ( .A1(n14397), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14400) );
  AOI22_X1 U17737 ( .A1(n19998), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n19996), .B2(P1_EBX_REG_29__SCAN_IN), .ZN(n14398) );
  OAI21_X1 U17738 ( .B1(n14617), .B2(n20002), .A(n14398), .ZN(n14399) );
  AOI211_X1 U17739 ( .C1(n14401), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14400), 
        .B(n14399), .ZN(n14402) );
  OAI211_X1 U17740 ( .C1(n20012), .C2(n14482), .A(n14403), .B(n14402), .ZN(
        P1_U2811) );
  OAI21_X1 U17741 ( .B1(n14405), .B2(n14418), .A(n10179), .ZN(n14789) );
  AOI21_X1 U17742 ( .B1(n14407), .B2(n14406), .A(n14218), .ZN(n14642) );
  NAND2_X1 U17743 ( .A1(n14642), .A2(n19965), .ZN(n14414) );
  INV_X1 U17744 ( .A(n14408), .ZN(n14421) );
  NOR2_X1 U17745 ( .A1(n14409), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14412) );
  AOI22_X1 U17746 ( .A1(n19998), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n19996), .B2(P1_EBX_REG_27__SCAN_IN), .ZN(n14410) );
  OAI21_X1 U17747 ( .B1(n14640), .B2(n20002), .A(n14410), .ZN(n14411) );
  AOI211_X1 U17748 ( .C1(n14421), .C2(P1_REIP_REG_27__SCAN_IN), .A(n14412), 
        .B(n14411), .ZN(n14413) );
  OAI211_X1 U17749 ( .C1(n20012), .C2(n14789), .A(n14414), .B(n14413), .ZN(
        P1_U2813) );
  OAI21_X1 U17750 ( .B1(n14415), .B2(n14416), .A(n14406), .ZN(n14648) );
  AND2_X1 U17751 ( .A1(n14431), .A2(n14417), .ZN(n14419) );
  OR2_X1 U17752 ( .A1(n14419), .A2(n14418), .ZN(n14802) );
  INV_X1 U17753 ( .A(n14802), .ZN(n14427) );
  INV_X1 U17754 ( .A(n14651), .ZN(n14425) );
  NAND2_X1 U17755 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14420) );
  NOR2_X1 U17756 ( .A1(n14451), .A2(n14420), .ZN(n14422) );
  OAI21_X1 U17757 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n14422), .A(n14421), 
        .ZN(n14424) );
  AOI22_X1 U17758 ( .A1(n19998), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n19996), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n14423) );
  OAI211_X1 U17759 ( .C1(n20002), .C2(n14425), .A(n14424), .B(n14423), .ZN(
        n14426) );
  AOI21_X1 U17760 ( .B1(n14427), .B2(n19988), .A(n14426), .ZN(n14428) );
  OAI21_X1 U17761 ( .B1(n14648), .B2(n19947), .A(n14428), .ZN(P1_U2814) );
  AOI21_X1 U17762 ( .B1(n14430), .B2(n14429), .A(n14415), .ZN(n14659) );
  INV_X1 U17763 ( .A(n14659), .ZN(n14552) );
  INV_X1 U17764 ( .A(n14431), .ZN(n14432) );
  AOI21_X1 U17765 ( .B1(n14433), .B2(n14456), .A(n14432), .ZN(n14811) );
  OAI22_X1 U17766 ( .A1(n14434), .A2(n19986), .B1(n20002), .B2(n14657), .ZN(
        n14440) );
  NAND2_X1 U17767 ( .A1(n19972), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14437) );
  NOR3_X1 U17768 ( .A1(n14451), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n20783), 
        .ZN(n14435) );
  AOI21_X1 U17769 ( .B1(P1_EBX_REG_25__SCAN_IN), .B2(n19996), .A(n14435), .ZN(
        n14436) );
  OAI21_X1 U17770 ( .B1(n14438), .B2(n14437), .A(n14436), .ZN(n14439) );
  AOI211_X1 U17771 ( .C1(n14811), .C2(n19988), .A(n14440), .B(n14439), .ZN(
        n14441) );
  OAI21_X1 U17772 ( .B1(n14552), .B2(n19947), .A(n14441), .ZN(P1_U2815) );
  OR2_X1 U17773 ( .A1(n14442), .A2(n14443), .ZN(n14444) );
  AND2_X1 U17774 ( .A1(n14429), .A2(n14444), .ZN(n14669) );
  INV_X1 U17775 ( .A(n14669), .ZN(n14560) );
  INV_X1 U17776 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14446) );
  INV_X1 U17777 ( .A(n14665), .ZN(n14445) );
  OAI22_X1 U17778 ( .A1(n14446), .A2(n19986), .B1(n20002), .B2(n14445), .ZN(
        n14453) );
  OR2_X1 U17779 ( .A1(n19984), .A2(n14489), .ZN(n14450) );
  INV_X1 U17780 ( .A(n14447), .ZN(n14448) );
  NOR2_X1 U17781 ( .A1(n15816), .A2(n14448), .ZN(n14467) );
  NAND2_X1 U17782 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14467), .ZN(n14449) );
  OAI211_X1 U17783 ( .C1(n14451), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14450), 
        .B(n14449), .ZN(n14452) );
  NOR2_X1 U17784 ( .A1(n14453), .A2(n14452), .ZN(n14458) );
  OR2_X1 U17785 ( .A1(n14461), .A2(n14454), .ZN(n14455) );
  AND2_X1 U17786 ( .A1(n14456), .A2(n14455), .ZN(n14818) );
  NAND2_X1 U17787 ( .A1(n14818), .A2(n19988), .ZN(n14457) );
  OAI211_X1 U17788 ( .C1(n14560), .C2(n19947), .A(n14458), .B(n14457), .ZN(
        P1_U2816) );
  NOR2_X1 U17789 ( .A1(n9895), .A2(n14459), .ZN(n14460) );
  OR2_X1 U17790 ( .A1(n14461), .A2(n14460), .ZN(n14823) );
  AOI21_X1 U17791 ( .B1(n14463), .B2(n14462), .A(n14442), .ZN(n14675) );
  NAND2_X1 U17792 ( .A1(n14675), .A2(n19965), .ZN(n14470) );
  INV_X1 U17793 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20779) );
  NAND2_X1 U17794 ( .A1(n15741), .A2(n14464), .ZN(n15744) );
  INV_X1 U17795 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20781) );
  OAI21_X1 U17796 ( .B1(n20779), .B2(n15744), .A(n20781), .ZN(n14468) );
  NOR2_X1 U17797 ( .A1(n20002), .A2(n14673), .ZN(n14466) );
  INV_X1 U17798 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14490) );
  OAI22_X1 U17799 ( .A1(n19986), .A2(n14117), .B1(n19984), .B2(n14490), .ZN(
        n14465) );
  AOI211_X1 U17800 ( .C1(n14468), .C2(n14467), .A(n14466), .B(n14465), .ZN(
        n14469) );
  OAI211_X1 U17801 ( .C1(n20012), .C2(n14823), .A(n14470), .B(n14469), .ZN(
        P1_U2817) );
  INV_X1 U17802 ( .A(n14471), .ZN(n14721) );
  INV_X1 U17803 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20767) );
  NAND2_X1 U17804 ( .A1(n14472), .A2(n15765), .ZN(n14473) );
  NOR2_X1 U17805 ( .A1(n20767), .A2(n14473), .ZN(n15794) );
  INV_X1 U17806 ( .A(n15794), .ZN(n14475) );
  NOR2_X1 U17807 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14473), .ZN(n15805) );
  NOR2_X1 U17808 ( .A1(n15805), .A2(n15799), .ZN(n14474) );
  MUX2_X1 U17809 ( .A(n14475), .B(n14474), .S(P1_REIP_REG_16__SCAN_IN), .Z(
        n14479) );
  AOI22_X1 U17810 ( .A1(n14718), .A2(n15809), .B1(n19996), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n14476) );
  OAI21_X1 U17811 ( .B1(n20012), .B2(n15899), .A(n14476), .ZN(n14477) );
  AOI211_X1 U17812 ( .C1(n19998), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n14477), .B(n12122), .ZN(n14478) );
  OAI211_X1 U17813 ( .C1(n14721), .C2(n19947), .A(n14479), .B(n14478), .ZN(
        P1_U2824) );
  OAI22_X1 U17814 ( .A1(n14756), .A2(n20015), .B1(n20029), .B2(n14480), .ZN(
        P1_U2841) );
  AOI22_X1 U17815 ( .A1(n14776), .A2(n20024), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n14527), .ZN(n14481) );
  OAI21_X1 U17816 ( .B1(n14534), .B2(n14529), .A(n14481), .ZN(P1_U2842) );
  INV_X1 U17817 ( .A(n14619), .ZN(n14540) );
  INV_X1 U17818 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14483) );
  OAI222_X1 U17819 ( .A1(n14529), .A2(n14540), .B1(n14483), .B2(n20029), .C1(
        n14482), .C2(n20015), .ZN(P1_U2843) );
  INV_X1 U17820 ( .A(n14642), .ZN(n14544) );
  INV_X1 U17821 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14484) );
  OAI222_X1 U17822 ( .A1(n14529), .A2(n14544), .B1(n14484), .B2(n20029), .C1(
        n14789), .C2(n20015), .ZN(P1_U2845) );
  OAI222_X1 U17823 ( .A1(n14529), .A2(n14648), .B1(n14485), .B2(n20029), .C1(
        n14802), .C2(n20015), .ZN(P1_U2846) );
  AOI22_X1 U17824 ( .A1(n14811), .A2(n20024), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n14527), .ZN(n14486) );
  OAI21_X1 U17825 ( .B1(n14552), .B2(n14529), .A(n14486), .ZN(P1_U2847) );
  NAND2_X1 U17826 ( .A1(n14669), .A2(n20025), .ZN(n14488) );
  NAND2_X1 U17827 ( .A1(n14818), .A2(n20024), .ZN(n14487) );
  OAI211_X1 U17828 ( .C1(n14489), .C2(n20029), .A(n14488), .B(n14487), .ZN(
        P1_U2848) );
  INV_X1 U17829 ( .A(n14675), .ZN(n14565) );
  OAI222_X1 U17830 ( .A1(n14529), .A2(n14565), .B1(n14490), .B2(n20029), .C1(
        n14823), .C2(n20015), .ZN(P1_U2849) );
  INV_X1 U17831 ( .A(n14462), .ZN(n14491) );
  AOI21_X1 U17832 ( .B1(n14492), .B2(n14495), .A(n14491), .ZN(n14683) );
  INV_X1 U17833 ( .A(n14683), .ZN(n15747) );
  AOI21_X1 U17834 ( .B1(n14493), .B2(n14497), .A(n9895), .ZN(n15745) );
  AOI22_X1 U17835 ( .A1(n15745), .A2(n20024), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14527), .ZN(n14494) );
  OAI21_X1 U17836 ( .B1(n15747), .B2(n14529), .A(n14494), .ZN(P1_U2850) );
  OAI21_X1 U17837 ( .B1(n14504), .B2(n14496), .A(n14495), .ZN(n14688) );
  INV_X1 U17838 ( .A(n14497), .ZN(n14498) );
  AOI21_X1 U17839 ( .B1(n14499), .B2(n14506), .A(n14498), .ZN(n15758) );
  AOI22_X1 U17840 ( .A1(n15758), .A2(n20024), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14527), .ZN(n14500) );
  OAI21_X1 U17841 ( .B1(n14688), .B2(n14529), .A(n14500), .ZN(P1_U2851) );
  NOR2_X1 U17842 ( .A1(n14501), .A2(n14502), .ZN(n14503) );
  OR2_X1 U17843 ( .A1(n14504), .A2(n14503), .ZN(n15767) );
  INV_X1 U17844 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14508) );
  OR2_X1 U17845 ( .A1(n14514), .A2(n14505), .ZN(n14507) );
  AND2_X1 U17846 ( .A1(n14507), .A2(n14506), .ZN(n14852) );
  INV_X1 U17847 ( .A(n14852), .ZN(n15766) );
  OAI222_X1 U17848 ( .A1(n14529), .A2(n15767), .B1(n20029), .B2(n14508), .C1(
        n15766), .C2(n20015), .ZN(P1_U2852) );
  AND2_X1 U17849 ( .A1(n10261), .A2(n14510), .ZN(n14511) );
  OR2_X1 U17850 ( .A1(n14511), .A2(n14501), .ZN(n15779) );
  AND2_X1 U17851 ( .A1(n14520), .A2(n14512), .ZN(n14513) );
  NOR2_X1 U17852 ( .A1(n14514), .A2(n14513), .ZN(n15877) );
  AOI22_X1 U17853 ( .A1(n15877), .A2(n20024), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14527), .ZN(n14515) );
  OAI21_X1 U17854 ( .B1(n15779), .B2(n14529), .A(n14515), .ZN(P1_U2853) );
  AOI21_X1 U17855 ( .B1(n14517), .B2(n14516), .A(n14509), .ZN(n14705) );
  INV_X1 U17856 ( .A(n14705), .ZN(n15785) );
  INV_X1 U17857 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14521) );
  NAND2_X1 U17858 ( .A1(n14523), .A2(n14518), .ZN(n14519) );
  NAND2_X1 U17859 ( .A1(n14520), .A2(n14519), .ZN(n15884) );
  OAI222_X1 U17860 ( .A1(n15785), .A2(n14529), .B1(n20029), .B2(n14521), .C1(
        n15884), .C2(n20015), .ZN(P1_U2854) );
  OAI21_X1 U17861 ( .B1(n13997), .B2(n14522), .A(n14516), .ZN(n15791) );
  INV_X1 U17862 ( .A(n14523), .ZN(n14524) );
  AOI21_X1 U17863 ( .B1(n14526), .B2(n14525), .A(n14524), .ZN(n15792) );
  AOI22_X1 U17864 ( .A1(n15792), .A2(n20024), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14527), .ZN(n14528) );
  OAI21_X1 U17865 ( .B1(n15791), .B2(n14529), .A(n14528), .ZN(P1_U2855) );
  OAI222_X1 U17866 ( .A1(n15919), .A2(n20015), .B1(n20029), .B2(n12072), .C1(
        n14747), .C2(n14529), .ZN(P1_U2859) );
  OAI22_X1 U17867 ( .A1(n14555), .A2(n20072), .B1(n14600), .B2(n14530), .ZN(
        n14531) );
  AOI21_X1 U17868 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n14557), .A(n14531), .ZN(
        n14533) );
  NAND2_X1 U17869 ( .A1(n14593), .A2(DATAI_30_), .ZN(n14532) );
  OAI211_X1 U17870 ( .C1(n14534), .C2(n14603), .A(n14533), .B(n14532), .ZN(
        P1_U2874) );
  NOR2_X1 U17871 ( .A1(n20144), .A2(n14535), .ZN(n14536) );
  AOI21_X1 U17872 ( .B1(DATAI_13_), .B2(n20144), .A(n14536), .ZN(n20069) );
  OAI22_X1 U17873 ( .A1(n14555), .A2(n20069), .B1(n14600), .B2(n13437), .ZN(
        n14537) );
  AOI21_X1 U17874 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14557), .A(n14537), .ZN(
        n14539) );
  NAND2_X1 U17875 ( .A1(n14593), .A2(DATAI_29_), .ZN(n14538) );
  OAI211_X1 U17876 ( .C1(n14540), .C2(n14603), .A(n14539), .B(n14538), .ZN(
        P1_U2875) );
  OAI22_X1 U17877 ( .A1(n14555), .A2(n20063), .B1(n14600), .B2(n13308), .ZN(
        n14541) );
  AOI21_X1 U17878 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14557), .A(n14541), .ZN(
        n14543) );
  NAND2_X1 U17879 ( .A1(n14593), .A2(DATAI_27_), .ZN(n14542) );
  OAI211_X1 U17880 ( .C1(n14544), .C2(n14603), .A(n14543), .B(n14542), .ZN(
        P1_U2877) );
  OAI22_X1 U17881 ( .A1(n14555), .A2(n20060), .B1(n14600), .B2(n13298), .ZN(
        n14545) );
  AOI21_X1 U17882 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n14557), .A(n14545), .ZN(
        n14547) );
  NAND2_X1 U17883 ( .A1(n14593), .A2(DATAI_26_), .ZN(n14546) );
  OAI211_X1 U17884 ( .C1(n14648), .C2(n14603), .A(n14547), .B(n14546), .ZN(
        P1_U2878) );
  INV_X1 U17885 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20168) );
  INV_X1 U17886 ( .A(n14555), .ZN(n14588) );
  AOI22_X1 U17887 ( .A1(n14588), .A2(n14548), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n14587), .ZN(n14549) );
  OAI21_X1 U17888 ( .B1(n20168), .B2(n14591), .A(n14549), .ZN(n14550) );
  AOI21_X1 U17889 ( .B1(n14593), .B2(DATAI_25_), .A(n14550), .ZN(n14551) );
  OAI21_X1 U17890 ( .B1(n14552), .B2(n14603), .A(n14551), .ZN(P1_U2879) );
  INV_X1 U17891 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14553) );
  OAI22_X1 U17892 ( .A1(n14555), .A2(n14554), .B1(n14600), .B2(n14553), .ZN(
        n14556) );
  AOI21_X1 U17893 ( .B1(BUF1_REG_24__SCAN_IN), .B2(n14557), .A(n14556), .ZN(
        n14559) );
  NAND2_X1 U17894 ( .A1(n14593), .A2(DATAI_24_), .ZN(n14558) );
  OAI211_X1 U17895 ( .C1(n14560), .C2(n14603), .A(n14559), .B(n14558), .ZN(
        P1_U2880) );
  INV_X1 U17896 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n14562) );
  AOI22_X1 U17897 ( .A1(n14588), .A2(n20217), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n14587), .ZN(n14561) );
  OAI21_X1 U17898 ( .B1(n14591), .B2(n14562), .A(n14561), .ZN(n14563) );
  AOI21_X1 U17899 ( .B1(n14593), .B2(DATAI_23_), .A(n14563), .ZN(n14564) );
  OAI21_X1 U17900 ( .B1(n14565), .B2(n14603), .A(n14564), .ZN(P1_U2881) );
  INV_X1 U17901 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14567) );
  AOI22_X1 U17902 ( .A1(n14588), .A2(n20206), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n14587), .ZN(n14566) );
  OAI21_X1 U17903 ( .B1(n14591), .B2(n14567), .A(n14566), .ZN(n14568) );
  AOI21_X1 U17904 ( .B1(n14593), .B2(DATAI_22_), .A(n14568), .ZN(n14569) );
  OAI21_X1 U17905 ( .B1(n15747), .B2(n14603), .A(n14569), .ZN(P1_U2882) );
  INV_X1 U17906 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n14571) );
  AOI22_X1 U17907 ( .A1(n14588), .A2(n20200), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n14587), .ZN(n14570) );
  OAI21_X1 U17908 ( .B1(n14591), .B2(n14571), .A(n14570), .ZN(n14572) );
  AOI21_X1 U17909 ( .B1(n14593), .B2(DATAI_21_), .A(n14572), .ZN(n14573) );
  OAI21_X1 U17910 ( .B1(n14688), .B2(n14603), .A(n14573), .ZN(P1_U2883) );
  AOI22_X1 U17911 ( .A1(n14588), .A2(n20193), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n14587), .ZN(n14574) );
  OAI21_X1 U17912 ( .B1(n14591), .B2(n20189), .A(n14574), .ZN(n14575) );
  AOI21_X1 U17913 ( .B1(n14593), .B2(DATAI_20_), .A(n14575), .ZN(n14576) );
  OAI21_X1 U17914 ( .B1(n15767), .B2(n14603), .A(n14576), .ZN(P1_U2884) );
  AOI22_X1 U17915 ( .A1(n14588), .A2(n20186), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n14587), .ZN(n14577) );
  OAI21_X1 U17916 ( .B1(n14591), .B2(n20181), .A(n14577), .ZN(n14578) );
  AOI21_X1 U17917 ( .B1(n14593), .B2(DATAI_19_), .A(n14578), .ZN(n14579) );
  OAI21_X1 U17918 ( .B1(n15779), .B2(n14603), .A(n14579), .ZN(P1_U2885) );
  AOI22_X1 U17919 ( .A1(n14588), .A2(n20178), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n14587), .ZN(n14580) );
  OAI21_X1 U17920 ( .B1(n14591), .B2(n20173), .A(n14580), .ZN(n14581) );
  AOI21_X1 U17921 ( .B1(n14593), .B2(DATAI_18_), .A(n14581), .ZN(n14582) );
  OAI21_X1 U17922 ( .B1(n15785), .B2(n14603), .A(n14582), .ZN(P1_U2886) );
  INV_X1 U17923 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14584) );
  AOI22_X1 U17924 ( .A1(n14588), .A2(n20170), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n14587), .ZN(n14583) );
  OAI21_X1 U17925 ( .B1(n14591), .B2(n14584), .A(n14583), .ZN(n14585) );
  AOI21_X1 U17926 ( .B1(n14593), .B2(DATAI_17_), .A(n14585), .ZN(n14586) );
  OAI21_X1 U17927 ( .B1(n15791), .B2(n14603), .A(n14586), .ZN(P1_U2887) );
  INV_X1 U17928 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14590) );
  AOI22_X1 U17929 ( .A1(n14588), .A2(n20159), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n14587), .ZN(n14589) );
  OAI21_X1 U17930 ( .B1(n14591), .B2(n14590), .A(n14589), .ZN(n14592) );
  AOI21_X1 U17931 ( .B1(n14593), .B2(DATAI_16_), .A(n14592), .ZN(n14594) );
  OAI21_X1 U17932 ( .B1(n14721), .B2(n14603), .A(n14594), .ZN(P1_U2888) );
  INV_X1 U17933 ( .A(n13961), .ZN(n14595) );
  AOI21_X1 U17934 ( .B1(n14597), .B2(n14596), .A(n14595), .ZN(n15841) );
  INV_X1 U17935 ( .A(n15841), .ZN(n14599) );
  OAI222_X1 U17936 ( .A1(n14603), .A2(n14599), .B1(n14600), .B2(n13384), .C1(
        n14602), .C2(n14598), .ZN(P1_U2889) );
  INV_X1 U17937 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14601) );
  OAI222_X1 U17938 ( .A1(n14603), .A2(n14747), .B1(n14602), .B2(n20069), .C1(
        n14601), .C2(n14600), .ZN(P1_U2891) );
  INV_X1 U17939 ( .A(n14604), .ZN(n14606) );
  NAND2_X1 U17940 ( .A1(n14606), .A2(n14605), .ZN(n14607) );
  NAND2_X1 U17941 ( .A1(n14608), .A2(n14607), .ZN(n14609) );
  XNOR2_X1 U17942 ( .A(n14609), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14778) );
  INV_X1 U17943 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20797) );
  NOR2_X1 U17944 ( .A1(n20135), .A2(n20797), .ZN(n14775) );
  AOI21_X1 U17945 ( .B1(n20090), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14775), .ZN(n14610) );
  OAI21_X1 U17946 ( .B1(n20101), .B2(n14611), .A(n14610), .ZN(n14612) );
  AOI21_X1 U17947 ( .B1(n14613), .B2(n20096), .A(n14612), .ZN(n14614) );
  OAI21_X1 U17948 ( .B1(n14778), .B2(n19922), .A(n14614), .ZN(P1_U2969) );
  AOI21_X1 U17949 ( .B1(n20090), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14615), .ZN(n14616) );
  OAI21_X1 U17950 ( .B1(n20101), .B2(n14617), .A(n14616), .ZN(n14618) );
  AOI21_X1 U17951 ( .B1(n14619), .B2(n20096), .A(n14618), .ZN(n14620) );
  OAI21_X1 U17952 ( .B1(n14621), .B2(n19922), .A(n14620), .ZN(P1_U2970) );
  NAND2_X1 U17953 ( .A1(n14622), .A2(n14798), .ZN(n14627) );
  NAND2_X1 U17954 ( .A1(n15852), .A2(n14624), .ZN(n14644) );
  NAND3_X1 U17955 ( .A1(n14623), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n14644), .ZN(n14626) );
  MUX2_X1 U17956 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n14798), .S(
        n15852), .Z(n14625) );
  AOI21_X1 U17957 ( .B1(n14627), .B2(n14626), .A(n14625), .ZN(n14628) );
  XNOR2_X1 U17958 ( .A(n14628), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14786) );
  NAND2_X1 U17959 ( .A1(n12122), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14780) );
  OAI21_X1 U17960 ( .B1(n14742), .B2(n14629), .A(n14780), .ZN(n14632) );
  NOR2_X1 U17961 ( .A1(n14630), .A2(n14748), .ZN(n14631) );
  OAI21_X1 U17962 ( .B1(n19922), .B2(n14786), .A(n14634), .ZN(P1_U2971) );
  MUX2_X1 U17963 ( .A(n14637), .B(n14636), .S(n10332), .Z(n14638) );
  XOR2_X1 U17964 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n14638), .Z(
        n14795) );
  NAND2_X1 U17965 ( .A1(n12122), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14787) );
  NAND2_X1 U17966 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14639) );
  OAI211_X1 U17967 ( .C1(n20101), .C2(n14640), .A(n14787), .B(n14639), .ZN(
        n14641) );
  AOI21_X1 U17968 ( .B1(n14642), .B2(n20096), .A(n14641), .ZN(n14643) );
  OAI21_X1 U17969 ( .B1(n19922), .B2(n14795), .A(n14643), .ZN(P1_U2972) );
  NOR2_X1 U17970 ( .A1(n14661), .A2(n10332), .ZN(n14645) );
  OAI21_X1 U17971 ( .B1(n14645), .B2(n14622), .A(n14644), .ZN(n14646) );
  XNOR2_X1 U17972 ( .A(n14646), .B(n14798), .ZN(n14806) );
  NAND2_X1 U17973 ( .A1(n12122), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14800) );
  OAI21_X1 U17974 ( .B1(n14742), .B2(n14647), .A(n14800), .ZN(n14650) );
  NOR2_X1 U17975 ( .A1(n14648), .A2(n14748), .ZN(n14649) );
  AOI211_X1 U17976 ( .C1(n15847), .C2(n14651), .A(n14650), .B(n14649), .ZN(
        n14652) );
  OAI21_X1 U17977 ( .B1(n19922), .B2(n14806), .A(n14652), .ZN(P1_U2973) );
  AND2_X1 U17978 ( .A1(n14654), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14662) );
  NAND2_X1 U17979 ( .A1(n14662), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14655) );
  NAND2_X1 U17980 ( .A1(n12122), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14807) );
  NAND2_X1 U17981 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14656) );
  OAI211_X1 U17982 ( .C1(n20101), .C2(n14657), .A(n14807), .B(n14656), .ZN(
        n14658) );
  AOI21_X1 U17983 ( .B1(n14659), .B2(n20096), .A(n14658), .ZN(n14660) );
  OAI21_X1 U17984 ( .B1(n19922), .B2(n14814), .A(n14660), .ZN(P1_U2974) );
  NAND2_X1 U17985 ( .A1(n14661), .A2(n10332), .ZN(n14663) );
  MUX2_X1 U17986 ( .A(n14663), .B(n10332), .S(n14662), .Z(n14664) );
  XNOR2_X1 U17987 ( .A(n14664), .B(n14819), .ZN(n14822) );
  NOR2_X1 U17988 ( .A1(n20135), .A2(n20783), .ZN(n14817) );
  AOI21_X1 U17989 ( .B1(n20090), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14817), .ZN(n14667) );
  NAND2_X1 U17990 ( .A1(n15847), .A2(n14665), .ZN(n14666) );
  NAND2_X1 U17991 ( .A1(n14667), .A2(n14666), .ZN(n14668) );
  AOI21_X1 U17992 ( .B1(n14669), .B2(n20096), .A(n14668), .ZN(n14670) );
  OAI21_X1 U17993 ( .B1(n14822), .B2(n19922), .A(n14670), .ZN(P1_U2975) );
  XNOR2_X1 U17994 ( .A(n15852), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14671) );
  XNOR2_X1 U17995 ( .A(n14623), .B(n14671), .ZN(n14831) );
  NAND2_X1 U17996 ( .A1(n12122), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14824) );
  NAND2_X1 U17997 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14672) );
  OAI211_X1 U17998 ( .C1(n20101), .C2(n14673), .A(n14824), .B(n14672), .ZN(
        n14674) );
  AOI21_X1 U17999 ( .B1(n14675), .B2(n20096), .A(n14674), .ZN(n14676) );
  OAI21_X1 U18000 ( .B1(n14831), .B2(n19922), .A(n14676), .ZN(P1_U2976) );
  NAND2_X1 U18001 ( .A1(n14678), .A2(n14677), .ZN(n14679) );
  XNOR2_X1 U18002 ( .A(n14679), .B(n14833), .ZN(n14838) );
  INV_X1 U18003 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14681) );
  NAND2_X1 U18004 ( .A1(n15847), .A2(n15742), .ZN(n14680) );
  NAND2_X1 U18005 ( .A1(n12122), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14832) );
  OAI211_X1 U18006 ( .C1(n14742), .C2(n14681), .A(n14680), .B(n14832), .ZN(
        n14682) );
  AOI21_X1 U18007 ( .B1(n14683), .B2(n20096), .A(n14682), .ZN(n14684) );
  OAI21_X1 U18008 ( .B1(n19922), .B2(n14838), .A(n14684), .ZN(P1_U2977) );
  NOR2_X1 U18009 ( .A1(n14685), .A2(n15852), .ZN(n14692) );
  NOR2_X1 U18010 ( .A1(n14686), .A2(n10332), .ZN(n14693) );
  MUX2_X1 U18011 ( .A(n14692), .B(n14693), .S(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n14687) );
  XNOR2_X1 U18012 ( .A(n14687), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14845) );
  INV_X1 U18013 ( .A(n14688), .ZN(n15759) );
  NAND2_X1 U18014 ( .A1(n12122), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14839) );
  NAND2_X1 U18015 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14689) );
  OAI211_X1 U18016 ( .C1(n20101), .C2(n15762), .A(n14839), .B(n14689), .ZN(
        n14690) );
  AOI21_X1 U18017 ( .B1(n15759), .B2(n20096), .A(n14690), .ZN(n14691) );
  OAI21_X1 U18018 ( .B1(n14845), .B2(n19922), .A(n14691), .ZN(P1_U2978) );
  NOR2_X1 U18019 ( .A1(n14693), .A2(n14692), .ZN(n14694) );
  XOR2_X1 U18020 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n14694), .Z(
        n14855) );
  NOR2_X1 U18021 ( .A1(n20135), .A2(n20776), .ZN(n14851) );
  NOR2_X1 U18022 ( .A1(n14742), .A2(n15773), .ZN(n14695) );
  AOI211_X1 U18023 ( .C1(n15847), .C2(n15763), .A(n14851), .B(n14695), .ZN(
        n14698) );
  INV_X1 U18024 ( .A(n15767), .ZN(n14696) );
  NAND2_X1 U18025 ( .A1(n14696), .A2(n20096), .ZN(n14697) );
  OAI211_X1 U18026 ( .C1(n14855), .C2(n19922), .A(n14698), .B(n14697), .ZN(
        P1_U2979) );
  OAI21_X1 U18027 ( .B1(n14701), .B2(n14700), .A(n14699), .ZN(n15885) );
  INV_X1 U18028 ( .A(n15788), .ZN(n14703) );
  AOI22_X1 U18029 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14702) );
  OAI21_X1 U18030 ( .B1(n14703), .B2(n20101), .A(n14702), .ZN(n14704) );
  AOI21_X1 U18031 ( .B1(n14705), .B2(n20096), .A(n14704), .ZN(n14706) );
  OAI21_X1 U18032 ( .B1(n19922), .B2(n15885), .A(n14706), .ZN(P1_U2981) );
  INV_X1 U18033 ( .A(n15851), .ZN(n14710) );
  INV_X1 U18034 ( .A(n14707), .ZN(n14709) );
  AOI21_X1 U18035 ( .B1(n14710), .B2(n14709), .A(n14708), .ZN(n14877) );
  INV_X1 U18036 ( .A(n14711), .ZN(n14712) );
  NAND3_X1 U18037 ( .A1(n14877), .A2(n14712), .A3(n14878), .ZN(n14879) );
  NAND2_X1 U18038 ( .A1(n14879), .A2(n14878), .ZN(n14714) );
  XNOR2_X1 U18039 ( .A(n14714), .B(n14713), .ZN(n15896) );
  NAND2_X1 U18040 ( .A1(n15896), .A2(n20097), .ZN(n14720) );
  INV_X1 U18041 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14715) );
  OAI22_X1 U18042 ( .A1(n14742), .A2(n14716), .B1(n20135), .B2(n14715), .ZN(
        n14717) );
  AOI21_X1 U18043 ( .B1(n14718), .B2(n15847), .A(n14717), .ZN(n14719) );
  OAI211_X1 U18044 ( .C1(n14748), .C2(n14721), .A(n14720), .B(n14719), .ZN(
        P1_U2983) );
  NAND2_X1 U18045 ( .A1(n15851), .A2(n14722), .ZN(n14859) );
  NAND3_X1 U18046 ( .A1(n14859), .A2(n14723), .A3(n14733), .ZN(n14725) );
  NAND2_X1 U18047 ( .A1(n14725), .A2(n14724), .ZN(n14727) );
  XNOR2_X1 U18048 ( .A(n15852), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14726) );
  XNOR2_X1 U18049 ( .A(n14727), .B(n14726), .ZN(n15900) );
  AOI22_X1 U18050 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14728) );
  OAI21_X1 U18051 ( .B1(n20101), .B2(n14729), .A(n14728), .ZN(n14730) );
  AOI21_X1 U18052 ( .B1(n14731), .B2(n20096), .A(n14730), .ZN(n14732) );
  OAI21_X1 U18053 ( .B1(n15900), .B2(n19922), .A(n14732), .ZN(P1_U2985) );
  INV_X1 U18054 ( .A(n14733), .ZN(n14735) );
  OAI22_X1 U18055 ( .A1(n15851), .A2(n14735), .B1(n14734), .B2(n15852), .ZN(
        n14891) );
  INV_X1 U18056 ( .A(n14738), .ZN(n14736) );
  OAI21_X1 U18057 ( .B1(n15852), .B2(n14737), .A(n14736), .ZN(n14890) );
  NOR2_X1 U18058 ( .A1(n14891), .A2(n14890), .ZN(n14889) );
  NOR2_X1 U18059 ( .A1(n14889), .A2(n14738), .ZN(n14740) );
  XNOR2_X1 U18060 ( .A(n14740), .B(n14739), .ZN(n15916) );
  NAND2_X1 U18061 ( .A1(n15916), .A2(n20097), .ZN(n14746) );
  INV_X1 U18062 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14741) );
  OAI22_X1 U18063 ( .A1(n14742), .A2(n14741), .B1(n20135), .B2(n20763), .ZN(
        n14743) );
  AOI21_X1 U18064 ( .B1(n15847), .B2(n14744), .A(n14743), .ZN(n14745) );
  OAI211_X1 U18065 ( .C1(n14748), .C2(n14747), .A(n14746), .B(n14745), .ZN(
        P1_U2986) );
  MUX2_X1 U18066 ( .A(n14749), .B(n15851), .S(n15852), .Z(n14750) );
  XNOR2_X1 U18067 ( .A(n14750), .B(n12061), .ZN(n15934) );
  AOI22_X1 U18068 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14751) );
  OAI21_X1 U18069 ( .B1(n20101), .B2(n14752), .A(n14751), .ZN(n14753) );
  AOI21_X1 U18070 ( .B1(n14754), .B2(n20096), .A(n14753), .ZN(n14755) );
  OAI21_X1 U18071 ( .B1(n15934), .B2(n19922), .A(n14755), .ZN(P1_U2989) );
  NOR2_X1 U18072 ( .A1(n14756), .A2(n15936), .ZN(n14767) );
  INV_X1 U18073 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14758) );
  NOR4_X1 U18074 ( .A1(n14770), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14758), .A4(n14757), .ZN(n14766) );
  OAI21_X1 U18075 ( .B1(n15952), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14759) );
  NOR2_X1 U18076 ( .A1(n14760), .A2(n14759), .ZN(n14772) );
  INV_X1 U18077 ( .A(n14761), .ZN(n14763) );
  NOR3_X1 U18078 ( .A1(n14772), .A2(n14763), .A3(n14762), .ZN(n14764) );
  OAI21_X1 U18079 ( .B1(n14769), .B2(n15935), .A(n14768), .ZN(P1_U3000) );
  INV_X1 U18080 ( .A(n14770), .ZN(n14771) );
  AOI21_X1 U18081 ( .B1(n14771), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14773) );
  NOR2_X1 U18082 ( .A1(n14773), .A2(n14772), .ZN(n14774) );
  AOI211_X1 U18083 ( .C1(n20126), .C2(n14776), .A(n14775), .B(n14774), .ZN(
        n14777) );
  OAI21_X1 U18084 ( .B1(n14778), .B2(n15935), .A(n14777), .ZN(P1_U3001) );
  XNOR2_X1 U18085 ( .A(n14782), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14784) );
  NAND2_X1 U18086 ( .A1(n14779), .A2(n20126), .ZN(n14781) );
  OAI211_X1 U18087 ( .C1(n14788), .C2(n14782), .A(n14781), .B(n14780), .ZN(
        n14783) );
  AOI21_X1 U18088 ( .B1(n14793), .B2(n14784), .A(n14783), .ZN(n14785) );
  OAI21_X1 U18089 ( .B1(n14786), .B2(n15935), .A(n14785), .ZN(P1_U3003) );
  INV_X1 U18090 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14792) );
  OAI21_X1 U18091 ( .B1(n14788), .B2(n14792), .A(n14787), .ZN(n14791) );
  NOR2_X1 U18092 ( .A1(n14789), .A2(n15936), .ZN(n14790) );
  AOI211_X1 U18093 ( .C1(n14793), .C2(n14792), .A(n14791), .B(n14790), .ZN(
        n14794) );
  OAI21_X1 U18094 ( .B1(n14795), .B2(n15935), .A(n14794), .ZN(P1_U3004) );
  NAND3_X1 U18095 ( .A1(n14829), .A2(n14797), .A3(n14808), .ZN(n14812) );
  AOI21_X1 U18096 ( .B1(n14812), .B2(n14809), .A(n14798), .ZN(n14804) );
  NAND3_X1 U18097 ( .A1(n14829), .A2(n14799), .A3(n14798), .ZN(n14801) );
  OAI211_X1 U18098 ( .C1(n15936), .C2(n14802), .A(n14801), .B(n14800), .ZN(
        n14803) );
  NOR2_X1 U18099 ( .A1(n14804), .A2(n14803), .ZN(n14805) );
  OAI21_X1 U18100 ( .B1(n14806), .B2(n15935), .A(n14805), .ZN(P1_U3005) );
  OAI21_X1 U18101 ( .B1(n14809), .B2(n14808), .A(n14807), .ZN(n14810) );
  AOI21_X1 U18102 ( .B1(n14811), .B2(n20126), .A(n14810), .ZN(n14813) );
  OAI211_X1 U18103 ( .C1(n14814), .C2(n15935), .A(n14813), .B(n14812), .ZN(
        P1_U3006) );
  INV_X1 U18104 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14828) );
  OAI21_X1 U18105 ( .B1(n14892), .B2(n14899), .A(n14828), .ZN(n14815) );
  AOI21_X1 U18106 ( .B1(n14825), .B2(n14815), .A(n14819), .ZN(n14816) );
  AOI211_X1 U18107 ( .C1(n14818), .C2(n20126), .A(n14817), .B(n14816), .ZN(
        n14821) );
  NAND3_X1 U18108 ( .A1(n14829), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14819), .ZN(n14820) );
  OAI211_X1 U18109 ( .C1(n14822), .C2(n15935), .A(n14821), .B(n14820), .ZN(
        P1_U3007) );
  NOR2_X1 U18110 ( .A1(n14823), .A2(n15936), .ZN(n14827) );
  OAI21_X1 U18111 ( .B1(n14825), .B2(n14828), .A(n14824), .ZN(n14826) );
  AOI211_X1 U18112 ( .C1(n14829), .C2(n14828), .A(n14827), .B(n14826), .ZN(
        n14830) );
  OAI21_X1 U18113 ( .B1(n14831), .B2(n15935), .A(n14830), .ZN(P1_U3008) );
  OAI21_X1 U18114 ( .B1(n14840), .B2(n14833), .A(n14832), .ZN(n14836) );
  XNOR2_X1 U18115 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14834) );
  NOR2_X1 U18116 ( .A1(n14841), .A2(n14834), .ZN(n14835) );
  AOI211_X1 U18117 ( .C1(n20126), .C2(n15745), .A(n14836), .B(n14835), .ZN(
        n14837) );
  OAI21_X1 U18118 ( .B1(n14838), .B2(n15935), .A(n14837), .ZN(P1_U3009) );
  OAI21_X1 U18119 ( .B1(n14840), .B2(n12416), .A(n14839), .ZN(n14843) );
  NOR2_X1 U18120 ( .A1(n14841), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14842) );
  AOI211_X1 U18121 ( .C1(n20126), .C2(n15758), .A(n14843), .B(n14842), .ZN(
        n14844) );
  OAI21_X1 U18122 ( .B1(n14845), .B2(n15935), .A(n14844), .ZN(P1_U3010) );
  OAI21_X1 U18123 ( .B1(n14847), .B2(n14846), .A(n21133), .ZN(n14849) );
  INV_X1 U18124 ( .A(n15880), .ZN(n14848) );
  AOI21_X1 U18125 ( .B1(n14849), .B2(n14848), .A(n12415), .ZN(n14850) );
  AOI211_X1 U18126 ( .C1(n20126), .C2(n14852), .A(n14851), .B(n14850), .ZN(
        n14854) );
  NAND3_X1 U18127 ( .A1(n15881), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n12415), .ZN(n14853) );
  OAI211_X1 U18128 ( .C1(n14855), .C2(n15935), .A(n14854), .B(n14853), .ZN(
        P1_U3011) );
  INV_X1 U18129 ( .A(n14856), .ZN(n14858) );
  OAI21_X1 U18130 ( .B1(n14859), .B2(n14858), .A(n14857), .ZN(n14862) );
  NAND2_X1 U18131 ( .A1(n14862), .A2(n14860), .ZN(n14861) );
  MUX2_X1 U18132 ( .A(n14862), .B(n14861), .S(n10332), .Z(n14864) );
  XNOR2_X1 U18133 ( .A(n14864), .B(n14863), .ZN(n15839) );
  NOR2_X1 U18134 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14865), .ZN(
        n15912) );
  NOR2_X1 U18135 ( .A1(n20132), .A2(n15931), .ZN(n14866) );
  NOR2_X1 U18136 ( .A1(n14868), .A2(n14867), .ZN(n15913) );
  INV_X1 U18137 ( .A(n14869), .ZN(n15914) );
  OAI22_X1 U18138 ( .A1(n14871), .A2(n20132), .B1(n14870), .B2(n15914), .ZN(
        n14872) );
  NOR2_X1 U18139 ( .A1(n15912), .A2(n15915), .ZN(n15904) );
  OAI21_X1 U18140 ( .B1(n15952), .B2(n14873), .A(n15904), .ZN(n15888) );
  OAI21_X1 U18141 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n14874), .A(
        n15888), .ZN(n14876) );
  AOI22_X1 U18142 ( .A1(n15792), .A2(n20126), .B1(n12122), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n14875) );
  OAI211_X1 U18143 ( .C1(n15839), .C2(n15935), .A(n14876), .B(n14875), .ZN(
        P1_U3014) );
  INV_X1 U18144 ( .A(n14877), .ZN(n14882) );
  OAI21_X1 U18145 ( .B1(n15892), .B2(n15852), .A(n14878), .ZN(n14881) );
  INV_X1 U18146 ( .A(n14879), .ZN(n14880) );
  AOI21_X1 U18147 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n15844) );
  OAI21_X1 U18148 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15952), .A(
        n15904), .ZN(n15895) );
  NOR2_X1 U18149 ( .A1(n9917), .A2(n14883), .ZN(n14884) );
  OR2_X1 U18150 ( .A1(n14885), .A2(n14884), .ZN(n15825) );
  NOR2_X1 U18151 ( .A1(n15825), .A2(n15936), .ZN(n14887) );
  OAI22_X1 U18152 ( .A1(n20135), .A2(n20767), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15891), .ZN(n14886) );
  AOI211_X1 U18153 ( .C1(n15895), .C2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n14887), .B(n14886), .ZN(n14888) );
  OAI21_X1 U18154 ( .B1(n15844), .B2(n15935), .A(n14888), .ZN(P1_U3016) );
  AOI21_X1 U18155 ( .B1(n14891), .B2(n14890), .A(n14889), .ZN(n15850) );
  NOR2_X1 U18156 ( .A1(n20135), .A2(n20760), .ZN(n14906) );
  NAND2_X1 U18157 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14892), .ZN(
        n20141) );
  NOR2_X1 U18158 ( .A1(n21116), .A2(n20141), .ZN(n14901) );
  INV_X1 U18159 ( .A(n14901), .ZN(n15955) );
  NAND2_X1 U18160 ( .A1(n20132), .A2(n15955), .ZN(n15901) );
  NAND2_X1 U18161 ( .A1(n15931), .A2(n15901), .ZN(n15979) );
  NOR2_X1 U18162 ( .A1(n14898), .A2(n15979), .ZN(n14904) );
  INV_X1 U18163 ( .A(n14895), .ZN(n14893) );
  NOR3_X1 U18164 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14894), .A3(
        n14893), .ZN(n15924) );
  AOI21_X1 U18165 ( .B1(n14896), .B2(n14895), .A(n15930), .ZN(n14897) );
  AOI211_X1 U18166 ( .C1(n14899), .C2(n14898), .A(n14897), .B(n15953), .ZN(
        n15929) );
  INV_X1 U18167 ( .A(n15929), .ZN(n14900) );
  AOI21_X1 U18168 ( .B1(n14901), .B2(n15924), .A(n14900), .ZN(n14902) );
  INV_X1 U18169 ( .A(n14902), .ZN(n14903) );
  MUX2_X1 U18170 ( .A(n14904), .B(n14903), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n14905) );
  AOI211_X1 U18171 ( .C1(n20126), .C2(n15808), .A(n14906), .B(n14905), .ZN(
        n14907) );
  OAI21_X1 U18172 ( .B1(n15850), .B2(n15935), .A(n14907), .ZN(P1_U3019) );
  NAND3_X1 U18173 ( .A1(n14908), .A2(n9815), .A3(n20123), .ZN(n14918) );
  NOR2_X1 U18174 ( .A1(n14910), .A2(n14909), .ZN(n14911) );
  NOR2_X1 U18175 ( .A1(n20122), .A2(n14911), .ZN(n14912) );
  AOI211_X1 U18176 ( .C1(n20126), .C2(n14914), .A(n14913), .B(n14912), .ZN(
        n14917) );
  OR3_X1 U18177 ( .A1(n15952), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n14915), .ZN(n14916) );
  NAND3_X1 U18178 ( .A1(n14918), .A2(n14917), .A3(n14916), .ZN(P1_U3030) );
  XNOR2_X1 U18179 ( .A(n9821), .B(P1_STATEBS16_REG_SCAN_IN), .ZN(n14920) );
  OAI22_X1 U18180 ( .A1(n14920), .A2(n20669), .B1(n13725), .B2(n14922), .ZN(
        n14921) );
  MUX2_X1 U18181 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14921), .S(
        n20142), .Z(P1_U3477) );
  NAND2_X1 U18182 ( .A1(n9821), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20665) );
  XNOR2_X1 U18183 ( .A(n14925), .B(n20665), .ZN(n14923) );
  OAI22_X1 U18184 ( .A1(n14923), .A2(n20669), .B1(n13091), .B2(n14922), .ZN(
        n14924) );
  MUX2_X1 U18185 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14924), .S(
        n20142), .Z(P1_U3476) );
  NOR2_X1 U18186 ( .A1(n20390), .A2(n20665), .ZN(n20394) );
  AOI211_X1 U18187 ( .C1(n20146), .C2(n20622), .A(n20515), .B(n20394), .ZN(
        n14930) );
  AOI21_X1 U18188 ( .B1(n14928), .B2(n20421), .A(n10331), .ZN(n14929) );
  OAI21_X1 U18189 ( .B1(n14930), .B2(n20669), .A(n14929), .ZN(n14931) );
  MUX2_X1 U18190 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n14931), .S(
        n20142), .Z(P1_U3475) );
  NOR2_X1 U18191 ( .A1(n14932), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14935) );
  NOR3_X1 U18192 ( .A1(n14933), .A2(n14937), .A3(n11832), .ZN(n14934) );
  AOI211_X1 U18193 ( .C1(n20625), .C2(n14936), .A(n14935), .B(n14934), .ZN(
        n15693) );
  NOR3_X1 U18194 ( .A1(n11832), .A2(n14937), .A3(n20805), .ZN(n14938) );
  AOI21_X1 U18195 ( .B1(n14940), .B2(n14939), .A(n14938), .ZN(n14941) );
  OAI21_X1 U18196 ( .B1(n15693), .B2(n20807), .A(n14941), .ZN(n14942) );
  MUX2_X1 U18197 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14942), .S(
        n20809), .Z(P1_U3473) );
  NAND2_X1 U18198 ( .A1(n14984), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14943) );
  OAI21_X1 U18199 ( .B1(n11783), .B2(n14984), .A(n14943), .ZN(P2_U2856) );
  NAND2_X1 U18200 ( .A1(n14945), .A2(n14944), .ZN(n14946) );
  XOR2_X1 U18201 ( .A(n14947), .B(n14946), .Z(n15047) );
  NOR2_X1 U18202 ( .A1(n15296), .A2(n14984), .ZN(n14948) );
  AOI21_X1 U18203 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n14984), .A(n14948), .ZN(
        n14949) );
  OAI21_X1 U18204 ( .B1(n15047), .B2(n15038), .A(n14949), .ZN(P2_U2859) );
  OAI21_X1 U18205 ( .B1(n14952), .B2(n14951), .A(n14950), .ZN(n15058) );
  NOR2_X1 U18206 ( .A1(n15119), .A2(n14984), .ZN(n14953) );
  AOI21_X1 U18207 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n14984), .A(n14953), .ZN(
        n14954) );
  OAI21_X1 U18208 ( .B1(n15058), .B2(n15038), .A(n14954), .ZN(P2_U2860) );
  OR2_X1 U18209 ( .A1(n14966), .A2(n14955), .ZN(n14956) );
  NAND2_X1 U18210 ( .A1(n12948), .A2(n14956), .ZN(n16031) );
  AOI21_X1 U18211 ( .B1(n14959), .B2(n14958), .A(n14957), .ZN(n15059) );
  NAND2_X1 U18212 ( .A1(n15059), .A2(n15021), .ZN(n14961) );
  NAND2_X1 U18213 ( .A1(n14984), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14960) );
  OAI211_X1 U18214 ( .C1(n16031), .C2(n14984), .A(n14961), .B(n14960), .ZN(
        P2_U2861) );
  OAI21_X1 U18215 ( .B1(n14962), .B2(n14964), .A(n14963), .ZN(n15078) );
  AND2_X1 U18216 ( .A1(n14975), .A2(n14965), .ZN(n14967) );
  OR2_X1 U18217 ( .A1(n14967), .A2(n14966), .ZN(n15143) );
  NOR2_X1 U18218 ( .A1(n15143), .A2(n14984), .ZN(n14968) );
  AOI21_X1 U18219 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n14984), .A(n14968), .ZN(
        n14969) );
  OAI21_X1 U18220 ( .B1(n15078), .B2(n15038), .A(n14969), .ZN(P2_U2862) );
  OAI21_X1 U18221 ( .B1(n14972), .B2(n14971), .A(n14970), .ZN(n14973) );
  XOR2_X1 U18222 ( .A(n14974), .B(n14973), .Z(n15086) );
  INV_X1 U18223 ( .A(n14975), .ZN(n14976) );
  AOI21_X1 U18224 ( .B1(n14978), .B2(n14977), .A(n14976), .ZN(n16050) );
  INV_X1 U18225 ( .A(n16050), .ZN(n15346) );
  NOR2_X1 U18226 ( .A1(n15346), .A2(n14984), .ZN(n14979) );
  AOI21_X1 U18227 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n14984), .A(n14979), .ZN(
        n14980) );
  OAI21_X1 U18228 ( .B1(n15086), .B2(n15038), .A(n14980), .ZN(P2_U2863) );
  OAI21_X1 U18229 ( .B1(n14983), .B2(n14982), .A(n14981), .ZN(n15091) );
  MUX2_X1 U18230 ( .A(n15352), .B(n14985), .S(n14984), .Z(n14986) );
  OAI21_X1 U18231 ( .B1(n15091), .B2(n15038), .A(n14986), .ZN(P2_U2864) );
  OAI21_X1 U18232 ( .B1(n14987), .B2(n14988), .A(n12677), .ZN(n16060) );
  INV_X1 U18233 ( .A(n14990), .ZN(n14991) );
  AOI21_X1 U18234 ( .B1(n10295), .B2(n14991), .A(n9899), .ZN(n15687) );
  NAND2_X1 U18235 ( .A1(n15687), .A2(n15036), .ZN(n14993) );
  NAND2_X1 U18236 ( .A1(n14984), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14992) );
  OAI211_X1 U18237 ( .C1(n16060), .C2(n15038), .A(n14993), .B(n14992), .ZN(
        P2_U2865) );
  AOI21_X1 U18238 ( .B1(n14995), .B2(n14994), .A(n14987), .ZN(n15092) );
  NAND2_X1 U18239 ( .A1(n15092), .A2(n15021), .ZN(n14997) );
  NAND2_X1 U18240 ( .A1(n14984), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14996) );
  OAI211_X1 U18241 ( .C1(n15387), .C2(n14984), .A(n14997), .B(n14996), .ZN(
        P2_U2866) );
  INV_X1 U18242 ( .A(n14999), .ZN(n15000) );
  AOI21_X1 U18243 ( .B1(n15001), .B2(n14998), .A(n15000), .ZN(n18856) );
  NAND2_X1 U18244 ( .A1(n18856), .A2(n15036), .ZN(n15006) );
  OR2_X1 U18245 ( .A1(n15002), .A2(n15003), .ZN(n15004) );
  AND2_X1 U18246 ( .A1(n14994), .A2(n15004), .ZN(n16067) );
  NAND2_X1 U18247 ( .A1(n16067), .A2(n15021), .ZN(n15005) );
  OAI211_X1 U18248 ( .C1(n15036), .C2(n15007), .A(n15006), .B(n15005), .ZN(
        P2_U2867) );
  OR2_X1 U18249 ( .A1(n15017), .A2(n15008), .ZN(n15009) );
  AND2_X1 U18250 ( .A1(n14998), .A2(n15009), .ZN(n18876) );
  INV_X1 U18251 ( .A(n18876), .ZN(n15014) );
  AOI21_X1 U18252 ( .B1(n15011), .B2(n15018), .A(n15002), .ZN(n15103) );
  NAND2_X1 U18253 ( .A1(n15103), .A2(n15021), .ZN(n15013) );
  NAND2_X1 U18254 ( .A1(n14984), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15012) );
  OAI211_X1 U18255 ( .C1(n15014), .C2(n14984), .A(n15013), .B(n15012), .ZN(
        P2_U2868) );
  NOR2_X1 U18256 ( .A1(n9896), .A2(n15015), .ZN(n15016) );
  OR2_X1 U18257 ( .A1(n15017), .A2(n15016), .ZN(n18889) );
  INV_X1 U18258 ( .A(n15018), .ZN(n15019) );
  AOI21_X1 U18259 ( .B1(n15020), .B2(n13757), .A(n15019), .ZN(n16072) );
  NAND2_X1 U18260 ( .A1(n16072), .A2(n15021), .ZN(n15023) );
  NAND2_X1 U18261 ( .A1(n14984), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15022) );
  OAI211_X1 U18262 ( .C1(n18889), .C2(n14984), .A(n15023), .B(n15022), .ZN(
        P2_U2869) );
  AOI21_X1 U18263 ( .B1(n15024), .B2(n15031), .A(n9896), .ZN(n18899) );
  NAND2_X1 U18264 ( .A1(n18899), .A2(n15036), .ZN(n15026) );
  NAND2_X1 U18265 ( .A1(n14984), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15025) );
  OAI211_X1 U18266 ( .C1(n15027), .C2(n15038), .A(n15026), .B(n15025), .ZN(
        P2_U2870) );
  AND2_X1 U18267 ( .A1(n15029), .A2(n15028), .ZN(n15030) );
  OR2_X1 U18268 ( .A1(n15030), .A2(n13756), .ZN(n19094) );
  INV_X1 U18269 ( .A(n15031), .ZN(n15032) );
  AOI21_X1 U18270 ( .B1(n15033), .B2(n13604), .A(n15032), .ZN(n18909) );
  INV_X1 U18271 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n15034) );
  NOR2_X1 U18272 ( .A1(n15036), .A2(n15034), .ZN(n15035) );
  AOI21_X1 U18273 ( .B1(n18909), .B2(n15036), .A(n15035), .ZN(n15037) );
  OAI21_X1 U18274 ( .B1(n15038), .B2(n19094), .A(n15037), .ZN(P2_U2871) );
  OR2_X1 U18275 ( .A1(n19100), .A2(n15039), .ZN(n15041) );
  NAND2_X1 U18276 ( .A1(n19100), .A2(BUF2_REG_12__SCAN_IN), .ZN(n15040) );
  AND2_X1 U18277 ( .A1(n15041), .A2(n15040), .ZN(n19228) );
  INV_X1 U18278 ( .A(n19228), .ZN(n15042) );
  AOI22_X1 U18279 ( .A1(n19088), .A2(n15042), .B1(n19125), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15043) );
  OAI21_X1 U18280 ( .B1(n15054), .B2(n17222), .A(n15043), .ZN(n15045) );
  NOR2_X1 U18281 ( .A1(n15301), .A2(n19092), .ZN(n15044) );
  AOI211_X1 U18282 ( .C1(n19089), .C2(BUF1_REG_28__SCAN_IN), .A(n15045), .B(
        n15044), .ZN(n15046) );
  OAI21_X1 U18283 ( .B1(n15047), .B2(n19093), .A(n15046), .ZN(P2_U2891) );
  INV_X1 U18284 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n15053) );
  OR2_X1 U18285 ( .A1(n19100), .A2(n15048), .ZN(n15050) );
  NAND2_X1 U18286 ( .A1(n19100), .A2(BUF2_REG_11__SCAN_IN), .ZN(n15049) );
  AND2_X1 U18287 ( .A1(n15050), .A2(n15049), .ZN(n19226) );
  INV_X1 U18288 ( .A(n19226), .ZN(n15051) );
  AOI22_X1 U18289 ( .A1(n19088), .A2(n15051), .B1(n19125), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15052) );
  OAI21_X1 U18290 ( .B1(n15054), .B2(n15053), .A(n15052), .ZN(n15056) );
  NOR2_X1 U18291 ( .A1(n15314), .A2(n19092), .ZN(n15055) );
  AOI211_X1 U18292 ( .C1(n19089), .C2(BUF1_REG_27__SCAN_IN), .A(n15056), .B(
        n15055), .ZN(n15057) );
  OAI21_X1 U18293 ( .B1(n15058), .B2(n19093), .A(n15057), .ZN(P2_U2892) );
  NAND2_X1 U18294 ( .A1(n15059), .A2(n19127), .ZN(n15066) );
  AOI22_X1 U18295 ( .A1(n19088), .A2(n19111), .B1(n19125), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15065) );
  AOI22_X1 U18296 ( .A1(n19089), .A2(BUF1_REG_26__SCAN_IN), .B1(n19090), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15064) );
  AND2_X1 U18297 ( .A1(n15069), .A2(n15060), .ZN(n15061) );
  NOR2_X1 U18298 ( .A1(n15062), .A2(n15061), .ZN(n16034) );
  NAND2_X1 U18299 ( .A1(n16034), .A2(n19099), .ZN(n15063) );
  NAND4_X1 U18300 ( .A1(n15066), .A2(n15065), .A3(n15064), .A4(n15063), .ZN(
        P2_U2893) );
  NAND2_X1 U18301 ( .A1(n15079), .A2(n15067), .ZN(n15068) );
  NAND2_X1 U18302 ( .A1(n15069), .A2(n15068), .ZN(n16042) );
  INV_X1 U18303 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n15070) );
  OR2_X1 U18304 ( .A1(n19100), .A2(n15070), .ZN(n15072) );
  NAND2_X1 U18305 ( .A1(n19100), .A2(BUF2_REG_9__SCAN_IN), .ZN(n15071) );
  AND2_X1 U18306 ( .A1(n15072), .A2(n15071), .ZN(n19224) );
  INV_X1 U18307 ( .A(n19224), .ZN(n15073) );
  AOI22_X1 U18308 ( .A1(n19088), .A2(n15073), .B1(n19125), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15075) );
  AOI22_X1 U18309 ( .A1(n19089), .A2(BUF1_REG_25__SCAN_IN), .B1(n19090), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15074) );
  OAI211_X1 U18310 ( .C1(n16042), .C2(n19092), .A(n15075), .B(n15074), .ZN(
        n15076) );
  INV_X1 U18311 ( .A(n15076), .ZN(n15077) );
  OAI21_X1 U18312 ( .B1(n15078), .B2(n19093), .A(n15077), .ZN(P2_U2894) );
  AOI21_X1 U18313 ( .B1(n15080), .B2(n12937), .A(n10138), .ZN(n16049) );
  INV_X1 U18314 ( .A(n19116), .ZN(n15081) );
  OAI22_X1 U18315 ( .A1(n15082), .A2(n15081), .B1(n19121), .B2(n19155), .ZN(
        n15083) );
  AOI21_X1 U18316 ( .B1(n16049), .B2(n19099), .A(n15083), .ZN(n15085) );
  AOI22_X1 U18317 ( .A1(n19089), .A2(BUF1_REG_24__SCAN_IN), .B1(n19090), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15084) );
  OAI211_X1 U18318 ( .C1(n15086), .C2(n19093), .A(n15085), .B(n15084), .ZN(
        P2_U2895) );
  AOI22_X1 U18319 ( .A1(n19089), .A2(BUF1_REG_23__SCAN_IN), .B1(n19090), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15088) );
  AOI22_X1 U18320 ( .A1(n19088), .A2(n15645), .B1(n19125), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15087) );
  OAI211_X1 U18321 ( .C1(n19092), .C2(n15355), .A(n15088), .B(n15087), .ZN(
        n15089) );
  INV_X1 U18322 ( .A(n15089), .ZN(n15090) );
  OAI21_X1 U18323 ( .B1(n15091), .B2(n19093), .A(n15090), .ZN(P2_U2896) );
  NAND2_X1 U18324 ( .A1(n15092), .A2(n19127), .ZN(n15096) );
  AOI22_X1 U18325 ( .A1(n19088), .A2(n19124), .B1(n19125), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U18326 ( .A1(n19089), .A2(BUF1_REG_21__SCAN_IN), .B1(n19090), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15094) );
  NAND2_X1 U18327 ( .A1(n19099), .A2(n15380), .ZN(n15093) );
  NAND4_X1 U18328 ( .A1(n15096), .A2(n15095), .A3(n15094), .A4(n15093), .ZN(
        P2_U2898) );
  AND2_X1 U18329 ( .A1(n15419), .A2(n15097), .ZN(n15098) );
  OR2_X1 U18330 ( .A1(n15098), .A2(n15393), .ZN(n18878) );
  AOI22_X1 U18331 ( .A1(n19089), .A2(BUF1_REG_19__SCAN_IN), .B1(n19090), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n15101) );
  AOI22_X1 U18332 ( .A1(n19088), .A2(n15099), .B1(n19125), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15100) );
  OAI211_X1 U18333 ( .C1(n19092), .C2(n18878), .A(n15101), .B(n15100), .ZN(
        n15102) );
  AOI21_X1 U18334 ( .B1(n15103), .B2(n19127), .A(n15102), .ZN(n15104) );
  INV_X1 U18335 ( .A(n15104), .ZN(P2_U2900) );
  NAND2_X1 U18336 ( .A1(n15106), .A2(n15105), .ZN(n15108) );
  XOR2_X1 U18337 ( .A(n15108), .B(n15107), .Z(n15294) );
  INV_X1 U18338 ( .A(n16024), .ZN(n15290) );
  NAND2_X1 U18339 ( .A1(n19236), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15287) );
  NAND2_X1 U18340 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15109) );
  OAI211_X1 U18341 ( .C1(n19247), .C2(n15110), .A(n15287), .B(n15109), .ZN(
        n15111) );
  AOI21_X1 U18342 ( .B1(n15290), .B2(n9787), .A(n15111), .ZN(n15115) );
  AOI21_X1 U18343 ( .B1(n15284), .B2(n15113), .A(n15112), .ZN(n15291) );
  NAND2_X1 U18344 ( .A1(n15291), .A2(n19241), .ZN(n15114) );
  OAI211_X1 U18345 ( .C1(n15294), .C2(n12452), .A(n15115), .B(n15114), .ZN(
        P2_U2985) );
  XNOR2_X1 U18346 ( .A(n15116), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15318) );
  INV_X1 U18347 ( .A(n15117), .ZN(n15118) );
  INV_X1 U18348 ( .A(n15119), .ZN(n15317) );
  NAND2_X1 U18349 ( .A1(n16143), .A2(n15120), .ZN(n15121) );
  NAND2_X1 U18350 ( .A1(n19236), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15310) );
  OAI211_X1 U18351 ( .C1(n16150), .C2(n15122), .A(n15121), .B(n15310), .ZN(
        n15123) );
  INV_X1 U18352 ( .A(n15123), .ZN(n15124) );
  OAI21_X1 U18353 ( .B1(n15318), .B2(n12452), .A(n15128), .ZN(P2_U2987) );
  OAI21_X1 U18354 ( .B1(n15129), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15117), .ZN(n15330) );
  AOI21_X1 U18355 ( .B1(n15130), .B2(n15139), .A(n15138), .ZN(n15132) );
  XNOR2_X1 U18356 ( .A(n15132), .B(n15131), .ZN(n15328) );
  NOR2_X1 U18357 ( .A1(n16031), .A2(n16130), .ZN(n15136) );
  NAND2_X1 U18358 ( .A1(n19236), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15319) );
  NAND2_X1 U18359 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15133) );
  OAI211_X1 U18360 ( .C1(n19247), .C2(n15134), .A(n15319), .B(n15133), .ZN(
        n15135) );
  AOI211_X1 U18361 ( .C1(n15328), .C2(n19242), .A(n15136), .B(n15135), .ZN(
        n15137) );
  OAI21_X1 U18362 ( .B1(n16145), .B2(n15330), .A(n15137), .ZN(P2_U2988) );
  NAND2_X1 U18363 ( .A1(n10304), .A2(n15139), .ZN(n15140) );
  XNOR2_X1 U18364 ( .A(n15130), .B(n15140), .ZN(n15339) );
  AOI21_X1 U18365 ( .B1(n15332), .B2(n15142), .A(n15129), .ZN(n15331) );
  NAND2_X1 U18366 ( .A1(n15331), .A2(n19241), .ZN(n15148) );
  INV_X1 U18367 ( .A(n15143), .ZN(n16045) );
  NAND2_X1 U18368 ( .A1(n16143), .A2(n16037), .ZN(n15144) );
  NAND2_X1 U18369 ( .A1(n19236), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15334) );
  OAI211_X1 U18370 ( .C1(n16150), .C2(n15145), .A(n15144), .B(n15334), .ZN(
        n15146) );
  AOI21_X1 U18371 ( .B1(n16045), .B2(n9787), .A(n15146), .ZN(n15147) );
  OAI211_X1 U18372 ( .C1(n12452), .C2(n15339), .A(n15148), .B(n15147), .ZN(
        P2_U2989) );
  OAI21_X1 U18373 ( .B1(n9861), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15142), .ZN(n15350) );
  XOR2_X1 U18374 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15149), .Z(
        n15150) );
  XNOR2_X1 U18375 ( .A(n15151), .B(n15150), .ZN(n15348) );
  NAND2_X1 U18376 ( .A1(n16050), .A2(n9787), .ZN(n15153) );
  NOR2_X1 U18377 ( .A1(n19034), .A2(n19820), .ZN(n15344) );
  AOI21_X1 U18378 ( .B1(n19237), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15344), .ZN(n15152) );
  OAI211_X1 U18379 ( .C1(n19247), .C2(n15154), .A(n15153), .B(n15152), .ZN(
        n15155) );
  AOI21_X1 U18380 ( .B1(n15348), .B2(n19242), .A(n15155), .ZN(n15156) );
  OAI21_X1 U18381 ( .B1(n15350), .B2(n16145), .A(n15156), .ZN(P2_U2990) );
  XNOR2_X1 U18382 ( .A(n15157), .B(n15158), .ZN(n15365) );
  AOI21_X1 U18383 ( .B1(n15359), .B2(n15159), .A(n9861), .ZN(n15351) );
  NAND2_X1 U18384 ( .A1(n15351), .A2(n19241), .ZN(n15165) );
  NAND2_X1 U18385 ( .A1(n19236), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15358) );
  OAI21_X1 U18386 ( .B1(n16150), .B2(n15160), .A(n15358), .ZN(n15162) );
  NOR2_X1 U18387 ( .A1(n15352), .A2(n16130), .ZN(n15161) );
  AOI211_X1 U18388 ( .C1(n16143), .C2(n15163), .A(n15162), .B(n15161), .ZN(
        n15164) );
  OAI211_X1 U18389 ( .C1(n15365), .C2(n12452), .A(n15165), .B(n15164), .ZN(
        P2_U2991) );
  OAI21_X1 U18390 ( .B1(n15166), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15159), .ZN(n15379) );
  NAND2_X1 U18391 ( .A1(n19236), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n15371) );
  NAND2_X1 U18392 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15167) );
  OAI211_X1 U18393 ( .C1(n19247), .C2(n15168), .A(n15371), .B(n15167), .ZN(
        n15174) );
  NAND2_X1 U18394 ( .A1(n10072), .A2(n15170), .ZN(n15171) );
  XNOR2_X1 U18395 ( .A(n15172), .B(n15171), .ZN(n15376) );
  NOR2_X1 U18396 ( .A1(n15376), .A2(n12452), .ZN(n15173) );
  AOI211_X1 U18397 ( .C1(n9787), .C2(n15687), .A(n15174), .B(n15173), .ZN(
        n15175) );
  OAI21_X1 U18398 ( .B1(n16145), .B2(n15379), .A(n15175), .ZN(P2_U2992) );
  AOI21_X1 U18399 ( .B1(n15176), .B2(n16084), .A(n16086), .ZN(n16079) );
  INV_X1 U18400 ( .A(n15177), .ZN(n16077) );
  INV_X1 U18401 ( .A(n16076), .ZN(n15178) );
  AOI21_X1 U18402 ( .B1(n16079), .B2(n16077), .A(n15178), .ZN(n15253) );
  AOI21_X1 U18403 ( .B1(n15253), .B2(n15250), .A(n15249), .ZN(n15241) );
  NAND2_X1 U18404 ( .A1(n15241), .A2(n15240), .ZN(n15239) );
  NAND2_X1 U18405 ( .A1(n15239), .A2(n15179), .ZN(n15232) );
  NOR2_X1 U18406 ( .A1(n15180), .A2(n15181), .ZN(n15231) );
  NAND3_X1 U18407 ( .A1(n15223), .A2(n15209), .A3(n15220), .ZN(n15198) );
  INV_X1 U18408 ( .A(n15197), .ZN(n15182) );
  NOR2_X1 U18409 ( .A1(n15182), .A2(n15196), .ZN(n15183) );
  AOI21_X1 U18410 ( .B1(n15198), .B2(n15183), .A(n15195), .ZN(n15187) );
  NAND2_X1 U18411 ( .A1(n15185), .A2(n15184), .ZN(n15186) );
  XNOR2_X1 U18412 ( .A(n15187), .B(n15186), .ZN(n15391) );
  AOI21_X1 U18413 ( .B1(n20968), .B2(n15188), .A(n15166), .ZN(n15389) );
  NAND2_X1 U18414 ( .A1(n19236), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15382) );
  OAI21_X1 U18415 ( .B1(n16150), .B2(n15189), .A(n15382), .ZN(n15190) );
  AOI21_X1 U18416 ( .B1(n16143), .B2(n15191), .A(n15190), .ZN(n15192) );
  OAI21_X1 U18417 ( .B1(n15387), .B2(n16130), .A(n15192), .ZN(n15193) );
  AOI21_X1 U18418 ( .B1(n15389), .B2(n19241), .A(n15193), .ZN(n15194) );
  OAI21_X1 U18419 ( .B1(n15391), .B2(n12452), .A(n15194), .ZN(P2_U2993) );
  NOR2_X1 U18420 ( .A1(n15196), .A2(n15195), .ZN(n15200) );
  NAND2_X1 U18421 ( .A1(n15198), .A2(n15197), .ZN(n15199) );
  XOR2_X1 U18422 ( .A(n15200), .B(n15199), .Z(n15403) );
  NOR2_X1 U18423 ( .A1(n19034), .A2(n15201), .ZN(n15395) );
  AOI21_X1 U18424 ( .B1(n19237), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15395), .ZN(n15202) );
  OAI21_X1 U18425 ( .B1(n19247), .B2(n15203), .A(n15202), .ZN(n15206) );
  OAI21_X1 U18426 ( .B1(n15204), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15188), .ZN(n15399) );
  NOR2_X1 U18427 ( .A1(n15399), .A2(n16145), .ZN(n15205) );
  AOI211_X1 U18428 ( .C1(n9787), .C2(n18856), .A(n15206), .B(n15205), .ZN(
        n15207) );
  OAI21_X1 U18429 ( .B1(n15403), .B2(n12452), .A(n15207), .ZN(P2_U2994) );
  NAND2_X1 U18430 ( .A1(n15209), .A2(n15208), .ZN(n15212) );
  INV_X1 U18431 ( .A(n15221), .ZN(n15210) );
  OAI21_X1 U18432 ( .B1(n15223), .B2(n15210), .A(n15220), .ZN(n15211) );
  XOR2_X1 U18433 ( .A(n15212), .B(n15211), .Z(n15415) );
  NAND2_X1 U18434 ( .A1(n18869), .A2(n16143), .ZN(n15213) );
  NAND2_X1 U18435 ( .A1(n19236), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15405) );
  OAI211_X1 U18436 ( .C1(n16150), .C2(n15214), .A(n15213), .B(n15405), .ZN(
        n15215) );
  AOI21_X1 U18437 ( .B1(n18876), .B2(n9787), .A(n15215), .ZN(n15219) );
  AND2_X1 U18438 ( .A1(n15216), .A2(n15404), .ZN(n15217) );
  NOR2_X1 U18439 ( .A1(n15204), .A2(n15217), .ZN(n15412) );
  NAND2_X1 U18440 ( .A1(n15412), .A2(n19241), .ZN(n15218) );
  OAI211_X1 U18441 ( .C1(n15415), .C2(n12452), .A(n15219), .B(n15218), .ZN(
        P2_U2995) );
  NAND2_X1 U18442 ( .A1(n15221), .A2(n15220), .ZN(n15222) );
  XNOR2_X1 U18443 ( .A(n15223), .B(n15222), .ZN(n15431) );
  NAND2_X1 U18444 ( .A1(n15224), .A2(n15425), .ZN(n15225) );
  AND2_X1 U18445 ( .A1(n15216), .A2(n15225), .ZN(n15429) );
  NOR2_X1 U18446 ( .A1(n18889), .A2(n16130), .ZN(n15229) );
  NAND2_X1 U18447 ( .A1(n19236), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15420) );
  NAND2_X1 U18448 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15226) );
  OAI211_X1 U18449 ( .C1(n15227), .C2(n19247), .A(n15420), .B(n15226), .ZN(
        n15228) );
  AOI211_X1 U18450 ( .C1(n15429), .C2(n19241), .A(n15229), .B(n15228), .ZN(
        n15230) );
  OAI21_X1 U18451 ( .B1(n15431), .B2(n12452), .A(n15230), .ZN(P2_U2996) );
  XNOR2_X1 U18452 ( .A(n15232), .B(n15231), .ZN(n15447) );
  NAND2_X1 U18453 ( .A1(n18892), .A2(n16143), .ZN(n15233) );
  NAND2_X1 U18454 ( .A1(n19236), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15432) );
  OAI211_X1 U18455 ( .C1(n16150), .C2(n15234), .A(n15233), .B(n15432), .ZN(
        n15235) );
  AOI21_X1 U18456 ( .B1(n18899), .B2(n9787), .A(n15235), .ZN(n15238) );
  OAI211_X1 U18457 ( .C1(n15236), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15224), .B(n19241), .ZN(n15237) );
  OAI211_X1 U18458 ( .C1(n15447), .C2(n12452), .A(n15238), .B(n15237), .ZN(
        P2_U2997) );
  OAI21_X1 U18459 ( .B1(n15241), .B2(n15240), .A(n15239), .ZN(n15458) );
  NOR2_X1 U18460 ( .A1(n15451), .A2(n19034), .ZN(n15244) );
  AOI22_X1 U18461 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16143), .B2(n18904), .ZN(n15242) );
  INV_X1 U18462 ( .A(n15242), .ZN(n15243) );
  AOI211_X1 U18463 ( .C1(n18909), .C2(n9787), .A(n15244), .B(n15243), .ZN(
        n15248) );
  NOR2_X1 U18464 ( .A1(n15245), .A2(n15466), .ZN(n15246) );
  INV_X1 U18465 ( .A(n15236), .ZN(n15438) );
  OAI211_X1 U18466 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15246), .A(
        n15438), .B(n19241), .ZN(n15247) );
  OAI211_X1 U18467 ( .C1(n15458), .C2(n12452), .A(n15248), .B(n15247), .ZN(
        P2_U2998) );
  INV_X1 U18468 ( .A(n15249), .ZN(n15251) );
  NAND2_X1 U18469 ( .A1(n15251), .A2(n15250), .ZN(n15252) );
  XNOR2_X1 U18470 ( .A(n15253), .B(n15252), .ZN(n15472) );
  XNOR2_X1 U18471 ( .A(n15245), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15470) );
  NAND2_X1 U18472 ( .A1(n19236), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n15463) );
  OAI21_X1 U18473 ( .B1(n16150), .B2(n21083), .A(n15463), .ZN(n15254) );
  AOI21_X1 U18474 ( .B1(n16143), .B2(n18920), .A(n15254), .ZN(n15255) );
  OAI21_X1 U18475 ( .B1(n18917), .B2(n16130), .A(n15255), .ZN(n15256) );
  AOI21_X1 U18476 ( .B1(n15470), .B2(n19241), .A(n15256), .ZN(n15257) );
  OAI21_X1 U18477 ( .B1(n15472), .B2(n12452), .A(n15257), .ZN(P2_U2999) );
  INV_X1 U18478 ( .A(n15258), .ZN(n16110) );
  NOR2_X1 U18479 ( .A1(n15259), .A2(n16110), .ZN(n15261) );
  XOR2_X1 U18480 ( .A(n15261), .B(n15260), .Z(n15517) );
  INV_X1 U18481 ( .A(n15262), .ZN(n15263) );
  INV_X1 U18482 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15508) );
  NAND2_X1 U18483 ( .A1(n15263), .A2(n15508), .ZN(n15507) );
  NAND2_X1 U18484 ( .A1(n15262), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16108) );
  NAND3_X1 U18485 ( .A1(n15507), .A2(n19241), .A3(n16108), .ZN(n15269) );
  OAI22_X1 U18486 ( .A1(n16150), .A2(n15264), .B1(n11324), .B2(n19034), .ZN(
        n15267) );
  NOR2_X1 U18487 ( .A1(n15265), .A2(n16130), .ZN(n15266) );
  AOI211_X1 U18488 ( .C1(n16143), .C2(n18981), .A(n15267), .B(n15266), .ZN(
        n15268) );
  OAI211_X1 U18489 ( .C1(n12452), .C2(n15517), .A(n15269), .B(n15268), .ZN(
        P2_U3005) );
  INV_X1 U18490 ( .A(n16124), .ZN(n15271) );
  NOR2_X1 U18491 ( .A1(n15271), .A2(n16123), .ZN(n15272) );
  XNOR2_X1 U18492 ( .A(n15270), .B(n15272), .ZN(n15530) );
  OR2_X1 U18493 ( .A1(n15274), .A2(n15273), .ZN(n15518) );
  NAND3_X1 U18494 ( .A1(n15518), .A2(n19241), .A3(n15275), .ZN(n15280) );
  OAI22_X1 U18495 ( .A1(n16150), .A2(n15276), .B1(n19794), .B2(n19034), .ZN(
        n15278) );
  NOR2_X1 U18496 ( .A1(n19002), .A2(n16130), .ZN(n15277) );
  AOI211_X1 U18497 ( .C1(n16143), .C2(n18997), .A(n15278), .B(n15277), .ZN(
        n15279) );
  OAI211_X1 U18498 ( .C1(n15530), .C2(n12452), .A(n15280), .B(n15279), .ZN(
        P2_U3007) );
  NOR2_X1 U18499 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15281), .ZN(
        n15308) );
  NOR2_X1 U18500 ( .A1(n15311), .A2(n15308), .ZN(n15298) );
  NAND3_X1 U18501 ( .A1(n15297), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15283), .ZN(n15299) );
  AOI21_X1 U18502 ( .B1(n15298), .B2(n15299), .A(n15284), .ZN(n15289) );
  INV_X1 U18503 ( .A(n15282), .ZN(n15285) );
  NAND3_X1 U18504 ( .A1(n15285), .A2(n15284), .A3(n15283), .ZN(n15286) );
  OAI211_X1 U18505 ( .C1(n16020), .C2(n16177), .A(n15287), .B(n15286), .ZN(
        n15288) );
  AOI211_X1 U18506 ( .C1(n15290), .C2(n16182), .A(n15289), .B(n15288), .ZN(
        n15293) );
  NAND2_X1 U18507 ( .A1(n15291), .A2(n16183), .ZN(n15292) );
  OAI211_X1 U18508 ( .C1(n15294), .C2(n16187), .A(n15293), .B(n15292), .ZN(
        P2_U3017) );
  NOR2_X1 U18509 ( .A1(n15295), .A2(n16199), .ZN(n15305) );
  NOR2_X1 U18510 ( .A1(n15296), .A2(n16194), .ZN(n15304) );
  NOR2_X1 U18511 ( .A1(n15298), .A2(n15297), .ZN(n15303) );
  OAI211_X1 U18512 ( .C1(n15301), .C2(n16177), .A(n15300), .B(n15299), .ZN(
        n15302) );
  NOR4_X2 U18513 ( .A1(n15305), .A2(n15304), .A3(n15303), .A4(n15302), .ZN(
        n15306) );
  OAI21_X1 U18514 ( .B1(n15307), .B2(n16187), .A(n15306), .ZN(P2_U3018) );
  INV_X1 U18515 ( .A(n15308), .ZN(n15309) );
  AND2_X1 U18516 ( .A1(n15310), .A2(n15309), .ZN(n15313) );
  NAND2_X1 U18517 ( .A1(n15311), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15312) );
  OAI211_X1 U18518 ( .C1(n15314), .C2(n16177), .A(n15313), .B(n15312), .ZN(
        n15316) );
  INV_X1 U18519 ( .A(n15319), .ZN(n15321) );
  NOR4_X1 U18520 ( .A1(n15342), .A2(n15332), .A3(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(n15341), .ZN(n15320) );
  AOI211_X1 U18521 ( .C1(n16034), .C2(n16192), .A(n15321), .B(n15320), .ZN(
        n15326) );
  NOR2_X1 U18522 ( .A1(n15342), .A2(n15322), .ZN(n15340) );
  INV_X1 U18523 ( .A(n15341), .ZN(n15323) );
  NAND3_X1 U18524 ( .A1(n15332), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15323), .ZN(n15333) );
  OAI21_X1 U18525 ( .B1(n15495), .B2(n15340), .A(n15333), .ZN(n15324) );
  NAND2_X1 U18526 ( .A1(n15324), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15325) );
  OAI211_X1 U18527 ( .C1(n16031), .C2(n16194), .A(n15326), .B(n15325), .ZN(
        n15327) );
  AOI21_X1 U18528 ( .B1(n15328), .B2(n16196), .A(n15327), .ZN(n15329) );
  OAI21_X1 U18529 ( .B1(n16199), .B2(n15330), .A(n15329), .ZN(P2_U3020) );
  NAND2_X1 U18530 ( .A1(n15331), .A2(n16183), .ZN(n15338) );
  NOR3_X1 U18531 ( .A1(n15495), .A2(n15340), .A3(n15332), .ZN(n15336) );
  OAI211_X1 U18532 ( .C1(n16042), .C2(n16177), .A(n15334), .B(n15333), .ZN(
        n15335) );
  AOI211_X1 U18533 ( .C1(n16045), .C2(n16182), .A(n15336), .B(n15335), .ZN(
        n15337) );
  OAI211_X1 U18534 ( .C1(n15339), .C2(n16187), .A(n15338), .B(n15337), .ZN(
        P2_U3021) );
  AOI21_X1 U18535 ( .B1(n15342), .B2(n15341), .A(n15340), .ZN(n15343) );
  AOI211_X1 U18536 ( .C1(n16049), .C2(n16192), .A(n15344), .B(n15343), .ZN(
        n15345) );
  OAI21_X1 U18537 ( .B1(n15346), .B2(n16194), .A(n15345), .ZN(n15347) );
  AOI21_X1 U18538 ( .B1(n15348), .B2(n16196), .A(n15347), .ZN(n15349) );
  OAI21_X1 U18539 ( .B1(n15350), .B2(n16199), .A(n15349), .ZN(P2_U3022) );
  NAND2_X1 U18540 ( .A1(n15351), .A2(n16183), .ZN(n15364) );
  INV_X1 U18541 ( .A(n15352), .ZN(n15362) );
  INV_X1 U18542 ( .A(n15353), .ZN(n15366) );
  AOI211_X1 U18543 ( .C1(n15359), .C2(n15372), .A(n15354), .B(n15366), .ZN(
        n15361) );
  INV_X1 U18544 ( .A(n15355), .ZN(n15356) );
  NAND2_X1 U18545 ( .A1(n15356), .A2(n16192), .ZN(n15357) );
  OAI211_X1 U18546 ( .C1(n15373), .C2(n15359), .A(n15358), .B(n15357), .ZN(
        n15360) );
  AOI211_X1 U18547 ( .C1(n15362), .C2(n16182), .A(n15361), .B(n15360), .ZN(
        n15363) );
  OAI211_X1 U18548 ( .C1(n15365), .C2(n16187), .A(n15364), .B(n15363), .ZN(
        P2_U3023) );
  NOR2_X1 U18549 ( .A1(n15366), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15375) );
  AOI21_X1 U18550 ( .B1(n15369), .B2(n15368), .A(n15367), .ZN(n16061) );
  NAND2_X1 U18551 ( .A1(n16061), .A2(n16192), .ZN(n15370) );
  OAI211_X1 U18552 ( .C1(n15373), .C2(n15372), .A(n15371), .B(n15370), .ZN(
        n15374) );
  AOI211_X1 U18553 ( .C1(n15687), .C2(n16182), .A(n15375), .B(n15374), .ZN(
        n15378) );
  OR2_X1 U18554 ( .A1(n15376), .A2(n16187), .ZN(n15377) );
  OAI211_X1 U18555 ( .C1(n15379), .C2(n16199), .A(n15378), .B(n15377), .ZN(
        P2_U3024) );
  NAND2_X1 U18556 ( .A1(n16192), .A2(n15380), .ZN(n15381) );
  OAI211_X1 U18557 ( .C1(n15383), .C2(n20968), .A(n15382), .B(n15381), .ZN(
        n15384) );
  AOI21_X1 U18558 ( .B1(n15385), .B2(n20968), .A(n15384), .ZN(n15386) );
  OAI21_X1 U18559 ( .B1(n15387), .B2(n16194), .A(n15386), .ZN(n15388) );
  AOI21_X1 U18560 ( .B1(n15389), .B2(n16183), .A(n15388), .ZN(n15390) );
  OAI21_X1 U18561 ( .B1(n15391), .B2(n16187), .A(n15390), .ZN(P2_U3025) );
  XNOR2_X1 U18562 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15398) );
  OR2_X1 U18563 ( .A1(n15393), .A2(n15392), .ZN(n15394) );
  AND2_X1 U18564 ( .A1(n12924), .A2(n15394), .ZN(n18855) );
  AOI21_X1 U18565 ( .B1(n16192), .B2(n18855), .A(n15395), .ZN(n15397) );
  NAND3_X1 U18566 ( .A1(n15408), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15440), .ZN(n15396) );
  OAI211_X1 U18567 ( .C1(n15410), .C2(n15398), .A(n15397), .B(n15396), .ZN(
        n15401) );
  NOR2_X1 U18568 ( .A1(n15399), .A2(n16199), .ZN(n15400) );
  AOI211_X1 U18569 ( .C1(n18856), .C2(n16182), .A(n15401), .B(n15400), .ZN(
        n15402) );
  OAI21_X1 U18570 ( .B1(n15403), .B2(n16187), .A(n15402), .ZN(P2_U3026) );
  NOR2_X1 U18571 ( .A1(n15495), .A2(n15404), .ZN(n15407) );
  OAI21_X1 U18572 ( .B1(n16177), .B2(n18878), .A(n15405), .ZN(n15406) );
  AOI21_X1 U18573 ( .B1(n15408), .B2(n15407), .A(n15406), .ZN(n15409) );
  OAI21_X1 U18574 ( .B1(n15410), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15409), .ZN(n15411) );
  AOI21_X1 U18575 ( .B1(n18876), .B2(n16182), .A(n15411), .ZN(n15414) );
  NAND2_X1 U18576 ( .A1(n15412), .A2(n16183), .ZN(n15413) );
  OAI211_X1 U18577 ( .C1(n15415), .C2(n16187), .A(n15414), .B(n15413), .ZN(
        P2_U3027) );
  NAND2_X1 U18578 ( .A1(n15417), .A2(n15416), .ZN(n15418) );
  AND2_X1 U18579 ( .A1(n15419), .A2(n15418), .ZN(n18887) );
  INV_X1 U18580 ( .A(n15420), .ZN(n15423) );
  NOR3_X1 U18581 ( .A1(n15421), .A2(n15495), .A3(n15425), .ZN(n15422) );
  AOI211_X1 U18582 ( .C1(n16192), .C2(n18887), .A(n15423), .B(n15422), .ZN(
        n15427) );
  NAND3_X1 U18583 ( .A1(n15467), .A2(n10314), .A3(n15425), .ZN(n15426) );
  OAI211_X1 U18584 ( .C1(n18889), .C2(n16194), .A(n15427), .B(n15426), .ZN(
        n15428) );
  AOI21_X1 U18585 ( .B1(n15429), .B2(n16183), .A(n15428), .ZN(n15430) );
  OAI21_X1 U18586 ( .B1(n15431), .B2(n16187), .A(n15430), .ZN(P2_U3028) );
  OAI21_X1 U18587 ( .B1(n16177), .B2(n18901), .A(n15432), .ZN(n15436) );
  AOI22_X1 U18588 ( .A1(n15236), .A2(n16183), .B1(n15433), .B2(n15467), .ZN(
        n15434) );
  NOR2_X1 U18589 ( .A1(n15434), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15435) );
  AOI211_X1 U18590 ( .C1(n18899), .C2(n16182), .A(n15436), .B(n15435), .ZN(
        n15446) );
  INV_X1 U18591 ( .A(n15437), .ZN(n15439) );
  OAI21_X1 U18592 ( .B1(n16183), .B2(n15439), .A(n15438), .ZN(n15442) );
  NAND2_X1 U18593 ( .A1(n15441), .A2(n15440), .ZN(n15459) );
  OAI211_X1 U18594 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15443), .A(
        n15442), .B(n15459), .ZN(n15455) );
  NOR2_X1 U18595 ( .A1(n15481), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15444) );
  OAI21_X1 U18596 ( .B1(n15455), .B2(n15444), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15445) );
  OAI211_X1 U18597 ( .C1(n15447), .C2(n16187), .A(n15446), .B(n15445), .ZN(
        P2_U3029) );
  NOR2_X1 U18598 ( .A1(n15448), .A2(n15460), .ZN(n15449) );
  OR2_X1 U18599 ( .A1(n15450), .A2(n15449), .ZN(n19091) );
  OAI22_X1 U18600 ( .A1(n16177), .A2(n19091), .B1(n15451), .B2(n19034), .ZN(
        n15454) );
  INV_X1 U18601 ( .A(n15245), .ZN(n16081) );
  AOI21_X1 U18602 ( .B1(n16081), .B2(n16183), .A(n15467), .ZN(n15452) );
  NOR3_X1 U18603 ( .A1(n15452), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15466), .ZN(n15453) );
  AOI211_X1 U18604 ( .C1(n18909), .C2(n16182), .A(n15454), .B(n15453), .ZN(
        n15457) );
  NAND2_X1 U18605 ( .A1(n15455), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15456) );
  OAI211_X1 U18606 ( .C1(n15458), .C2(n16187), .A(n15457), .B(n15456), .ZN(
        P2_U3030) );
  NOR2_X1 U18607 ( .A1(n15459), .A2(n15466), .ZN(n15465) );
  NOR2_X1 U18608 ( .A1(n16152), .A2(n16164), .ZN(n16151) );
  INV_X1 U18609 ( .A(n15460), .ZN(n15461) );
  OAI21_X1 U18610 ( .B1(n15462), .B2(n16151), .A(n15461), .ZN(n19102) );
  OAI21_X1 U18611 ( .B1(n16177), .B2(n19102), .A(n15463), .ZN(n15464) );
  AOI211_X1 U18612 ( .C1(n15467), .C2(n15466), .A(n15465), .B(n15464), .ZN(
        n15468) );
  OAI21_X1 U18613 ( .B1(n16194), .B2(n18917), .A(n15468), .ZN(n15469) );
  AOI21_X1 U18614 ( .B1(n15470), .B2(n16183), .A(n15469), .ZN(n15471) );
  OAI21_X1 U18615 ( .B1(n15472), .B2(n16187), .A(n15471), .ZN(P2_U3031) );
  INV_X1 U18616 ( .A(n15496), .ZN(n15473) );
  OR2_X1 U18617 ( .A1(n16108), .A2(n15473), .ZN(n15491) );
  NAND2_X1 U18618 ( .A1(n15491), .A2(n11191), .ZN(n15475) );
  NAND2_X1 U18619 ( .A1(n15475), .A2(n15474), .ZN(n16097) );
  OR2_X1 U18620 ( .A1(n15477), .A2(n15476), .ZN(n15478) );
  NAND2_X1 U18621 ( .A1(n15479), .A2(n15478), .ZN(n16094) );
  AOI21_X1 U18622 ( .B1(n15480), .B2(n9894), .A(n16165), .ZN(n19108) );
  NAND2_X1 U18623 ( .A1(n16154), .A2(n16153), .ZN(n15484) );
  INV_X1 U18624 ( .A(n15484), .ZN(n15483) );
  OAI21_X1 U18625 ( .B1(n16154), .B2(n15481), .A(n15513), .ZN(n15482) );
  AOI21_X1 U18626 ( .B1(n15483), .B2(n11191), .A(n15482), .ZN(n16167) );
  AOI21_X1 U18627 ( .B1(n11191), .B2(n15484), .A(n16167), .ZN(n15486) );
  NOR2_X1 U18628 ( .A1(n19034), .A2(n11333), .ZN(n15485) );
  AOI211_X1 U18629 ( .C1(n16192), .C2(n19108), .A(n15486), .B(n15485), .ZN(
        n15487) );
  OAI21_X1 U18630 ( .B1(n15488), .B2(n16194), .A(n15487), .ZN(n15489) );
  AOI21_X1 U18631 ( .B1(n16094), .B2(n16196), .A(n15489), .ZN(n15490) );
  OAI21_X1 U18632 ( .B1(n16199), .B2(n16097), .A(n15490), .ZN(P2_U3034) );
  NOR2_X1 U18633 ( .A1(n16108), .A2(n16109), .ZN(n16107) );
  OAI21_X1 U18634 ( .B1(n16107), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15491), .ZN(n16102) );
  NOR2_X1 U18635 ( .A1(n9923), .A2(n15493), .ZN(n15494) );
  XNOR2_X1 U18636 ( .A(n15492), .B(n15494), .ZN(n16101) );
  AOI21_X1 U18637 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15513), .A(
        n15495), .ZN(n16180) );
  INV_X1 U18638 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19800) );
  NOR2_X1 U18639 ( .A1(n19800), .A2(n19034), .ZN(n15499) );
  NAND2_X1 U18640 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16153), .ZN(
        n16176) );
  AOI211_X1 U18641 ( .C1(n15497), .C2(n16109), .A(n15496), .B(n16176), .ZN(
        n15498) );
  AOI211_X1 U18642 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16180), .A(
        n15499), .B(n15498), .ZN(n15504) );
  OAI21_X1 U18643 ( .B1(n15501), .B2(n15500), .A(n9894), .ZN(n19110) );
  INV_X1 U18644 ( .A(n19110), .ZN(n15502) );
  AOI22_X1 U18645 ( .A1(n18961), .A2(n16182), .B1(n16192), .B2(n15502), .ZN(
        n15503) );
  OAI211_X1 U18646 ( .C1(n16101), .C2(n16187), .A(n15504), .B(n15503), .ZN(
        n15505) );
  INV_X1 U18647 ( .A(n15505), .ZN(n15506) );
  OAI21_X1 U18648 ( .B1(n16102), .B2(n16199), .A(n15506), .ZN(P2_U3035) );
  NAND3_X1 U18649 ( .A1(n15507), .A2(n16183), .A3(n16108), .ZN(n15516) );
  NAND2_X1 U18650 ( .A1(n16153), .A2(n15508), .ZN(n15512) );
  OAI21_X1 U18651 ( .B1(n15509), .B2(n16190), .A(n16174), .ZN(n19114) );
  INV_X1 U18652 ( .A(n19114), .ZN(n15510) );
  AOI22_X1 U18653 ( .A1(n16192), .A2(n15510), .B1(n16202), .B2(
        P2_REIP_REG_9__SCAN_IN), .ZN(n15511) );
  OAI211_X1 U18654 ( .C1(n15513), .C2(n15508), .A(n15512), .B(n15511), .ZN(
        n15514) );
  AOI21_X1 U18655 ( .B1(n16182), .B2(n18982), .A(n15514), .ZN(n15515) );
  OAI211_X1 U18656 ( .C1(n15517), .C2(n16187), .A(n15516), .B(n15515), .ZN(
        P2_U3037) );
  NAND3_X1 U18657 ( .A1(n15518), .A2(n16183), .A3(n15275), .ZN(n15529) );
  INV_X1 U18658 ( .A(n15519), .ZN(n16204) );
  OAI21_X1 U18659 ( .B1(n15522), .B2(n15521), .A(n15520), .ZN(n19119) );
  INV_X1 U18660 ( .A(n19119), .ZN(n15524) );
  OAI22_X1 U18661 ( .A1(n16189), .A2(n15527), .B1(n19794), .B2(n19034), .ZN(
        n15523) );
  AOI21_X1 U18662 ( .B1(n15524), .B2(n16192), .A(n15523), .ZN(n15525) );
  OAI21_X1 U18663 ( .B1(n16194), .B2(n19002), .A(n15525), .ZN(n15526) );
  AOI21_X1 U18664 ( .B1(n16204), .B2(n15527), .A(n15526), .ZN(n15528) );
  OAI211_X1 U18665 ( .C1(n15530), .C2(n16187), .A(n15529), .B(n15528), .ZN(
        P2_U3039) );
  OAI21_X1 U18666 ( .B1(n15531), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15532), .ZN(n16139) );
  INV_X1 U18667 ( .A(n15533), .ZN(n15535) );
  NAND3_X1 U18668 ( .A1(n13628), .A2(n15535), .A3(n15534), .ZN(n15536) );
  NAND2_X1 U18669 ( .A1(n15537), .A2(n15536), .ZN(n19122) );
  NOR2_X1 U18670 ( .A1(n11312), .A2(n19034), .ZN(n15538) );
  AOI21_X1 U18671 ( .B1(n15540), .B2(n15539), .A(n15538), .ZN(n15543) );
  NAND2_X1 U18672 ( .A1(n15541), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15542) );
  OAI211_X1 U18673 ( .C1(n19122), .C2(n16177), .A(n15543), .B(n15542), .ZN(
        n15547) );
  XNOR2_X1 U18674 ( .A(n15544), .B(n15545), .ZN(n16136) );
  NOR2_X1 U18675 ( .A1(n16136), .A2(n16187), .ZN(n15546) );
  AOI211_X1 U18676 ( .C1(n19015), .C2(n16182), .A(n15547), .B(n15546), .ZN(
        n15548) );
  OAI21_X1 U18677 ( .B1(n16199), .B2(n16139), .A(n15548), .ZN(P2_U3040) );
  OAI22_X1 U18678 ( .A1(n16187), .A2(n15549), .B1(n16194), .B2(n9968), .ZN(
        n15550) );
  AOI21_X1 U18679 ( .B1(n15551), .B2(n13015), .A(n15550), .ZN(n15558) );
  INV_X1 U18680 ( .A(n15552), .ZN(n15554) );
  AOI22_X1 U18681 ( .A1(n15554), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n16183), .B2(n15553), .ZN(n15557) );
  NAND2_X1 U18682 ( .A1(n16192), .A2(n19065), .ZN(n15555) );
  NAND4_X1 U18683 ( .A1(n15558), .A2(n15557), .A3(n15556), .A4(n15555), .ZN(
        P2_U3046) );
  INV_X1 U18684 ( .A(n16252), .ZN(n15593) );
  INV_X1 U18685 ( .A(n15559), .ZN(n15561) );
  NAND2_X1 U18686 ( .A1(n15561), .A2(n15560), .ZN(n15569) );
  MUX2_X1 U18687 ( .A(n11464), .B(n15569), .S(n15562), .Z(n15563) );
  AOI21_X1 U18688 ( .B1(n12485), .B2(n15576), .A(n15563), .ZN(n16213) );
  INV_X1 U18689 ( .A(n15564), .ZN(n15565) );
  OAI222_X1 U18690 ( .A1(n15593), .A2(n12494), .B1(n15592), .B2(n16213), .C1(
        n11393), .C2(n15565), .ZN(n15566) );
  MUX2_X1 U18691 ( .A(n15566), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15594), .Z(P2_U3601) );
  NAND2_X1 U18692 ( .A1(n12489), .A2(n15576), .ZN(n15571) );
  NOR2_X1 U18693 ( .A1(n10856), .A2(n15567), .ZN(n15568) );
  AOI22_X1 U18694 ( .A1(n15569), .A2(n15568), .B1(n11464), .B2(n10795), .ZN(
        n15570) );
  AND2_X1 U18695 ( .A1(n15571), .A2(n15570), .ZN(n16214) );
  INV_X1 U18696 ( .A(n15572), .ZN(n15574) );
  OAI222_X1 U18697 ( .A1(n19868), .A2(n15593), .B1(n15592), .B2(n16214), .C1(
        n15574), .C2(n15573), .ZN(n15575) );
  MUX2_X1 U18698 ( .A(n15575), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15594), .Z(P2_U3600) );
  INV_X1 U18699 ( .A(n15576), .ZN(n15577) );
  OR2_X1 U18700 ( .A1(n15578), .A2(n15577), .ZN(n15591) );
  INV_X1 U18701 ( .A(n9799), .ZN(n15580) );
  INV_X1 U18702 ( .A(n15584), .ZN(n15579) );
  AOI21_X1 U18703 ( .B1(n11464), .B2(n15580), .A(n15579), .ZN(n15581) );
  OAI21_X1 U18704 ( .B1(n15582), .B2(n10867), .A(n15581), .ZN(n15583) );
  INV_X1 U18705 ( .A(n15583), .ZN(n15587) );
  AOI22_X1 U18706 ( .A1(n15585), .A2(n15584), .B1(n9799), .B2(n11464), .ZN(
        n15586) );
  MUX2_X1 U18707 ( .A(n15587), .B(n15586), .S(n10676), .Z(n15589) );
  AND2_X1 U18708 ( .A1(n15589), .A2(n15588), .ZN(n15590) );
  AND2_X1 U18709 ( .A1(n15591), .A2(n15590), .ZN(n16220) );
  OAI22_X1 U18710 ( .A1(n19846), .A2(n15593), .B1(n15592), .B2(n16220), .ZN(
        n15595) );
  MUX2_X1 U18711 ( .A(n15595), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15594), .Z(P2_U3596) );
  INV_X1 U18712 ( .A(n15596), .ZN(n19648) );
  NAND2_X1 U18713 ( .A1(n19275), .A2(n19648), .ZN(n15597) );
  OR2_X1 U18714 ( .A1(n15596), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19651) );
  OAI21_X1 U18715 ( .B1(n19698), .B2(n15597), .A(n19651), .ZN(n15604) );
  INV_X1 U18716 ( .A(n15598), .ZN(n15599) );
  AND2_X1 U18717 ( .A1(n15599), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19751) );
  INV_X1 U18718 ( .A(n19751), .ZN(n15600) );
  NAND2_X1 U18719 ( .A1(n15604), .A2(n15600), .ZN(n15601) );
  OAI211_X1 U18720 ( .C1(n15603), .C2(n19654), .A(n15601), .B(n19469), .ZN(
        n15602) );
  AND2_X1 U18721 ( .A1(n19466), .A2(n16209), .ZN(n15605) );
  INV_X1 U18722 ( .A(n15605), .ZN(n15647) );
  INV_X1 U18723 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18166) );
  OAI22_X2 U18724 ( .A1(n14590), .A2(n15651), .B1(n18166), .B2(n15650), .ZN(
        n19662) );
  OAI21_X1 U18725 ( .B1(n15603), .B2(n15605), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15607) );
  OAI21_X1 U18726 ( .B1(n19751), .B2(n15605), .A(n15604), .ZN(n15606) );
  NAND2_X1 U18727 ( .A1(n19204), .A2(n19707), .ZN(n19665) );
  NAND2_X1 U18728 ( .A1(n16231), .A2(n15646), .ZN(n19248) );
  OAI22_X1 U18729 ( .A1(n15648), .A2(n19665), .B1(n15647), .B2(n19248), .ZN(
        n15609) );
  AOI21_X1 U18730 ( .B1(n19662), .B2(n19265), .A(n15609), .ZN(n15611) );
  INV_X1 U18731 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20149) );
  INV_X1 U18732 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n21086) );
  OAI22_X2 U18733 ( .A1(n20149), .A2(n15651), .B1(n21086), .B2(n15650), .ZN(
        n19710) );
  NAND2_X1 U18734 ( .A1(n19710), .A2(n19698), .ZN(n15610) );
  OAI211_X1 U18735 ( .C1(n15655), .C2(n15612), .A(n15611), .B(n15610), .ZN(
        P2_U3048) );
  INV_X1 U18736 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n15613) );
  OAI22_X2 U18737 ( .A1(n14584), .A2(n15651), .B1(n15613), .B2(n15650), .ZN(
        n19666) );
  NOR2_X1 U18738 ( .A1(n19214), .A2(n19536), .ZN(n19715) );
  INV_X1 U18739 ( .A(n19715), .ZN(n19669) );
  NAND2_X1 U18740 ( .A1(n15614), .A2(n15646), .ZN(n19251) );
  OAI22_X1 U18741 ( .A1(n15648), .A2(n19669), .B1(n15647), .B2(n19251), .ZN(
        n15615) );
  AOI21_X1 U18742 ( .B1(n19666), .B2(n19265), .A(n15615), .ZN(n15617) );
  INV_X1 U18743 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18175) );
  OAI22_X2 U18744 ( .A1(n20168), .A2(n15651), .B1(n18175), .B2(n15650), .ZN(
        n19716) );
  NAND2_X1 U18745 ( .A1(n19716), .A2(n19698), .ZN(n15616) );
  OAI211_X1 U18746 ( .C1(n15655), .C2(n15618), .A(n15617), .B(n15616), .ZN(
        P2_U3049) );
  INV_X1 U18747 ( .A(n19720), .ZN(n15619) );
  OAI22_X1 U18748 ( .A1(n15648), .A2(n19673), .B1(n15647), .B2(n15619), .ZN(
        n15620) );
  AOI21_X1 U18749 ( .B1(n19670), .B2(n19265), .A(n15620), .ZN(n15622) );
  NAND2_X1 U18750 ( .A1(n19722), .A2(n19698), .ZN(n15621) );
  OAI211_X1 U18751 ( .C1(n15655), .C2(n15623), .A(n15622), .B(n15621), .ZN(
        P2_U3050) );
  INV_X1 U18752 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20181) );
  INV_X1 U18753 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15624) );
  OAI22_X2 U18754 ( .A1(n20181), .A2(n15651), .B1(n15624), .B2(n15650), .ZN(
        n19674) );
  NOR2_X1 U18755 ( .A1(n19216), .A2(n19536), .ZN(n19727) );
  INV_X1 U18756 ( .A(n19727), .ZN(n19677) );
  NAND2_X1 U18757 ( .A1(n15625), .A2(n15646), .ZN(n19256) );
  OAI22_X1 U18758 ( .A1(n15648), .A2(n19677), .B1(n15647), .B2(n19256), .ZN(
        n15626) );
  AOI21_X1 U18759 ( .B1(n19674), .B2(n19265), .A(n15626), .ZN(n15628) );
  INV_X1 U18760 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20184) );
  OAI22_X2 U18761 ( .A1(n20184), .A2(n15651), .B1(n15053), .B2(n15650), .ZN(
        n19728) );
  NAND2_X1 U18762 ( .A1(n19728), .A2(n19698), .ZN(n15627) );
  OAI211_X1 U18763 ( .C1(n15655), .C2(n15629), .A(n15628), .B(n15627), .ZN(
        P2_U3051) );
  INV_X1 U18764 ( .A(n19732), .ZN(n15630) );
  OAI22_X1 U18765 ( .A1(n15648), .A2(n19681), .B1(n15647), .B2(n15630), .ZN(
        n15631) );
  AOI21_X1 U18766 ( .B1(n19678), .B2(n19265), .A(n15631), .ZN(n15633) );
  NAND2_X1 U18767 ( .A1(n19734), .A2(n19698), .ZN(n15632) );
  OAI211_X1 U18768 ( .C1(n15655), .C2(n15634), .A(n15633), .B(n15632), .ZN(
        P2_U3052) );
  INV_X1 U18769 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18193) );
  OAI22_X2 U18770 ( .A1(n14571), .A2(n15651), .B1(n18193), .B2(n15650), .ZN(
        n19682) );
  NOR2_X1 U18771 ( .A1(n19218), .A2(n19536), .ZN(n19739) );
  INV_X1 U18772 ( .A(n19739), .ZN(n19685) );
  NAND2_X1 U18773 ( .A1(n15635), .A2(n15646), .ZN(n19261) );
  OAI22_X1 U18774 ( .A1(n15648), .A2(n19685), .B1(n15647), .B2(n19261), .ZN(
        n15636) );
  AOI21_X1 U18775 ( .B1(n19682), .B2(n19265), .A(n15636), .ZN(n15638) );
  INV_X1 U18776 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20198) );
  OAI22_X2 U18777 ( .A1(n12820), .A2(n15650), .B1(n20198), .B2(n15651), .ZN(
        n19740) );
  NAND2_X1 U18778 ( .A1(n19740), .A2(n19698), .ZN(n15637) );
  OAI211_X1 U18779 ( .C1(n15655), .C2(n15639), .A(n15638), .B(n15637), .ZN(
        P2_U3053) );
  INV_X1 U18780 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15644) );
  INV_X1 U18781 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18197) );
  OAI22_X2 U18782 ( .A1(n14567), .A2(n15651), .B1(n18197), .B2(n15650), .ZN(
        n19686) );
  INV_X1 U18783 ( .A(n19745), .ZN(n19689) );
  NAND2_X1 U18784 ( .A1(n15640), .A2(n15646), .ZN(n19264) );
  OAI22_X1 U18785 ( .A1(n15648), .A2(n19689), .B1(n15647), .B2(n19264), .ZN(
        n15641) );
  AOI21_X1 U18786 ( .B1(n19686), .B2(n19265), .A(n15641), .ZN(n15643) );
  INV_X1 U18787 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20205) );
  OAI22_X2 U18788 ( .A1(n14324), .A2(n15650), .B1(n20205), .B2(n15651), .ZN(
        n19746) );
  NAND2_X1 U18789 ( .A1(n19746), .A2(n19698), .ZN(n15642) );
  OAI211_X1 U18790 ( .C1(n15655), .C2(n15644), .A(n15643), .B(n15642), .ZN(
        P2_U3054) );
  INV_X1 U18791 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18202) );
  OAI22_X2 U18792 ( .A1(n18202), .A2(n15650), .B1(n14562), .B2(n15651), .ZN(
        n19692) );
  INV_X1 U18793 ( .A(n15645), .ZN(n19222) );
  NOR2_X1 U18794 ( .A1(n19222), .A2(n19536), .ZN(n19752) );
  INV_X1 U18795 ( .A(n19752), .ZN(n19696) );
  OAI22_X1 U18796 ( .A1(n15648), .A2(n19696), .B1(n15647), .B2(n19269), .ZN(
        n15649) );
  AOI21_X1 U18797 ( .B1(n19692), .B2(n19265), .A(n15649), .ZN(n15653) );
  INV_X1 U18798 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n16403) );
  OAI22_X2 U18799 ( .A1(n20213), .A2(n15651), .B1(n16403), .B2(n15650), .ZN(
        n19754) );
  NAND2_X1 U18800 ( .A1(n19754), .A2(n19698), .ZN(n15652) );
  OAI211_X1 U18801 ( .C1(n15655), .C2(n15654), .A(n15653), .B(n15652), .ZN(
        P2_U3055) );
  INV_X1 U18802 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17433) );
  INV_X1 U18803 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17365) );
  INV_X1 U18804 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17286) );
  NAND3_X1 U18805 ( .A1(n18172), .A2(n18813), .A3(n16817), .ZN(n15658) );
  INV_X1 U18806 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17406) );
  NAND4_X1 U18807 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(P3_EAX_REG_5__SCAN_IN), .ZN(n15660) );
  NOR2_X1 U18808 ( .A1(n17406), .A2(n15660), .ZN(n17326) );
  NAND4_X1 U18809 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_1__SCAN_IN), .A4(n17326), .ZN(n17290) );
  INV_X1 U18810 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n21142) );
  INV_X1 U18811 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17463) );
  INV_X1 U18812 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17397) );
  NAND2_X1 U18813 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .ZN(n17296) );
  NOR4_X1 U18814 ( .A1(n21142), .A2(n17463), .A3(n17397), .A4(n17296), .ZN(
        n15661) );
  NAND3_X1 U18815 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .ZN(n17249) );
  NAND3_X1 U18816 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .ZN(n15662) );
  NAND2_X1 U18817 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17244), .ZN(n17243) );
  NAND2_X1 U18818 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17239), .ZN(n17238) );
  NAND2_X1 U18819 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17218), .ZN(n17214) );
  NAND2_X1 U18820 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17209), .ZN(n17208) );
  NAND3_X1 U18821 ( .A1(n17350), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n17208), 
        .ZN(n15665) );
  NAND2_X1 U18822 ( .A1(n15663), .A2(n17321), .ZN(n17250) );
  NAND2_X1 U18823 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17279), .ZN(n15664) );
  OAI211_X1 U18824 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n17208), .A(n15665), .B(
        n15664), .ZN(P3_U2704) );
  NAND2_X1 U18825 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18387) );
  AOI221_X1 U18826 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18387), .C1(n15667), 
        .C2(n18387), .A(n15666), .ZN(n18164) );
  NOR2_X1 U18827 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18168), .ZN(
        n18252) );
  AOI211_X1 U18828 ( .C1(n18512), .C2(n15668), .A(n18161), .B(n18252), .ZN(
        n15669) );
  INV_X1 U18829 ( .A(n15669), .ZN(n18162) );
  AOI22_X1 U18830 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18164), .B1(
        n18162), .B2(n18650), .ZN(P3_U2865) );
  AOI21_X1 U18831 ( .B1(n15670), .B2(n17490), .A(n9878), .ZN(n15671) );
  XNOR2_X1 U18832 ( .A(n16284), .B(n15671), .ZN(n16299) );
  OAI21_X1 U18833 ( .B1(n18052), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15672), .ZN(n16319) );
  AOI21_X1 U18834 ( .B1(n18076), .B2(n17467), .A(n16319), .ZN(n15674) );
  OAI211_X1 U18835 ( .C1(n15674), .C2(n18142), .A(n15673), .B(n18109), .ZN(
        n15677) );
  NOR3_X1 U18836 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16295), .A3(
        n15675), .ZN(n15676) );
  AOI21_X1 U18837 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15677), .A(
        n15676), .ZN(n15678) );
  NAND2_X1 U18838 ( .A1(n9790), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16289) );
  OAI211_X1 U18839 ( .C1(n16299), .C2(n10104), .A(n15678), .B(n16289), .ZN(
        P3_U2833) );
  AOI211_X1 U18840 ( .C1(n15681), .C2(n15679), .A(n15680), .B(n19061), .ZN(
        n15686) );
  INV_X1 U18841 ( .A(n15682), .ZN(n15684) );
  AOI22_X1 U18842 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19080), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19049), .ZN(n15683) );
  OAI21_X1 U18843 ( .B1(n15684), .B2(n19070), .A(n15683), .ZN(n15685) );
  AOI211_X1 U18844 ( .C1(P2_EBX_REG_22__SCAN_IN), .C2(n19063), .A(n15686), .B(
        n15685), .ZN(n15689) );
  AOI22_X1 U18845 ( .A1(n15687), .A2(n19062), .B1(n16061), .B2(n19064), .ZN(
        n15688) );
  NAND2_X1 U18846 ( .A1(n15689), .A2(n15688), .ZN(P2_U2833) );
  AOI21_X1 U18847 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15691), .A(
        n15690), .ZN(n15697) );
  AOI211_X1 U18848 ( .C1(n15694), .C2(n15697), .A(n15693), .B(n15692), .ZN(
        n15695) );
  INV_X1 U18849 ( .A(n15695), .ZN(n15696) );
  OAI211_X1 U18850 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n15697), .A(
        n15696), .B(n20545), .ZN(n15699) );
  INV_X1 U18851 ( .A(n15699), .ZN(n15701) );
  AOI21_X1 U18852 ( .B1(n15699), .B2(n20420), .A(n15698), .ZN(n15700) );
  AOI21_X1 U18853 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15701), .A(
        n15700), .ZN(n15703) );
  INV_X1 U18854 ( .A(n15703), .ZN(n15706) );
  INV_X1 U18855 ( .A(n15702), .ZN(n15705) );
  OAI21_X1 U18856 ( .B1(n15703), .B2(n15702), .A(n20618), .ZN(n15704) );
  OAI21_X1 U18857 ( .B1(n15706), .B2(n15705), .A(n15704), .ZN(n15715) );
  INV_X1 U18858 ( .A(n15707), .ZN(n15711) );
  OAI21_X1 U18859 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15708), .ZN(n15709) );
  NAND4_X1 U18860 ( .A1(n15712), .A2(n15711), .A3(n15710), .A4(n15709), .ZN(
        n15713) );
  AOI211_X1 U18861 ( .C1(n15715), .C2(n20143), .A(n15714), .B(n15713), .ZN(
        n15716) );
  INV_X1 U18862 ( .A(n15716), .ZN(n15725) );
  NAND2_X1 U18863 ( .A1(n15718), .A2(n15717), .ZN(n15720) );
  AOI21_X1 U18864 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATE2_REG_1__SCAN_IN), .A(n13230), .ZN(n20726) );
  NOR2_X1 U18865 ( .A1(n15722), .A2(n15730), .ZN(n15996) );
  INV_X1 U18866 ( .A(n15996), .ZN(n15719) );
  OAI211_X1 U18867 ( .C1(n15721), .C2(n15720), .A(n20726), .B(n15719), .ZN(
        n16001) );
  AOI221_X1 U18868 ( .B1(n20824), .B2(n15722), .C1(n15725), .C2(n15722), .A(
        n16001), .ZN(n15729) );
  NOR2_X1 U18869 ( .A1(n20823), .A2(n20805), .ZN(n15728) );
  OAI21_X1 U18870 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n15730), .A(n13230), 
        .ZN(n15999) );
  NOR2_X1 U18871 ( .A1(n15729), .A2(n20824), .ZN(n16004) );
  OAI211_X1 U18872 ( .C1(n15996), .C2(n15999), .A(n16004), .B(n15723), .ZN(
        n15724) );
  AOI21_X1 U18873 ( .B1(n15726), .B2(n15725), .A(n15724), .ZN(n15727) );
  AOI221_X1 U18874 ( .B1(n15729), .B2(n20824), .C1(n15728), .C2(n20824), .A(
        n15727), .ZN(P1_U3161) );
  INV_X1 U18875 ( .A(HOLD), .ZN(n20740) );
  NOR2_X1 U18876 ( .A1(n11841), .A2(n20740), .ZN(n20730) );
  AOI22_X1 U18877 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15732) );
  NAND2_X1 U18878 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15730), .ZN(n20728) );
  OAI211_X1 U18879 ( .C1(n20730), .C2(n15732), .A(n15731), .B(n20728), .ZN(
        P1_U3195) );
  INV_X1 U18880 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16405) );
  NOR2_X1 U18881 ( .A1(n20045), .A2(n16405), .ZN(P1_U2905) );
  NOR3_X1 U18882 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15733) );
  INV_X1 U18883 ( .A(n19900), .ZN(n16253) );
  NOR2_X1 U18884 ( .A1(n19901), .A2(n19762), .ZN(n16248) );
  NOR4_X1 U18885 ( .A1(n15733), .A2(n16253), .A3(n16259), .A4(n16248), .ZN(
        P2_U3178) );
  INV_X1 U18886 ( .A(n15734), .ZN(n19890) );
  OAI221_X1 U18887 ( .B1(n15736), .B2(n15735), .C1(n19890), .C2(n15735), .A(
        n19536), .ZN(n19882) );
  NOR2_X1 U18888 ( .A1(n16246), .A2(n19882), .ZN(P2_U3047) );
  NAND2_X1 U18889 ( .A1(n18206), .A2(n15738), .ZN(n17324) );
  INV_X1 U18890 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17415) );
  AOI22_X1 U18891 ( .A1(n17354), .A2(BUF2_REG_0__SCAN_IN), .B1(n17353), .B2(
        n17844), .ZN(n15737) );
  OAI221_X1 U18892 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17324), .C1(n17415), 
        .C2(n15738), .A(n15737), .ZN(P3_U2735) );
  AOI21_X1 U18893 ( .B1(n15740), .B2(n15739), .A(n15816), .ZN(n15770) );
  INV_X1 U18894 ( .A(n15770), .ZN(n15751) );
  NAND2_X1 U18895 ( .A1(n15741), .A2(n20948), .ZN(n15753) );
  AOI22_X1 U18896 ( .A1(n15809), .A2(n15742), .B1(n19996), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n15743) );
  OAI21_X1 U18897 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15744), .A(n15743), 
        .ZN(n15749) );
  INV_X1 U18898 ( .A(n15745), .ZN(n15746) );
  OAI22_X1 U18899 ( .A1(n15747), .A2(n19947), .B1(n15746), .B2(n20012), .ZN(
        n15748) );
  AOI211_X1 U18900 ( .C1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n19998), .A(
        n15749), .B(n15748), .ZN(n15750) );
  OAI221_X1 U18901 ( .B1(n20779), .B2(n15751), .C1(n20779), .C2(n15753), .A(
        n15750), .ZN(P1_U2818) );
  NOR2_X1 U18902 ( .A1(n20948), .A2(n15751), .ZN(n15757) );
  NOR2_X1 U18903 ( .A1(n15753), .A2(n15752), .ZN(n15756) );
  INV_X1 U18904 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15754) );
  OAI22_X1 U18905 ( .A1(n19986), .A2(n14069), .B1(n19984), .B2(n15754), .ZN(
        n15755) );
  NOR3_X1 U18906 ( .A1(n15757), .A2(n15756), .A3(n15755), .ZN(n15761) );
  AOI22_X1 U18907 ( .A1(n15759), .A2(n19965), .B1(n15758), .B2(n19988), .ZN(
        n15760) );
  OAI211_X1 U18908 ( .C1(n15762), .C2(n20002), .A(n15761), .B(n15760), .ZN(
        P1_U2819) );
  AOI22_X1 U18909 ( .A1(n15809), .A2(n15763), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n19996), .ZN(n15772) );
  INV_X1 U18910 ( .A(n15764), .ZN(n15776) );
  NAND2_X1 U18911 ( .A1(n15776), .A2(n15765), .ZN(n15790) );
  OAI21_X1 U18912 ( .B1(n15774), .B2(n15790), .A(n20776), .ZN(n15769) );
  OAI22_X1 U18913 ( .A1(n15767), .A2(n19947), .B1(n15766), .B2(n20012), .ZN(
        n15768) );
  AOI21_X1 U18914 ( .B1(n15770), .B2(n15769), .A(n15768), .ZN(n15771) );
  OAI211_X1 U18915 ( .C1(n15773), .C2(n19986), .A(n15772), .B(n15771), .ZN(
        P1_U2820) );
  OAI21_X1 U18916 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n15774), .ZN(n15782) );
  OAI21_X1 U18917 ( .B1(n15816), .B2(n15776), .A(n15775), .ZN(n15793) );
  AOI22_X1 U18918 ( .A1(n15793), .A2(P1_REIP_REG_19__SCAN_IN), .B1(n19996), 
        .B2(P1_EBX_REG_19__SCAN_IN), .ZN(n15777) );
  OAI21_X1 U18919 ( .B1(n15834), .B2(n20002), .A(n15777), .ZN(n15778) );
  AOI211_X1 U18920 ( .C1(n19998), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n12122), .B(n15778), .ZN(n15781) );
  INV_X1 U18921 ( .A(n15779), .ZN(n15831) );
  AOI22_X1 U18922 ( .A1(n15831), .A2(n19965), .B1(n15877), .B2(n19988), .ZN(
        n15780) );
  OAI211_X1 U18923 ( .C1(n15790), .C2(n15782), .A(n15781), .B(n15780), .ZN(
        P1_U2821) );
  AOI22_X1 U18924 ( .A1(n15793), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_EBX_REG_18__SCAN_IN), .B2(n19996), .ZN(n15783) );
  OAI211_X1 U18925 ( .C1(n19986), .C2(n15784), .A(n15783), .B(n20135), .ZN(
        n15787) );
  OAI22_X1 U18926 ( .A1(n15785), .A2(n19947), .B1(n20012), .B2(n15884), .ZN(
        n15786) );
  AOI211_X1 U18927 ( .C1(n15788), .C2(n15809), .A(n15787), .B(n15786), .ZN(
        n15789) );
  OAI21_X1 U18928 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n15790), .A(n15789), 
        .ZN(P1_U2822) );
  AOI22_X1 U18929 ( .A1(n19998), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n19996), .B2(P1_EBX_REG_17__SCAN_IN), .ZN(n15798) );
  AOI21_X1 U18930 ( .B1(n15809), .B2(n15835), .A(n12122), .ZN(n15797) );
  INV_X1 U18931 ( .A(n15791), .ZN(n15836) );
  AOI22_X1 U18932 ( .A1(n15836), .A2(n19965), .B1(n15792), .B2(n19988), .ZN(
        n15796) );
  OAI221_X1 U18933 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(P1_REIP_REG_16__SCAN_IN), .C1(P1_REIP_REG_17__SCAN_IN), .C2(n15794), .A(n15793), .ZN(n15795) );
  NAND4_X1 U18934 ( .A1(n15798), .A2(n15797), .A3(n15796), .A4(n15795), .ZN(
        P1_U2823) );
  AOI22_X1 U18935 ( .A1(n15841), .A2(n19965), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n15799), .ZN(n15807) );
  OAI22_X1 U18936 ( .A1(n15825), .A2(n20012), .B1(n15800), .B2(n19984), .ZN(
        n15801) );
  INV_X1 U18937 ( .A(n15801), .ZN(n15802) );
  OAI211_X1 U18938 ( .C1(n19986), .C2(n15803), .A(n15802), .B(n20135), .ZN(
        n15804) );
  AOI211_X1 U18939 ( .C1(n15809), .C2(n15840), .A(n15805), .B(n15804), .ZN(
        n15806) );
  NAND2_X1 U18940 ( .A1(n15807), .A2(n15806), .ZN(P1_U2825) );
  AOI22_X1 U18941 ( .A1(n19998), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19996), .B2(P1_EBX_REG_12__SCAN_IN), .ZN(n15814) );
  AOI21_X1 U18942 ( .B1(n15808), .B2(n19988), .A(n12122), .ZN(n15813) );
  AOI22_X1 U18943 ( .A1(n15846), .A2(n15809), .B1(n19965), .B2(n15845), .ZN(
        n15812) );
  NOR2_X1 U18944 ( .A1(n20758), .A2(n15817), .ZN(n15815) );
  OAI21_X1 U18945 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(n15815), .A(n15810), 
        .ZN(n15811) );
  NAND4_X1 U18946 ( .A1(n15814), .A2(n15813), .A3(n15812), .A4(n15811), .ZN(
        P1_U2828) );
  AOI211_X1 U18947 ( .C1(n15817), .C2(n20758), .A(n15816), .B(n15815), .ZN(
        n15823) );
  INV_X1 U18948 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15821) );
  OAI22_X1 U18949 ( .A1(n15920), .A2(n20012), .B1(n19984), .B2(n15818), .ZN(
        n15819) );
  INV_X1 U18950 ( .A(n15819), .ZN(n15820) );
  OAI211_X1 U18951 ( .C1(n19986), .C2(n15821), .A(n15820), .B(n20135), .ZN(
        n15822) );
  AOI211_X1 U18952 ( .C1(n15856), .C2(n19965), .A(n15823), .B(n15822), .ZN(
        n15824) );
  OAI21_X1 U18953 ( .B1(n15859), .B2(n20002), .A(n15824), .ZN(P1_U2829) );
  INV_X1 U18954 ( .A(n15825), .ZN(n15826) );
  AOI22_X1 U18955 ( .A1(n15841), .A2(n20025), .B1(n20024), .B2(n15826), .ZN(
        n15827) );
  OAI21_X1 U18956 ( .B1(n20029), .B2(n15800), .A(n15827), .ZN(P1_U2857) );
  AOI22_X1 U18957 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15833) );
  OAI21_X1 U18958 ( .B1(n15852), .B2(n15828), .A(n14699), .ZN(n15830) );
  XNOR2_X1 U18959 ( .A(n15852), .B(n21133), .ZN(n15829) );
  XNOR2_X1 U18960 ( .A(n15830), .B(n15829), .ZN(n15878) );
  AOI22_X1 U18961 ( .A1(n15878), .A2(n20097), .B1(n20096), .B2(n15831), .ZN(
        n15832) );
  OAI211_X1 U18962 ( .C1(n20101), .C2(n15834), .A(n15833), .B(n15832), .ZN(
        P1_U2980) );
  AOI22_X1 U18963 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15838) );
  AOI22_X1 U18964 ( .A1(n15836), .A2(n20096), .B1(n15835), .B2(n15847), .ZN(
        n15837) );
  OAI211_X1 U18965 ( .C1(n15839), .C2(n19922), .A(n15838), .B(n15837), .ZN(
        P1_U2982) );
  AOI22_X1 U18966 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15843) );
  AOI22_X1 U18967 ( .A1(n15841), .A2(n20096), .B1(n15840), .B2(n15847), .ZN(
        n15842) );
  OAI211_X1 U18968 ( .C1(n15844), .C2(n19922), .A(n15843), .B(n15842), .ZN(
        P1_U2984) );
  AOI22_X1 U18969 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15849) );
  AOI22_X1 U18970 ( .A1(n15847), .A2(n15846), .B1(n20096), .B2(n15845), .ZN(
        n15848) );
  OAI211_X1 U18971 ( .C1(n15850), .C2(n19922), .A(n15849), .B(n15848), .ZN(
        P1_U2987) );
  AOI22_X1 U18972 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15858) );
  NOR2_X1 U18973 ( .A1(n14749), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15854) );
  NOR2_X1 U18974 ( .A1(n15851), .A2(n12061), .ZN(n15853) );
  MUX2_X1 U18975 ( .A(n15854), .B(n15853), .S(n15852), .Z(n15855) );
  XOR2_X1 U18976 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n15855), .Z(
        n15925) );
  AOI22_X1 U18977 ( .A1(n20097), .A2(n15925), .B1(n20096), .B2(n15856), .ZN(
        n15857) );
  OAI211_X1 U18978 ( .C1(n20101), .C2(n15859), .A(n15858), .B(n15857), .ZN(
        P1_U2988) );
  AOI22_X1 U18979 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15865) );
  NAND2_X1 U18980 ( .A1(n15862), .A2(n15861), .ZN(n15863) );
  XNOR2_X1 U18981 ( .A(n15860), .B(n15863), .ZN(n15970) );
  AOI22_X1 U18982 ( .A1(n15970), .A2(n20097), .B1(n20096), .B2(n20020), .ZN(
        n15864) );
  OAI211_X1 U18983 ( .C1(n20101), .C2(n19960), .A(n15865), .B(n15864), .ZN(
        P1_U2992) );
  AOI22_X1 U18984 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15870) );
  XNOR2_X1 U18985 ( .A(n15867), .B(n15961), .ZN(n15868) );
  XNOR2_X1 U18986 ( .A(n15866), .B(n15868), .ZN(n15976) );
  AOI22_X1 U18987 ( .A1(n15976), .A2(n20097), .B1(n20096), .B2(n19966), .ZN(
        n15869) );
  OAI211_X1 U18988 ( .C1(n20101), .C2(n19970), .A(n15870), .B(n15869), .ZN(
        P1_U2993) );
  AOI22_X1 U18989 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15876) );
  OAI21_X1 U18990 ( .B1(n15873), .B2(n15872), .A(n15871), .ZN(n15874) );
  INV_X1 U18991 ( .A(n15874), .ZN(n15985) );
  AOI22_X1 U18992 ( .A1(n15985), .A2(n20097), .B1(n20096), .B2(n20026), .ZN(
        n15875) );
  OAI211_X1 U18993 ( .C1(n20101), .C2(n19978), .A(n15876), .B(n15875), .ZN(
        P1_U2994) );
  AOI22_X1 U18994 ( .A1(n15878), .A2(n20123), .B1(n20126), .B2(n15877), .ZN(
        n15883) );
  INV_X1 U18995 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21098) );
  NOR2_X1 U18996 ( .A1(n20135), .A2(n21098), .ZN(n15879) );
  AOI221_X1 U18997 ( .B1(n15881), .B2(n21133), .C1(n15880), .C2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15879), .ZN(n15882) );
  NAND2_X1 U18998 ( .A1(n15883), .A2(n15882), .ZN(P1_U3012) );
  INV_X1 U18999 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20773) );
  NOR2_X1 U19000 ( .A1(n20135), .A2(n20773), .ZN(n15887) );
  OAI22_X1 U19001 ( .A1(n15885), .A2(n15935), .B1(n15936), .B2(n15884), .ZN(
        n15886) );
  AOI211_X1 U19002 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15888), .A(
        n15887), .B(n15886), .ZN(n15889) );
  OAI21_X1 U19003 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15890), .A(
        n15889), .ZN(P1_U3013) );
  AOI21_X1 U19004 ( .B1(n15892), .B2(n14860), .A(n15891), .ZN(n15894) );
  AOI22_X1 U19005 ( .A1(n12122), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n15894), 
        .B2(n15893), .ZN(n15898) );
  AOI22_X1 U19006 ( .A1(n15896), .A2(n20123), .B1(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15895), .ZN(n15897) );
  OAI211_X1 U19007 ( .C1(n15936), .C2(n15899), .A(n15898), .B(n15897), .ZN(
        P1_U3015) );
  INV_X1 U19008 ( .A(n15900), .ZN(n15907) );
  INV_X1 U19009 ( .A(n15901), .ZN(n15922) );
  NAND2_X1 U19010 ( .A1(n15902), .A2(n15903), .ZN(n15905) );
  OAI22_X1 U19011 ( .A1(n15922), .A2(n15905), .B1(n15904), .B2(n15903), .ZN(
        n15906) );
  AOI21_X1 U19012 ( .B1(n15907), .B2(n20123), .A(n15906), .ZN(n15909) );
  NAND2_X1 U19013 ( .A1(n12122), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n15908) );
  OAI211_X1 U19014 ( .C1(n15936), .C2(n15910), .A(n15909), .B(n15908), .ZN(
        P1_U3017) );
  NOR2_X1 U19015 ( .A1(n20135), .A2(n20763), .ZN(n15911) );
  AOI211_X1 U19016 ( .C1(n15914), .C2(n15913), .A(n15912), .B(n15911), .ZN(
        n15918) );
  AOI22_X1 U19017 ( .A1(n15916), .A2(n20123), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15915), .ZN(n15917) );
  OAI211_X1 U19018 ( .C1(n15936), .C2(n15919), .A(n15918), .B(n15917), .ZN(
        P1_U3018) );
  INV_X1 U19019 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15928) );
  INV_X1 U19020 ( .A(n15920), .ZN(n15921) );
  AOI22_X1 U19021 ( .A1(n12122), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20126), 
        .B2(n15921), .ZN(n15927) );
  NOR2_X1 U19022 ( .A1(n15923), .A2(n15922), .ZN(n20115) );
  AOI22_X1 U19023 ( .A1(n15925), .A2(n20123), .B1(n20115), .B2(n15924), .ZN(
        n15926) );
  OAI211_X1 U19024 ( .C1(n15929), .C2(n15928), .A(n15927), .B(n15926), .ZN(
        P1_U3020) );
  INV_X1 U19025 ( .A(n15930), .ZN(n20121) );
  AOI21_X1 U19026 ( .B1(n20121), .B2(n20128), .A(n20120), .ZN(n20102) );
  NAND2_X1 U19027 ( .A1(n15931), .A2(n20102), .ZN(n15933) );
  OAI21_X1 U19028 ( .B1(n15939), .B2(n15933), .A(n15932), .ZN(n15950) );
  INV_X1 U19029 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20756) );
  OAI222_X1 U19030 ( .A1(n15937), .A2(n15936), .B1(n20135), .B2(n20756), .C1(
        n15935), .C2(n15934), .ZN(n15938) );
  INV_X1 U19031 ( .A(n15938), .ZN(n15941) );
  NOR2_X1 U19032 ( .A1(n15939), .A2(n15979), .ZN(n15946) );
  OAI221_X1 U19033 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n12061), .C2(n15951), .A(
        n15946), .ZN(n15940) );
  OAI211_X1 U19034 ( .C1(n12061), .C2(n15950), .A(n15941), .B(n15940), .ZN(
        P1_U3021) );
  NAND2_X1 U19035 ( .A1(n15943), .A2(n15942), .ZN(n15944) );
  AND2_X1 U19036 ( .A1(n15945), .A2(n15944), .ZN(n20013) );
  AOI22_X1 U19037 ( .A1(n12122), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n20126), 
        .B2(n20013), .ZN(n15949) );
  AOI22_X1 U19038 ( .A1(n15947), .A2(n20123), .B1(n15951), .B2(n15946), .ZN(
        n15948) );
  OAI211_X1 U19039 ( .C1(n15951), .C2(n15950), .A(n15949), .B(n15948), .ZN(
        P1_U3022) );
  INV_X1 U19040 ( .A(n15952), .ZN(n15956) );
  NOR2_X1 U19041 ( .A1(n20106), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15984) );
  INV_X1 U19042 ( .A(n15984), .ZN(n15954) );
  AOI221_X1 U19043 ( .B1(n20128), .B2(n20121), .C1(n20106), .C2(n20121), .A(
        n15953), .ZN(n15989) );
  OAI21_X1 U19044 ( .B1(n15955), .B2(n15954), .A(n15989), .ZN(n15975) );
  AOI21_X1 U19045 ( .B1(n15961), .B2(n15956), .A(n15975), .ZN(n15974) );
  INV_X1 U19046 ( .A(n15957), .ZN(n15960) );
  INV_X1 U19047 ( .A(n15958), .ZN(n15959) );
  AOI222_X1 U19048 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n12122), .B1(n20126), 
        .B2(n15960), .C1(n20123), .C2(n15959), .ZN(n15963) );
  INV_X1 U19049 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15973) );
  NOR2_X1 U19050 ( .A1(n15961), .A2(n15979), .ZN(n15969) );
  OAI221_X1 U19051 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n12400), .C2(n15973), .A(
        n15969), .ZN(n15962) );
  OAI211_X1 U19052 ( .C1(n15974), .C2(n12400), .A(n15963), .B(n15962), .ZN(
        P1_U3023) );
  INV_X1 U19053 ( .A(n15983), .ZN(n15966) );
  AOI21_X1 U19054 ( .B1(n15966), .B2(n15965), .A(n15964), .ZN(n15968) );
  AOI22_X1 U19055 ( .A1(n12122), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n20126), 
        .B2(n10345), .ZN(n15972) );
  AOI22_X1 U19056 ( .A1(n15970), .A2(n20123), .B1(n15969), .B2(n15973), .ZN(
        n15971) );
  OAI211_X1 U19057 ( .C1(n15974), .C2(n15973), .A(n15972), .B(n15971), .ZN(
        P1_U3024) );
  AOI22_X1 U19058 ( .A1(n12122), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20126), 
        .B2(n19964), .ZN(n15978) );
  AOI22_X1 U19059 ( .A1(n15976), .A2(n20123), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15975), .ZN(n15977) );
  OAI211_X1 U19060 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15979), .A(
        n15978), .B(n15977), .ZN(P1_U3025) );
  NAND2_X1 U19061 ( .A1(n15981), .A2(n15980), .ZN(n15982) );
  AND2_X1 U19062 ( .A1(n15983), .A2(n15982), .ZN(n20023) );
  AOI22_X1 U19063 ( .A1(n12122), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n20126), 
        .B2(n20023), .ZN(n15987) );
  AOI22_X1 U19064 ( .A1(n15985), .A2(n20123), .B1(n20115), .B2(n15984), .ZN(
        n15986) );
  OAI211_X1 U19065 ( .C1(n15989), .C2(n15988), .A(n15987), .B(n15986), .ZN(
        P1_U3026) );
  INV_X1 U19066 ( .A(n19991), .ZN(n15993) );
  INV_X1 U19067 ( .A(n12428), .ZN(n15991) );
  NAND4_X1 U19068 ( .A1(n15993), .A2(n15992), .A3(n15991), .A4(n15990), .ZN(
        n15994) );
  OAI21_X1 U19069 ( .B1(n20809), .B2(n15995), .A(n15994), .ZN(P1_U3468) );
  NAND3_X1 U19070 ( .A1(n13230), .A2(n15996), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n15998) );
  NAND2_X1 U19071 ( .A1(n15998), .A2(n15997), .ZN(n20725) );
  AOI21_X1 U19072 ( .B1(n16004), .B2(n15999), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n16000) );
  AOI221_X1 U19073 ( .B1(n16002), .B2(n16001), .C1(n20725), .C2(n16001), .A(
        n16000), .ZN(P1_U3162) );
  OAI21_X1 U19074 ( .B1(n16004), .B2(n20551), .A(n16003), .ZN(P1_U3466) );
  INV_X1 U19075 ( .A(n16005), .ZN(n16008) );
  NAND3_X1 U19076 ( .A1(n19231), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n16006), 
        .ZN(n16007) );
  OAI21_X1 U19077 ( .B1(n16008), .B2(n19070), .A(n16007), .ZN(n16010) );
  INV_X1 U19078 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19836) );
  OAI22_X1 U19079 ( .A1(n11424), .A2(n19035), .B1(n19836), .B2(n19069), .ZN(
        n16009) );
  AOI211_X1 U19080 ( .C1(n19064), .C2(n19085), .A(n16010), .B(n16009), .ZN(
        n16014) );
  NAND4_X1 U19081 ( .A1(n19764), .A2(n16011), .A3(n16012), .A4(n9925), .ZN(
        n16013) );
  OAI211_X1 U19082 ( .C1(n11783), .C2(n19047), .A(n16014), .B(n16013), .ZN(
        P2_U2824) );
  AOI21_X1 U19083 ( .B1(n16015), .B2(n16016), .A(n16011), .ZN(n16022) );
  INV_X1 U19084 ( .A(n19070), .ZN(n18999) );
  AOI22_X1 U19085 ( .A1(n16017), .A2(n18999), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19080), .ZN(n16019) );
  AOI22_X1 U19086 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19063), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19049), .ZN(n16018) );
  OAI211_X1 U19087 ( .C1(n16020), .C2(n19053), .A(n16019), .B(n16018), .ZN(
        n16021) );
  AOI21_X1 U19088 ( .B1(n19764), .B2(n16022), .A(n16021), .ZN(n16023) );
  OAI21_X1 U19089 ( .B1(n16024), .B2(n19047), .A(n16023), .ZN(P2_U2826) );
  AOI211_X1 U19090 ( .C1(n16027), .C2(n16025), .A(n16026), .B(n19061), .ZN(
        n16033) );
  AOI22_X1 U19091 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19080), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19049), .ZN(n16030) );
  AOI22_X1 U19092 ( .A1(n16028), .A2(n18999), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n19063), .ZN(n16029) );
  OAI211_X1 U19093 ( .C1(n16031), .C2(n19047), .A(n16030), .B(n16029), .ZN(
        n16032) );
  AOI211_X1 U19094 ( .C1(n19064), .C2(n16034), .A(n16033), .B(n16032), .ZN(
        n16035) );
  INV_X1 U19095 ( .A(n16035), .ZN(P2_U2829) );
  AOI211_X1 U19096 ( .C1(n16037), .C2(n16036), .A(n9910), .B(n19061), .ZN(
        n16044) );
  INV_X1 U19097 ( .A(n16038), .ZN(n16039) );
  AOI22_X1 U19098 ( .A1(n16039), .A2(n18999), .B1(P2_REIP_REG_25__SCAN_IN), 
        .B2(n19049), .ZN(n16041) );
  AOI22_X1 U19099 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19063), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19080), .ZN(n16040) );
  OAI211_X1 U19100 ( .C1(n16042), .C2(n19053), .A(n16041), .B(n16040), .ZN(
        n16043) );
  AOI211_X1 U19101 ( .C1(n19062), .C2(n16045), .A(n16044), .B(n16043), .ZN(
        n16046) );
  INV_X1 U19102 ( .A(n16046), .ZN(P2_U2830) );
  OAI22_X1 U19103 ( .A1(n16047), .A2(n19070), .B1(n19820), .B2(n19069), .ZN(
        n16048) );
  INV_X1 U19104 ( .A(n16048), .ZN(n16058) );
  AOI22_X1 U19105 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19063), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19080), .ZN(n16057) );
  AOI22_X1 U19106 ( .A1(n16050), .A2(n19062), .B1(n16049), .B2(n19064), .ZN(
        n16056) );
  AOI21_X1 U19107 ( .B1(n16053), .B2(n16051), .A(n16052), .ZN(n16054) );
  NAND2_X1 U19108 ( .A1(n19764), .A2(n16054), .ZN(n16055) );
  NAND4_X1 U19109 ( .A1(n16058), .A2(n16057), .A3(n16056), .A4(n16055), .ZN(
        P2_U2831) );
  INV_X1 U19110 ( .A(n19220), .ZN(n16059) );
  AOI22_X1 U19111 ( .A1(n19088), .A2(n16059), .B1(n19125), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16065) );
  AOI22_X1 U19112 ( .A1(n19090), .A2(BUF2_REG_22__SCAN_IN), .B1(n19089), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16064) );
  INV_X1 U19113 ( .A(n16060), .ZN(n16062) );
  AOI22_X1 U19114 ( .A1(n16062), .A2(n19127), .B1(n19099), .B2(n16061), .ZN(
        n16063) );
  NAND3_X1 U19115 ( .A1(n16065), .A2(n16064), .A3(n16063), .ZN(P2_U2897) );
  AOI22_X1 U19116 ( .A1(n19088), .A2(n16066), .B1(n19125), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16070) );
  AOI22_X1 U19117 ( .A1(n19090), .A2(BUF2_REG_20__SCAN_IN), .B1(n19089), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16069) );
  AOI22_X1 U19118 ( .A1(n16067), .A2(n19127), .B1(n19099), .B2(n18855), .ZN(
        n16068) );
  NAND3_X1 U19119 ( .A1(n16070), .A2(n16069), .A3(n16068), .ZN(P2_U2899) );
  AOI22_X1 U19120 ( .A1(n19088), .A2(n16071), .B1(n19125), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16075) );
  AOI22_X1 U19121 ( .A1(n19090), .A2(BUF2_REG_18__SCAN_IN), .B1(n19089), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16074) );
  AOI22_X1 U19122 ( .A1(n16072), .A2(n19127), .B1(n19099), .B2(n18887), .ZN(
        n16073) );
  NAND3_X1 U19123 ( .A1(n16075), .A2(n16074), .A3(n16073), .ZN(P2_U2901) );
  AOI22_X1 U19124 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n16202), .ZN(n16083) );
  NAND2_X1 U19125 ( .A1(n16077), .A2(n16076), .ZN(n16078) );
  XNOR2_X1 U19126 ( .A(n16079), .B(n16078), .ZN(n16160) );
  AOI21_X1 U19127 ( .B1(n16155), .B2(n16080), .A(n16081), .ZN(n16159) );
  AOI222_X1 U19128 ( .A1(n16160), .A2(n19242), .B1(n19241), .B2(n16159), .C1(
        n9787), .C2(n16158), .ZN(n16082) );
  OAI211_X1 U19129 ( .C1(n19247), .C2(n18927), .A(n16083), .B(n16082), .ZN(
        P2_U3000) );
  AOI22_X1 U19130 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n16202), .B1(n16143), 
        .B2(n18941), .ZN(n16093) );
  INV_X1 U19131 ( .A(n16084), .ZN(n16085) );
  NOR2_X1 U19132 ( .A1(n16086), .A2(n16085), .ZN(n16087) );
  XNOR2_X1 U19133 ( .A(n15176), .B(n16087), .ZN(n16170) );
  INV_X1 U19134 ( .A(n16080), .ZN(n16088) );
  AOI21_X1 U19135 ( .B1(n15474), .B2(n16089), .A(n16088), .ZN(n16169) );
  AOI22_X1 U19136 ( .A1(n16170), .A2(n19242), .B1(n19241), .B2(n16169), .ZN(
        n16090) );
  INV_X1 U19137 ( .A(n16090), .ZN(n16091) );
  AOI21_X1 U19138 ( .B1(n9787), .B2(n18940), .A(n16091), .ZN(n16092) );
  OAI211_X1 U19139 ( .C1(n16150), .C2(n10216), .A(n16093), .B(n16092), .ZN(
        P2_U3001) );
  AOI22_X1 U19140 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19236), .ZN(n16100) );
  NAND2_X1 U19141 ( .A1(n16094), .A2(n19242), .ZN(n16096) );
  NAND2_X1 U19142 ( .A1(n18950), .A2(n9787), .ZN(n16095) );
  OAI211_X1 U19143 ( .C1(n16097), .C2(n16145), .A(n16096), .B(n16095), .ZN(
        n16098) );
  INV_X1 U19144 ( .A(n16098), .ZN(n16099) );
  OAI211_X1 U19145 ( .C1(n19247), .C2(n18945), .A(n16100), .B(n16099), .ZN(
        P2_U3002) );
  AOI22_X1 U19146 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n16202), .B1(n16143), 
        .B2(n18960), .ZN(n16105) );
  OAI22_X1 U19147 ( .A1(n16102), .A2(n16145), .B1(n16101), .B2(n12452), .ZN(
        n16103) );
  AOI21_X1 U19148 ( .B1(n9787), .B2(n18961), .A(n16103), .ZN(n16104) );
  OAI211_X1 U19149 ( .C1(n16150), .C2(n16106), .A(n16105), .B(n16104), .ZN(
        P2_U3003) );
  AOI22_X1 U19150 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n16202), .ZN(n16118) );
  AOI21_X1 U19151 ( .B1(n16109), .B2(n16108), .A(n16107), .ZN(n16184) );
  NOR2_X1 U19152 ( .A1(n16111), .A2(n16110), .ZN(n16115) );
  NAND2_X1 U19153 ( .A1(n16113), .A2(n16112), .ZN(n16114) );
  XNOR2_X1 U19154 ( .A(n16115), .B(n16114), .ZN(n16188) );
  OAI22_X1 U19155 ( .A1(n16188), .A2(n12452), .B1(n16130), .B2(n18970), .ZN(
        n16116) );
  AOI21_X1 U19156 ( .B1(n16184), .B2(n19241), .A(n16116), .ZN(n16117) );
  OAI211_X1 U19157 ( .C1(n19247), .C2(n18967), .A(n16118), .B(n16117), .ZN(
        P2_U3004) );
  AOI22_X1 U19158 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19236), .ZN(n16135) );
  OR2_X1 U19159 ( .A1(n16121), .A2(n16120), .ZN(n16122) );
  NAND2_X1 U19160 ( .A1(n16119), .A2(n16122), .ZN(n16200) );
  AOI21_X1 U19161 ( .B1(n15270), .B2(n16124), .A(n16123), .ZN(n16129) );
  INV_X1 U19162 ( .A(n16125), .ZN(n16127) );
  NOR2_X1 U19163 ( .A1(n16127), .A2(n16126), .ZN(n16128) );
  XNOR2_X1 U19164 ( .A(n16129), .B(n16128), .ZN(n16197) );
  NOR2_X1 U19165 ( .A1(n18995), .A2(n16130), .ZN(n16131) );
  AOI21_X1 U19166 ( .B1(n16197), .B2(n19242), .A(n16131), .ZN(n16132) );
  OAI21_X1 U19167 ( .B1(n16200), .B2(n16145), .A(n16132), .ZN(n16133) );
  INV_X1 U19168 ( .A(n16133), .ZN(n16134) );
  OAI211_X1 U19169 ( .C1(n19247), .C2(n18990), .A(n16135), .B(n16134), .ZN(
        P2_U3006) );
  AOI22_X1 U19170 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n16202), .ZN(n16142) );
  NAND2_X1 U19171 ( .A1(n19015), .A2(n9787), .ZN(n16138) );
  OR2_X1 U19172 ( .A1(n16136), .A2(n12452), .ZN(n16137) );
  OAI211_X1 U19173 ( .C1(n16139), .C2(n16145), .A(n16138), .B(n16137), .ZN(
        n16140) );
  INV_X1 U19174 ( .A(n16140), .ZN(n16141) );
  OAI211_X1 U19175 ( .C1(n19247), .C2(n19013), .A(n16142), .B(n16141), .ZN(
        P2_U3008) );
  AOI22_X1 U19176 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19236), .B1(n16143), 
        .B2(n19026), .ZN(n16149) );
  OAI22_X1 U19177 ( .A1(n16146), .A2(n12452), .B1(n16145), .B2(n16144), .ZN(
        n16147) );
  AOI21_X1 U19178 ( .B1(n9787), .B2(n19027), .A(n16147), .ZN(n16148) );
  OAI211_X1 U19179 ( .C1(n16150), .C2(n19019), .A(n16149), .B(n16148), .ZN(
        P2_U3009) );
  AOI21_X1 U19180 ( .B1(n16152), .B2(n16164), .A(n16151), .ZN(n19103) );
  NOR2_X1 U19181 ( .A1(n19034), .A2(n11341), .ZN(n16157) );
  NAND3_X1 U19182 ( .A1(n16154), .A2(n16153), .A3(n16089), .ZN(n16173) );
  AOI21_X1 U19183 ( .B1(n16167), .B2(n16173), .A(n16155), .ZN(n16156) );
  AOI211_X1 U19184 ( .C1(n16192), .C2(n19103), .A(n16157), .B(n16156), .ZN(
        n16162) );
  AOI222_X1 U19185 ( .A1(n16160), .A2(n16196), .B1(n16183), .B2(n16159), .C1(
        n16182), .C2(n16158), .ZN(n16161) );
  OAI211_X1 U19186 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16163), .A(
        n16162), .B(n16161), .ZN(P2_U3032) );
  OAI21_X1 U19187 ( .B1(n16166), .B2(n16165), .A(n16164), .ZN(n19107) );
  OAI22_X1 U19188 ( .A1(n16167), .A2(n16089), .B1(n19107), .B2(n16177), .ZN(
        n16168) );
  AOI21_X1 U19189 ( .B1(P2_REIP_REG_13__SCAN_IN), .B2(n19236), .A(n16168), 
        .ZN(n16172) );
  AOI222_X1 U19190 ( .A1(n16170), .A2(n16196), .B1(n16169), .B2(n16183), .C1(
        n16182), .C2(n18940), .ZN(n16171) );
  OAI211_X1 U19191 ( .C1(n11191), .C2(n16173), .A(n16172), .B(n16171), .ZN(
        P2_U3033) );
  INV_X1 U19192 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19798) );
  NOR2_X1 U19193 ( .A1(n19798), .A2(n19034), .ZN(n16179) );
  XNOR2_X1 U19194 ( .A(n16175), .B(n16174), .ZN(n19113) );
  OAI22_X1 U19195 ( .A1(n16177), .A2(n19113), .B1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16176), .ZN(n16178) );
  AOI211_X1 U19196 ( .C1(n16180), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16179), .B(n16178), .ZN(n16186) );
  INV_X1 U19197 ( .A(n18970), .ZN(n16181) );
  AOI22_X1 U19198 ( .A1(n16184), .A2(n16183), .B1(n16182), .B2(n16181), .ZN(
        n16185) );
  OAI211_X1 U19199 ( .C1(n16188), .C2(n16187), .A(n16186), .B(n16185), .ZN(
        P2_U3036) );
  INV_X1 U19200 ( .A(n16189), .ZN(n16193) );
  AOI21_X1 U19201 ( .B1(n16191), .B2(n15520), .A(n16190), .ZN(n19115) );
  AOI22_X1 U19202 ( .A1(n16193), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16192), .B2(n19115), .ZN(n16208) );
  NOR2_X1 U19203 ( .A1(n18995), .A2(n16194), .ZN(n16195) );
  AOI21_X1 U19204 ( .B1(n16197), .B2(n16196), .A(n16195), .ZN(n16198) );
  OAI21_X1 U19205 ( .B1(n16200), .B2(n16199), .A(n16198), .ZN(n16201) );
  INV_X1 U19206 ( .A(n16201), .ZN(n16207) );
  NAND2_X1 U19207 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n16202), .ZN(n16206) );
  OAI211_X1 U19208 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16204), .B(n16203), .ZN(n16205) );
  NAND4_X1 U19209 ( .A1(n16208), .A2(n16207), .A3(n16206), .A4(n16205), .ZN(
        P2_U3038) );
  INV_X1 U19210 ( .A(n16209), .ZN(n19311) );
  INV_X1 U19211 ( .A(n16210), .ZN(n16219) );
  MUX2_X1 U19212 ( .A(n16211), .B(n16219), .S(n16239), .Z(n16241) );
  AOI21_X1 U19213 ( .B1(n16214), .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n16212), .ZN(n16217) );
  INV_X1 U19214 ( .A(n16213), .ZN(n16216) );
  NAND2_X1 U19215 ( .A1(n16214), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n16215) );
  OAI211_X1 U19216 ( .C1(n16217), .C2(n16216), .A(n16239), .B(n16215), .ZN(
        n16218) );
  AOI21_X1 U19217 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16219), .A(
        n16218), .ZN(n16222) );
  INV_X1 U19218 ( .A(n16220), .ZN(n16221) );
  MUX2_X1 U19219 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16221), .S(
        n16239), .Z(n16238) );
  AOI222_X1 U19220 ( .A1(n16222), .A2(n16238), .B1(n16222), .B2(n19858), .C1(
        n16238), .C2(n19858), .ZN(n16223) );
  OAI21_X1 U19221 ( .B1(n19311), .B2(n16241), .A(n16223), .ZN(n16245) );
  INV_X1 U19222 ( .A(n16224), .ZN(n16225) );
  OAI22_X1 U19223 ( .A1(n16230), .A2(n16227), .B1(n16226), .B2(n16225), .ZN(
        n16228) );
  AOI21_X1 U19224 ( .B1(n16230), .B2(n16229), .A(n16228), .ZN(n19889) );
  AOI22_X1 U19225 ( .A1(n16234), .A2(n16233), .B1(n16232), .B2(n16231), .ZN(
        n16237) );
  OAI21_X1 U19226 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n16235), .ZN(n16236) );
  NAND3_X1 U19227 ( .A1(n19889), .A2(n16237), .A3(n16236), .ZN(n16244) );
  INV_X1 U19228 ( .A(n16238), .ZN(n16242) );
  OAI22_X1 U19229 ( .A1(n16242), .A2(n16241), .B1(n16240), .B2(n16239), .ZN(
        n16243) );
  AOI211_X1 U19230 ( .C1(n16246), .C2(n16245), .A(n16244), .B(n16243), .ZN(
        n16258) );
  AOI211_X1 U19231 ( .C1(n16259), .C2(n19890), .A(n16248), .B(n16247), .ZN(
        n16257) );
  INV_X1 U19232 ( .A(n19901), .ZN(n19899) );
  NAND3_X1 U19233 ( .A1(n11721), .A2(n19903), .A3(n16249), .ZN(n16251) );
  AND3_X1 U19234 ( .A1(n16251), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n16250), 
        .ZN(n16254) );
  AOI22_X1 U19235 ( .A1(n19899), .A2(n16254), .B1(n16253), .B2(n16252), .ZN(
        n16255) );
  OAI221_X1 U19236 ( .B1(n19904), .B2(n16258), .C1(n19904), .C2(n11393), .A(
        n16254), .ZN(n19766) );
  NAND2_X1 U19237 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19766), .ZN(n16260) );
  OAI21_X1 U19238 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16255), .A(n16260), 
        .ZN(n16256) );
  OAI211_X1 U19239 ( .C1(n16258), .C2(n19134), .A(n16257), .B(n16256), .ZN(
        P2_U3176) );
  AOI21_X1 U19240 ( .B1(n16260), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16259), 
        .ZN(n16261) );
  INV_X1 U19241 ( .A(n16261), .ZN(P2_U3593) );
  NOR2_X1 U19242 ( .A1(n17754), .A2(n16262), .ZN(n16271) );
  OAI21_X1 U19243 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17754), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16263) );
  OAI221_X1 U19244 ( .B1(n16265), .B2(n16264), .C1(n17754), .C2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n16263), .ZN(n16270) );
  OAI21_X1 U19245 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16265), .A(
        n16264), .ZN(n16268) );
  NAND2_X1 U19246 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17754), .ZN(
        n16266) );
  OAI22_X1 U19247 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17754), .B1(
        n16266), .B2(n16265), .ZN(n16267) );
  OAI21_X1 U19248 ( .B1(n16271), .B2(n16268), .A(n16267), .ZN(n16269) );
  OAI21_X1 U19249 ( .B1(n16271), .B2(n16270), .A(n16269), .ZN(n16307) );
  INV_X1 U19250 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16463) );
  INV_X1 U19251 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18753) );
  NOR2_X1 U19252 ( .A1(n9796), .A2(n18753), .ZN(n16305) );
  XNOR2_X1 U19253 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16274) );
  OAI22_X1 U19254 ( .A1(n16275), .A2(n16274), .B1(n16273), .B2(n16463), .ZN(
        n16276) );
  AOI211_X1 U19255 ( .C1(n17604), .C2(n10009), .A(n16305), .B(n16276), .ZN(
        n16281) );
  NAND2_X1 U19256 ( .A1(n16277), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16278) );
  INV_X1 U19257 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18778) );
  XOR2_X1 U19258 ( .A(n16278), .B(n18778), .Z(n16302) );
  NAND2_X1 U19259 ( .A1(n16282), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16279) );
  XOR2_X1 U19260 ( .A(n16279), .B(n18778), .Z(n16301) );
  AOI22_X1 U19261 ( .A1(n17834), .A2(n16302), .B1(n17715), .B2(n16301), .ZN(
        n16280) );
  OAI211_X1 U19262 ( .C1(n17733), .C2(n16307), .A(n16281), .B(n16280), .ZN(
        P3_U2799) );
  NOR2_X1 U19263 ( .A1(n16295), .A2(n17855), .ZN(n16322) );
  INV_X1 U19264 ( .A(n16322), .ZN(n16283) );
  AOI211_X1 U19265 ( .C1(n16284), .C2(n16283), .A(n16282), .B(n17759), .ZN(
        n16293) );
  INV_X1 U19266 ( .A(n16285), .ZN(n16438) );
  AOI21_X1 U19267 ( .B1(n10015), .B2(n16438), .A(n16286), .ZN(n16487) );
  OAI21_X1 U19268 ( .B1(n16287), .B2(n17604), .A(n16487), .ZN(n16288) );
  OAI211_X1 U19269 ( .C1(n16291), .C2(n16290), .A(n16289), .B(n16288), .ZN(
        n16292) );
  AOI211_X1 U19270 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16294), .A(
        n16293), .B(n16292), .ZN(n16298) );
  NOR2_X1 U19271 ( .A1(n17858), .A2(n16295), .ZN(n16323) );
  OAI211_X1 U19272 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16323), .A(
        n17834), .B(n16296), .ZN(n16297) );
  OAI211_X1 U19273 ( .C1(n16299), .C2(n17733), .A(n16298), .B(n16297), .ZN(
        P3_U2801) );
  OAI21_X1 U19274 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18110), .A(
        n16300), .ZN(n16306) );
  AOI22_X1 U19275 ( .A1(n18066), .A2(n16309), .B1(n16308), .B2(n18068), .ZN(
        n17966) );
  OR2_X1 U19276 ( .A1(n17620), .A2(n17967), .ZN(n16311) );
  NOR2_X1 U19277 ( .A1(n17620), .A2(n18125), .ZN(n16310) );
  AOI22_X1 U19278 ( .A1(n18635), .A2(n17956), .B1(n17957), .B2(n16310), .ZN(
        n17883) );
  OAI21_X1 U19279 ( .B1(n17966), .B2(n16311), .A(n17883), .ZN(n17931) );
  NAND2_X1 U19280 ( .A1(n16312), .A2(n17931), .ZN(n17907) );
  NOR2_X1 U19281 ( .A1(n18142), .A2(n17907), .ZN(n17869) );
  NOR2_X1 U19282 ( .A1(n17685), .A2(n17491), .ZN(n16313) );
  AOI22_X1 U19283 ( .A1(n16314), .A2(n17869), .B1(n16313), .B2(n18141), .ZN(
        n16329) );
  AOI21_X1 U19284 ( .B1(n17754), .B2(n17491), .A(n17490), .ZN(n17469) );
  NAND2_X1 U19285 ( .A1(n16316), .A2(n16315), .ZN(n17468) );
  NOR2_X1 U19286 ( .A1(n17469), .A2(n17468), .ZN(n17470) );
  OAI211_X1 U19287 ( .C1(n16318), .C2(n17491), .A(n18609), .B(n16317), .ZN(
        n16321) );
  INV_X1 U19288 ( .A(n16319), .ZN(n16320) );
  OAI211_X1 U19289 ( .C1(n17470), .C2(n16321), .A(n16320), .B(n18109), .ZN(
        n16325) );
  OAI22_X1 U19290 ( .A1(n16323), .A2(n18611), .B1(n16322), .B2(n18015), .ZN(
        n16324) );
  OAI21_X1 U19291 ( .B1(n16325), .B2(n16324), .A(n9796), .ZN(n16328) );
  AND2_X1 U19292 ( .A1(n17468), .A2(n18078), .ZN(n16326) );
  AOI22_X1 U19293 ( .A1(n17490), .A2(n16326), .B1(n9790), .B2(
        P3_REIP_REG_28__SCAN_IN), .ZN(n16327) );
  OAI221_X1 U19294 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n16329), 
        .C1(n17467), .C2(n16328), .A(n16327), .ZN(P3_U2834) );
  NOR3_X1 U19295 ( .A1(P3_BE_N_REG_3__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n16331) );
  NOR4_X1 U19296 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16330) );
  NAND4_X1 U19297 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16331), .A3(n16330), .A4(
        U215), .ZN(U213) );
  INV_X1 U19298 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19141) );
  INV_X2 U19299 ( .A(U214), .ZN(n16370) );
  NOR2_X1 U19300 ( .A1(n16370), .A2(n16332), .ZN(n16367) );
  OAI222_X1 U19301 ( .A1(U212), .A2(n19141), .B1(n16372), .B2(n20213), .C1(
        U214), .C2(n16405), .ZN(U216) );
  AOI222_X1 U19302 ( .A1(n16369), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16367), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16370), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n16333) );
  INV_X1 U19303 ( .A(n16333), .ZN(U217) );
  AOI22_X1 U19304 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16369), .ZN(n16334) );
  OAI21_X1 U19305 ( .B1(n20198), .B2(n16372), .A(n16334), .ZN(U218) );
  AOI22_X1 U19306 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16369), .ZN(n16335) );
  OAI21_X1 U19307 ( .B1(n20191), .B2(n16372), .A(n16335), .ZN(U219) );
  AOI22_X1 U19308 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16369), .ZN(n16336) );
  OAI21_X1 U19309 ( .B1(n20184), .B2(n16372), .A(n16336), .ZN(U220) );
  AOI22_X1 U19310 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16369), .ZN(n16337) );
  OAI21_X1 U19311 ( .B1(n20176), .B2(n16372), .A(n16337), .ZN(U221) );
  AOI222_X1 U19312 ( .A1(n16369), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(n16367), 
        .B2(BUF1_REG_25__SCAN_IN), .C1(n16370), .C2(P1_DATAO_REG_25__SCAN_IN), 
        .ZN(n16338) );
  INV_X1 U19313 ( .A(n16338), .ZN(U222) );
  AOI22_X1 U19314 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16369), .ZN(n16339) );
  OAI21_X1 U19315 ( .B1(n20149), .B2(n16372), .A(n16339), .ZN(U223) );
  AOI22_X1 U19316 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16369), .ZN(n16340) );
  OAI21_X1 U19317 ( .B1(n14562), .B2(n16372), .A(n16340), .ZN(U224) );
  INV_X1 U19318 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16396) );
  OAI222_X1 U19319 ( .A1(U212), .A2(n16396), .B1(n16372), .B2(n14567), .C1(
        U214), .C2(n16341), .ZN(U225) );
  AOI22_X1 U19320 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16369), .ZN(n16342) );
  OAI21_X1 U19321 ( .B1(n14571), .B2(n16372), .A(n16342), .ZN(U226) );
  AOI22_X1 U19322 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16369), .ZN(n16343) );
  OAI21_X1 U19323 ( .B1(n20189), .B2(n16372), .A(n16343), .ZN(U227) );
  AOI22_X1 U19324 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16369), .ZN(n16344) );
  OAI21_X1 U19325 ( .B1(n20181), .B2(n16372), .A(n16344), .ZN(U228) );
  AOI22_X1 U19326 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16369), .ZN(n16345) );
  OAI21_X1 U19327 ( .B1(n20173), .B2(n16372), .A(n16345), .ZN(U229) );
  AOI22_X1 U19328 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16369), .ZN(n16346) );
  OAI21_X1 U19329 ( .B1(n14584), .B2(n16372), .A(n16346), .ZN(U230) );
  AOI222_X1 U19330 ( .A1(n16370), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n16367), 
        .B2(BUF1_REG_16__SCAN_IN), .C1(n16369), .C2(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n16347) );
  INV_X1 U19331 ( .A(n16347), .ZN(U231) );
  AOI22_X1 U19332 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16369), .ZN(n16348) );
  OAI21_X1 U19333 ( .B1(n13379), .B2(n16372), .A(n16348), .ZN(U232) );
  AOI22_X1 U19334 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16369), .ZN(n16349) );
  OAI21_X1 U19335 ( .B1(n13909), .B2(n16372), .A(n16349), .ZN(U233) );
  AOI22_X1 U19336 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16369), .ZN(n16350) );
  OAI21_X1 U19337 ( .B1(n14535), .B2(n16372), .A(n16350), .ZN(U234) );
  AOI22_X1 U19338 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16369), .ZN(n16351) );
  OAI21_X1 U19339 ( .B1(n15039), .B2(n16372), .A(n16351), .ZN(U235) );
  AOI22_X1 U19340 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16369), .ZN(n16352) );
  OAI21_X1 U19341 ( .B1(n15048), .B2(n16372), .A(n16352), .ZN(U236) );
  AOI22_X1 U19342 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16369), .ZN(n16353) );
  OAI21_X1 U19343 ( .B1(n16354), .B2(n16372), .A(n16353), .ZN(U237) );
  AOI22_X1 U19344 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16369), .ZN(n16355) );
  OAI21_X1 U19345 ( .B1(n15070), .B2(n16372), .A(n16355), .ZN(U238) );
  AOI22_X1 U19346 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16369), .ZN(n16356) );
  OAI21_X1 U19347 ( .B1(n16357), .B2(n16372), .A(n16356), .ZN(U239) );
  AOI22_X1 U19348 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16369), .ZN(n16358) );
  OAI21_X1 U19349 ( .B1(n16359), .B2(n16372), .A(n16358), .ZN(U240) );
  AOI222_X1 U19350 ( .A1(n16369), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n16367), 
        .B2(BUF1_REG_6__SCAN_IN), .C1(n16370), .C2(P1_DATAO_REG_6__SCAN_IN), 
        .ZN(n16360) );
  INV_X1 U19351 ( .A(n16360), .ZN(U241) );
  INV_X1 U19352 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n20044) );
  AOI22_X1 U19353 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16367), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16369), .ZN(n16361) );
  OAI21_X1 U19354 ( .B1(n20044), .B2(U214), .A(n16361), .ZN(U242) );
  AOI22_X1 U19355 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16369), .ZN(n16362) );
  OAI21_X1 U19356 ( .B1(n16363), .B2(n16372), .A(n16362), .ZN(U243) );
  INV_X1 U19357 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16377) );
  AOI22_X1 U19358 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16367), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16370), .ZN(n16364) );
  OAI21_X1 U19359 ( .B1(n16377), .B2(U212), .A(n16364), .ZN(U244) );
  AOI22_X1 U19360 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16369), .ZN(n16365) );
  OAI21_X1 U19361 ( .B1(n16366), .B2(n16372), .A(n16365), .ZN(U245) );
  INV_X1 U19362 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16375) );
  AOI22_X1 U19363 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16367), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16370), .ZN(n16368) );
  OAI21_X1 U19364 ( .B1(n16375), .B2(U212), .A(n16368), .ZN(U246) );
  AOI22_X1 U19365 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16370), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16369), .ZN(n16371) );
  OAI21_X1 U19366 ( .B1(n16373), .B2(n16372), .A(n16371), .ZN(U247) );
  OAI22_X1 U19367 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16404), .ZN(n16374) );
  INV_X1 U19368 ( .A(n16374), .ZN(U251) );
  INV_X1 U19369 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18176) );
  AOI22_X1 U19370 ( .A1(n16404), .A2(n16375), .B1(n18176), .B2(U215), .ZN(U252) );
  OAI22_X1 U19371 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16390), .ZN(n16376) );
  INV_X1 U19372 ( .A(n16376), .ZN(U253) );
  INV_X1 U19373 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18184) );
  AOI22_X1 U19374 ( .A1(n16404), .A2(n16377), .B1(n18184), .B2(U215), .ZN(U254) );
  OAI22_X1 U19375 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16390), .ZN(n16378) );
  INV_X1 U19376 ( .A(n16378), .ZN(U255) );
  OAI22_X1 U19377 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16390), .ZN(n16379) );
  INV_X1 U19378 ( .A(n16379), .ZN(U256) );
  INV_X1 U19379 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16380) );
  INV_X1 U19380 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18198) );
  AOI22_X1 U19381 ( .A1(n16404), .A2(n16380), .B1(n18198), .B2(U215), .ZN(U257) );
  OAI22_X1 U19382 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16390), .ZN(n16381) );
  INV_X1 U19383 ( .A(n16381), .ZN(U258) );
  OAI22_X1 U19384 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16390), .ZN(n16382) );
  INV_X1 U19385 ( .A(n16382), .ZN(U259) );
  OAI22_X1 U19386 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16390), .ZN(n16383) );
  INV_X1 U19387 ( .A(n16383), .ZN(U260) );
  OAI22_X1 U19388 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16390), .ZN(n16384) );
  INV_X1 U19389 ( .A(n16384), .ZN(U261) );
  OAI22_X1 U19390 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16404), .ZN(n16385) );
  INV_X1 U19391 ( .A(n16385), .ZN(U262) );
  OAI22_X1 U19392 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16390), .ZN(n16386) );
  INV_X1 U19393 ( .A(n16386), .ZN(U263) );
  OAI22_X1 U19394 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16404), .ZN(n16387) );
  INV_X1 U19395 ( .A(n16387), .ZN(U264) );
  OAI22_X1 U19396 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16390), .ZN(n16388) );
  INV_X1 U19397 ( .A(n16388), .ZN(U265) );
  OAI22_X1 U19398 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16404), .ZN(n16389) );
  INV_X1 U19399 ( .A(n16389), .ZN(U266) );
  INV_X1 U19400 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n21146) );
  AOI22_X1 U19401 ( .A1(n16404), .A2(n21146), .B1(n18166), .B2(U215), .ZN(U267) );
  OAI22_X1 U19402 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16390), .ZN(n16391) );
  INV_X1 U19403 ( .A(n16391), .ZN(U268) );
  OAI22_X1 U19404 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16404), .ZN(n16392) );
  INV_X1 U19405 ( .A(n16392), .ZN(U269) );
  OAI22_X1 U19406 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16404), .ZN(n16393) );
  INV_X1 U19407 ( .A(n16393), .ZN(U270) );
  OAI22_X1 U19408 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16404), .ZN(n16394) );
  INV_X1 U19409 ( .A(n16394), .ZN(U271) );
  OAI22_X1 U19410 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16404), .ZN(n16395) );
  INV_X1 U19411 ( .A(n16395), .ZN(U272) );
  AOI22_X1 U19412 ( .A1(n16404), .A2(n16396), .B1(n18197), .B2(U215), .ZN(U273) );
  OAI22_X1 U19413 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16404), .ZN(n16397) );
  INV_X1 U19414 ( .A(n16397), .ZN(U274) );
  OAI22_X1 U19415 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16404), .ZN(n16398) );
  INV_X1 U19416 ( .A(n16398), .ZN(U275) );
  INV_X1 U19417 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n19152) );
  AOI22_X1 U19418 ( .A1(n16404), .A2(n19152), .B1(n18175), .B2(U215), .ZN(U276) );
  OAI22_X1 U19419 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16404), .ZN(n16399) );
  INV_X1 U19420 ( .A(n16399), .ZN(U277) );
  OAI22_X1 U19421 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16404), .ZN(n16400) );
  INV_X1 U19422 ( .A(n16400), .ZN(U278) );
  OAI22_X1 U19423 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16404), .ZN(n16401) );
  INV_X1 U19424 ( .A(n16401), .ZN(U279) );
  OAI22_X1 U19425 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16404), .ZN(n16402) );
  INV_X1 U19426 ( .A(n16402), .ZN(U280) );
  INV_X1 U19427 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n21031) );
  AOI22_X1 U19428 ( .A1(n16404), .A2(n21031), .B1(n14324), .B2(U215), .ZN(U281) );
  AOI22_X1 U19429 ( .A1(n16404), .A2(n19141), .B1(n16403), .B2(U215), .ZN(U282) );
  INV_X1 U19430 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17359) );
  AOI222_X1 U19431 ( .A1(n16405), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19141), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17359), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16406) );
  INV_X2 U19432 ( .A(n16408), .ZN(n16407) );
  INV_X1 U19433 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18717) );
  INV_X1 U19434 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19799) );
  AOI22_X1 U19435 ( .A1(n16407), .A2(n18717), .B1(n19799), .B2(n16408), .ZN(
        U347) );
  INV_X1 U19436 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18715) );
  INV_X1 U19437 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19797) );
  AOI22_X1 U19438 ( .A1(n16407), .A2(n18715), .B1(n19797), .B2(n16408), .ZN(
        U348) );
  INV_X1 U19439 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18714) );
  INV_X1 U19440 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19796) );
  AOI22_X1 U19441 ( .A1(n16407), .A2(n18714), .B1(n19796), .B2(n16408), .ZN(
        U349) );
  INV_X1 U19442 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18712) );
  INV_X1 U19443 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19795) );
  AOI22_X1 U19444 ( .A1(n16407), .A2(n18712), .B1(n19795), .B2(n16408), .ZN(
        U350) );
  INV_X1 U19445 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18710) );
  INV_X1 U19446 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19793) );
  AOI22_X1 U19447 ( .A1(n16407), .A2(n18710), .B1(n19793), .B2(n16408), .ZN(
        U351) );
  INV_X1 U19448 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18708) );
  INV_X1 U19449 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19792) );
  AOI22_X1 U19450 ( .A1(n16407), .A2(n18708), .B1(n19792), .B2(n16408), .ZN(
        U352) );
  INV_X1 U19451 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18706) );
  INV_X1 U19452 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19791) );
  AOI22_X1 U19453 ( .A1(n16407), .A2(n18706), .B1(n19791), .B2(n16408), .ZN(
        U353) );
  INV_X1 U19454 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18704) );
  AOI22_X1 U19455 ( .A1(n16407), .A2(n18704), .B1(n19790), .B2(n16408), .ZN(
        U354) );
  INV_X1 U19456 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18755) );
  INV_X1 U19457 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19835) );
  AOI22_X1 U19458 ( .A1(n16407), .A2(n18755), .B1(n19835), .B2(n16408), .ZN(
        U355) );
  INV_X1 U19459 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18751) );
  INV_X1 U19460 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19831) );
  AOI22_X1 U19461 ( .A1(n16407), .A2(n18751), .B1(n19831), .B2(n16408), .ZN(
        U356) );
  INV_X1 U19462 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n21151) );
  INV_X1 U19463 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19829) );
  AOI22_X1 U19464 ( .A1(n16407), .A2(n21151), .B1(n19829), .B2(n16408), .ZN(
        U357) );
  INV_X1 U19465 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18748) );
  INV_X1 U19466 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19826) );
  AOI22_X1 U19467 ( .A1(n16407), .A2(n18748), .B1(n19826), .B2(n16408), .ZN(
        U358) );
  INV_X1 U19468 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18747) );
  INV_X1 U19469 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19825) );
  AOI22_X1 U19470 ( .A1(n16407), .A2(n18747), .B1(n19825), .B2(n16408), .ZN(
        U359) );
  INV_X1 U19471 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18745) );
  INV_X1 U19472 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19823) );
  AOI22_X1 U19473 ( .A1(n16407), .A2(n18745), .B1(n19823), .B2(n16408), .ZN(
        U360) );
  INV_X1 U19474 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18742) );
  INV_X1 U19475 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19821) );
  AOI22_X1 U19476 ( .A1(n16407), .A2(n18742), .B1(n19821), .B2(n16408), .ZN(
        U361) );
  INV_X1 U19477 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18741) );
  INV_X1 U19478 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19819) );
  AOI22_X1 U19479 ( .A1(n16407), .A2(n18741), .B1(n19819), .B2(n16408), .ZN(
        U362) );
  INV_X1 U19480 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18740) );
  INV_X1 U19481 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19817) );
  AOI22_X1 U19482 ( .A1(n16407), .A2(n18740), .B1(n19817), .B2(n16408), .ZN(
        U363) );
  INV_X1 U19483 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18738) );
  INV_X1 U19484 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19815) );
  AOI22_X1 U19485 ( .A1(n16407), .A2(n18738), .B1(n19815), .B2(n16408), .ZN(
        U364) );
  INV_X1 U19486 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18702) );
  INV_X1 U19487 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U19488 ( .A1(n16407), .A2(n18702), .B1(n19788), .B2(n16408), .ZN(
        U365) );
  INV_X1 U19489 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18735) );
  INV_X1 U19490 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19813) );
  AOI22_X1 U19491 ( .A1(n16407), .A2(n18735), .B1(n19813), .B2(n16408), .ZN(
        U366) );
  INV_X1 U19492 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18734) );
  INV_X1 U19493 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19812) );
  AOI22_X1 U19494 ( .A1(n16407), .A2(n18734), .B1(n19812), .B2(n16408), .ZN(
        U367) );
  INV_X1 U19495 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18732) );
  INV_X1 U19496 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19810) );
  AOI22_X1 U19497 ( .A1(n16407), .A2(n18732), .B1(n19810), .B2(n16408), .ZN(
        U368) );
  INV_X1 U19498 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18730) );
  INV_X1 U19499 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n21075) );
  AOI22_X1 U19500 ( .A1(n16407), .A2(n18730), .B1(n21075), .B2(n16408), .ZN(
        U369) );
  INV_X1 U19501 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18729) );
  INV_X1 U19502 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19807) );
  AOI22_X1 U19503 ( .A1(n16407), .A2(n18729), .B1(n19807), .B2(n16408), .ZN(
        U370) );
  INV_X1 U19504 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18727) );
  INV_X1 U19505 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19806) );
  AOI22_X1 U19506 ( .A1(n16407), .A2(n18727), .B1(n19806), .B2(n16408), .ZN(
        U371) );
  INV_X1 U19507 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18724) );
  INV_X1 U19508 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19804) );
  AOI22_X1 U19509 ( .A1(n16407), .A2(n18724), .B1(n19804), .B2(n16408), .ZN(
        U372) );
  INV_X1 U19510 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18723) );
  INV_X1 U19511 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19803) );
  AOI22_X1 U19512 ( .A1(n16407), .A2(n18723), .B1(n19803), .B2(n16408), .ZN(
        U373) );
  INV_X1 U19513 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18720) );
  INV_X1 U19514 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19802) );
  AOI22_X1 U19515 ( .A1(n16407), .A2(n18720), .B1(n19802), .B2(n16408), .ZN(
        U374) );
  INV_X1 U19516 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18719) );
  INV_X1 U19517 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19801) );
  AOI22_X1 U19518 ( .A1(n16407), .A2(n18719), .B1(n19801), .B2(n16408), .ZN(
        U375) );
  INV_X1 U19519 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18700) );
  INV_X1 U19520 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19787) );
  AOI22_X1 U19521 ( .A1(n16407), .A2(n18700), .B1(n19787), .B2(n16408), .ZN(
        U376) );
  INV_X1 U19522 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18699) );
  NAND2_X1 U19523 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18699), .ZN(n18688) );
  NOR2_X1 U19524 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n18685) );
  INV_X1 U19525 ( .A(n18685), .ZN(n16409) );
  OAI21_X1 U19526 ( .B1(n18688), .B2(n16410), .A(n16409), .ZN(n18767) );
  AOI21_X1 U19527 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18767), .ZN(n16411) );
  INV_X1 U19528 ( .A(n16411), .ZN(P3_U2633) );
  NAND2_X1 U19529 ( .A1(n18779), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n16456) );
  INV_X1 U19530 ( .A(n17416), .ZN(n17418) );
  OAI21_X1 U19531 ( .B1(n16417), .B2(n17418), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16412) );
  OAI21_X1 U19532 ( .B1(n16456), .B2(n16413), .A(n16412), .ZN(P3_U2634) );
  AOI22_X1 U19533 ( .A1(n18685), .A2(n18699), .B1(P3_D_C_N_REG_SCAN_IN), .B2(
        n18822), .ZN(n16414) );
  OAI21_X1 U19534 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n18822), .A(n16414), 
        .ZN(P3_U2635) );
  OAI21_X1 U19535 ( .B1(n16415), .B2(BS16), .A(n18767), .ZN(n18765) );
  OAI21_X1 U19536 ( .B1(n18767), .B2(n18812), .A(n18765), .ZN(P3_U2636) );
  NOR3_X1 U19537 ( .A1(n16417), .A2(n16416), .A3(n18607), .ZN(n18614) );
  NOR2_X1 U19538 ( .A1(n18614), .A2(n18669), .ZN(n18806) );
  OAI21_X1 U19539 ( .B1(n18806), .B2(n16419), .A(n16418), .ZN(P3_U2637) );
  NOR4_X1 U19540 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16423) );
  NOR4_X1 U19541 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16422) );
  NOR4_X1 U19542 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16421) );
  NOR4_X1 U19543 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16420) );
  NAND4_X1 U19544 ( .A1(n16423), .A2(n16422), .A3(n16421), .A4(n16420), .ZN(
        n16429) );
  NOR4_X1 U19545 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16427) );
  AOI211_X1 U19546 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_10__SCAN_IN), .B(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16426) );
  NOR4_X1 U19547 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16425) );
  NOR4_X1 U19548 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16424) );
  NAND4_X1 U19549 ( .A1(n16427), .A2(n16426), .A3(n16425), .A4(n16424), .ZN(
        n16428) );
  NOR2_X1 U19550 ( .A1(n16429), .A2(n16428), .ZN(n18804) );
  INV_X1 U19551 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16431) );
  NOR3_X1 U19552 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16432) );
  OAI21_X1 U19553 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16432), .A(n18804), .ZN(
        n16430) );
  OAI21_X1 U19554 ( .B1(n18804), .B2(n16431), .A(n16430), .ZN(P3_U2638) );
  INV_X1 U19555 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18798) );
  INV_X1 U19556 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18766) );
  AOI21_X1 U19557 ( .B1(n18798), .B2(n18766), .A(n16432), .ZN(n16433) );
  INV_X1 U19558 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18758) );
  INV_X1 U19559 ( .A(n18804), .ZN(n18800) );
  AOI22_X1 U19560 ( .A1(n18804), .A2(n16433), .B1(n18758), .B2(n18800), .ZN(
        P3_U2639) );
  INV_X1 U19561 ( .A(n16434), .ZN(n16435) );
  NAND2_X1 U19562 ( .A1(n16436), .A2(n16435), .ZN(n18606) );
  NAND2_X1 U19563 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16819), .ZN(n16437) );
  AOI211_X4 U19564 ( .C1(n18812), .C2(n18814), .A(n16459), .B(n16437), .ZN(
        n16775) );
  INV_X1 U19565 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16944) );
  NOR3_X1 U19566 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16786) );
  NAND2_X1 U19567 ( .A1(n16786), .A2(n17195), .ZN(n16774) );
  NOR2_X1 U19568 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16774), .ZN(n16758) );
  INV_X1 U19569 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17183) );
  NAND2_X1 U19570 ( .A1(n16758), .A2(n17183), .ZN(n16751) );
  INV_X1 U19571 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17174) );
  NAND2_X1 U19572 ( .A1(n16733), .A2(n17174), .ZN(n16730) );
  INV_X1 U19573 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16707) );
  NAND2_X1 U19574 ( .A1(n16717), .A2(n16707), .ZN(n16704) );
  INV_X1 U19575 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16688) );
  NAND2_X1 U19576 ( .A1(n16691), .A2(n16688), .ZN(n16685) );
  INV_X1 U19577 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16656) );
  NAND2_X1 U19578 ( .A1(n16671), .A2(n16656), .ZN(n16655) );
  INV_X1 U19579 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16637) );
  NAND2_X1 U19580 ( .A1(n16641), .A2(n16637), .ZN(n16634) );
  INV_X1 U19581 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16617) );
  NAND2_X1 U19582 ( .A1(n16620), .A2(n16617), .ZN(n16616) );
  INV_X1 U19583 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16593) );
  NAND2_X1 U19584 ( .A1(n16602), .A2(n16593), .ZN(n16592) );
  INV_X1 U19585 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n21069) );
  NAND2_X1 U19586 ( .A1(n16576), .A2(n21069), .ZN(n16570) );
  NOR2_X1 U19587 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16570), .ZN(n16559) );
  INV_X1 U19588 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16933) );
  NAND2_X1 U19589 ( .A1(n16559), .A2(n16933), .ZN(n16551) );
  NOR2_X1 U19590 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16551), .ZN(n16536) );
  INV_X1 U19591 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16532) );
  NAND2_X1 U19592 ( .A1(n16536), .A2(n16532), .ZN(n16531) );
  NOR2_X1 U19593 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16531), .ZN(n16513) );
  INV_X1 U19594 ( .A(n16513), .ZN(n16505) );
  NOR2_X1 U19595 ( .A1(n16505), .A2(P3_EBX_REG_27__SCAN_IN), .ZN(n16504) );
  NAND2_X1 U19596 ( .A1(n16944), .A2(n16504), .ZN(n16499) );
  OR2_X1 U19597 ( .A1(n16499), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n16475) );
  NOR2_X1 U19598 ( .A1(n16809), .A2(n16475), .ZN(n16478) );
  INV_X1 U19599 ( .A(n16478), .ZN(n16472) );
  AOI211_X1 U19600 ( .C1(n18811), .C2(n18813), .A(n18693), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16458) );
  AOI211_X4 U19601 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16819), .A(n16458), .B(
        n16459), .ZN(n16767) );
  INV_X1 U19602 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17494) );
  NOR2_X1 U19603 ( .A1(n17841), .A2(n17517), .ZN(n16451) );
  INV_X1 U19604 ( .A(n16451), .ZN(n16450) );
  NOR2_X1 U19605 ( .A1(n17520), .A2(n16450), .ZN(n17475) );
  NAND2_X1 U19606 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17475), .ZN(
        n16454) );
  NOR2_X1 U19607 ( .A1(n17494), .A2(n16454), .ZN(n16439) );
  OAI21_X1 U19608 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16439), .A(
        n16438), .ZN(n17474) );
  INV_X1 U19609 ( .A(n17474), .ZN(n16496) );
  AOI21_X1 U19610 ( .B1(n17494), .B2(n16454), .A(n16439), .ZN(n17488) );
  INV_X1 U19611 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17522) );
  NAND2_X1 U19612 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16451), .ZN(
        n16440) );
  AOI21_X1 U19613 ( .B1(n17522), .B2(n16440), .A(n17475), .ZN(n17530) );
  INV_X1 U19614 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17519) );
  NAND2_X1 U19615 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9893), .ZN(
        n16446) );
  INV_X1 U19616 ( .A(n16446), .ZN(n16447) );
  NAND2_X1 U19617 ( .A1(n17567), .A2(n16447), .ZN(n17516) );
  AOI21_X1 U19618 ( .B1(n17519), .B2(n17516), .A(n16451), .ZN(n17548) );
  NOR2_X1 U19619 ( .A1(n17577), .A2(n16446), .ZN(n16441) );
  OAI21_X1 U19620 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16441), .A(
        n17516), .ZN(n17565) );
  INV_X1 U19621 ( .A(n17565), .ZN(n16558) );
  INV_X1 U19622 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n21027) );
  INV_X1 U19623 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17601) );
  NAND2_X1 U19624 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17599), .ZN(
        n17598) );
  NOR3_X1 U19625 ( .A1(n21027), .A2(n17601), .A3(n17598), .ZN(n16444) );
  INV_X1 U19626 ( .A(n16444), .ZN(n17563) );
  AOI21_X1 U19627 ( .B1(n17588), .B2(n17563), .A(n16447), .ZN(n17592) );
  INV_X1 U19628 ( .A(n17598), .ZN(n16443) );
  OAI22_X1 U19629 ( .A1(n21027), .A2(n17598), .B1(n16443), .B2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17612) );
  INV_X1 U19630 ( .A(n17612), .ZN(n16601) );
  NOR2_X1 U19631 ( .A1(n17841), .A2(n9891), .ZN(n17639) );
  NAND3_X1 U19632 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(n17639), .ZN(n16621) );
  AOI21_X1 U19633 ( .B1(n21007), .B2(n16621), .A(n16443), .ZN(n17627) );
  INV_X1 U19634 ( .A(n17624), .ZN(n16442) );
  NOR3_X1 U19635 ( .A1(n17841), .A2(n17781), .A3(n17775), .ZN(n16679) );
  NAND2_X1 U19636 ( .A1(n17677), .A2(n16679), .ZN(n17674) );
  NOR2_X1 U19637 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17674), .ZN(
        n16665) );
  NAND2_X1 U19638 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16443), .ZN(
        n16445) );
  AOI21_X1 U19639 ( .B1(n17601), .B2(n16445), .A(n16444), .ZN(n17603) );
  NOR2_X1 U19640 ( .A1(n17592), .A2(n16580), .ZN(n16579) );
  NOR2_X1 U19641 ( .A1(n16579), .A2(n9890), .ZN(n16569) );
  AOI22_X1 U19642 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16447), .B1(
        n16446), .B2(n17577), .ZN(n17574) );
  NAND2_X1 U19643 ( .A1(n16449), .A2(n16448), .ZN(n16567) );
  NOR2_X1 U19644 ( .A1(n16556), .A2(n9890), .ZN(n16547) );
  NOR2_X1 U19645 ( .A1(n17548), .A2(n16547), .ZN(n16546) );
  NOR2_X1 U19646 ( .A1(n16546), .A2(n9890), .ZN(n16541) );
  INV_X1 U19647 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17538) );
  AOI22_X1 U19648 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16451), .B1(
        n16450), .B2(n17538), .ZN(n17535) );
  NOR2_X1 U19649 ( .A1(n17530), .A2(n16526), .ZN(n16525) );
  OR2_X1 U19650 ( .A1(n16525), .A2(n9890), .ZN(n16515) );
  OAI21_X1 U19651 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17475), .A(
        n16454), .ZN(n16455) );
  INV_X1 U19652 ( .A(n16455), .ZN(n17503) );
  NAND2_X1 U19653 ( .A1(n16515), .A2(n16455), .ZN(n16516) );
  NOR2_X1 U19654 ( .A1(n16506), .A2(n9890), .ZN(n16495) );
  NOR2_X1 U19655 ( .A1(n16496), .A2(n16495), .ZN(n16494) );
  NOR2_X1 U19656 ( .A1(n16494), .A2(n9890), .ZN(n16486) );
  NOR3_X1 U19657 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18682) );
  NAND2_X1 U19658 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18682), .ZN(n18679) );
  INV_X1 U19659 ( .A(n18679), .ZN(n16737) );
  NAND2_X1 U19660 ( .A1(n10009), .A2(n16737), .ZN(n16799) );
  NAND2_X1 U19661 ( .A1(n18661), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18674) );
  INV_X1 U19662 ( .A(n18674), .ZN(n18509) );
  INV_X1 U19663 ( .A(n16456), .ZN(n18675) );
  AOI211_X1 U19664 ( .C1(n18509), .C2(n18675), .A(n9790), .B(n16737), .ZN(
        n16457) );
  INV_X1 U19665 ( .A(n16458), .ZN(n18664) );
  INV_X1 U19666 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18721) );
  INV_X1 U19667 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18716) );
  INV_X1 U19668 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18713) );
  INV_X1 U19669 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18709) );
  INV_X1 U19670 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18705) );
  NAND3_X1 U19671 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16755) );
  NOR2_X1 U19672 ( .A1(n18705), .A2(n16755), .ZN(n16745) );
  NAND2_X1 U19673 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16745), .ZN(n16742) );
  NOR2_X1 U19674 ( .A1(n18709), .A2(n16742), .ZN(n16725) );
  NAND2_X1 U19675 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16725), .ZN(n16716) );
  NOR2_X1 U19676 ( .A1(n18713), .A2(n16716), .ZN(n16690) );
  NAND2_X1 U19677 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16690), .ZN(n16697) );
  NOR2_X1 U19678 ( .A1(n18716), .A2(n16697), .ZN(n16678) );
  NAND2_X1 U19679 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16678), .ZN(n16673) );
  NOR2_X1 U19680 ( .A1(n18721), .A2(n16673), .ZN(n16466) );
  NAND2_X1 U19681 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16460) );
  NAND4_X1 U19682 ( .A1(n16639), .A2(P3_REIP_REG_17__SCAN_IN), .A3(
        P3_REIP_REG_16__SCAN_IN), .A4(P3_REIP_REG_15__SCAN_IN), .ZN(n16607) );
  NAND2_X1 U19683 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n16461) );
  NAND3_X1 U19684 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(P3_REIP_REG_21__SCAN_IN), .ZN(n16468) );
  NAND2_X1 U19685 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16543), .ZN(n16535) );
  NAND2_X1 U19686 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n16469) );
  NAND4_X1 U19687 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16498), .ZN(n16465) );
  NAND2_X1 U19688 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18753), .ZN(n16462) );
  OAI22_X1 U19689 ( .A1(n16463), .A2(n16798), .B1(n16465), .B2(n16462), .ZN(
        n16464) );
  INV_X1 U19690 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18750) );
  NAND2_X1 U19691 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16483) );
  NOR2_X1 U19692 ( .A1(n18750), .A2(n16483), .ZN(n16470) );
  NAND3_X1 U19693 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16467) );
  NAND4_X1 U19694 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16466), .A3(
        P3_REIP_REG_13__SCAN_IN), .A4(n16800), .ZN(n16644) );
  NOR2_X1 U19695 ( .A1(n16467), .A2(n16644), .ZN(n16597) );
  NAND4_X1 U19696 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(P3_REIP_REG_19__SCAN_IN), .A4(n16597), .ZN(n16555) );
  NOR2_X1 U19697 ( .A1(n16468), .A2(n16555), .ZN(n16538) );
  NAND2_X1 U19698 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16538), .ZN(n16527) );
  NOR2_X1 U19699 ( .A1(n16469), .A2(n16527), .ZN(n16493) );
  NAND2_X1 U19700 ( .A1(n16756), .A2(n16800), .ZN(n16815) );
  AOI21_X1 U19701 ( .B1(n16470), .B2(n16493), .A(n16598), .ZN(n16482) );
  OAI21_X1 U19702 ( .B1(n16477), .B2(n16482), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16471) );
  XNOR2_X1 U19703 ( .A(n16474), .B(n16473), .ZN(n16481) );
  NAND2_X1 U19704 ( .A1(n16775), .A2(n16475), .ZN(n16484) );
  OAI22_X1 U19705 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16484), .B1(n21077), 
        .B2(n16798), .ZN(n16476) );
  AOI211_X1 U19706 ( .C1(P3_REIP_REG_30__SCAN_IN), .C2(n16482), .A(n16477), 
        .B(n16476), .ZN(n16480) );
  OAI21_X1 U19707 ( .B1(n16767), .B2(n16478), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16479) );
  OAI211_X1 U19708 ( .C1(n18679), .C2(n16481), .A(n16480), .B(n16479), .ZN(
        P3_U2641) );
  AOI22_X1 U19709 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16482), .B1(n16767), 
        .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n16492) );
  NOR2_X1 U19710 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16483), .ZN(n16490) );
  AOI21_X1 U19711 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16499), .A(n16484), .ZN(
        n16489) );
  AOI211_X1 U19712 ( .C1(n16487), .C2(n16486), .A(n16485), .B(n18679), .ZN(
        n16488) );
  OAI211_X1 U19713 ( .C1(n10015), .C2(n16798), .A(n16492), .B(n16491), .ZN(
        P3_U2642) );
  AOI22_X1 U19714 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16796), .B1(
        n16767), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16503) );
  NOR2_X1 U19715 ( .A1(n16598), .A2(n16493), .ZN(n16521) );
  INV_X1 U19716 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n21068) );
  AND2_X1 U19717 ( .A1(n21068), .A2(n16498), .ZN(n16510) );
  AOI211_X1 U19718 ( .C1(n16496), .C2(n16495), .A(n16494), .B(n18679), .ZN(
        n16497) );
  AOI221_X1 U19719 ( .B1(n16521), .B2(P3_REIP_REG_28__SCAN_IN), .C1(n16510), 
        .C2(P3_REIP_REG_28__SCAN_IN), .A(n16497), .ZN(n16502) );
  INV_X1 U19720 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18749) );
  NAND3_X1 U19721 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16498), .A3(n18749), 
        .ZN(n16501) );
  OAI211_X1 U19722 ( .C1(n16504), .C2(n16944), .A(n16775), .B(n16499), .ZN(
        n16500) );
  NAND4_X1 U19723 ( .A1(n16503), .A2(n16502), .A3(n16501), .A4(n16500), .ZN(
        P3_U2643) );
  AOI22_X1 U19724 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16521), .B1(n16767), 
        .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n16512) );
  AOI211_X1 U19725 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16505), .A(n16504), .B(
        n16809), .ZN(n16509) );
  AOI211_X1 U19726 ( .C1(n17488), .C2(n16507), .A(n16506), .B(n18679), .ZN(
        n16508) );
  NOR3_X1 U19727 ( .A1(n16510), .A2(n16509), .A3(n16508), .ZN(n16511) );
  OAI211_X1 U19728 ( .C1(n17494), .C2(n16798), .A(n16512), .B(n16511), .ZN(
        P3_U2644) );
  INV_X1 U19729 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16524) );
  AOI211_X1 U19730 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16531), .A(n16513), .B(
        n16809), .ZN(n16514) );
  AOI21_X1 U19731 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n16767), .A(n16514), .ZN(
        n16523) );
  INV_X1 U19732 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18744) );
  NOR3_X1 U19733 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16535), .A3(n18744), 
        .ZN(n16520) );
  INV_X1 U19734 ( .A(n16515), .ZN(n16518) );
  INV_X1 U19735 ( .A(n16516), .ZN(n16517) );
  AOI211_X1 U19736 ( .C1(n17503), .C2(n16518), .A(n16517), .B(n18679), .ZN(
        n16519) );
  AOI211_X1 U19737 ( .C1(n16521), .C2(P3_REIP_REG_26__SCAN_IN), .A(n16520), 
        .B(n16519), .ZN(n16522) );
  OAI211_X1 U19738 ( .C1(n16524), .C2(n16798), .A(n16523), .B(n16522), .ZN(
        P3_U2645) );
  AOI211_X1 U19739 ( .C1(n17530), .C2(n16526), .A(n16525), .B(n18679), .ZN(
        n16530) );
  NAND2_X1 U19740 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16527), .ZN(n16528) );
  OAI22_X1 U19741 ( .A1(n16598), .A2(n16528), .B1(n17522), .B2(n16798), .ZN(
        n16529) );
  AOI211_X1 U19742 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n16767), .A(n16530), .B(
        n16529), .ZN(n16534) );
  OAI211_X1 U19743 ( .C1(n16536), .C2(n16532), .A(n16775), .B(n16531), .ZN(
        n16533) );
  OAI211_X1 U19744 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16535), .A(n16534), 
        .B(n16533), .ZN(P3_U2646) );
  AOI211_X1 U19745 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16551), .A(n16536), .B(
        n16809), .ZN(n16537) );
  AOI21_X1 U19746 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16767), .A(n16537), .ZN(
        n16545) );
  NOR2_X1 U19747 ( .A1(n16598), .A2(n16538), .ZN(n16550) );
  INV_X1 U19748 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18743) );
  INV_X1 U19749 ( .A(n16539), .ZN(n16540) );
  AOI211_X1 U19750 ( .C1(n17535), .C2(n16541), .A(n16540), .B(n18679), .ZN(
        n16542) );
  AOI221_X1 U19751 ( .B1(n16550), .B2(P3_REIP_REG_24__SCAN_IN), .C1(n16543), 
        .C2(n18743), .A(n16542), .ZN(n16544) );
  OAI211_X1 U19752 ( .C1(n17538), .C2(n16798), .A(n16545), .B(n16544), .ZN(
        P3_U2647) );
  AOI22_X1 U19753 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16796), .B1(
        n16767), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n16554) );
  NAND2_X1 U19754 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16563) );
  NOR2_X1 U19755 ( .A1(n16575), .A2(n16563), .ZN(n16549) );
  INV_X1 U19756 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n21127) );
  AOI211_X1 U19757 ( .C1(n17548), .C2(n16547), .A(n16546), .B(n18679), .ZN(
        n16548) );
  AOI221_X1 U19758 ( .B1(n16550), .B2(P3_REIP_REG_23__SCAN_IN), .C1(n16549), 
        .C2(n21127), .A(n16548), .ZN(n16553) );
  OAI211_X1 U19759 ( .C1(n16559), .C2(n16933), .A(n16775), .B(n16551), .ZN(
        n16552) );
  NAND3_X1 U19760 ( .A1(n16554), .A2(n16553), .A3(n16552), .ZN(P3_U2648) );
  INV_X1 U19761 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18739) );
  NAND2_X1 U19762 ( .A1(n16815), .A2(n16555), .ZN(n16578) );
  AOI211_X1 U19763 ( .C1(n16558), .C2(n16557), .A(n16556), .B(n18679), .ZN(
        n16562) );
  AOI211_X1 U19764 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16570), .A(n16559), .B(
        n16809), .ZN(n16561) );
  OAI22_X1 U19765 ( .A1(n20966), .A2(n16798), .B1(n16810), .B2(n10110), .ZN(
        n16560) );
  NOR3_X1 U19766 ( .A1(n16562), .A2(n16561), .A3(n16560), .ZN(n16566) );
  INV_X1 U19767 ( .A(n16575), .ZN(n16564) );
  OAI211_X1 U19768 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16564), .B(n16563), .ZN(n16565) );
  OAI211_X1 U19769 ( .C1(n18739), .C2(n16578), .A(n16566), .B(n16565), .ZN(
        P3_U2649) );
  INV_X1 U19770 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18737) );
  INV_X1 U19771 ( .A(n16567), .ZN(n16568) );
  AOI211_X1 U19772 ( .C1(n17574), .C2(n16569), .A(n16568), .B(n18679), .ZN(
        n16573) );
  OAI211_X1 U19773 ( .C1(n16576), .C2(n21069), .A(n16775), .B(n16570), .ZN(
        n16571) );
  OAI21_X1 U19774 ( .B1(n21069), .B2(n16810), .A(n16571), .ZN(n16572) );
  AOI211_X1 U19775 ( .C1(n16796), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16573), .B(n16572), .ZN(n16574) );
  OAI221_X1 U19776 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16575), .C1(n18737), 
        .C2(n16578), .A(n16574), .ZN(P3_U2650) );
  AOI211_X1 U19777 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16592), .A(n16576), .B(
        n16809), .ZN(n16577) );
  AOI21_X1 U19778 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16767), .A(n16577), .ZN(
        n16585) );
  INV_X1 U19779 ( .A(n16578), .ZN(n16583) );
  INV_X1 U19780 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18736) );
  AOI211_X1 U19781 ( .C1(n17592), .C2(n16580), .A(n16579), .B(n18679), .ZN(
        n16581) );
  AOI221_X1 U19782 ( .B1(n16583), .B2(P3_REIP_REG_20__SCAN_IN), .C1(n16582), 
        .C2(n18736), .A(n16581), .ZN(n16584) );
  OAI211_X1 U19783 ( .C1(n17588), .C2(n16798), .A(n16585), .B(n16584), .ZN(
        P3_U2651) );
  AOI22_X1 U19784 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16796), .B1(
        n16767), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16596) );
  OAI22_X1 U19785 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16607), .B1(n16598), 
        .B2(n16597), .ZN(n16591) );
  INV_X1 U19786 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21167) );
  NOR3_X1 U19787 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n21167), .A3(n16607), 
        .ZN(n16590) );
  INV_X1 U19788 ( .A(n16586), .ZN(n16587) );
  AOI211_X1 U19789 ( .C1(n17603), .C2(n16588), .A(n16587), .B(n18679), .ZN(
        n16589) );
  AOI211_X1 U19790 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n16591), .A(n16590), 
        .B(n16589), .ZN(n16595) );
  OAI211_X1 U19791 ( .C1(n16602), .C2(n16593), .A(n16775), .B(n16592), .ZN(
        n16594) );
  NAND4_X1 U19792 ( .A1(n16596), .A2(n16595), .A3(n9796), .A4(n16594), .ZN(
        P3_U2652) );
  OR2_X1 U19793 ( .A1(n16598), .A2(n16597), .ZN(n16610) );
  AOI211_X1 U19794 ( .C1(n16601), .C2(n16600), .A(n16599), .B(n18679), .ZN(
        n16605) );
  AOI211_X1 U19795 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16616), .A(n16602), .B(
        n16809), .ZN(n16604) );
  INV_X1 U19796 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16821) );
  OAI22_X1 U19797 ( .A1(n21027), .A2(n16798), .B1(n16810), .B2(n16821), .ZN(
        n16603) );
  NOR4_X1 U19798 ( .A1(n9790), .A2(n16605), .A3(n16604), .A4(n16603), .ZN(
        n16606) );
  OAI221_X1 U19799 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16607), .C1(n21167), 
        .C2(n16610), .A(n16606), .ZN(P3_U2653) );
  AOI211_X1 U19800 ( .C1(n17627), .C2(n16609), .A(n16608), .B(n18679), .ZN(
        n16615) );
  OAI21_X1 U19801 ( .B1(n16810), .B2(n16617), .A(n9796), .ZN(n16614) );
  INV_X1 U19802 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18728) );
  NAND2_X1 U19803 ( .A1(n16639), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n16629) );
  NOR2_X1 U19804 ( .A1(n18728), .A2(n16629), .ZN(n16612) );
  INV_X1 U19805 ( .A(n16610), .ZN(n16611) );
  MUX2_X1 U19806 ( .A(n16612), .B(n16611), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n16613) );
  NOR3_X1 U19807 ( .A1(n16615), .A2(n16614), .A3(n16613), .ZN(n16619) );
  OAI211_X1 U19808 ( .C1(n16620), .C2(n16617), .A(n16775), .B(n16616), .ZN(
        n16618) );
  OAI211_X1 U19809 ( .C1(n16798), .C2(n21007), .A(n16619), .B(n16618), .ZN(
        P3_U2654) );
  INV_X1 U19810 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18726) );
  AOI22_X1 U19811 ( .A1(n16639), .A2(n18726), .B1(n16815), .B2(n16644), .ZN(
        n16628) );
  AOI211_X1 U19812 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16634), .A(n16620), .B(
        n16809), .ZN(n16626) );
  INV_X1 U19813 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16820) );
  NAND2_X1 U19814 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17639), .ZN(
        n16630) );
  INV_X1 U19815 ( .A(n16630), .ZN(n16622) );
  OAI21_X1 U19816 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16622), .A(
        n16621), .ZN(n17643) );
  OAI21_X1 U19817 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16630), .A(
        n10009), .ZN(n16631) );
  AOI21_X1 U19818 ( .B1(n17643), .B2(n16631), .A(n18679), .ZN(n16623) );
  OAI21_X1 U19819 ( .B1(n17643), .B2(n16631), .A(n16623), .ZN(n16624) );
  OAI211_X1 U19820 ( .C1(n16810), .C2(n16820), .A(n9796), .B(n16624), .ZN(
        n16625) );
  AOI211_X1 U19821 ( .C1(n16796), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16626), .B(n16625), .ZN(n16627) );
  OAI221_X1 U19822 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16629), .C1(n18728), 
        .C2(n16628), .A(n16627), .ZN(P3_U2655) );
  NAND2_X1 U19823 ( .A1(n16815), .A2(n16644), .ZN(n16648) );
  OAI21_X1 U19824 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17639), .A(
        n16630), .ZN(n17648) );
  INV_X1 U19825 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16811) );
  NAND2_X1 U19826 ( .A1(n16811), .A2(n16737), .ZN(n16773) );
  INV_X1 U19827 ( .A(n16773), .ZN(n16667) );
  AOI22_X1 U19828 ( .A1(n16737), .A2(n17648), .B1(n17639), .B2(n16667), .ZN(
        n16632) );
  NOR2_X1 U19829 ( .A1(n18679), .A2(n10009), .ZN(n16668) );
  INV_X1 U19830 ( .A(n16668), .ZN(n16785) );
  AOI22_X1 U19831 ( .A1(n16632), .A2(n16785), .B1(n17648), .B2(n16631), .ZN(
        n16633) );
  AOI211_X1 U19832 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16796), .A(
        n9790), .B(n16633), .ZN(n16636) );
  OAI211_X1 U19833 ( .C1(n16641), .C2(n16637), .A(n16775), .B(n16634), .ZN(
        n16635) );
  OAI211_X1 U19834 ( .C1(n16637), .C2(n16810), .A(n16636), .B(n16635), .ZN(
        n16638) );
  AOI21_X1 U19835 ( .B1(n16639), .B2(n18726), .A(n16638), .ZN(n16640) );
  OAI21_X1 U19836 ( .B1(n16648), .B2(n18726), .A(n16640), .ZN(P3_U2656) );
  INV_X1 U19837 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17084) );
  AOI211_X1 U19838 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16655), .A(n16641), .B(
        n16809), .ZN(n16650) );
  INV_X1 U19839 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18725) );
  INV_X1 U19840 ( .A(n17674), .ZN(n16666) );
  NAND2_X1 U19841 ( .A1(n17682), .A2(n16666), .ZN(n16652) );
  AOI21_X1 U19842 ( .B1(n17663), .B2(n16652), .A(n17639), .ZN(n17666) );
  INV_X1 U19843 ( .A(n16652), .ZN(n16642) );
  AOI21_X1 U19844 ( .B1(n16642), .B2(n16811), .A(n9890), .ZN(n16654) );
  AOI21_X1 U19845 ( .B1(n17666), .B2(n16654), .A(n18679), .ZN(n16643) );
  OAI21_X1 U19846 ( .B1(n17666), .B2(n16654), .A(n16643), .ZN(n16647) );
  INV_X1 U19847 ( .A(n16664), .ZN(n16645) );
  NAND3_X1 U19848 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16645), .A3(n16644), 
        .ZN(n16646) );
  OAI211_X1 U19849 ( .C1(n16648), .C2(n18725), .A(n16647), .B(n16646), .ZN(
        n16649) );
  AOI211_X1 U19850 ( .C1(n16796), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16650), .B(n16649), .ZN(n16651) );
  OAI211_X1 U19851 ( .C1(n16810), .C2(n17084), .A(n16651), .B(n9796), .ZN(
        P3_U2657) );
  AOI22_X1 U19852 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16796), .B1(
        n16767), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n16663) );
  AOI21_X1 U19853 ( .B1(n16790), .B2(n16673), .A(n16812), .ZN(n16682) );
  OAI21_X1 U19854 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16756), .A(n16682), 
        .ZN(n16661) );
  AOI21_X1 U19855 ( .B1(n16667), .B2(n21066), .A(n16668), .ZN(n16659) );
  NOR2_X1 U19856 ( .A1(n17699), .A2(n17674), .ZN(n16653) );
  OAI21_X1 U19857 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16653), .A(
        n16652), .ZN(n17680) );
  NAND3_X1 U19858 ( .A1(n16737), .A2(n16654), .A3(n17680), .ZN(n16658) );
  OAI211_X1 U19859 ( .C1(n16671), .C2(n16656), .A(n16775), .B(n16655), .ZN(
        n16657) );
  OAI211_X1 U19860 ( .C1(n16659), .C2(n17680), .A(n16658), .B(n16657), .ZN(
        n16660) );
  AOI211_X1 U19861 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16661), .A(n9790), .B(
        n16660), .ZN(n16662) );
  OAI211_X1 U19862 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16664), .A(n16663), 
        .B(n16662), .ZN(P3_U2658) );
  INV_X1 U19863 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17111) );
  NOR2_X1 U19864 ( .A1(n16665), .A2(n16799), .ZN(n16670) );
  AOI22_X1 U19865 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17674), .B1(
        n16666), .B2(n17699), .ZN(n17695) );
  NOR2_X1 U19866 ( .A1(n16668), .A2(n16667), .ZN(n16807) );
  AOI211_X1 U19867 ( .C1(n10009), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16807), .B(n17695), .ZN(n16669) );
  AOI211_X1 U19868 ( .C1(n16670), .C2(n17695), .A(n9790), .B(n16669), .ZN(
        n16677) );
  AOI211_X1 U19869 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16685), .A(n16671), .B(
        n16809), .ZN(n16675) );
  NAND2_X1 U19870 ( .A1(n16790), .A2(n18721), .ZN(n16672) );
  OAI22_X1 U19871 ( .A1(n18721), .A2(n16682), .B1(n16673), .B2(n16672), .ZN(
        n16674) );
  AOI211_X1 U19872 ( .C1(n16796), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16675), .B(n16674), .ZN(n16676) );
  OAI211_X1 U19873 ( .C1(n16810), .C2(n17111), .A(n16677), .B(n16676), .ZN(
        P3_U2659) );
  AOI21_X1 U19874 ( .B1(n16790), .B2(n16678), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16683) );
  INV_X1 U19875 ( .A(n16679), .ZN(n16734) );
  NOR2_X1 U19876 ( .A1(n17746), .A2(n16734), .ZN(n16712) );
  NAND2_X1 U19877 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16712), .ZN(
        n16701) );
  NOR2_X1 U19878 ( .A1(n16693), .A2(n16701), .ZN(n16692) );
  AOI21_X1 U19879 ( .B1(n16692), .B2(n16811), .A(n9890), .ZN(n16680) );
  OAI21_X1 U19880 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16692), .A(
        n17674), .ZN(n17721) );
  XOR2_X1 U19881 ( .A(n16680), .B(n17721), .Z(n16681) );
  OAI22_X1 U19882 ( .A1(n16683), .A2(n16682), .B1(n18679), .B2(n16681), .ZN(
        n16684) );
  AOI211_X1 U19883 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n16796), .A(
        n9790), .B(n16684), .ZN(n16687) );
  OAI211_X1 U19884 ( .C1(n16691), .C2(n16688), .A(n16775), .B(n16685), .ZN(
        n16686) );
  OAI211_X1 U19885 ( .C1(n16688), .C2(n16810), .A(n16687), .B(n16686), .ZN(
        P3_U2660) );
  NOR2_X1 U19886 ( .A1(n16690), .A2(n16756), .ZN(n16689) );
  NOR2_X1 U19887 ( .A1(n16812), .A2(n16689), .ZN(n16715) );
  INV_X1 U19888 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n21076) );
  NAND3_X1 U19889 ( .A1(n16790), .A2(n16690), .A3(n21076), .ZN(n16706) );
  AOI211_X1 U19890 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16704), .A(n16691), .B(
        n16809), .ZN(n16699) );
  NAND2_X1 U19891 ( .A1(n16790), .A2(n18716), .ZN(n16696) );
  AOI21_X1 U19892 ( .B1(n16693), .B2(n16701), .A(n16692), .ZN(n17729) );
  OAI21_X1 U19893 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16701), .A(
        n10009), .ZN(n16703) );
  XNOR2_X1 U19894 ( .A(n17729), .B(n16703), .ZN(n16694) );
  AOI22_X1 U19895 ( .A1(n16767), .A2(P3_EBX_REG_10__SCAN_IN), .B1(n16737), 
        .B2(n16694), .ZN(n16695) );
  OAI211_X1 U19896 ( .C1(n16697), .C2(n16696), .A(n16695), .B(n9796), .ZN(
        n16698) );
  AOI211_X1 U19897 ( .C1(n16796), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16699), .B(n16698), .ZN(n16700) );
  OAI221_X1 U19898 ( .B1(n18716), .B2(n16715), .C1(n18716), .C2(n16706), .A(
        n16700), .ZN(P3_U2661) );
  OAI21_X1 U19899 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16712), .A(
        n16701), .ZN(n17738) );
  OAI221_X1 U19900 ( .B1(n17738), .B2(n17709), .C1(n17738), .C2(n16811), .A(
        n16737), .ZN(n16702) );
  AOI22_X1 U19901 ( .A1(n17738), .A2(n16703), .B1(n16785), .B2(n16702), .ZN(
        n16710) );
  OAI211_X1 U19902 ( .C1(n16717), .C2(n16707), .A(n16775), .B(n16704), .ZN(
        n16705) );
  OAI21_X1 U19903 ( .B1(n16798), .B2(n17709), .A(n16705), .ZN(n16709) );
  OAI21_X1 U19904 ( .B1(n16707), .B2(n16810), .A(n16706), .ZN(n16708) );
  NOR4_X1 U19905 ( .A1(n9790), .A2(n16710), .A3(n16709), .A4(n16708), .ZN(
        n16711) );
  OAI21_X1 U19906 ( .B1(n16715), .B2(n21076), .A(n16711), .ZN(P3_U2662) );
  AND2_X1 U19907 ( .A1(n17708), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17747) );
  NOR2_X1 U19908 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17841), .ZN(
        n16789) );
  AOI21_X1 U19909 ( .B1(n17747), .B2(n16789), .A(n9890), .ZN(n16714) );
  INV_X1 U19910 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17763) );
  NOR2_X1 U19911 ( .A1(n17763), .A2(n16734), .ZN(n16723) );
  INV_X1 U19912 ( .A(n16712), .ZN(n16713) );
  OAI21_X1 U19913 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16723), .A(
        n16713), .ZN(n17749) );
  XOR2_X1 U19914 ( .A(n16714), .B(n17749), .Z(n16722) );
  AOI21_X1 U19915 ( .B1(n16767), .B2(P3_EBX_REG_8__SCAN_IN), .A(n9790), .ZN(
        n16721) );
  AOI221_X1 U19916 ( .B1(n16756), .B2(n18713), .C1(n16716), .C2(n18713), .A(
        n16715), .ZN(n16719) );
  AOI211_X1 U19917 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16730), .A(n16717), .B(
        n16809), .ZN(n16718) );
  AOI211_X1 U19918 ( .C1(n16796), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16719), .B(n16718), .ZN(n16720) );
  OAI211_X1 U19919 ( .C1(n18679), .C2(n16722), .A(n16721), .B(n16720), .ZN(
        P3_U2663) );
  AOI21_X1 U19920 ( .B1(n17763), .B2(n16734), .A(n16723), .ZN(n17768) );
  AOI21_X1 U19921 ( .B1(n17708), .B2(n16789), .A(n9890), .ZN(n16736) );
  OAI21_X1 U19922 ( .B1(n17768), .B2(n16736), .A(n16737), .ZN(n16724) );
  AOI21_X1 U19923 ( .B1(n17768), .B2(n16736), .A(n16724), .ZN(n16729) );
  NAND2_X1 U19924 ( .A1(n16790), .A2(n16725), .ZN(n16727) );
  INV_X1 U19925 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18711) );
  AOI221_X1 U19926 ( .B1(n18709), .B2(n16790), .C1(n16742), .C2(n16790), .A(
        n16812), .ZN(n16726) );
  OAI221_X1 U19927 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n16727), .C1(n18711), 
        .C2(n16726), .A(n9796), .ZN(n16728) );
  AOI211_X1 U19928 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16767), .A(n16729), .B(
        n16728), .ZN(n16732) );
  OAI211_X1 U19929 ( .C1(n16733), .C2(n17174), .A(n16775), .B(n16730), .ZN(
        n16731) );
  OAI211_X1 U19930 ( .C1(n16798), .C2(n17763), .A(n16732), .B(n16731), .ZN(
        P3_U2664) );
  AOI211_X1 U19931 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16751), .A(n16733), .B(
        n16809), .ZN(n16741) );
  AOI21_X1 U19932 ( .B1(n16790), .B2(n16742), .A(n16812), .ZN(n16749) );
  NOR2_X1 U19933 ( .A1(n17841), .A2(n17781), .ZN(n16746) );
  OAI21_X1 U19934 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16746), .A(
        n16734), .ZN(n17780) );
  AOI211_X1 U19935 ( .C1(n10009), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16807), .B(n17780), .ZN(n16735) );
  NOR2_X1 U19936 ( .A1(n9790), .A2(n16735), .ZN(n16739) );
  NAND3_X1 U19937 ( .A1(n16737), .A2(n16736), .A3(n17780), .ZN(n16738) );
  OAI211_X1 U19938 ( .C1(n16749), .C2(n18709), .A(n16739), .B(n16738), .ZN(
        n16740) );
  AOI211_X1 U19939 ( .C1(n16796), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16741), .B(n16740), .ZN(n16744) );
  OR3_X1 U19940 ( .A1(n16756), .A2(n16742), .A3(P3_REIP_REG_6__SCAN_IN), .ZN(
        n16743) );
  OAI211_X1 U19941 ( .C1(n10120), .C2(n16810), .A(n16744), .B(n16743), .ZN(
        P3_U2665) );
  INV_X1 U19942 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16754) );
  AOI21_X1 U19943 ( .B1(n16790), .B2(n16745), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16748) );
  NAND2_X1 U19944 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17783), .ZN(
        n16759) );
  AOI21_X1 U19945 ( .B1(n16754), .B2(n16759), .A(n16746), .ZN(n17791) );
  OAI21_X1 U19946 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16759), .A(
        n10009), .ZN(n16760) );
  XOR2_X1 U19947 ( .A(n17791), .B(n16760), .Z(n16747) );
  OAI22_X1 U19948 ( .A1(n16749), .A2(n16748), .B1(n18679), .B2(n16747), .ZN(
        n16750) );
  AOI211_X1 U19949 ( .C1(n16767), .C2(P3_EBX_REG_5__SCAN_IN), .A(n9790), .B(
        n16750), .ZN(n16753) );
  OAI211_X1 U19950 ( .C1(n16758), .C2(n17183), .A(n16775), .B(n16751), .ZN(
        n16752) );
  OAI211_X1 U19951 ( .C1(n16798), .C2(n16754), .A(n16753), .B(n16752), .ZN(
        P3_U2666) );
  AOI21_X1 U19952 ( .B1(n16790), .B2(n16755), .A(n16812), .ZN(n16777) );
  NOR3_X1 U19953 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16756), .A3(n16755), .ZN(
        n16757) );
  AOI21_X1 U19954 ( .B1(n16796), .B2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16757), .ZN(n16769) );
  AOI211_X1 U19955 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16774), .A(n16758), .B(
        n16809), .ZN(n16766) );
  OAI21_X1 U19956 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16770), .A(
        n16759), .ZN(n17805) );
  INV_X1 U19957 ( .A(n17805), .ZN(n16761) );
  AOI22_X1 U19958 ( .A1(n16761), .A2(n10009), .B1(n16760), .B2(n17805), .ZN(
        n16762) );
  AOI21_X1 U19959 ( .B1(n17799), .B2(n16789), .A(n16762), .ZN(n16764) );
  NOR2_X1 U19960 ( .A1(n16818), .A2(n18826), .ZN(n16783) );
  OAI21_X1 U19961 ( .B1(n16916), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16783), .ZN(n16763) );
  OAI211_X1 U19962 ( .C1(n16764), .C2(n18679), .A(n9796), .B(n16763), .ZN(
        n16765) );
  AOI211_X1 U19963 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16767), .A(n16766), .B(
        n16765), .ZN(n16768) );
  OAI211_X1 U19964 ( .C1(n18705), .C2(n16777), .A(n16769), .B(n16768), .ZN(
        P3_U2667) );
  NOR2_X1 U19965 ( .A1(n18796), .A2(n13971), .ZN(n18626) );
  OAI21_X1 U19966 ( .B1(n18626), .B2(n18775), .A(n16859), .ZN(n18772) );
  NAND2_X1 U19967 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16784) );
  INV_X1 U19968 ( .A(n16784), .ZN(n16772) );
  AOI21_X1 U19969 ( .B1(n16772), .B2(n16811), .A(n16799), .ZN(n16788) );
  INV_X1 U19970 ( .A(n16770), .ZN(n16771) );
  OAI21_X1 U19971 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16772), .A(
        n16771), .ZN(n17822) );
  AOI22_X1 U19972 ( .A1(n16783), .A2(n18772), .B1(n16788), .B2(n17822), .ZN(
        n16782) );
  AOI221_X1 U19973 ( .B1(n16784), .B2(n16785), .C1(n16773), .C2(n16785), .A(
        n17822), .ZN(n16780) );
  NAND3_X1 U19974 ( .A1(n16790), .A2(P3_REIP_REG_1__SCAN_IN), .A3(
        P3_REIP_REG_2__SCAN_IN), .ZN(n16778) );
  INV_X1 U19975 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18703) );
  OAI211_X1 U19976 ( .C1(n16786), .C2(n17195), .A(n16775), .B(n16774), .ZN(
        n16776) );
  OAI221_X1 U19977 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(n16778), .C1(n18703), 
        .C2(n16777), .A(n16776), .ZN(n16779) );
  AOI211_X1 U19978 ( .C1(n16796), .C2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n16780), .B(n16779), .ZN(n16781) );
  OAI211_X1 U19979 ( .C1(n16810), .C2(n17195), .A(n16782), .B(n16781), .ZN(
        P3_U2668) );
  INV_X1 U19980 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18701) );
  NAND2_X1 U19981 ( .A1(n16790), .A2(n18798), .ZN(n16805) );
  NAND2_X1 U19982 ( .A1(n18641), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n18630) );
  NAND2_X1 U19983 ( .A1(n10497), .A2(n18630), .ZN(n18624) );
  OAI21_X1 U19984 ( .B1(n13971), .B2(n18796), .A(n18624), .ZN(n18780) );
  INV_X1 U19985 ( .A(n16783), .ZN(n18828) );
  OAI21_X1 U19986 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16784), .ZN(n17828) );
  OAI22_X1 U19987 ( .A1(n18780), .A2(n18828), .B1(n17828), .B2(n16785), .ZN(
        n16795) );
  INV_X1 U19988 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16793) );
  INV_X1 U19989 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n16808) );
  INV_X1 U19990 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17201) );
  NAND2_X1 U19991 ( .A1(n16808), .A2(n17201), .ZN(n16801) );
  AOI211_X1 U19992 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16801), .A(n16786), .B(
        n16809), .ZN(n16787) );
  AOI221_X1 U19993 ( .B1(n16789), .B2(n16788), .C1(n17828), .C2(n16788), .A(
        n16787), .ZN(n16792) );
  NAND3_X1 U19994 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16790), .A3(n18701), 
        .ZN(n16791) );
  OAI211_X1 U19995 ( .C1(n16793), .C2(n16810), .A(n16792), .B(n16791), .ZN(
        n16794) );
  AOI211_X1 U19996 ( .C1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n16796), .A(
        n16795), .B(n16794), .ZN(n16797) );
  OAI221_X1 U19997 ( .B1(n18701), .B2(n16800), .C1(n18701), .C2(n16805), .A(
        n16797), .ZN(P3_U2669) );
  OAI21_X1 U19998 ( .B1(n16811), .B2(n16799), .A(n16798), .ZN(n16804) );
  OAI22_X1 U19999 ( .A1(n10495), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n18796), .B2(n18641), .ZN(n18788) );
  INV_X1 U20000 ( .A(n18788), .ZN(n18642) );
  OAI22_X1 U20001 ( .A1(n18798), .A2(n16800), .B1(n18642), .B2(n18828), .ZN(
        n16803) );
  OAI21_X1 U20002 ( .B1(n17201), .B2(n16808), .A(n16801), .ZN(n17203) );
  OAI22_X1 U20003 ( .A1(n16810), .A2(n17201), .B1(n16809), .B2(n17203), .ZN(
        n16802) );
  AOI211_X1 U20004 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n16804), .A(
        n16803), .B(n16802), .ZN(n16806) );
  OAI211_X1 U20005 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n16807), .A(
        n16806), .B(n16805), .ZN(P3_U2670) );
  AOI21_X1 U20006 ( .B1(n16810), .B2(n16809), .A(n16808), .ZN(n16814) );
  INV_X1 U20007 ( .A(n18824), .ZN(n18793) );
  NOR3_X1 U20008 ( .A1(n18793), .A2(n16812), .A3(n16811), .ZN(n16813) );
  AOI211_X1 U20009 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(n16815), .A(n16814), .B(
        n16813), .ZN(n16816) );
  OAI21_X1 U20010 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18828), .A(
        n16816), .ZN(P3_U2671) );
  INV_X1 U20011 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n21021) );
  NAND2_X1 U20012 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16936) );
  INV_X1 U20013 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16822) );
  INV_X1 U20014 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17177) );
  NOR2_X1 U20015 ( .A1(n16822), .A2(n17017), .ZN(n16980) );
  NAND4_X1 U20016 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .A4(n16980), .ZN(n16823) );
  NOR4_X1 U20017 ( .A1(n10110), .A2(n21069), .A3(n16936), .A4(n16823), .ZN(
        n16824) );
  NAND3_X1 U20018 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(n16824), .ZN(n16930) );
  NAND2_X1 U20019 ( .A1(n9793), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16826) );
  NAND2_X1 U20020 ( .A1(n16929), .A2(n18206), .ZN(n16825) );
  OAI22_X1 U20021 ( .A1(n16929), .A2(n16826), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16825), .ZN(P3_U2672) );
  AOI22_X1 U20022 ( .A1(n10396), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16830) );
  AOI22_X1 U20023 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16829) );
  AOI22_X1 U20024 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16828) );
  AOI22_X1 U20025 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16827) );
  NAND4_X1 U20026 ( .A1(n16830), .A2(n16829), .A3(n16828), .A4(n16827), .ZN(
        n16836) );
  AOI22_X1 U20027 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16834) );
  AOI22_X1 U20028 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16833) );
  AOI22_X1 U20029 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16832) );
  AOI22_X1 U20030 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16831) );
  NAND4_X1 U20031 ( .A1(n16834), .A2(n16833), .A3(n16832), .A4(n16831), .ZN(
        n16835) );
  NOR2_X1 U20032 ( .A1(n16836), .A2(n16835), .ZN(n16941) );
  AOI22_X1 U20033 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16840) );
  AOI22_X1 U20034 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16839) );
  AOI22_X1 U20035 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16838) );
  AOI22_X1 U20036 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16837) );
  NAND4_X1 U20037 ( .A1(n16840), .A2(n16839), .A3(n16838), .A4(n16837), .ZN(
        n16846) );
  AOI22_X1 U20038 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16882), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16844) );
  AOI22_X1 U20039 ( .A1(n10396), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16843) );
  AOI22_X1 U20040 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16842) );
  AOI22_X1 U20041 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10387), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16841) );
  NAND4_X1 U20042 ( .A1(n16844), .A2(n16843), .A3(n16842), .A4(n16841), .ZN(
        n16845) );
  NOR2_X1 U20043 ( .A1(n16846), .A2(n16845), .ZN(n16951) );
  AOI22_X1 U20044 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17138), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16850) );
  AOI22_X1 U20045 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17162), .B1(
        n9792), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16849) );
  AOI22_X1 U20046 ( .A1(n10396), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16848) );
  AOI22_X1 U20047 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n10414), .ZN(n16847) );
  NAND4_X1 U20048 ( .A1(n16850), .A2(n16849), .A3(n16848), .A4(n16847), .ZN(
        n16856) );
  AOI22_X1 U20049 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n16916), .ZN(n16854) );
  AOI22_X1 U20050 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17158), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17144), .ZN(n16853) );
  AOI22_X1 U20051 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n9795), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17057), .ZN(n16852) );
  AOI22_X1 U20052 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16851) );
  NAND4_X1 U20053 ( .A1(n16854), .A2(n16853), .A3(n16852), .A4(n16851), .ZN(
        n16855) );
  NOR2_X1 U20054 ( .A1(n16856), .A2(n16855), .ZN(n16961) );
  AOI22_X1 U20055 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16868) );
  AOI22_X1 U20056 ( .A1(n16878), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16867) );
  AOI22_X1 U20057 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9788), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16857) );
  OAI21_X1 U20058 ( .B1(n16858), .B2(n17207), .A(n16857), .ZN(n16865) );
  AOI22_X1 U20059 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16863) );
  AOI22_X1 U20060 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16862) );
  AOI22_X1 U20061 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16861) );
  AOI22_X1 U20062 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16860) );
  NAND4_X1 U20063 ( .A1(n16863), .A2(n16862), .A3(n16861), .A4(n16860), .ZN(
        n16864) );
  AOI211_X1 U20064 ( .C1(n17161), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n16865), .B(n16864), .ZN(n16866) );
  NAND3_X1 U20065 ( .A1(n16868), .A2(n16867), .A3(n16866), .ZN(n16965) );
  AOI22_X1 U20066 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16882), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16881) );
  AOI22_X1 U20067 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16880) );
  AOI22_X1 U20068 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16869) );
  OAI21_X1 U20069 ( .B1(n16871), .B2(n16870), .A(n16869), .ZN(n16877) );
  AOI22_X1 U20070 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9792), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16875) );
  AOI22_X1 U20071 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16874) );
  AOI22_X1 U20072 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16873) );
  AOI22_X1 U20073 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16872) );
  NAND4_X1 U20074 ( .A1(n16875), .A2(n16874), .A3(n16873), .A4(n16872), .ZN(
        n16876) );
  AOI211_X1 U20075 ( .C1(n16878), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n16877), .B(n16876), .ZN(n16879) );
  NAND3_X1 U20076 ( .A1(n16881), .A2(n16880), .A3(n16879), .ZN(n16966) );
  NAND2_X1 U20077 ( .A1(n16965), .A2(n16966), .ZN(n16964) );
  NOR2_X1 U20078 ( .A1(n16961), .A2(n16964), .ZN(n16958) );
  AOI22_X1 U20079 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16894) );
  AOI22_X1 U20080 ( .A1(n16878), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16882), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16893) );
  AOI22_X1 U20081 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16883) );
  OAI21_X1 U20082 ( .B1(n16884), .B2(n21128), .A(n16883), .ZN(n16891) );
  AOI22_X1 U20083 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U20084 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16885), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16888) );
  AOI22_X1 U20085 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16887) );
  AOI22_X1 U20086 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16886) );
  NAND4_X1 U20087 ( .A1(n16889), .A2(n16888), .A3(n16887), .A4(n16886), .ZN(
        n16890) );
  AOI211_X1 U20088 ( .C1(n9792), .C2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n16891), .B(n16890), .ZN(n16892) );
  NAND3_X1 U20089 ( .A1(n16894), .A2(n16893), .A3(n16892), .ZN(n16957) );
  NAND2_X1 U20090 ( .A1(n16958), .A2(n16957), .ZN(n16956) );
  NOR2_X1 U20091 ( .A1(n16951), .A2(n16956), .ZN(n16950) );
  AOI22_X1 U20092 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10416), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16904) );
  AOI22_X1 U20093 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16903) );
  AOI22_X1 U20094 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16895) );
  OAI21_X1 U20095 ( .B1(n10511), .B2(n20970), .A(n16895), .ZN(n16901) );
  AOI22_X1 U20096 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16899) );
  AOI22_X1 U20097 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16898) );
  AOI22_X1 U20098 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16897) );
  AOI22_X1 U20099 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16896) );
  NAND4_X1 U20100 ( .A1(n16899), .A2(n16898), .A3(n16897), .A4(n16896), .ZN(
        n16900) );
  AOI211_X1 U20101 ( .C1(n16885), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n16901), .B(n16900), .ZN(n16902) );
  NAND3_X1 U20102 ( .A1(n16904), .A2(n16903), .A3(n16902), .ZN(n16947) );
  NAND2_X1 U20103 ( .A1(n16950), .A2(n16947), .ZN(n16946) );
  NOR2_X1 U20104 ( .A1(n16941), .A2(n16946), .ZN(n16940) );
  INV_X1 U20105 ( .A(n16940), .ZN(n16935) );
  AOI22_X1 U20106 ( .A1(n16878), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16909) );
  AOI22_X1 U20107 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16908) );
  AOI22_X1 U20108 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16907) );
  AOI22_X1 U20109 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16906) );
  NAND4_X1 U20110 ( .A1(n16909), .A2(n16908), .A3(n16907), .A4(n16906), .ZN(
        n16915) );
  AOI22_X1 U20111 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20112 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20113 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16911) );
  AOI22_X1 U20114 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16910) );
  NAND4_X1 U20115 ( .A1(n16913), .A2(n16912), .A3(n16911), .A4(n16910), .ZN(
        n16914) );
  NOR2_X1 U20116 ( .A1(n16915), .A2(n16914), .ZN(n16934) );
  NOR2_X1 U20117 ( .A1(n16935), .A2(n16934), .ZN(n16928) );
  AOI22_X1 U20118 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16920) );
  AOI22_X1 U20119 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16919) );
  AOI22_X1 U20120 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16916), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16918) );
  AOI22_X1 U20121 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16917) );
  NAND4_X1 U20122 ( .A1(n16920), .A2(n16919), .A3(n16918), .A4(n16917), .ZN(
        n16926) );
  AOI22_X1 U20123 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16924) );
  AOI22_X1 U20124 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16923) );
  AOI22_X1 U20125 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16922) );
  AOI22_X1 U20126 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16921) );
  NAND4_X1 U20127 ( .A1(n16924), .A2(n16923), .A3(n16922), .A4(n16921), .ZN(
        n16925) );
  NOR2_X1 U20128 ( .A1(n16926), .A2(n16925), .ZN(n16927) );
  XOR2_X1 U20129 ( .A(n16928), .B(n16927), .Z(n17212) );
  AOI21_X1 U20130 ( .B1(n16930), .B2(n21021), .A(n16929), .ZN(n16931) );
  NAND2_X1 U20131 ( .A1(n9793), .A2(n16931), .ZN(n16932) );
  OAI21_X1 U20132 ( .B1(n17212), .B2(n9793), .A(n16932), .ZN(P3_U2673) );
  NAND2_X1 U20133 ( .A1(n18206), .A2(n9826), .ZN(n17202) );
  INV_X1 U20134 ( .A(n17202), .ZN(n17205) );
  NAND2_X1 U20135 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17005), .ZN(n16993) );
  NOR2_X1 U20136 ( .A1(n17193), .A2(n16955), .ZN(n16952) );
  AOI21_X1 U20137 ( .B1(n17205), .B2(n16936), .A(n16952), .ZN(n16943) );
  INV_X1 U20138 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16939) );
  XOR2_X1 U20139 ( .A(n16935), .B(n16934), .Z(n17213) );
  NOR3_X1 U20140 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16949), .A3(n16936), .ZN(
        n16937) );
  AOI21_X1 U20141 ( .B1(n17193), .B2(n17213), .A(n16937), .ZN(n16938) );
  OAI21_X1 U20142 ( .B1(n16943), .B2(n16939), .A(n16938), .ZN(P3_U2674) );
  NAND2_X1 U20143 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16955), .ZN(n16945) );
  AOI21_X1 U20144 ( .B1(n16941), .B2(n16946), .A(n16940), .ZN(n17217) );
  NAND2_X1 U20145 ( .A1(n17193), .A2(n17217), .ZN(n16942) );
  OAI221_X1 U20146 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16945), .C1(n16944), 
        .C2(n16943), .A(n16942), .ZN(P3_U2675) );
  OAI21_X1 U20147 ( .B1(n16950), .B2(n16947), .A(n16946), .ZN(n17226) );
  NAND3_X1 U20148 ( .A1(n16949), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n9793), .ZN(
        n16948) );
  OAI221_X1 U20149 ( .B1(n16949), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n9793), 
        .C2(n17226), .A(n16948), .ZN(P3_U2676) );
  NAND2_X1 U20150 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16963), .ZN(n16954) );
  AOI21_X1 U20151 ( .B1(n16951), .B2(n16956), .A(n16950), .ZN(n17227) );
  AOI22_X1 U20152 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16952), .B1(n17193), 
        .B2(n17227), .ZN(n16953) );
  OAI21_X1 U20153 ( .B1(n16955), .B2(n16954), .A(n16953), .ZN(P3_U2677) );
  OAI21_X1 U20154 ( .B1(n16958), .B2(n16957), .A(n16956), .ZN(n17237) );
  NAND3_X1 U20155 ( .A1(n16960), .A2(P3_EBX_REG_25__SCAN_IN), .A3(n9793), .ZN(
        n16959) );
  OAI221_X1 U20156 ( .B1(n16960), .B2(P3_EBX_REG_25__SCAN_IN), .C1(n9793), 
        .C2(n17237), .A(n16959), .ZN(P3_U2678) );
  AOI21_X1 U20157 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n9793), .A(n9897), .ZN(
        n16962) );
  XNOR2_X1 U20158 ( .A(n16961), .B(n16964), .ZN(n17242) );
  OAI22_X1 U20159 ( .A1(n16963), .A2(n16962), .B1(n9793), .B2(n17242), .ZN(
        P3_U2679) );
  AOI21_X1 U20160 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n9793), .A(n9898), .ZN(
        n16967) );
  OAI21_X1 U20161 ( .B1(n16966), .B2(n16965), .A(n16964), .ZN(n17247) );
  OAI22_X1 U20162 ( .A1(n9897), .A2(n16967), .B1(n9793), .B2(n17247), .ZN(
        P3_U2680) );
  AOI21_X1 U20163 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n9793), .A(n16968), .ZN(
        n16979) );
  AOI22_X1 U20164 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10397), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20165 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U20166 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16970) );
  AOI22_X1 U20167 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16969) );
  NAND4_X1 U20168 ( .A1(n16972), .A2(n16971), .A3(n16970), .A4(n16969), .ZN(
        n16978) );
  AOI22_X1 U20169 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16976) );
  AOI22_X1 U20170 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9792), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16975) );
  AOI22_X1 U20171 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20172 ( .A1(n16878), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16973) );
  NAND4_X1 U20173 ( .A1(n16976), .A2(n16975), .A3(n16974), .A4(n16973), .ZN(
        n16977) );
  NOR2_X1 U20174 ( .A1(n16978), .A2(n16977), .ZN(n17251) );
  OAI22_X1 U20175 ( .A1(n9898), .A2(n16979), .B1(n17251), .B2(n9793), .ZN(
        P3_U2681) );
  NOR2_X1 U20176 ( .A1(n17193), .A2(n16980), .ZN(n17004) );
  AOI22_X1 U20177 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16991) );
  AOI22_X1 U20178 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16990) );
  INV_X1 U20179 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n21049) );
  AOI22_X1 U20180 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16981) );
  OAI21_X1 U20181 ( .B1(n16982), .B2(n21049), .A(n16981), .ZN(n16988) );
  AOI22_X1 U20182 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16986) );
  AOI22_X1 U20183 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U20184 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16916), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16984) );
  AOI22_X1 U20185 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16983) );
  NAND4_X1 U20186 ( .A1(n16986), .A2(n16985), .A3(n16984), .A4(n16983), .ZN(
        n16987) );
  AOI211_X1 U20187 ( .C1(n9792), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n16988), .B(n16987), .ZN(n16989) );
  NAND3_X1 U20188 ( .A1(n16991), .A2(n16990), .A3(n16989), .ZN(n17255) );
  AOI22_X1 U20189 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17004), .B1(n17193), 
        .B2(n17255), .ZN(n16992) );
  OAI21_X1 U20190 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16993), .A(n16992), .ZN(
        P3_U2682) );
  AOI22_X1 U20191 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16997) );
  AOI22_X1 U20192 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16996) );
  AOI22_X1 U20193 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20194 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16994) );
  NAND4_X1 U20195 ( .A1(n16997), .A2(n16996), .A3(n16995), .A4(n16994), .ZN(
        n17003) );
  AOI22_X1 U20196 ( .A1(n16878), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20197 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20198 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20199 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16998) );
  NAND4_X1 U20200 ( .A1(n17001), .A2(n17000), .A3(n16999), .A4(n16998), .ZN(
        n17002) );
  NOR2_X1 U20201 ( .A1(n17003), .A2(n17002), .ZN(n17263) );
  OAI21_X1 U20202 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17005), .A(n17004), .ZN(
        n17006) );
  OAI21_X1 U20203 ( .B1(n17263), .B2(n9793), .A(n17006), .ZN(P3_U2683) );
  AOI22_X1 U20204 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20205 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17009) );
  AOI22_X1 U20206 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10397), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20207 ( .A1(n16878), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17007) );
  NAND4_X1 U20208 ( .A1(n17010), .A2(n17009), .A3(n17008), .A4(n17007), .ZN(
        n17016) );
  AOI22_X1 U20209 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20210 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20211 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U20212 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17011) );
  NAND4_X1 U20213 ( .A1(n17014), .A2(n17013), .A3(n17012), .A4(n17011), .ZN(
        n17015) );
  NOR2_X1 U20214 ( .A1(n17016), .A2(n17015), .ZN(n17268) );
  OAI21_X1 U20215 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n9900), .A(n17017), .ZN(
        n17018) );
  AOI22_X1 U20216 ( .A1(n17193), .A2(n17268), .B1(n17018), .B2(n9793), .ZN(
        P3_U2684) );
  NOR2_X1 U20217 ( .A1(n17248), .A2(n17019), .ZN(n17041) );
  OAI21_X1 U20218 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17041), .A(n9793), .ZN(
        n17030) );
  AOI22_X1 U20219 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20220 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20221 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17021) );
  AOI22_X1 U20222 ( .A1(n10396), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17020) );
  NAND4_X1 U20223 ( .A1(n17023), .A2(n17022), .A3(n17021), .A4(n17020), .ZN(
        n17029) );
  AOI22_X1 U20224 ( .A1(n16878), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16916), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20225 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20226 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U20227 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17024) );
  NAND4_X1 U20228 ( .A1(n17027), .A2(n17026), .A3(n17025), .A4(n17024), .ZN(
        n17028) );
  NOR2_X1 U20229 ( .A1(n17029), .A2(n17028), .ZN(n17272) );
  OAI22_X1 U20230 ( .A1(n9900), .A2(n17030), .B1(n17272), .B2(n9793), .ZN(
        P3_U2685) );
  AOI22_X1 U20231 ( .A1(n10396), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17057), .ZN(n17034) );
  AOI22_X1 U20232 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20233 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n16916), .ZN(n17032) );
  AOI22_X1 U20234 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17144), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n10414), .ZN(n17031) );
  NAND4_X1 U20235 ( .A1(n17034), .A2(n17033), .A3(n17032), .A4(n17031), .ZN(
        n17040) );
  AOI22_X1 U20236 ( .A1(n16878), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20237 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17162), .ZN(n17037) );
  AOI22_X1 U20238 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17163), .ZN(n17036) );
  AOI22_X1 U20239 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17158), .ZN(n17035) );
  NAND4_X1 U20240 ( .A1(n17038), .A2(n17037), .A3(n17036), .A4(n17035), .ZN(
        n17039) );
  NOR2_X1 U20241 ( .A1(n17040), .A2(n17039), .ZN(n17278) );
  NOR3_X1 U20242 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17193), .A3(n17053), .ZN(
        n17042) );
  AOI211_X1 U20243 ( .C1(n17193), .C2(n17278), .A(n17042), .B(n17041), .ZN(
        P3_U2686) );
  AOI22_X1 U20244 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17046) );
  AOI22_X1 U20245 ( .A1(n16878), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20246 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20247 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17043) );
  NAND4_X1 U20248 ( .A1(n17046), .A2(n17045), .A3(n17044), .A4(n17043), .ZN(
        n17052) );
  AOI22_X1 U20249 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17050) );
  AOI22_X1 U20250 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20251 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20252 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17047) );
  NAND4_X1 U20253 ( .A1(n17050), .A2(n17049), .A3(n17048), .A4(n17047), .ZN(
        n17051) );
  NOR2_X1 U20254 ( .A1(n17052), .A2(n17051), .ZN(n17284) );
  INV_X1 U20255 ( .A(n17068), .ZN(n17055) );
  NOR2_X1 U20256 ( .A1(n17193), .A2(n17053), .ZN(n17054) );
  OAI21_X1 U20257 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17055), .A(n17054), .ZN(
        n17056) );
  OAI21_X1 U20258 ( .B1(n17284), .B2(n9793), .A(n17056), .ZN(P3_U2687) );
  AOI22_X1 U20259 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U20260 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17060) );
  AOI22_X1 U20261 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10416), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17059) );
  AOI22_X1 U20262 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17058) );
  NAND4_X1 U20263 ( .A1(n17061), .A2(n17060), .A3(n17059), .A4(n17058), .ZN(
        n17067) );
  AOI22_X1 U20264 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U20265 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17064) );
  AOI22_X1 U20266 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17063) );
  AOI22_X1 U20267 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17062) );
  NAND4_X1 U20268 ( .A1(n17065), .A2(n17064), .A3(n17063), .A4(n17062), .ZN(
        n17066) );
  NOR2_X1 U20269 ( .A1(n17067), .A2(n17066), .ZN(n17289) );
  OAI21_X1 U20270 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17069), .A(n17068), .ZN(
        n17070) );
  AOI22_X1 U20271 ( .A1(n17193), .A2(n17289), .B1(n17070), .B2(n9793), .ZN(
        P3_U2688) );
  NAND2_X1 U20272 ( .A1(n9793), .A2(n17081), .ZN(n17096) );
  AOI22_X1 U20273 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17080) );
  AOI22_X1 U20274 ( .A1(n16878), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U20275 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17071) );
  OAI21_X1 U20276 ( .B1(n10435), .B2(n21159), .A(n17071), .ZN(n17077) );
  AOI22_X1 U20277 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17075) );
  AOI22_X1 U20278 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17074) );
  AOI22_X1 U20279 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20280 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17072) );
  NAND4_X1 U20281 ( .A1(n17075), .A2(n17074), .A3(n17073), .A4(n17072), .ZN(
        n17076) );
  AOI211_X1 U20282 ( .C1(n9792), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17077), .B(n17076), .ZN(n17078) );
  NAND3_X1 U20283 ( .A1(n17080), .A2(n17079), .A3(n17078), .ZN(n17291) );
  NOR3_X1 U20284 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17248), .A3(n17081), .ZN(
        n17082) );
  AOI21_X1 U20285 ( .B1(n17193), .B2(n17291), .A(n17082), .ZN(n17083) );
  OAI21_X1 U20286 ( .B1(n17084), .B2(n17096), .A(n17083), .ZN(P3_U2689) );
  AOI22_X1 U20287 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20288 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9795), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17087) );
  AOI22_X1 U20289 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10416), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20290 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17085) );
  NAND4_X1 U20291 ( .A1(n17088), .A2(n17087), .A3(n17086), .A4(n17085), .ZN(
        n17095) );
  AOI22_X1 U20292 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17093) );
  AOI22_X1 U20293 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U20294 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17091) );
  AOI22_X1 U20295 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17090) );
  NAND4_X1 U20296 ( .A1(n17093), .A2(n17092), .A3(n17091), .A4(n17090), .ZN(
        n17094) );
  NOR2_X1 U20297 ( .A1(n17095), .A2(n17094), .ZN(n17297) );
  NOR2_X1 U20298 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n9924), .ZN(n17097) );
  OAI22_X1 U20299 ( .A1(n17297), .A2(n9793), .B1(n17097), .B2(n17096), .ZN(
        P3_U2690) );
  NAND2_X1 U20300 ( .A1(n9793), .A2(n17108), .ZN(n17122) );
  AOI22_X1 U20301 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10416), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17107) );
  AOI22_X1 U20302 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17106) );
  AOI22_X1 U20303 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17098) );
  OAI21_X1 U20304 ( .B1(n10435), .B2(n21164), .A(n17098), .ZN(n17104) );
  AOI22_X1 U20305 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U20306 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U20307 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20308 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17099) );
  NAND4_X1 U20309 ( .A1(n17102), .A2(n17101), .A3(n17100), .A4(n17099), .ZN(
        n17103) );
  AOI211_X1 U20310 ( .C1(n9797), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17104), .B(n17103), .ZN(n17105) );
  NAND3_X1 U20311 ( .A1(n17107), .A2(n17106), .A3(n17105), .ZN(n17303) );
  NOR3_X1 U20312 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17248), .A3(n17108), .ZN(
        n17109) );
  AOI21_X1 U20313 ( .B1(n17193), .B2(n17303), .A(n17109), .ZN(n17110) );
  OAI21_X1 U20314 ( .B1(n17111), .B2(n17122), .A(n17110), .ZN(P3_U2691) );
  AOI22_X1 U20315 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10396), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20316 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20317 ( .A1(n16878), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17113) );
  AOI22_X1 U20318 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17112) );
  NAND4_X1 U20319 ( .A1(n17115), .A2(n17114), .A3(n17113), .A4(n17112), .ZN(
        n17121) );
  AOI22_X1 U20320 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U20321 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17118) );
  AOI22_X1 U20322 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17117) );
  AOI22_X1 U20323 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17116) );
  NAND4_X1 U20324 ( .A1(n17119), .A2(n17118), .A3(n17117), .A4(n17116), .ZN(
        n17120) );
  NOR2_X1 U20325 ( .A1(n17121), .A2(n17120), .ZN(n17307) );
  NOR2_X1 U20326 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17136), .ZN(n17123) );
  OAI22_X1 U20327 ( .A1(n17307), .A2(n9793), .B1(n17123), .B2(n17122), .ZN(
        P3_U2692) );
  OAI21_X1 U20328 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17124), .A(n9793), .ZN(
        n17135) );
  AOI22_X1 U20329 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20330 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20331 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10414), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20332 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17125) );
  NAND4_X1 U20333 ( .A1(n17128), .A2(n17127), .A3(n17126), .A4(n17125), .ZN(
        n17134) );
  AOI22_X1 U20334 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17132) );
  AOI22_X1 U20335 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9792), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20336 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20337 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17129) );
  NAND4_X1 U20338 ( .A1(n17132), .A2(n17131), .A3(n17130), .A4(n17129), .ZN(
        n17133) );
  NOR2_X1 U20339 ( .A1(n17134), .A2(n17133), .ZN(n17311) );
  OAI22_X1 U20340 ( .A1(n17136), .A2(n17135), .B1(n17311), .B2(n9793), .ZN(
        P3_U2693) );
  AOI22_X1 U20341 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17138), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20342 ( .A1(n9797), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20343 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n9795), .ZN(n17140) );
  AOI22_X1 U20344 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10414), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17162), .ZN(n17139) );
  NAND4_X1 U20345 ( .A1(n17142), .A2(n17141), .A3(n17140), .A4(n17139), .ZN(
        n17151) );
  AOI22_X1 U20346 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9792), .ZN(n17149) );
  AOI22_X1 U20347 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17143), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n9788), .ZN(n17148) );
  AOI22_X1 U20348 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17144), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U20349 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10396), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17146) );
  NAND4_X1 U20350 ( .A1(n17149), .A2(n17148), .A3(n17147), .A4(n17146), .ZN(
        n17150) );
  NOR2_X1 U20351 ( .A1(n17151), .A2(n17150), .ZN(n17316) );
  OAI21_X1 U20352 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17153), .A(n17152), .ZN(
        n17154) );
  AOI22_X1 U20353 ( .A1(n17193), .A2(n17316), .B1(n17154), .B2(n9793), .ZN(
        P3_U2694) );
  NAND2_X1 U20354 ( .A1(n9793), .A2(n17155), .ZN(n17179) );
  AOI22_X1 U20355 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17173) );
  AOI22_X1 U20356 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17172) );
  AOI22_X1 U20357 ( .A1(n16885), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17159) );
  OAI21_X1 U20358 ( .B1(n17160), .B2(n17207), .A(n17159), .ZN(n17170) );
  AOI22_X1 U20359 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17168) );
  AOI22_X1 U20360 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10565), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17167) );
  AOI22_X1 U20361 ( .A1(n9792), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17166) );
  AOI22_X1 U20362 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17165) );
  NAND4_X1 U20363 ( .A1(n17168), .A2(n17167), .A3(n17166), .A4(n17165), .ZN(
        n17169) );
  AOI211_X1 U20364 ( .C1(n9797), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n17170), .B(n17169), .ZN(n17171) );
  NAND3_X1 U20365 ( .A1(n17173), .A2(n17172), .A3(n17171), .ZN(n17319) );
  NOR2_X1 U20366 ( .A1(n17248), .A2(n9916), .ZN(n17181) );
  NOR3_X1 U20367 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17174), .A3(n10120), .ZN(
        n17175) );
  AOI22_X1 U20368 ( .A1(n17193), .A2(n17319), .B1(n17181), .B2(n17175), .ZN(
        n17176) );
  OAI21_X1 U20369 ( .B1(n17177), .B2(n17179), .A(n17176), .ZN(P3_U2695) );
  AOI21_X1 U20370 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17181), .A(
        P3_EBX_REG_7__SCAN_IN), .ZN(n17180) );
  INV_X1 U20371 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17178) );
  OAI22_X1 U20372 ( .A1(n17180), .A2(n17179), .B1(n17178), .B2(n9793), .ZN(
        P3_U2696) );
  NAND2_X1 U20373 ( .A1(n9793), .A2(n9916), .ZN(n17185) );
  AOI22_X1 U20374 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17193), .B1(
        n17181), .B2(n10120), .ZN(n17182) );
  OAI21_X1 U20375 ( .B1(n10120), .B2(n17185), .A(n17182), .ZN(P3_U2697) );
  AND2_X1 U20376 ( .A1(n17183), .A2(n17187), .ZN(n17186) );
  INV_X1 U20377 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17184) );
  OAI22_X1 U20378 ( .A1(n17186), .A2(n17185), .B1(n17184), .B2(n9793), .ZN(
        P3_U2698) );
  INV_X1 U20379 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17190) );
  OAI21_X1 U20380 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17188), .A(n17187), .ZN(
        n17189) );
  AOI22_X1 U20381 ( .A1(n17193), .A2(n17190), .B1(n17189), .B2(n9793), .ZN(
        P3_U2699) );
  NAND2_X1 U20382 ( .A1(n9793), .A2(n17191), .ZN(n17198) );
  NOR3_X1 U20383 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17248), .A3(n17191), .ZN(
        n17192) );
  AOI21_X1 U20384 ( .B1(n17193), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n17192), .ZN(n17194) );
  OAI21_X1 U20385 ( .B1(n17195), .B2(n17198), .A(n17194), .ZN(P3_U2700) );
  NOR2_X1 U20386 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17196), .ZN(n17199) );
  INV_X1 U20387 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17197) );
  OAI22_X1 U20388 ( .A1(n17199), .A2(n17198), .B1(n17197), .B2(n9793), .ZN(
        P3_U2701) );
  OAI222_X1 U20389 ( .A1(n17203), .A2(n17202), .B1(n17201), .B2(n9826), .C1(
        n17200), .C2(n9793), .ZN(P3_U2702) );
  OAI21_X1 U20390 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17205), .A(n17204), .ZN(
        n17206) );
  OAI21_X1 U20391 ( .B1(n9793), .B2(n17207), .A(n17206), .ZN(P3_U2703) );
  NAND2_X1 U20392 ( .A1(n18194), .A2(n17321), .ZN(n17254) );
  AOI22_X1 U20393 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17280), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17279), .ZN(n17211) );
  OAI211_X1 U20394 ( .C1(n17209), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17350), .B(
        n17208), .ZN(n17210) );
  OAI211_X1 U20395 ( .C1(n17212), .C2(n17345), .A(n17211), .B(n17210), .ZN(
        P3_U2705) );
  AOI22_X1 U20396 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17280), .B1(n17213), .B2(
        n17353), .ZN(n17216) );
  OAI211_X1 U20397 ( .C1(n17218), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17350), .B(
        n17214), .ZN(n17215) );
  OAI211_X1 U20398 ( .C1(n17250), .C2(n12820), .A(n17216), .B(n17215), .ZN(
        P3_U2706) );
  AOI22_X1 U20399 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17280), .B1(n17217), .B2(
        n17353), .ZN(n17221) );
  AOI211_X1 U20400 ( .C1(n17433), .C2(n17223), .A(n17218), .B(n17321), .ZN(
        n17219) );
  INV_X1 U20401 ( .A(n17219), .ZN(n17220) );
  OAI211_X1 U20402 ( .C1(n17250), .C2(n17222), .A(n17221), .B(n17220), .ZN(
        P3_U2707) );
  AOI22_X1 U20403 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17280), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17279), .ZN(n17225) );
  OAI211_X1 U20404 ( .C1(n17228), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17350), .B(
        n17223), .ZN(n17224) );
  OAI211_X1 U20405 ( .C1(n17345), .C2(n17226), .A(n17225), .B(n17224), .ZN(
        P3_U2708) );
  AOI22_X1 U20406 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17280), .B1(n17227), .B2(
        n17353), .ZN(n17231) );
  AOI211_X1 U20407 ( .C1(n17365), .C2(n17233), .A(n17228), .B(n17321), .ZN(
        n17229) );
  INV_X1 U20408 ( .A(n17229), .ZN(n17230) );
  OAI211_X1 U20409 ( .C1(n17250), .C2(n17232), .A(n17231), .B(n17230), .ZN(
        P3_U2709) );
  AOI22_X1 U20410 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17280), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17279), .ZN(n17236) );
  OAI211_X1 U20411 ( .C1(n17234), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17350), .B(
        n17233), .ZN(n17235) );
  OAI211_X1 U20412 ( .C1(n17345), .C2(n17237), .A(n17236), .B(n17235), .ZN(
        P3_U2710) );
  AOI22_X1 U20413 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17280), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17279), .ZN(n17241) );
  OAI211_X1 U20414 ( .C1(n17239), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17350), .B(
        n17238), .ZN(n17240) );
  OAI211_X1 U20415 ( .C1(n17345), .C2(n17242), .A(n17241), .B(n17240), .ZN(
        P3_U2711) );
  AOI22_X1 U20416 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17280), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17279), .ZN(n17246) );
  OAI211_X1 U20417 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17244), .A(n17350), .B(
        n17243), .ZN(n17245) );
  OAI211_X1 U20418 ( .C1(n17345), .C2(n17247), .A(n17246), .B(n17245), .ZN(
        P3_U2712) );
  INV_X1 U20419 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n21033) );
  NOR3_X1 U20420 ( .A1(n17248), .A2(n21033), .A3(n17281), .ZN(n17273) );
  NAND2_X1 U20421 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17273), .ZN(n17269) );
  NOR2_X1 U20422 ( .A1(n17249), .A2(n17269), .ZN(n17259) );
  NOR2_X1 U20423 ( .A1(n17321), .A2(n17259), .ZN(n17256) );
  INV_X1 U20424 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17372) );
  OAI22_X1 U20425 ( .A1(n17251), .A2(n17345), .B1(n18197), .B2(n17250), .ZN(
        n17252) );
  AOI221_X1 U20426 ( .B1(n17256), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17259), 
        .C2(n17372), .A(n17252), .ZN(n17253) );
  OAI21_X1 U20427 ( .B1(n18198), .B2(n17254), .A(n17253), .ZN(P3_U2713) );
  INV_X1 U20428 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17376) );
  INV_X1 U20429 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17378) );
  OR3_X1 U20430 ( .A1(n17376), .A2(n17378), .A3(n17269), .ZN(n17260) );
  AOI22_X1 U20431 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17279), .B1(n17353), .B2(
        n17255), .ZN(n17258) );
  AOI22_X1 U20432 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17280), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n17256), .ZN(n17257) );
  OAI211_X1 U20433 ( .C1(n17259), .C2(n17260), .A(n17258), .B(n17257), .ZN(
        P3_U2714) );
  AOI22_X1 U20434 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17280), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17279), .ZN(n17262) );
  NOR2_X1 U20435 ( .A1(n17378), .A2(n17269), .ZN(n17264) );
  OAI211_X1 U20436 ( .C1(n17264), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17350), .B(
        n17260), .ZN(n17261) );
  OAI211_X1 U20437 ( .C1(n17263), .C2(n17345), .A(n17262), .B(n17261), .ZN(
        P3_U2715) );
  AOI22_X1 U20438 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17280), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17279), .ZN(n17267) );
  AOI211_X1 U20439 ( .C1(n17378), .C2(n17269), .A(n17264), .B(n17321), .ZN(
        n17265) );
  INV_X1 U20440 ( .A(n17265), .ZN(n17266) );
  OAI211_X1 U20441 ( .C1(n17268), .C2(n17345), .A(n17267), .B(n17266), .ZN(
        P3_U2716) );
  AOI22_X1 U20442 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17280), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17279), .ZN(n17271) );
  OAI211_X1 U20443 ( .C1(n17273), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17350), .B(
        n17269), .ZN(n17270) );
  OAI211_X1 U20444 ( .C1(n17272), .C2(n17345), .A(n17271), .B(n17270), .ZN(
        P3_U2717) );
  AOI22_X1 U20445 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17280), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17279), .ZN(n17277) );
  INV_X1 U20446 ( .A(n17281), .ZN(n17275) );
  INV_X1 U20447 ( .A(n17273), .ZN(n17274) );
  OAI211_X1 U20448 ( .C1(n17275), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17350), .B(
        n17274), .ZN(n17276) );
  OAI211_X1 U20449 ( .C1(n17278), .C2(n17345), .A(n17277), .B(n17276), .ZN(
        P3_U2718) );
  AOI22_X1 U20450 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17280), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17279), .ZN(n17283) );
  OAI211_X1 U20451 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17285), .A(n17281), .B(
        n17350), .ZN(n17282) );
  OAI211_X1 U20452 ( .C1(n17284), .C2(n17345), .A(n17283), .B(n17282), .ZN(
        P3_U2719) );
  AOI211_X1 U20453 ( .C1(n17286), .C2(n17292), .A(n17321), .B(n17285), .ZN(
        n17287) );
  AOI21_X1 U20454 ( .B1(n17354), .B2(BUF2_REG_15__SCAN_IN), .A(n17287), .ZN(
        n17288) );
  OAI21_X1 U20455 ( .B1(n17289), .B2(n17345), .A(n17288), .ZN(P3_U2720) );
  INV_X1 U20456 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17455) );
  INV_X1 U20457 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17395) );
  NOR2_X1 U20458 ( .A1(n17290), .A2(n17324), .ZN(n17329) );
  NAND2_X1 U20459 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17329), .ZN(n17314) );
  NOR2_X1 U20460 ( .A1(n17395), .A2(n17314), .ZN(n17318) );
  NAND2_X1 U20461 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17318), .ZN(n17310) );
  NOR2_X1 U20462 ( .A1(n17455), .A2(n17310), .ZN(n17302) );
  NAND2_X1 U20463 ( .A1(n17302), .A2(n17463), .ZN(n17295) );
  AOI22_X1 U20464 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17354), .B1(n17353), .B2(
        n17291), .ZN(n17294) );
  NAND3_X1 U20465 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17350), .A3(n17292), 
        .ZN(n17293) );
  OAI211_X1 U20466 ( .C1(n17296), .C2(n17295), .A(n17294), .B(n17293), .ZN(
        P3_U2721) );
  NAND2_X1 U20467 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17302), .ZN(n17301) );
  NAND2_X1 U20468 ( .A1(n17301), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n17300) );
  INV_X1 U20469 ( .A(n17297), .ZN(n17298) );
  AOI22_X1 U20470 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17354), .B1(n17353), .B2(
        n17298), .ZN(n17299) );
  OAI221_X1 U20471 ( .B1(n17301), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n17300), 
        .C2(n17321), .A(n17299), .ZN(P3_U2722) );
  INV_X1 U20472 ( .A(n17301), .ZN(n17306) );
  AOI21_X1 U20473 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17350), .A(n17302), .ZN(
        n17305) );
  AOI22_X1 U20474 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17354), .B1(n17353), .B2(
        n17303), .ZN(n17304) );
  OAI21_X1 U20475 ( .B1(n17306), .B2(n17305), .A(n17304), .ZN(P3_U2723) );
  NAND2_X1 U20476 ( .A1(n17350), .A2(n17310), .ZN(n17313) );
  INV_X1 U20477 ( .A(n17307), .ZN(n17308) );
  AOI22_X1 U20478 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17354), .B1(n17353), .B2(
        n17308), .ZN(n17309) );
  OAI221_X1 U20479 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17310), .C1(n17455), 
        .C2(n17313), .A(n17309), .ZN(P3_U2724) );
  INV_X1 U20480 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17453) );
  NOR2_X1 U20481 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17318), .ZN(n17312) );
  OAI222_X1 U20482 ( .A1(n17348), .A2(n17453), .B1(n17313), .B2(n17312), .C1(
        n17345), .C2(n17311), .ZN(P3_U2725) );
  INV_X1 U20483 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17449) );
  OAI21_X1 U20484 ( .B1(n17395), .B2(n17321), .A(n17314), .ZN(n17315) );
  INV_X1 U20485 ( .A(n17315), .ZN(n17317) );
  OAI222_X1 U20486 ( .A1(n17348), .A2(n17449), .B1(n17318), .B2(n17317), .C1(
        n17345), .C2(n17316), .ZN(P3_U2726) );
  INV_X1 U20487 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17447) );
  AOI22_X1 U20488 ( .A1(n17353), .A2(n17319), .B1(n17329), .B2(n17397), .ZN(
        n17323) );
  OR3_X1 U20489 ( .A1(n17321), .A2(n17320), .A3(n17397), .ZN(n17322) );
  OAI211_X1 U20490 ( .C1(n17348), .C2(n17447), .A(n17323), .B(n17322), .ZN(
        P3_U2727) );
  NAND2_X1 U20491 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .ZN(n17325) );
  NOR2_X1 U20492 ( .A1(n17325), .A2(n17324), .ZN(n17357) );
  AND2_X1 U20493 ( .A1(n17326), .A2(n17357), .ZN(n17331) );
  AOI21_X1 U20494 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17350), .A(n17331), .ZN(
        n17328) );
  OAI222_X1 U20495 ( .A1(n17348), .A2(n18203), .B1(n17329), .B2(n17328), .C1(
        n17345), .C2(n17327), .ZN(P3_U2728) );
  INV_X1 U20496 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17404) );
  INV_X1 U20497 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17408) );
  NAND2_X1 U20498 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17357), .ZN(n17340) );
  NOR2_X1 U20499 ( .A1(n17408), .A2(n17340), .ZN(n17343) );
  NAND2_X1 U20500 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17343), .ZN(n17333) );
  NOR2_X1 U20501 ( .A1(n17404), .A2(n17333), .ZN(n17335) );
  AOI21_X1 U20502 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17350), .A(n17335), .ZN(
        n17332) );
  OAI222_X1 U20503 ( .A1(n17348), .A2(n18198), .B1(n17332), .B2(n17331), .C1(
        n17345), .C2(n17330), .ZN(P3_U2729) );
  INV_X1 U20504 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21119) );
  INV_X1 U20505 ( .A(n17333), .ZN(n17339) );
  AOI21_X1 U20506 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17350), .A(n17339), .ZN(
        n17336) );
  OAI222_X1 U20507 ( .A1(n17348), .A2(n21119), .B1(n17336), .B2(n17335), .C1(
        n17345), .C2(n17334), .ZN(P3_U2730) );
  AOI21_X1 U20508 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17350), .A(n17343), .ZN(
        n17338) );
  OAI222_X1 U20509 ( .A1(n18189), .A2(n17348), .B1(n17339), .B2(n17338), .C1(
        n17345), .C2(n17337), .ZN(P3_U2731) );
  INV_X1 U20510 ( .A(n17340), .ZN(n17347) );
  AOI21_X1 U20511 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17350), .A(n17347), .ZN(
        n17342) );
  OAI222_X1 U20512 ( .A1(n18184), .A2(n17348), .B1(n17343), .B2(n17342), .C1(
        n17345), .C2(n17341), .ZN(P3_U2732) );
  AOI21_X1 U20513 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17350), .A(n17357), .ZN(
        n17346) );
  OAI222_X1 U20514 ( .A1(n18180), .A2(n17348), .B1(n17347), .B2(n17346), .C1(
        n17345), .C2(n17344), .ZN(P3_U2733) );
  NOR2_X1 U20515 ( .A1(n17415), .A2(n17349), .ZN(n17351) );
  OAI21_X1 U20516 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17351), .A(n17350), .ZN(
        n17356) );
  AOI22_X1 U20517 ( .A1(n17354), .A2(BUF2_REG_1__SCAN_IN), .B1(n17353), .B2(
        n17352), .ZN(n17355) );
  OAI21_X1 U20518 ( .B1(n17357), .B2(n17356), .A(n17355), .ZN(P3_U2734) );
  NAND2_X1 U20519 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17675), .ZN(n17388) );
  NOR2_X1 U20520 ( .A1(n17385), .A2(n17359), .ZN(P3_U2736) );
  INV_X1 U20521 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n21082) );
  NOR2_X1 U20522 ( .A1(n17414), .A2(n18172), .ZN(n17383) );
  INV_X2 U20523 ( .A(n17388), .ZN(n17412) );
  AOI22_X1 U20524 ( .A1(n17412), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17360) );
  OAI21_X1 U20525 ( .B1(n21082), .B2(n17382), .A(n17360), .ZN(P3_U2737) );
  INV_X1 U20526 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17435) );
  AOI22_X1 U20527 ( .A1(n17412), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17361) );
  OAI21_X1 U20528 ( .B1(n17435), .B2(n17382), .A(n17361), .ZN(P3_U2738) );
  AOI22_X1 U20529 ( .A1(n17412), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17362) );
  OAI21_X1 U20530 ( .B1(n17433), .B2(n17382), .A(n17362), .ZN(P3_U2739) );
  INV_X1 U20531 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17431) );
  AOI22_X1 U20532 ( .A1(n17412), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17363) );
  OAI21_X1 U20533 ( .B1(n17431), .B2(n17382), .A(n17363), .ZN(P3_U2740) );
  AOI22_X1 U20534 ( .A1(n17412), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17364) );
  OAI21_X1 U20535 ( .B1(n17365), .B2(n17382), .A(n17364), .ZN(P3_U2741) );
  INV_X1 U20536 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17367) );
  AOI22_X1 U20537 ( .A1(n17412), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17366) );
  OAI21_X1 U20538 ( .B1(n17367), .B2(n17382), .A(n17366), .ZN(P3_U2742) );
  INV_X1 U20539 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U20540 ( .A1(n17412), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17368) );
  OAI21_X1 U20541 ( .B1(n17369), .B2(n17382), .A(n17368), .ZN(P3_U2743) );
  INV_X1 U20542 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n21060) );
  AOI22_X1 U20543 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17383), .B1(n17412), 
        .B2(P3_UWORD_REG_7__SCAN_IN), .ZN(n17370) );
  OAI21_X1 U20544 ( .B1(n21060), .B2(n17385), .A(n17370), .ZN(P3_U2744) );
  AOI22_X1 U20545 ( .A1(n17412), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17371) );
  OAI21_X1 U20546 ( .B1(n17372), .B2(n17382), .A(n17371), .ZN(P3_U2745) );
  INV_X1 U20547 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17374) );
  AOI22_X1 U20548 ( .A1(n17412), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17373) );
  OAI21_X1 U20549 ( .B1(n17374), .B2(n17382), .A(n17373), .ZN(P3_U2746) );
  AOI22_X1 U20550 ( .A1(n17412), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17375) );
  OAI21_X1 U20551 ( .B1(n17376), .B2(n17382), .A(n17375), .ZN(P3_U2747) );
  AOI22_X1 U20552 ( .A1(n17412), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17377) );
  OAI21_X1 U20553 ( .B1(n17378), .B2(n17382), .A(n17377), .ZN(P3_U2748) );
  INV_X1 U20554 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17380) );
  AOI22_X1 U20555 ( .A1(n17412), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17379) );
  OAI21_X1 U20556 ( .B1(n17380), .B2(n17382), .A(n17379), .ZN(P3_U2749) );
  AOI22_X1 U20557 ( .A1(n17412), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17381) );
  OAI21_X1 U20558 ( .B1(n21033), .B2(n17382), .A(n17381), .ZN(P3_U2750) );
  INV_X1 U20559 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n20949) );
  AOI22_X1 U20560 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17383), .B1(n17412), 
        .B2(P3_UWORD_REG_0__SCAN_IN), .ZN(n17384) );
  OAI21_X1 U20561 ( .B1(n20949), .B2(n17385), .A(n17384), .ZN(P3_U2751) );
  INV_X1 U20562 ( .A(P3_LWORD_REG_15__SCAN_IN), .ZN(n20958) );
  INV_X1 U20563 ( .A(n17414), .ZN(n17386) );
  AOI22_X1 U20564 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n17386), .B1(n17402), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17387) );
  OAI21_X1 U20565 ( .B1(n20958), .B2(n17388), .A(n17387), .ZN(P3_U2752) );
  AOI22_X1 U20566 ( .A1(n17412), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17389) );
  OAI21_X1 U20567 ( .B1(n17463), .B2(n17414), .A(n17389), .ZN(P3_U2753) );
  INV_X1 U20568 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U20569 ( .A1(n17412), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17390) );
  OAI21_X1 U20570 ( .B1(n17460), .B2(n17414), .A(n17390), .ZN(P3_U2754) );
  INV_X1 U20571 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17458) );
  AOI22_X1 U20572 ( .A1(n17412), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17391) );
  OAI21_X1 U20573 ( .B1(n17458), .B2(n17414), .A(n17391), .ZN(P3_U2755) );
  AOI22_X1 U20574 ( .A1(n17412), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17392) );
  OAI21_X1 U20575 ( .B1(n17455), .B2(n17414), .A(n17392), .ZN(P3_U2756) );
  AOI22_X1 U20576 ( .A1(n17412), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17393) );
  OAI21_X1 U20577 ( .B1(n21142), .B2(n17414), .A(n17393), .ZN(P3_U2757) );
  AOI22_X1 U20578 ( .A1(n17412), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17394) );
  OAI21_X1 U20579 ( .B1(n17395), .B2(n17414), .A(n17394), .ZN(P3_U2758) );
  AOI22_X1 U20580 ( .A1(n17412), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17396) );
  OAI21_X1 U20581 ( .B1(n17397), .B2(n17414), .A(n17396), .ZN(P3_U2759) );
  INV_X1 U20582 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U20583 ( .A1(n17412), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17398) );
  OAI21_X1 U20584 ( .B1(n17399), .B2(n17414), .A(n17398), .ZN(P3_U2760) );
  INV_X1 U20585 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17401) );
  AOI22_X1 U20586 ( .A1(n17412), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17400) );
  OAI21_X1 U20587 ( .B1(n17401), .B2(n17414), .A(n17400), .ZN(P3_U2761) );
  AOI22_X1 U20588 ( .A1(n17412), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17403) );
  OAI21_X1 U20589 ( .B1(n17404), .B2(n17414), .A(n17403), .ZN(P3_U2762) );
  AOI22_X1 U20590 ( .A1(n17412), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17405) );
  OAI21_X1 U20591 ( .B1(n17406), .B2(n17414), .A(n17405), .ZN(P3_U2763) );
  AOI22_X1 U20592 ( .A1(n17412), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17407) );
  OAI21_X1 U20593 ( .B1(n17408), .B2(n17414), .A(n17407), .ZN(P3_U2764) );
  INV_X1 U20594 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U20595 ( .A1(n17412), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17409) );
  OAI21_X1 U20596 ( .B1(n17410), .B2(n17414), .A(n17409), .ZN(P3_U2765) );
  INV_X1 U20597 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17439) );
  AOI22_X1 U20598 ( .A1(n17412), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17411) );
  OAI21_X1 U20599 ( .B1(n17439), .B2(n17414), .A(n17411), .ZN(P3_U2766) );
  AOI22_X1 U20600 ( .A1(n17412), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17402), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17413) );
  OAI21_X1 U20601 ( .B1(n17415), .B2(n17414), .A(n17413), .ZN(P3_U2767) );
  OAI211_X1 U20602 ( .C1(n18814), .C2(n18813), .A(n17417), .B(n17416), .ZN(
        n17456) );
  AOI22_X1 U20603 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17450), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17465), .ZN(n17419) );
  OAI21_X1 U20604 ( .B1(n18167), .B2(n17452), .A(n17419), .ZN(P3_U2768) );
  AOI22_X1 U20605 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17464), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17465), .ZN(n17420) );
  OAI21_X1 U20606 ( .B1(n21033), .B2(n17462), .A(n17420), .ZN(P3_U2769) );
  AOI22_X1 U20607 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17450), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17465), .ZN(n17421) );
  OAI21_X1 U20608 ( .B1(n18180), .B2(n17452), .A(n17421), .ZN(P3_U2770) );
  AOI22_X1 U20609 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17450), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17465), .ZN(n17422) );
  OAI21_X1 U20610 ( .B1(n18184), .B2(n17452), .A(n17422), .ZN(P3_U2771) );
  AOI22_X1 U20611 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17450), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17465), .ZN(n17423) );
  OAI21_X1 U20612 ( .B1(n18189), .B2(n17452), .A(n17423), .ZN(P3_U2772) );
  AOI22_X1 U20613 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17450), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17465), .ZN(n17424) );
  OAI21_X1 U20614 ( .B1(n21119), .B2(n17452), .A(n17424), .ZN(P3_U2773) );
  AOI22_X1 U20615 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17450), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17465), .ZN(n17425) );
  OAI21_X1 U20616 ( .B1(n18198), .B2(n17452), .A(n17425), .ZN(P3_U2774) );
  AOI22_X1 U20617 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17450), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17465), .ZN(n17426) );
  OAI21_X1 U20618 ( .B1(n18203), .B2(n17452), .A(n17426), .ZN(P3_U2775) );
  AOI22_X1 U20619 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17450), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17465), .ZN(n17427) );
  OAI21_X1 U20620 ( .B1(n17447), .B2(n17452), .A(n17427), .ZN(P3_U2776) );
  AOI22_X1 U20621 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17450), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17465), .ZN(n17428) );
  OAI21_X1 U20622 ( .B1(n17449), .B2(n17452), .A(n17428), .ZN(P3_U2777) );
  AOI22_X1 U20623 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17450), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17465), .ZN(n17429) );
  OAI21_X1 U20624 ( .B1(n17453), .B2(n17452), .A(n17429), .ZN(P3_U2778) );
  AOI22_X1 U20625 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17464), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17465), .ZN(n17430) );
  OAI21_X1 U20626 ( .B1(n17431), .B2(n17462), .A(n17430), .ZN(P3_U2779) );
  AOI22_X1 U20627 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17464), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17465), .ZN(n17432) );
  OAI21_X1 U20628 ( .B1(n17433), .B2(n17462), .A(n17432), .ZN(P3_U2780) );
  AOI22_X1 U20629 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17464), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17465), .ZN(n17434) );
  OAI21_X1 U20630 ( .B1(n17435), .B2(n17462), .A(n17434), .ZN(P3_U2781) );
  AOI22_X1 U20631 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17464), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17465), .ZN(n17436) );
  OAI21_X1 U20632 ( .B1(n21082), .B2(n17462), .A(n17436), .ZN(P3_U2782) );
  AOI22_X1 U20633 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17450), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17465), .ZN(n17437) );
  OAI21_X1 U20634 ( .B1(n18167), .B2(n17452), .A(n17437), .ZN(P3_U2783) );
  AOI22_X1 U20635 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17465), .ZN(n17438) );
  OAI21_X1 U20636 ( .B1(n17439), .B2(n17462), .A(n17438), .ZN(P3_U2784) );
  AOI22_X1 U20637 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17450), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17465), .ZN(n17440) );
  OAI21_X1 U20638 ( .B1(n18180), .B2(n17452), .A(n17440), .ZN(P3_U2785) );
  AOI22_X1 U20639 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17450), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17456), .ZN(n17441) );
  OAI21_X1 U20640 ( .B1(n18184), .B2(n17452), .A(n17441), .ZN(P3_U2786) );
  AOI22_X1 U20641 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17450), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17456), .ZN(n17442) );
  OAI21_X1 U20642 ( .B1(n18189), .B2(n17452), .A(n17442), .ZN(P3_U2787) );
  AOI22_X1 U20643 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17450), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17456), .ZN(n17443) );
  OAI21_X1 U20644 ( .B1(n21119), .B2(n17452), .A(n17443), .ZN(P3_U2788) );
  AOI22_X1 U20645 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17450), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17456), .ZN(n17444) );
  OAI21_X1 U20646 ( .B1(n18198), .B2(n17452), .A(n17444), .ZN(P3_U2789) );
  AOI22_X1 U20647 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17450), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17456), .ZN(n17445) );
  OAI21_X1 U20648 ( .B1(n18203), .B2(n17452), .A(n17445), .ZN(P3_U2790) );
  AOI22_X1 U20649 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17450), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17456), .ZN(n17446) );
  OAI21_X1 U20650 ( .B1(n17447), .B2(n17452), .A(n17446), .ZN(P3_U2791) );
  AOI22_X1 U20651 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17450), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17456), .ZN(n17448) );
  OAI21_X1 U20652 ( .B1(n17449), .B2(n17452), .A(n17448), .ZN(P3_U2792) );
  AOI22_X1 U20653 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17450), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17456), .ZN(n17451) );
  OAI21_X1 U20654 ( .B1(n17453), .B2(n17452), .A(n17451), .ZN(P3_U2793) );
  AOI22_X1 U20655 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17456), .ZN(n17454) );
  OAI21_X1 U20656 ( .B1(n17455), .B2(n17462), .A(n17454), .ZN(P3_U2794) );
  AOI22_X1 U20657 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17456), .ZN(n17457) );
  OAI21_X1 U20658 ( .B1(n17458), .B2(n17462), .A(n17457), .ZN(P3_U2795) );
  AOI22_X1 U20659 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17465), .ZN(n17459) );
  OAI21_X1 U20660 ( .B1(n17460), .B2(n17462), .A(n17459), .ZN(P3_U2796) );
  AOI22_X1 U20661 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17465), .ZN(n17461) );
  OAI21_X1 U20662 ( .B1(n17463), .B2(n17462), .A(n17461), .ZN(P3_U2797) );
  INV_X1 U20663 ( .A(n17466), .ZN(P3_U2798) );
  NAND2_X1 U20664 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17467), .ZN(
        n17487) );
  AOI21_X1 U20665 ( .B1(n17469), .B2(n17468), .A(n17733), .ZN(n17484) );
  NOR2_X1 U20666 ( .A1(n17694), .A2(n17477), .ZN(n17495) );
  OAI211_X1 U20667 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17495), .B(n17471), .ZN(n17473) );
  NAND2_X1 U20668 ( .A1(n9790), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17472) );
  OAI211_X1 U20669 ( .C1(n17696), .C2(n17474), .A(n17473), .B(n17472), .ZN(
        n17481) );
  OAI21_X1 U20670 ( .B1(n17475), .B2(n17846), .A(n17845), .ZN(n17476) );
  AOI21_X1 U20671 ( .B1(n17803), .B2(n17477), .A(n17476), .ZN(n17513) );
  OAI21_X1 U20672 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17564), .A(
        n17513), .ZN(n17489) );
  INV_X1 U20673 ( .A(n17489), .ZN(n17479) );
  INV_X1 U20674 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17478) );
  NOR2_X1 U20675 ( .A1(n17479), .A2(n17478), .ZN(n17480) );
  AOI22_X1 U20676 ( .A1(n17834), .A2(n17858), .B1(n17715), .B2(n17855), .ZN(
        n17508) );
  NAND2_X1 U20677 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17508), .ZN(
        n17497) );
  OAI211_X1 U20678 ( .C1(n17834), .C2(n17715), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17497), .ZN(n17485) );
  OAI211_X1 U20679 ( .C1(n17496), .C2(n17487), .A(n17486), .B(n17485), .ZN(
        P3_U2802) );
  AOI22_X1 U20680 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17489), .B1(
        n17604), .B2(n17488), .ZN(n17501) );
  INV_X1 U20681 ( .A(n17490), .ZN(n17492) );
  NAND2_X1 U20682 ( .A1(n17492), .A2(n17491), .ZN(n17493) );
  XOR2_X1 U20683 ( .A(n17754), .B(n17493), .Z(n17866) );
  AOI22_X1 U20684 ( .A1(n17755), .A2(n17866), .B1(n17495), .B2(n17494), .ZN(
        n17500) );
  INV_X1 U20685 ( .A(n17496), .ZN(n17498) );
  OAI21_X1 U20686 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17498), .A(
        n17497), .ZN(n17499) );
  NAND2_X1 U20687 ( .A1(n9790), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17867) );
  NAND4_X1 U20688 ( .A1(n17501), .A2(n17500), .A3(n17499), .A4(n17867), .ZN(
        P3_U2803) );
  AOI21_X1 U20689 ( .B1(n18552), .B2(n17502), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17512) );
  NAND2_X1 U20690 ( .A1(n17696), .A2(n17564), .ZN(n17837) );
  AOI22_X1 U20691 ( .A1(n9790), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n17503), 
        .B2(n17837), .ZN(n17511) );
  INV_X1 U20692 ( .A(n17633), .ZN(n17647) );
  NOR2_X1 U20693 ( .A1(n17523), .A2(n17647), .ZN(n17541) );
  NAND2_X1 U20694 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17514) );
  NOR2_X1 U20695 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17514), .ZN(
        n17870) );
  AOI21_X1 U20696 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17506), .A(
        n17505), .ZN(n17877) );
  OAI22_X1 U20697 ( .A1(n17508), .A2(n17507), .B1(n17877), .B2(n17733), .ZN(
        n17509) );
  AOI21_X1 U20698 ( .B1(n17541), .B2(n17870), .A(n17509), .ZN(n17510) );
  OAI211_X1 U20699 ( .C1(n17513), .C2(n17512), .A(n17511), .B(n17510), .ZN(
        P3_U2804) );
  INV_X1 U20700 ( .A(n17982), .ZN(n17915) );
  NOR2_X1 U20701 ( .A1(n17893), .A2(n17899), .ZN(n17515) );
  OAI22_X1 U20702 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17515), .B1(
        n17514), .B2(n17899), .ZN(n17888) );
  AOI22_X1 U20703 ( .A1(n18552), .A2(n17517), .B1(n17675), .B2(n17516), .ZN(
        n17518) );
  NAND2_X1 U20704 ( .A1(n17518), .A2(n17845), .ZN(n17553) );
  AOI21_X1 U20705 ( .B1(n17675), .B2(n17519), .A(n17553), .ZN(n17539) );
  AND2_X1 U20706 ( .A1(n17678), .A2(n9893), .ZN(n17578) );
  NAND2_X1 U20707 ( .A1(n17567), .A2(n17578), .ZN(n17550) );
  NOR2_X1 U20708 ( .A1(n17519), .A2(n17550), .ZN(n17534) );
  OAI211_X1 U20709 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17534), .B(n17520), .ZN(n17521) );
  NAND2_X1 U20710 ( .A1(n9790), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17890) );
  OAI211_X1 U20711 ( .C1(n17539), .C2(n17522), .A(n17521), .B(n17890), .ZN(
        n17529) );
  NOR2_X1 U20712 ( .A1(n17988), .A2(n17523), .ZN(n17896) );
  NAND2_X1 U20713 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17896), .ZN(
        n17524) );
  XOR2_X1 U20714 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17524), .Z(
        n17885) );
  OAI21_X1 U20715 ( .B1(n17685), .B2(n17526), .A(n17525), .ZN(n17527) );
  XOR2_X1 U20716 ( .A(n17527), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17892) );
  OAI22_X1 U20717 ( .A1(n17850), .A2(n17885), .B1(n17733), .B2(n17892), .ZN(
        n17528) );
  AOI211_X1 U20718 ( .C1(n17604), .C2(n17530), .A(n17529), .B(n17528), .ZN(
        n17531) );
  OAI21_X1 U20719 ( .B1(n17759), .B2(n17888), .A(n17531), .ZN(P3_U2805) );
  OAI21_X1 U20720 ( .B1(n17533), .B2(n17893), .A(n17532), .ZN(n17895) );
  INV_X1 U20721 ( .A(n17895), .ZN(n17543) );
  NAND2_X1 U20722 ( .A1(n17899), .A2(n17715), .ZN(n17544) );
  OAI21_X1 U20723 ( .B1(n17896), .B2(n17850), .A(n17544), .ZN(n17558) );
  AOI22_X1 U20724 ( .A1(n17535), .A2(n17604), .B1(n17534), .B2(n17538), .ZN(
        n17537) );
  NAND2_X1 U20725 ( .A1(n9790), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17536) );
  OAI211_X1 U20726 ( .C1(n17539), .C2(n17538), .A(n17537), .B(n17536), .ZN(
        n17540) );
  AOI221_X1 U20727 ( .B1(n17541), .B2(n17893), .C1(n17558), .C2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n17540), .ZN(n17542) );
  OAI21_X1 U20728 ( .B1(n17543), .B2(n17733), .A(n17542), .ZN(P3_U2806) );
  NOR2_X1 U20729 ( .A1(n17896), .A2(n17850), .ZN(n17546) );
  INV_X1 U20730 ( .A(n17544), .ZN(n17545) );
  AOI22_X1 U20731 ( .A1(n17547), .A2(n17546), .B1(n17982), .B2(n17545), .ZN(
        n17561) );
  NAND2_X1 U20732 ( .A1(n9790), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17911) );
  INV_X1 U20733 ( .A(n17911), .ZN(n17552) );
  INV_X1 U20734 ( .A(n17548), .ZN(n17549) );
  OAI22_X1 U20735 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17550), .B1(
        n17549), .B2(n17696), .ZN(n17551) );
  AOI211_X1 U20736 ( .C1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n17553), .A(
        n17552), .B(n17551), .ZN(n17560) );
  OAI22_X1 U20737 ( .A1(n17754), .A2(n17930), .B1(n17569), .B2(n17554), .ZN(
        n17556) );
  NOR2_X1 U20738 ( .A1(n17556), .A2(n17555), .ZN(n17557) );
  XOR2_X1 U20739 ( .A(n17557), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n17910) );
  AOI22_X1 U20740 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17558), .B1(
        n17755), .B2(n17910), .ZN(n17559) );
  OAI211_X1 U20741 ( .C1(n17561), .C2(n17853), .A(n17560), .B(n17559), .ZN(
        P3_U2807) );
  INV_X1 U20742 ( .A(n17803), .ZN(n17817) );
  OAI21_X1 U20743 ( .B1(n9893), .B2(n17817), .A(n17845), .ZN(n17562) );
  AOI21_X1 U20744 ( .B1(n17675), .B2(n17563), .A(n17562), .ZN(n17587) );
  OAI21_X1 U20745 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17564), .A(
        n17587), .ZN(n17576) );
  OAI21_X1 U20746 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17578), .ZN(n17566) );
  OAI22_X1 U20747 ( .A1(n17567), .A2(n17566), .B1(n17565), .B2(n17696), .ZN(
        n17568) );
  AOI21_X1 U20748 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17576), .A(
        n17568), .ZN(n17573) );
  NOR2_X1 U20749 ( .A1(n17834), .A2(n17715), .ZN(n17593) );
  NOR2_X1 U20750 ( .A1(n17620), .A2(n17914), .ZN(n17919) );
  AOI22_X1 U20751 ( .A1(n17834), .A2(n17988), .B1(n17715), .B2(n17915), .ZN(
        n17646) );
  OAI21_X1 U20752 ( .B1(n17593), .B2(n17919), .A(n17646), .ZN(n17584) );
  OAI221_X1 U20753 ( .B1(n17569), .B2(n17637), .C1(n17569), .C2(n17919), .A(
        n10475), .ZN(n17570) );
  XOR2_X1 U20754 ( .A(n17930), .B(n17570), .Z(n17927) );
  AOI22_X1 U20755 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17584), .B1(
        n17755), .B2(n17927), .ZN(n17572) );
  NAND2_X1 U20756 ( .A1(n9790), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17928) );
  NAND3_X1 U20757 ( .A1(n17633), .A2(n17919), .A3(n17930), .ZN(n17571) );
  NAND4_X1 U20758 ( .A1(n17573), .A2(n17572), .A3(n17928), .A4(n17571), .ZN(
        P3_U2808) );
  OR2_X1 U20759 ( .A1(n17582), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17943) );
  NOR2_X1 U20760 ( .A1(n17620), .A2(n17623), .ZN(n17933) );
  NAND2_X1 U20761 ( .A1(n17633), .A2(n17933), .ZN(n17610) );
  OAI22_X1 U20762 ( .A1(n9796), .A2(n18737), .B1(n17696), .B2(n16448), .ZN(
        n17575) );
  AOI221_X1 U20763 ( .B1(n17578), .B2(n17577), .C1(n17576), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17575), .ZN(n17586) );
  NAND3_X1 U20764 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17754), .A3(
        n17579), .ZN(n17605) );
  INV_X1 U20765 ( .A(n17580), .ZN(n17618) );
  OAI22_X1 U20766 ( .A1(n17582), .A2(n17605), .B1(n17581), .B2(n17618), .ZN(
        n17583) );
  XOR2_X1 U20767 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17583), .Z(
        n17932) );
  AOI22_X1 U20768 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17584), .B1(
        n17755), .B2(n17932), .ZN(n17585) );
  OAI211_X1 U20769 ( .C1(n17943), .C2(n17610), .A(n17586), .B(n17585), .ZN(
        P3_U2809) );
  NAND2_X1 U20770 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21062), .ZN(
        n17950) );
  AOI221_X1 U20771 ( .B1(n17589), .B2(n17588), .C1(n18464), .C2(n17588), .A(
        n17587), .ZN(n17591) );
  NOR2_X1 U20772 ( .A1(n9796), .A2(n18736), .ZN(n17590) );
  AOI211_X1 U20773 ( .C1(n17592), .C2(n17837), .A(n17591), .B(n17590), .ZN(
        n17597) );
  NAND2_X1 U20774 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17933), .ZN(
        n17916) );
  INV_X1 U20775 ( .A(n17916), .ZN(n17945) );
  OAI21_X1 U20776 ( .B1(n17593), .B2(n17945), .A(n17646), .ZN(n17607) );
  INV_X1 U20777 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17594) );
  AOI221_X1 U20778 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17605), 
        .C1(n17594), .C2(n17617), .A(n17555), .ZN(n17595) );
  XOR2_X1 U20779 ( .A(n17595), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n17944) );
  AOI22_X1 U20780 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17607), .B1(
        n17755), .B2(n17944), .ZN(n17596) );
  OAI211_X1 U20781 ( .C1(n17950), .C2(n17610), .A(n17597), .B(n17596), .ZN(
        P3_U2810) );
  OAI21_X1 U20782 ( .B1(n17599), .B2(n17817), .A(n17845), .ZN(n17626) );
  AOI21_X1 U20783 ( .B1(n17675), .B2(n17598), .A(n17626), .ZN(n17613) );
  AND2_X1 U20784 ( .A1(n17678), .A2(n17599), .ZN(n17616) );
  OAI221_X1 U20785 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(n21027), .C2(n17601), .A(
        n17616), .ZN(n17600) );
  NAND2_X1 U20786 ( .A1(n9790), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17953) );
  OAI211_X1 U20787 ( .C1(n17613), .C2(n17601), .A(n17600), .B(n17953), .ZN(
        n17602) );
  AOI21_X1 U20788 ( .B1(n17604), .B2(n17603), .A(n17602), .ZN(n17609) );
  OAI21_X1 U20789 ( .B1(n17617), .B2(n17618), .A(n17605), .ZN(n17606) );
  XOR2_X1 U20790 ( .A(n17606), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n17951) );
  AOI22_X1 U20791 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17607), .B1(
        n17755), .B2(n17951), .ZN(n17608) );
  OAI211_X1 U20792 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17610), .A(
        n17609), .B(n17608), .ZN(P3_U2811) );
  INV_X1 U20793 ( .A(n17646), .ZN(n17611) );
  AOI21_X1 U20794 ( .B1(n17633), .B2(n17620), .A(n17611), .ZN(n17631) );
  NOR2_X1 U20795 ( .A1(n9796), .A2(n21167), .ZN(n17615) );
  OAI22_X1 U20796 ( .A1(n17613), .A2(n21027), .B1(n17696), .B2(n17612), .ZN(
        n17614) );
  AOI211_X1 U20797 ( .C1(n17616), .C2(n21027), .A(n17615), .B(n17614), .ZN(
        n17622) );
  OAI21_X1 U20798 ( .B1(n17623), .B2(n17685), .A(n17617), .ZN(n17619) );
  XOR2_X1 U20799 ( .A(n17619), .B(n17618), .Z(n17969) );
  NOR2_X1 U20800 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17620), .ZN(
        n17968) );
  AOI22_X1 U20801 ( .A1(n17755), .A2(n17969), .B1(n17633), .B2(n17968), .ZN(
        n17621) );
  OAI211_X1 U20802 ( .C1(n17631), .C2(n17623), .A(n17622), .B(n17621), .ZN(
        P3_U2812) );
  INV_X1 U20803 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18731) );
  OAI21_X1 U20804 ( .B1(n18464), .B2(n17624), .A(n21007), .ZN(n17625) );
  AOI22_X1 U20805 ( .A1(n17627), .A2(n17837), .B1(n17626), .B2(n17625), .ZN(
        n17635) );
  NOR2_X1 U20806 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17978), .ZN(
        n21220) );
  AOI21_X1 U20807 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17630), .A(
        n17629), .ZN(n21224) );
  OAI22_X1 U20808 ( .A1(n21224), .A2(n17733), .B1(n17631), .B2(n17963), .ZN(
        n17632) );
  AOI21_X1 U20809 ( .B1(n17633), .B2(n21220), .A(n17632), .ZN(n17634) );
  OAI211_X1 U20810 ( .C1(n9796), .C2(n18731), .A(n17635), .B(n17634), .ZN(
        P3_U2813) );
  OAI21_X1 U20811 ( .B1(n17685), .B2(n17637), .A(n17636), .ZN(n17638) );
  XOR2_X1 U20812 ( .A(n17638), .B(n17978), .Z(n17979) );
  AOI21_X1 U20813 ( .B1(n17803), .B2(n9891), .A(n17818), .ZN(n17662) );
  OAI21_X1 U20814 ( .B1(n17639), .B2(n17846), .A(n17662), .ZN(n17650) );
  AOI22_X1 U20815 ( .A1(n9790), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17650), .ZN(n17642) );
  NOR2_X1 U20816 ( .A1(n17694), .A2(n9891), .ZN(n17652) );
  OAI211_X1 U20817 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17652), .B(n17640), .ZN(n17641) );
  OAI211_X1 U20818 ( .C1(n17643), .C2(n17696), .A(n17642), .B(n17641), .ZN(
        n17644) );
  AOI21_X1 U20819 ( .B1(n17755), .B2(n17979), .A(n17644), .ZN(n17645) );
  OAI221_X1 U20820 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17647), 
        .C1(n17978), .C2(n17646), .A(n17645), .ZN(P3_U2814) );
  INV_X1 U20821 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17651) );
  NAND2_X1 U20822 ( .A1(n9790), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17995) );
  OAI21_X1 U20823 ( .B1(n17696), .B2(n17648), .A(n17995), .ZN(n17649) );
  AOI221_X1 U20824 ( .B1(n17652), .B2(n17651), .C1(n17650), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17649), .ZN(n17660) );
  NOR2_X1 U20825 ( .A1(n17702), .A2(n17653), .ZN(n17686) );
  NOR4_X1 U20826 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n17754), .A4(n17735), .ZN(
        n17713) );
  INV_X1 U20827 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17717) );
  NAND2_X1 U20828 ( .A1(n17713), .A2(n17717), .ZN(n17701) );
  NOR2_X1 U20829 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17701), .ZN(
        n17668) );
  AOI21_X1 U20830 ( .B1(n17654), .B2(n17686), .A(n17668), .ZN(n17655) );
  AOI221_X1 U20831 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18032), 
        .C1(n17685), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17655), .ZN(
        n17656) );
  XOR2_X1 U20832 ( .A(n17656), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n17994) );
  NOR2_X1 U20833 ( .A1(n17982), .A2(n17759), .ZN(n17657) );
  NAND2_X1 U20834 ( .A1(n17989), .A2(n17661), .ZN(n17985) );
  AOI22_X1 U20835 ( .A1(n17755), .A2(n17994), .B1(n17657), .B2(n17985), .ZN(
        n17659) );
  OAI211_X1 U20836 ( .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n17667), .A(
        n17834), .B(n17988), .ZN(n17658) );
  NAND3_X1 U20837 ( .A1(n17660), .A2(n17659), .A3(n17658), .ZN(P3_U2815) );
  OAI221_X1 U20838 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18016), .A(n17661), .ZN(
        n18003) );
  INV_X1 U20839 ( .A(n17693), .ZN(n17679) );
  NAND2_X1 U20840 ( .A1(n18552), .A2(n17679), .ZN(n17712) );
  AOI221_X1 U20841 ( .B1(n17664), .B2(n17663), .C1(n17712), .C2(n17663), .A(
        n17662), .ZN(n17665) );
  NOR2_X1 U20842 ( .A1(n9796), .A2(n18725), .ZN(n18008) );
  AOI211_X1 U20843 ( .C1(n17666), .C2(n17837), .A(n17665), .B(n18008), .ZN(
        n17672) );
  NOR2_X1 U20844 ( .A1(n17690), .A2(n17999), .ZN(n17669) );
  INV_X1 U20845 ( .A(n17669), .ZN(n18002) );
  AOI221_X1 U20846 ( .B1(n18037), .B2(n18006), .C1(n18002), .C2(n18006), .A(
        n17667), .ZN(n18009) );
  NOR2_X1 U20847 ( .A1(n17685), .A2(n18036), .ZN(n17723) );
  AOI22_X1 U20848 ( .A1(n17723), .A2(n17669), .B1(n17668), .B2(n18032), .ZN(
        n17670) );
  XOR2_X1 U20849 ( .A(n18006), .B(n17670), .Z(n18010) );
  AOI22_X1 U20850 ( .A1(n17834), .A2(n18009), .B1(n17755), .B2(n18010), .ZN(
        n17671) );
  OAI211_X1 U20851 ( .C1(n17759), .C2(n18003), .A(n17672), .B(n17671), .ZN(
        P3_U2816) );
  NAND2_X1 U20852 ( .A1(n17673), .A2(n17690), .ZN(n18023) );
  OAI21_X1 U20853 ( .B1(n17708), .B2(n17817), .A(n17845), .ZN(n17765) );
  AOI21_X1 U20854 ( .B1(n17675), .B2(n17674), .A(n17765), .ZN(n17676) );
  OAI21_X1 U20855 ( .B1(n17677), .B2(n17817), .A(n17676), .ZN(n17698) );
  INV_X1 U20856 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18722) );
  NOR2_X1 U20857 ( .A1(n9796), .A2(n18722), .ZN(n17684) );
  OAI211_X1 U20858 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17679), .B(n17678), .ZN(n17681) );
  OAI22_X1 U20859 ( .A1(n17682), .A2(n17681), .B1(n17680), .B2(n17696), .ZN(
        n17683) );
  AOI211_X1 U20860 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17698), .A(
        n17684), .B(n17683), .ZN(n17692) );
  OAI22_X1 U20861 ( .A1(n18017), .A2(n17850), .B1(n18016), .B2(n17759), .ZN(
        n17704) );
  NOR2_X1 U20862 ( .A1(n18032), .A2(n17685), .ZN(n17688) );
  INV_X1 U20863 ( .A(n17701), .ZN(n17687) );
  OAI22_X1 U20864 ( .A1(n17688), .A2(n17687), .B1(n17686), .B2(n18032), .ZN(
        n17689) );
  XOR2_X1 U20865 ( .A(n17690), .B(n17689), .Z(n18014) );
  AOI22_X1 U20866 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17704), .B1(
        n17755), .B2(n18014), .ZN(n17691) );
  OAI211_X1 U20867 ( .C1(n17745), .C2(n18023), .A(n17692), .B(n17691), .ZN(
        P3_U2817) );
  INV_X1 U20868 ( .A(n17702), .ZN(n18025) );
  NAND2_X1 U20869 ( .A1(n18025), .A2(n18032), .ZN(n17707) );
  NOR2_X1 U20870 ( .A1(n17694), .A2(n17693), .ZN(n17700) );
  NAND2_X1 U20871 ( .A1(n9790), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18030) );
  OAI21_X1 U20872 ( .B1(n17696), .B2(n17695), .A(n18030), .ZN(n17697) );
  AOI221_X1 U20873 ( .B1(n17700), .B2(n17699), .C1(n17698), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17697), .ZN(n17706) );
  INV_X1 U20874 ( .A(n17723), .ZN(n17734) );
  OAI21_X1 U20875 ( .B1(n17702), .B2(n17734), .A(n17701), .ZN(n17703) );
  XOR2_X1 U20876 ( .A(n17703), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18029) );
  AOI22_X1 U20877 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17704), .B1(
        n17755), .B2(n18029), .ZN(n17705) );
  OAI211_X1 U20878 ( .C1(n17745), .C2(n17707), .A(n17706), .B(n17705), .ZN(
        P3_U2818) );
  NAND2_X1 U20879 ( .A1(n18552), .A2(n17708), .ZN(n17777) );
  NOR3_X1 U20880 ( .A1(n17746), .A2(n17709), .A3(n17777), .ZN(n17740) );
  NAND2_X1 U20881 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17740), .ZN(
        n17730) );
  OAI21_X1 U20882 ( .B1(n17842), .B2(n17710), .A(n17730), .ZN(n17711) );
  AOI22_X1 U20883 ( .A1(n16272), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17712), 
        .B2(n17711), .ZN(n17720) );
  AOI21_X1 U20884 ( .B1(n18034), .B2(n17723), .A(n17713), .ZN(n17714) );
  XOR2_X1 U20885 ( .A(n17717), .B(n17714), .Z(n18033) );
  NAND2_X1 U20886 ( .A1(n18034), .A2(n17717), .ZN(n18048) );
  AOI22_X1 U20887 ( .A1(n18036), .A2(n17715), .B1(n17834), .B2(n18037), .ZN(
        n17744) );
  OAI21_X1 U20888 ( .B1(n18034), .B2(n17745), .A(n17744), .ZN(n17716) );
  INV_X1 U20889 ( .A(n17716), .ZN(n17725) );
  OAI22_X1 U20890 ( .A1(n17745), .A2(n18048), .B1(n17725), .B2(n17717), .ZN(
        n17718) );
  AOI21_X1 U20891 ( .B1(n17755), .B2(n18033), .A(n17718), .ZN(n17719) );
  OAI211_X1 U20892 ( .C1(n17829), .C2(n17721), .A(n17720), .B(n17719), .ZN(
        P3_U2819) );
  NOR3_X1 U20893 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17754), .A3(
        n17735), .ZN(n17722) );
  AOI21_X1 U20894 ( .B1(n17723), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17722), .ZN(n17724) );
  XNOR2_X1 U20895 ( .A(n17726), .B(n17724), .ZN(n18056) );
  AOI221_X1 U20896 ( .B1(n17745), .B2(n17726), .C1(n18063), .C2(n17726), .A(
        n17725), .ZN(n17728) );
  NOR2_X1 U20897 ( .A1(n9796), .A2(n18716), .ZN(n17727) );
  AOI211_X1 U20898 ( .C1(n17729), .C2(n17837), .A(n17728), .B(n17727), .ZN(
        n17732) );
  INV_X1 U20899 ( .A(n17842), .ZN(n17782) );
  OAI211_X1 U20900 ( .C1(n17740), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17782), .B(n17730), .ZN(n17731) );
  OAI211_X1 U20901 ( .C1(n18056), .C2(n17733), .A(n17732), .B(n17731), .ZN(
        P3_U2820) );
  OAI21_X1 U20902 ( .B1(n17735), .B2(n17754), .A(n17734), .ZN(n17736) );
  XOR2_X1 U20903 ( .A(n17736), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18060) );
  NOR2_X1 U20904 ( .A1(n9796), .A2(n21076), .ZN(n17742) );
  NOR2_X1 U20905 ( .A1(n17746), .A2(n17777), .ZN(n17737) );
  AOI21_X1 U20906 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17782), .A(
        n17737), .ZN(n17739) );
  OAI22_X1 U20907 ( .A1(n17740), .A2(n17739), .B1(n17829), .B2(n17738), .ZN(
        n17741) );
  AOI211_X1 U20908 ( .C1(n17755), .C2(n18060), .A(n17742), .B(n17741), .ZN(
        n17743) );
  OAI221_X1 U20909 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17745), .C1(
        n18063), .C2(n17744), .A(n17743), .ZN(P3_U2821) );
  OAI211_X1 U20910 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17747), .A(
        n18552), .B(n17746), .ZN(n17748) );
  NAND2_X1 U20911 ( .A1(n9790), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18080) );
  OAI211_X1 U20912 ( .C1(n17829), .C2(n17749), .A(n17748), .B(n18080), .ZN(
        n17750) );
  AOI21_X1 U20913 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17765), .A(
        n17750), .ZN(n17757) );
  AOI21_X1 U20914 ( .B1(n17752), .B2(n18070), .A(n17751), .ZN(n18065) );
  OAI21_X1 U20915 ( .B1(n17754), .B2(n18067), .A(n17753), .ZN(n18077) );
  AOI22_X1 U20916 ( .A1(n17834), .A2(n18065), .B1(n17755), .B2(n18077), .ZN(
        n17756) );
  OAI211_X1 U20917 ( .C1(n17759), .C2(n17758), .A(n17757), .B(n17756), .ZN(
        P3_U2822) );
  NAND2_X1 U20918 ( .A1(n17761), .A2(n17760), .ZN(n17762) );
  XOR2_X1 U20919 ( .A(n17762), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18090) );
  INV_X1 U20920 ( .A(n17777), .ZN(n17764) );
  NOR2_X1 U20921 ( .A1(n9796), .A2(n18711), .ZN(n18083) );
  AOI221_X1 U20922 ( .B1(n17765), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n17764), .C2(n17763), .A(n18083), .ZN(n17770) );
  AOI21_X1 U20923 ( .B1(n18085), .B2(n17767), .A(n17766), .ZN(n18086) );
  AOI22_X1 U20924 ( .A1(n17838), .A2(n18086), .B1(n17768), .B2(n17837), .ZN(
        n17769) );
  OAI211_X1 U20925 ( .C1(n17850), .C2(n18090), .A(n17770), .B(n17769), .ZN(
        P3_U2823) );
  AOI21_X1 U20926 ( .B1(n17772), .B2(n17771), .A(n9926), .ZN(n18094) );
  AOI22_X1 U20927 ( .A1(n17838), .A2(n18094), .B1(n9790), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n17779) );
  AOI21_X1 U20928 ( .B1(n18091), .B2(n17774), .A(n17773), .ZN(n18093) );
  OAI22_X1 U20929 ( .A1(n17842), .A2(n17775), .B1(n18464), .B2(n17781), .ZN(
        n17776) );
  AOI22_X1 U20930 ( .A1(n17834), .A2(n18093), .B1(n17777), .B2(n17776), .ZN(
        n17778) );
  OAI211_X1 U20931 ( .C1(n17829), .C2(n17780), .A(n17779), .B(n17778), .ZN(
        P3_U2824) );
  NOR2_X1 U20932 ( .A1(n18464), .A2(n17781), .ZN(n17795) );
  OAI221_X1 U20933 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17783), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n17845), .A(n17782), .ZN(n17794) );
  AOI21_X1 U20934 ( .B1(n17786), .B2(n17785), .A(n17784), .ZN(n18099) );
  AOI22_X1 U20935 ( .A1(n17834), .A2(n18099), .B1(n9790), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17793) );
  AOI21_X1 U20936 ( .B1(n17789), .B2(n17788), .A(n17787), .ZN(n17790) );
  XOR2_X1 U20937 ( .A(n17790), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18100) );
  AOI22_X1 U20938 ( .A1(n17838), .A2(n18100), .B1(n17791), .B2(n17837), .ZN(
        n17792) );
  OAI211_X1 U20939 ( .C1(n17795), .C2(n17794), .A(n17793), .B(n17792), .ZN(
        P3_U2825) );
  AOI21_X1 U20940 ( .B1(n17798), .B2(n17797), .A(n17796), .ZN(n18105) );
  AOI22_X1 U20941 ( .A1(n17834), .A2(n18105), .B1(n18552), .B2(n17799), .ZN(
        n17808) );
  AOI21_X1 U20942 ( .B1(n17802), .B2(n17801), .A(n17800), .ZN(n18111) );
  OAI22_X1 U20943 ( .A1(n17829), .A2(n17805), .B1(n17812), .B2(n17804), .ZN(
        n17806) );
  AOI21_X1 U20944 ( .B1(n17838), .B2(n18111), .A(n17806), .ZN(n17807) );
  OAI211_X1 U20945 ( .C1(n9796), .C2(n18705), .A(n17808), .B(n17807), .ZN(
        P3_U2826) );
  AOI21_X1 U20946 ( .B1(n17811), .B2(n17810), .A(n17809), .ZN(n18119) );
  INV_X1 U20947 ( .A(n17812), .ZN(n17813) );
  AOI22_X1 U20948 ( .A1(n17838), .A2(n18119), .B1(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17813), .ZN(n17821) );
  AOI21_X1 U20949 ( .B1(n17816), .B2(n17815), .A(n17814), .ZN(n18118) );
  NOR2_X1 U20950 ( .A1(n9796), .A2(n18703), .ZN(n18117) );
  INV_X1 U20951 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17832) );
  NOR4_X1 U20952 ( .A1(n17818), .A2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        n17832), .A4(n17817), .ZN(n17819) );
  AOI211_X1 U20953 ( .C1(n17834), .C2(n18118), .A(n18117), .B(n17819), .ZN(
        n17820) );
  OAI211_X1 U20954 ( .C1(n17829), .C2(n17822), .A(n17821), .B(n17820), .ZN(
        P3_U2827) );
  AOI21_X1 U20955 ( .B1(n17825), .B2(n17824), .A(n17823), .ZN(n18132) );
  NOR2_X1 U20956 ( .A1(n9796), .A2(n18701), .ZN(n18124) );
  XNOR2_X1 U20957 ( .A(n17827), .B(n17826), .ZN(n18137) );
  OAI22_X1 U20958 ( .A1(n17829), .A2(n17828), .B1(n17850), .B2(n18137), .ZN(
        n17830) );
  AOI211_X1 U20959 ( .C1(n17838), .C2(n18132), .A(n18124), .B(n17830), .ZN(
        n17831) );
  OAI221_X1 U20960 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18464), .C1(
        n17832), .C2(n17845), .A(n17831), .ZN(P3_U2828) );
  NOR2_X1 U20961 ( .A1(n17844), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17833) );
  XNOR2_X1 U20962 ( .A(n17833), .B(n17836), .ZN(n18138) );
  AOI22_X1 U20963 ( .A1(n17834), .A2(n18138), .B1(n9790), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17840) );
  AOI21_X1 U20964 ( .B1(n17836), .B2(n17843), .A(n17835), .ZN(n18140) );
  AOI22_X1 U20965 ( .A1(n17838), .A2(n18140), .B1(n17841), .B2(n17837), .ZN(
        n17839) );
  OAI211_X1 U20966 ( .C1(n17842), .C2(n17841), .A(n17840), .B(n17839), .ZN(
        P3_U2829) );
  OAI21_X1 U20967 ( .B1(n17844), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17843), .ZN(n18155) );
  INV_X1 U20968 ( .A(n18155), .ZN(n18157) );
  NAND3_X1 U20969 ( .A1(n18779), .A2(n17846), .A3(n17845), .ZN(n17847) );
  AOI22_X1 U20970 ( .A1(n9790), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17847), .ZN(n17848) );
  OAI221_X1 U20971 ( .B1(n18157), .B2(n17850), .C1(n18155), .C2(n17849), .A(
        n17848), .ZN(P3_U2830) );
  OAI21_X1 U20972 ( .B1(n17851), .B2(n17907), .A(n17862), .ZN(n17865) );
  NOR2_X1 U20973 ( .A1(n18637), .A2(n18635), .ZN(n18143) );
  INV_X1 U20974 ( .A(n18143), .ZN(n17861) );
  NOR2_X1 U20975 ( .A1(n17852), .A2(n18612), .ZN(n17872) );
  NOR2_X1 U20976 ( .A1(n18043), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18126) );
  INV_X1 U20977 ( .A(n17957), .ZN(n17917) );
  NOR3_X1 U20978 ( .A1(n18126), .A2(n17917), .A3(n17853), .ZN(n17897) );
  NAND2_X1 U20979 ( .A1(n18639), .A2(n18043), .ZN(n18128) );
  INV_X1 U20980 ( .A(n18128), .ZN(n18072) );
  AOI21_X1 U20981 ( .B1(n17854), .B2(n17897), .A(n18072), .ZN(n17880) );
  AOI22_X1 U20982 ( .A1(n17855), .A2(n18068), .B1(n18623), .B2(n17871), .ZN(
        n17856) );
  INV_X1 U20983 ( .A(n17856), .ZN(n17857) );
  AOI211_X1 U20984 ( .C1(n18066), .C2(n17858), .A(n17880), .B(n17857), .ZN(
        n17873) );
  OAI211_X1 U20985 ( .C1(n18639), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17873), .ZN(n17859) );
  AOI211_X1 U20986 ( .C1(n17861), .C2(n17860), .A(n17872), .B(n17859), .ZN(
        n17863) );
  OAI22_X1 U20987 ( .A1(n17863), .A2(n18142), .B1(n17862), .B2(n18109), .ZN(
        n17864) );
  AOI22_X1 U20988 ( .A1(n18078), .A2(n17866), .B1(n17865), .B2(n17864), .ZN(
        n17868) );
  NAND2_X1 U20989 ( .A1(n17868), .A2(n17867), .ZN(P3_U2835) );
  AND2_X1 U20990 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17869), .ZN(
        n17894) );
  AOI22_X1 U20991 ( .A1(n9790), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n17870), 
        .B2(n17894), .ZN(n17876) );
  NOR2_X1 U20992 ( .A1(n17872), .A2(n17871), .ZN(n17878) );
  OAI211_X1 U20993 ( .C1(n18143), .C2(n17878), .A(n17873), .B(n18150), .ZN(
        n17874) );
  NAND3_X1 U20994 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n9796), .A3(
        n17874), .ZN(n17875) );
  OAI211_X1 U20995 ( .C1(n17877), .C2(n10104), .A(n17876), .B(n17875), .ZN(
        P3_U2836) );
  INV_X1 U20996 ( .A(n17878), .ZN(n17879) );
  NOR2_X1 U20997 ( .A1(n17880), .A2(n17879), .ZN(n17887) );
  NOR3_X1 U20998 ( .A1(n17883), .A2(n17882), .A3(n17881), .ZN(n17884) );
  NOR2_X1 U20999 ( .A1(n17884), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17886) );
  OAI222_X1 U21000 ( .A1(n17888), .A2(n18015), .B1(n17887), .B2(n17886), .C1(
        n18611), .C2(n17885), .ZN(n17889) );
  AOI22_X1 U21001 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18144), .B1(
        n18150), .B2(n17889), .ZN(n17891) );
  OAI211_X1 U21002 ( .C1(n17892), .C2(n10104), .A(n17891), .B(n17890), .ZN(
        P3_U2837) );
  AOI22_X1 U21003 ( .A1(n18078), .A2(n17895), .B1(n17894), .B2(n17893), .ZN(
        n17905) );
  OAI22_X1 U21004 ( .A1(n18072), .A2(n17897), .B1(n17896), .B2(n18611), .ZN(
        n17898) );
  AOI211_X1 U21005 ( .C1(n18068), .C2(n17899), .A(n18144), .B(n17898), .ZN(
        n17902) );
  INV_X1 U21006 ( .A(n17902), .ZN(n17903) );
  AOI21_X1 U21007 ( .B1(n18635), .B2(n17900), .A(n17906), .ZN(n17901) );
  AOI21_X1 U21008 ( .B1(n17902), .B2(n17901), .A(n9790), .ZN(n17909) );
  OAI211_X1 U21009 ( .C1(n18076), .C2(n17903), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17909), .ZN(n17904) );
  OAI211_X1 U21010 ( .C1(n18743), .C2(n9796), .A(n17905), .B(n17904), .ZN(
        P3_U2838) );
  OAI21_X1 U21011 ( .B1(n18144), .B2(n17907), .A(n17906), .ZN(n17908) );
  AOI22_X1 U21012 ( .A1(n18078), .A2(n17910), .B1(n17909), .B2(n17908), .ZN(
        n17912) );
  NAND2_X1 U21013 ( .A1(n17912), .A2(n17911), .ZN(P3_U2839) );
  NAND2_X1 U21014 ( .A1(n18150), .A2(n17931), .ZN(n17913) );
  OAI22_X1 U21015 ( .A1(n17914), .A2(n17913), .B1(n17930), .B2(n18142), .ZN(
        n17926) );
  NOR2_X1 U21016 ( .A1(n18637), .A2(n17930), .ZN(n17923) );
  AOI22_X1 U21017 ( .A1(n18066), .A2(n17988), .B1(n18068), .B2(n17915), .ZN(
        n17935) );
  INV_X1 U21018 ( .A(n18052), .ZN(n17921) );
  OAI21_X1 U21019 ( .B1(n17917), .B2(n17916), .A(n18623), .ZN(n17918) );
  OAI221_X1 U21020 ( .B1(n18612), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), 
        .C1(n18612), .C2(n17956), .A(n17918), .ZN(n17936) );
  NAND2_X1 U21021 ( .A1(n18611), .A2(n18015), .ZN(n18041) );
  INV_X1 U21022 ( .A(n18041), .ZN(n17961) );
  OAI22_X1 U21023 ( .A1(n18639), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17961), .B2(n17919), .ZN(n17940) );
  AOI211_X1 U21024 ( .C1(n17921), .C2(n17920), .A(n17936), .B(n17940), .ZN(
        n17922) );
  OAI211_X1 U21025 ( .C1(n17924), .C2(n17923), .A(n17935), .B(n17922), .ZN(
        n17925) );
  AOI22_X1 U21026 ( .A1(n18078), .A2(n17927), .B1(n17926), .B2(n17925), .ZN(
        n17929) );
  OAI211_X1 U21027 ( .C1(n18109), .C2(n17930), .A(n17929), .B(n17928), .ZN(
        P3_U2840) );
  NAND3_X1 U21028 ( .A1(n18134), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17931), .ZN(n17955) );
  AOI22_X1 U21029 ( .A1(n16272), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18078), 
        .B2(n17932), .ZN(n17942) );
  AOI21_X1 U21030 ( .B1(n17934), .B2(n17933), .A(n18043), .ZN(n17937) );
  NAND2_X1 U21031 ( .A1(n18150), .A2(n17935), .ZN(n17977) );
  NOR3_X1 U21032 ( .A1(n17937), .A2(n17977), .A3(n17936), .ZN(n17946) );
  OAI21_X1 U21033 ( .B1(n17938), .B2(n18143), .A(n17946), .ZN(n17939) );
  OAI211_X1 U21034 ( .C1(n17940), .C2(n17939), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n9796), .ZN(n17941) );
  OAI211_X1 U21035 ( .C1(n17943), .C2(n17955), .A(n17942), .B(n17941), .ZN(
        P3_U2841) );
  AOI22_X1 U21036 ( .A1(n16272), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18078), 
        .B2(n17944), .ZN(n17949) );
  AOI221_X1 U21037 ( .B1(n17961), .B2(n17946), .C1(n17945), .C2(n17946), .A(
        n9790), .ZN(n17952) );
  NOR3_X1 U21038 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18143), .A3(
        n18661), .ZN(n17947) );
  OAI21_X1 U21039 ( .B1(n17952), .B2(n17947), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17948) );
  OAI211_X1 U21040 ( .C1(n17950), .C2(n17955), .A(n17949), .B(n17948), .ZN(
        P3_U2842) );
  AOI22_X1 U21041 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17952), .B1(
        n18078), .B2(n17951), .ZN(n17954) );
  OAI211_X1 U21042 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17955), .A(
        n17954), .B(n17953), .ZN(P3_U2843) );
  NOR2_X1 U21043 ( .A1(n17956), .A2(n18612), .ZN(n17959) );
  AOI21_X1 U21044 ( .B1(n17957), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n18072), .ZN(n17958) );
  NOR4_X1 U21045 ( .A1(n18126), .A2(n17959), .A3(n17958), .A4(n17977), .ZN(
        n17960) );
  OAI21_X1 U21046 ( .B1(n17962), .B2(n17961), .A(n17960), .ZN(n21221) );
  OAI221_X1 U21047 ( .B1(n21221), .B2(n17963), .C1(n21221), .C2(n18128), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17971) );
  INV_X1 U21048 ( .A(n17964), .ZN(n17965) );
  OAI22_X1 U21049 ( .A1(n18106), .A2(n18612), .B1(n18108), .B2(n18125), .ZN(
        n18116) );
  NAND2_X1 U21050 ( .A1(n17965), .A2(n18116), .ZN(n18098) );
  NOR3_X1 U21051 ( .A1(n18085), .A2(n18091), .A3(n18098), .ZN(n18069) );
  NAND2_X1 U21052 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18069), .ZN(
        n17998) );
  NAND2_X1 U21053 ( .A1(n17966), .A2(n17998), .ZN(n18024) );
  NAND2_X1 U21054 ( .A1(n18134), .A2(n18024), .ZN(n18064) );
  NOR2_X1 U21055 ( .A1(n17967), .A2(n18064), .ZN(n21219) );
  AOI22_X1 U21056 ( .A1(n18078), .A2(n17969), .B1(n21219), .B2(n17968), .ZN(
        n17970) );
  OAI221_X1 U21057 ( .B1(n9790), .B2(n17971), .C1(n9796), .C2(n21167), .A(
        n17970), .ZN(P3_U2844) );
  NAND2_X1 U21058 ( .A1(n18623), .A2(n17972), .ZN(n18050) );
  NAND2_X1 U21059 ( .A1(n18043), .A2(n18050), .ZN(n18057) );
  NAND2_X1 U21060 ( .A1(n18635), .A2(n17973), .ZN(n18038) );
  INV_X1 U21061 ( .A(n18038), .ZN(n17974) );
  AOI211_X1 U21062 ( .C1(n17975), .C2(n18057), .A(n17989), .B(n17974), .ZN(
        n17983) );
  OAI21_X1 U21063 ( .B1(n18052), .B2(n17976), .A(n17983), .ZN(n17987) );
  OAI221_X1 U21064 ( .B1(n17977), .B2(n18076), .C1(n17977), .C2(n17987), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17981) );
  AOI22_X1 U21065 ( .A1(n17979), .A2(n18078), .B1(n21219), .B2(n17978), .ZN(
        n17980) );
  OAI221_X1 U21066 ( .B1(n9790), .B2(n17981), .C1(n9796), .C2(n18728), .A(
        n17980), .ZN(P3_U2846) );
  NOR2_X1 U21067 ( .A1(n17982), .A2(n18015), .ZN(n17986) );
  NOR4_X1 U21068 ( .A1(n17983), .A2(n17998), .A3(n18006), .A4(n18002), .ZN(
        n17984) );
  AOI21_X1 U21069 ( .B1(n17986), .B2(n17985), .A(n17984), .ZN(n17997) );
  AOI211_X1 U21070 ( .C1(n18066), .C2(n17988), .A(n18142), .B(n17987), .ZN(
        n17990) );
  NOR3_X1 U21071 ( .A1(n9790), .A2(n17990), .A3(n17989), .ZN(n17993) );
  NOR3_X1 U21072 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17991), .A3(
        n18156), .ZN(n17992) );
  AOI211_X1 U21073 ( .C1(n17994), .C2(n18078), .A(n17993), .B(n17992), .ZN(
        n17996) );
  OAI211_X1 U21074 ( .C1(n17997), .C2(n18142), .A(n17996), .B(n17995), .ZN(
        P3_U2847) );
  NOR2_X1 U21075 ( .A1(n17998), .A2(n18002), .ZN(n18007) );
  INV_X1 U21076 ( .A(n18050), .ZN(n18001) );
  OAI21_X1 U21077 ( .B1(n17999), .B2(n18058), .A(n18637), .ZN(n18000) );
  NAND2_X1 U21078 ( .A1(n18038), .A2(n18000), .ZN(n18019) );
  AOI211_X1 U21079 ( .C1(n18076), .C2(n18002), .A(n18001), .B(n18019), .ZN(
        n18004) );
  OAI22_X1 U21080 ( .A1(n18004), .A2(n18006), .B1(n18015), .B2(n18003), .ZN(
        n18005) );
  AOI21_X1 U21081 ( .B1(n18007), .B2(n18006), .A(n18005), .ZN(n18013) );
  AOI21_X1 U21082 ( .B1(n18144), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18008), .ZN(n18012) );
  AOI22_X1 U21083 ( .A1(n18078), .A2(n18010), .B1(n18139), .B2(n18009), .ZN(
        n18011) );
  OAI211_X1 U21084 ( .C1(n18013), .C2(n18142), .A(n18012), .B(n18011), .ZN(
        P3_U2848) );
  AOI22_X1 U21085 ( .A1(n16272), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18078), 
        .B2(n18014), .ZN(n18022) );
  AOI21_X1 U21086 ( .B1(n18025), .B2(n18050), .A(n18052), .ZN(n18045) );
  OAI22_X1 U21087 ( .A1(n18017), .A2(n18611), .B1(n18016), .B2(n18015), .ZN(
        n18018) );
  NOR3_X1 U21088 ( .A1(n18045), .A2(n18019), .A3(n18018), .ZN(n18027) );
  OAI211_X1 U21089 ( .C1(n18052), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18150), .B(n18027), .ZN(n18020) );
  NAND3_X1 U21090 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n9796), .A3(
        n18020), .ZN(n18021) );
  OAI211_X1 U21091 ( .C1(n18023), .C2(n18064), .A(n18022), .B(n18021), .ZN(
        P3_U2849) );
  NAND3_X1 U21092 ( .A1(n18025), .A2(n18024), .A3(n18032), .ZN(n18026) );
  OAI21_X1 U21093 ( .B1(n18027), .B2(n18032), .A(n18026), .ZN(n18028) );
  AOI22_X1 U21094 ( .A1(n18078), .A2(n18029), .B1(n18150), .B2(n18028), .ZN(
        n18031) );
  OAI211_X1 U21095 ( .C1(n18109), .C2(n18032), .A(n18031), .B(n18030), .ZN(
        P3_U2850) );
  AOI22_X1 U21096 ( .A1(n9790), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18078), 
        .B2(n18033), .ZN(n18047) );
  INV_X1 U21097 ( .A(n18034), .ZN(n18042) );
  AOI21_X1 U21098 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18035), .A(
        n18043), .ZN(n18040) );
  AOI22_X1 U21099 ( .A1(n18066), .A2(n18037), .B1(n18068), .B2(n18036), .ZN(
        n18039) );
  NAND3_X1 U21100 ( .A1(n18134), .A2(n18039), .A3(n18038), .ZN(n18059) );
  AOI211_X1 U21101 ( .C1(n18042), .C2(n18041), .A(n18040), .B(n18059), .ZN(
        n18051) );
  OAI21_X1 U21102 ( .B1(n18043), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18051), .ZN(n18044) );
  OAI211_X1 U21103 ( .C1(n18045), .C2(n18044), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n9796), .ZN(n18046) );
  OAI211_X1 U21104 ( .C1(n18048), .C2(n18064), .A(n18047), .B(n18046), .ZN(
        P3_U2851) );
  NOR2_X1 U21105 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18064), .ZN(
        n18049) );
  AOI22_X1 U21106 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18049), .B1(
        n9790), .B2(P3_REIP_REG_10__SCAN_IN), .ZN(n18055) );
  OAI211_X1 U21107 ( .C1(n18052), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18051), .B(n18050), .ZN(n18053) );
  NAND3_X1 U21108 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n9796), .A3(
        n18053), .ZN(n18054) );
  OAI211_X1 U21109 ( .C1(n18056), .C2(n10104), .A(n18055), .B(n18054), .ZN(
        P3_U2852) );
  OAI221_X1 U21110 ( .B1(n18059), .B2(n18058), .C1(n18059), .C2(n18057), .A(
        n9796), .ZN(n18062) );
  AOI22_X1 U21111 ( .A1(n9790), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18078), .B2(
        n18060), .ZN(n18061) );
  OAI221_X1 U21112 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18064), .C1(
        n18063), .C2(n18062), .A(n18061), .ZN(P3_U2853) );
  AOI222_X1 U21113 ( .A1(n18070), .A2(n18069), .B1(n18068), .B2(n18067), .C1(
        n18066), .C2(n18065), .ZN(n18082) );
  OAI22_X1 U21114 ( .A1(n18073), .A2(n18072), .B1(n18071), .B2(n18612), .ZN(
        n18074) );
  NOR2_X1 U21115 ( .A1(n18126), .A2(n18074), .ZN(n18092) );
  INV_X1 U21116 ( .A(n18092), .ZN(n18075) );
  AOI211_X1 U21117 ( .C1(n18076), .C2(n18091), .A(n18085), .B(n18075), .ZN(
        n18084) );
  OAI21_X1 U21118 ( .B1(n18084), .B2(n18110), .A(n18109), .ZN(n18079) );
  AOI22_X1 U21119 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18079), .B1(
        n18078), .B2(n18077), .ZN(n18081) );
  OAI211_X1 U21120 ( .C1(n18082), .C2(n18142), .A(n18081), .B(n18080), .ZN(
        P3_U2854) );
  AOI21_X1 U21121 ( .B1(n18144), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18083), .ZN(n18089) );
  AOI221_X1 U21122 ( .B1(n18091), .B2(n18085), .C1(n18098), .C2(n18085), .A(
        n18084), .ZN(n18087) );
  AOI22_X1 U21123 ( .A1(n18134), .A2(n18087), .B1(n18141), .B2(n18086), .ZN(
        n18088) );
  OAI211_X1 U21124 ( .C1(n18156), .C2(n18090), .A(n18089), .B(n18088), .ZN(
        P3_U2855) );
  NAND2_X1 U21125 ( .A1(n18134), .A2(n18091), .ZN(n18097) );
  OAI21_X1 U21126 ( .B1(n18092), .B2(n18142), .A(n18109), .ZN(n18101) );
  AOI22_X1 U21127 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18101), .B1(
        n9790), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n18096) );
  AOI22_X1 U21128 ( .A1(n18141), .A2(n18094), .B1(n18139), .B2(n18093), .ZN(
        n18095) );
  OAI211_X1 U21129 ( .C1(n18098), .C2(n18097), .A(n18096), .B(n18095), .ZN(
        P3_U2856) );
  NAND4_X1 U21130 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n18134), .A4(n18116), .ZN(
        n18104) );
  AOI22_X1 U21131 ( .A1(n9790), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18139), .B2(
        n18099), .ZN(n18103) );
  AOI22_X1 U21132 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18101), .B1(
        n18141), .B2(n18100), .ZN(n18102) );
  OAI211_X1 U21133 ( .C1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n18104), .A(
        n18103), .B(n18102), .ZN(P3_U2857) );
  NAND3_X1 U21134 ( .A1(n18150), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18116), .ZN(n18115) );
  AOI22_X1 U21135 ( .A1(n9790), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18139), .B2(
        n18105), .ZN(n18114) );
  NAND2_X1 U21136 ( .A1(n18635), .A2(n18106), .ZN(n18129) );
  NAND2_X1 U21137 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18129), .ZN(
        n18107) );
  AOI211_X1 U21138 ( .C1(n18108), .C2(n18128), .A(n18126), .B(n18107), .ZN(
        n18123) );
  OAI21_X1 U21139 ( .B1(n18123), .B2(n18110), .A(n18109), .ZN(n18112) );
  AOI22_X1 U21140 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18112), .B1(
        n18141), .B2(n18111), .ZN(n18113) );
  OAI211_X1 U21141 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n18115), .A(
        n18114), .B(n18113), .ZN(P3_U2858) );
  OAI21_X1 U21142 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18116), .A(
        n18150), .ZN(n18122) );
  AOI21_X1 U21143 ( .B1(n18144), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n18117), .ZN(n18121) );
  AOI22_X1 U21144 ( .A1(n18141), .A2(n18119), .B1(n18139), .B2(n18118), .ZN(
        n18120) );
  OAI211_X1 U21145 ( .C1(n18123), .C2(n18122), .A(n18121), .B(n18120), .ZN(
        P3_U2859) );
  AOI21_X1 U21146 ( .B1(n18144), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18124), .ZN(n18136) );
  OR2_X1 U21147 ( .A1(n10446), .A2(n18125), .ZN(n18131) );
  NOR3_X1 U21148 ( .A1(n18612), .A2(n10446), .A3(n21150), .ZN(n18127) );
  AOI211_X1 U21149 ( .C1(n10446), .C2(n18128), .A(n18127), .B(n18126), .ZN(
        n18130) );
  OAI221_X1 U21150 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18131), .C1(
        n10459), .C2(n18130), .A(n18129), .ZN(n18133) );
  AOI22_X1 U21151 ( .A1(n18134), .A2(n18133), .B1(n18141), .B2(n18132), .ZN(
        n18135) );
  OAI211_X1 U21152 ( .C1(n18156), .C2(n18137), .A(n18136), .B(n18135), .ZN(
        P3_U2860) );
  AOI22_X1 U21153 ( .A1(n18141), .A2(n18140), .B1(n18139), .B2(n18138), .ZN(
        n18149) );
  NAND2_X1 U21154 ( .A1(n9790), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18148) );
  NOR3_X1 U21155 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18143), .A3(
        n18142), .ZN(n18151) );
  OAI21_X1 U21156 ( .B1(n18144), .B2(n18151), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18147) );
  OAI211_X1 U21157 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18623), .A(
        n18145), .B(n10446), .ZN(n18146) );
  NAND4_X1 U21158 ( .A1(n18149), .A2(n18148), .A3(n18147), .A4(n18146), .ZN(
        P3_U2861) );
  AOI21_X1 U21159 ( .B1(n18639), .B2(n18150), .A(n21150), .ZN(n18152) );
  AOI221_X1 U21160 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n9790), .C1(n18152), 
        .C2(n9796), .A(n18151), .ZN(n18153) );
  OAI221_X1 U21161 ( .B1(n18157), .B2(n18156), .C1(n18155), .C2(n18154), .A(
        n18153), .ZN(P3_U2862) );
  OAI211_X1 U21162 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18158), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18662)
         );
  OAI21_X1 U21163 ( .B1(n18161), .B2(n18159), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18160) );
  OAI221_X1 U21164 ( .B1(n18161), .B2(n18662), .C1(n18161), .C2(n18210), .A(
        n18160), .ZN(P3_U2863) );
  INV_X1 U21165 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18653) );
  NOR2_X1 U21166 ( .A1(n18650), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18341) );
  INV_X1 U21167 ( .A(n18341), .ZN(n18343) );
  NAND2_X1 U21168 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18650), .ZN(
        n18438) );
  AND2_X1 U21169 ( .A1(n18343), .A2(n18438), .ZN(n18163) );
  OAI22_X1 U21170 ( .A1(n18164), .A2(n18653), .B1(n18163), .B2(n18162), .ZN(
        P3_U2866) );
  NOR2_X1 U21171 ( .A1(n18654), .A2(n18165), .ZN(P3_U2867) );
  NOR2_X1 U21172 ( .A1(n18464), .A2(n18166), .ZN(n18548) );
  INV_X1 U21173 ( .A(n18548), .ZN(n18418) );
  NOR2_X1 U21174 ( .A1(n18653), .A2(n18387), .ZN(n18550) );
  NAND2_X1 U21175 ( .A1(n18550), .A2(n18412), .ZN(n18510) );
  NOR3_X1 U21176 ( .A1(n18650), .A2(n18653), .A3(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18551) );
  NAND2_X1 U21177 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18551), .ZN(
        n18605) );
  INV_X1 U21178 ( .A(n18605), .ZN(n18589) );
  NAND2_X1 U21179 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18552), .ZN(n18556) );
  INV_X1 U21180 ( .A(n18556), .ZN(n18413) );
  NOR2_X2 U21181 ( .A1(n18251), .A2(n18167), .ZN(n18547) );
  NAND2_X1 U21182 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18644) );
  NAND2_X1 U21183 ( .A1(n18412), .A2(n18645), .ZN(n18646) );
  NOR2_X1 U21184 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18253) );
  INV_X1 U21185 ( .A(n18253), .ZN(n18211) );
  NOR2_X2 U21186 ( .A1(n18646), .A2(n18211), .ZN(n18267) );
  NOR2_X1 U21187 ( .A1(n18600), .A2(n18267), .ZN(n18230) );
  NOR2_X1 U21188 ( .A1(n18509), .A2(n18230), .ZN(n18204) );
  AOI22_X1 U21189 ( .A1(n18589), .A2(n18413), .B1(n18547), .B2(n18204), .ZN(
        n18174) );
  INV_X1 U21190 ( .A(n18251), .ZN(n18463) );
  AOI21_X1 U21191 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18230), .ZN(n18169) );
  AOI21_X1 U21192 ( .B1(n18510), .B2(n18605), .A(n18251), .ZN(n18514) );
  AOI22_X1 U21193 ( .A1(n18463), .A2(n18169), .B1(n18168), .B2(n18514), .ZN(
        n18207) );
  NAND2_X1 U21194 ( .A1(n18171), .A2(n18170), .ZN(n18205) );
  NOR2_X2 U21195 ( .A1(n18172), .A2(n18205), .ZN(n18553) );
  AOI22_X1 U21196 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18207), .B1(
        n18267), .B2(n18553), .ZN(n18173) );
  OAI211_X1 U21197 ( .C1(n18418), .C2(n18510), .A(n18174), .B(n18173), .ZN(
        P3_U2868) );
  NOR2_X1 U21198 ( .A1(n18175), .A2(n18464), .ZN(n18558) );
  INV_X1 U21199 ( .A(n18558), .ZN(n18444) );
  INV_X1 U21200 ( .A(n18510), .ZN(n18541) );
  NAND2_X1 U21201 ( .A1(n18552), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18562) );
  INV_X1 U21202 ( .A(n18562), .ZN(n18441) );
  NOR2_X2 U21203 ( .A1(n18251), .A2(n18176), .ZN(n18557) );
  AOI22_X1 U21204 ( .A1(n18541), .A2(n18441), .B1(n18204), .B2(n18557), .ZN(
        n18178) );
  NOR2_X2 U21205 ( .A1(n18813), .A2(n18205), .ZN(n18559) );
  AOI22_X1 U21206 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18207), .B1(
        n18267), .B2(n18559), .ZN(n18177) );
  OAI211_X1 U21207 ( .C1(n18605), .C2(n18444), .A(n18178), .B(n18177), .ZN(
        P3_U2869) );
  NOR2_X1 U21208 ( .A1(n18464), .A2(n18179), .ZN(n18520) );
  INV_X1 U21209 ( .A(n18520), .ZN(n18568) );
  NAND2_X1 U21210 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18552), .ZN(n18523) );
  INV_X1 U21211 ( .A(n18523), .ZN(n18564) );
  NOR2_X2 U21212 ( .A1(n18251), .A2(n18180), .ZN(n18563) );
  AOI22_X1 U21213 ( .A1(n18589), .A2(n18564), .B1(n18204), .B2(n18563), .ZN(
        n18183) );
  NOR2_X2 U21214 ( .A1(n18181), .A2(n18205), .ZN(n18565) );
  AOI22_X1 U21215 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18207), .B1(
        n18267), .B2(n18565), .ZN(n18182) );
  OAI211_X1 U21216 ( .C1(n18510), .C2(n18568), .A(n18183), .B(n18182), .ZN(
        P3_U2870) );
  NOR2_X1 U21217 ( .A1(n15053), .A2(n18464), .ZN(n18524) );
  INV_X1 U21218 ( .A(n18524), .ZN(n18574) );
  NAND2_X1 U21219 ( .A1(n18552), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18527) );
  INV_X1 U21220 ( .A(n18527), .ZN(n18570) );
  NOR2_X2 U21221 ( .A1(n18251), .A2(n18184), .ZN(n18569) );
  AOI22_X1 U21222 ( .A1(n18541), .A2(n18570), .B1(n18204), .B2(n18569), .ZN(
        n18187) );
  NOR2_X2 U21223 ( .A1(n18185), .A2(n18205), .ZN(n18571) );
  AOI22_X1 U21224 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18207), .B1(
        n18267), .B2(n18571), .ZN(n18186) );
  OAI211_X1 U21225 ( .C1(n18605), .C2(n18574), .A(n18187), .B(n18186), .ZN(
        P3_U2871) );
  NOR2_X1 U21226 ( .A1(n18464), .A2(n18188), .ZN(n18576) );
  INV_X1 U21227 ( .A(n18576), .ZN(n18452) );
  NAND2_X1 U21228 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18552), .ZN(n18580) );
  INV_X1 U21229 ( .A(n18580), .ZN(n18449) );
  NOR2_X2 U21230 ( .A1(n18251), .A2(n18189), .ZN(n18575) );
  AOI22_X1 U21231 ( .A1(n18589), .A2(n18449), .B1(n18204), .B2(n18575), .ZN(
        n18192) );
  NOR2_X2 U21232 ( .A1(n18190), .A2(n18205), .ZN(n18577) );
  AOI22_X1 U21233 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18207), .B1(
        n18267), .B2(n18577), .ZN(n18191) );
  OAI211_X1 U21234 ( .C1(n18510), .C2(n18452), .A(n18192), .B(n18191), .ZN(
        P3_U2872) );
  NOR2_X1 U21235 ( .A1(n18193), .A2(n18464), .ZN(n18582) );
  INV_X1 U21236 ( .A(n18582), .ZN(n18533) );
  NAND2_X1 U21237 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18552), .ZN(n18586) );
  INV_X1 U21238 ( .A(n18586), .ZN(n18530) );
  NOR2_X2 U21239 ( .A1(n21119), .A2(n18251), .ZN(n18581) );
  AOI22_X1 U21240 ( .A1(n18589), .A2(n18530), .B1(n18204), .B2(n18581), .ZN(
        n18196) );
  NOR2_X2 U21241 ( .A1(n18194), .A2(n18205), .ZN(n18583) );
  AOI22_X1 U21242 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18207), .B1(
        n18267), .B2(n18583), .ZN(n18195) );
  OAI211_X1 U21243 ( .C1(n18510), .C2(n18533), .A(n18196), .B(n18195), .ZN(
        P3_U2873) );
  NOR2_X1 U21244 ( .A1(n18197), .A2(n18464), .ZN(n18588) );
  INV_X1 U21245 ( .A(n18588), .ZN(n18538) );
  NAND2_X1 U21246 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18552), .ZN(n18594) );
  INV_X1 U21247 ( .A(n18594), .ZN(n18535) );
  NOR2_X2 U21248 ( .A1(n18198), .A2(n18251), .ZN(n18587) );
  AOI22_X1 U21249 ( .A1(n18589), .A2(n18535), .B1(n18204), .B2(n18587), .ZN(
        n18201) );
  NOR2_X2 U21250 ( .A1(n18199), .A2(n18205), .ZN(n18590) );
  AOI22_X1 U21251 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18207), .B1(
        n18267), .B2(n18590), .ZN(n18200) );
  OAI211_X1 U21252 ( .C1(n18510), .C2(n18538), .A(n18201), .B(n18200), .ZN(
        P3_U2874) );
  NOR2_X1 U21253 ( .A1(n18202), .A2(n18464), .ZN(n18540) );
  INV_X1 U21254 ( .A(n18540), .ZN(n18604) );
  NAND2_X1 U21255 ( .A1(n18552), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18546) );
  INV_X1 U21256 ( .A(n18546), .ZN(n18598) );
  NOR2_X2 U21257 ( .A1(n18203), .A2(n18251), .ZN(n18596) );
  AOI22_X1 U21258 ( .A1(n18589), .A2(n18598), .B1(n18204), .B2(n18596), .ZN(
        n18209) );
  NOR2_X2 U21259 ( .A1(n18206), .A2(n18205), .ZN(n18599) );
  AOI22_X1 U21260 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18207), .B1(
        n18267), .B2(n18599), .ZN(n18208) );
  OAI211_X1 U21261 ( .C1(n18510), .C2(n18604), .A(n18209), .B(n18208), .ZN(
        P3_U2875) );
  INV_X1 U21262 ( .A(n18600), .ZN(n18250) );
  NAND2_X1 U21263 ( .A1(n18645), .A2(n18674), .ZN(n18386) );
  NOR2_X1 U21264 ( .A1(n18211), .A2(n18386), .ZN(n18226) );
  AOI22_X1 U21265 ( .A1(n18541), .A2(n18413), .B1(n18547), .B2(n18226), .ZN(
        n18213) );
  NAND2_X1 U21266 ( .A1(n18463), .A2(n18210), .ZN(n18388) );
  NOR2_X1 U21267 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18388), .ZN(
        n18297) );
  AOI22_X1 U21268 ( .A1(n18552), .A2(n18550), .B1(n18253), .B2(n18297), .ZN(
        n18227) );
  NAND2_X1 U21269 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18645), .ZN(
        n18390) );
  NOR2_X2 U21270 ( .A1(n18211), .A2(n18390), .ZN(n18293) );
  AOI22_X1 U21271 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18227), .B1(
        n18553), .B2(n18293), .ZN(n18212) );
  OAI211_X1 U21272 ( .C1(n18418), .C2(n18250), .A(n18213), .B(n18212), .ZN(
        P3_U2876) );
  AOI22_X1 U21273 ( .A1(n18541), .A2(n18558), .B1(n18557), .B2(n18226), .ZN(
        n18215) );
  AOI22_X1 U21274 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18227), .B1(
        n18559), .B2(n18293), .ZN(n18214) );
  OAI211_X1 U21275 ( .C1(n18250), .C2(n18562), .A(n18215), .B(n18214), .ZN(
        P3_U2877) );
  AOI22_X1 U21276 ( .A1(n18600), .A2(n18520), .B1(n18563), .B2(n18226), .ZN(
        n18217) );
  AOI22_X1 U21277 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18227), .B1(
        n18565), .B2(n18293), .ZN(n18216) );
  OAI211_X1 U21278 ( .C1(n18510), .C2(n18523), .A(n18217), .B(n18216), .ZN(
        P3_U2878) );
  AOI22_X1 U21279 ( .A1(n18600), .A2(n18570), .B1(n18569), .B2(n18226), .ZN(
        n18219) );
  AOI22_X1 U21280 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18227), .B1(
        n18571), .B2(n18293), .ZN(n18218) );
  OAI211_X1 U21281 ( .C1(n18510), .C2(n18574), .A(n18219), .B(n18218), .ZN(
        P3_U2879) );
  AOI22_X1 U21282 ( .A1(n18600), .A2(n18576), .B1(n18575), .B2(n18226), .ZN(
        n18221) );
  AOI22_X1 U21283 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18227), .B1(
        n18577), .B2(n18293), .ZN(n18220) );
  OAI211_X1 U21284 ( .C1(n18510), .C2(n18580), .A(n18221), .B(n18220), .ZN(
        P3_U2880) );
  AOI22_X1 U21285 ( .A1(n18600), .A2(n18582), .B1(n18581), .B2(n18226), .ZN(
        n18223) );
  AOI22_X1 U21286 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18227), .B1(
        n18583), .B2(n18293), .ZN(n18222) );
  OAI211_X1 U21287 ( .C1(n18510), .C2(n18586), .A(n18223), .B(n18222), .ZN(
        P3_U2881) );
  AOI22_X1 U21288 ( .A1(n18600), .A2(n18588), .B1(n18587), .B2(n18226), .ZN(
        n18225) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18227), .B1(
        n18590), .B2(n18293), .ZN(n18224) );
  OAI211_X1 U21290 ( .C1(n18510), .C2(n18594), .A(n18225), .B(n18224), .ZN(
        P3_U2882) );
  AOI22_X1 U21291 ( .A1(n18541), .A2(n18598), .B1(n18596), .B2(n18226), .ZN(
        n18229) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18227), .B1(
        n18599), .B2(n18293), .ZN(n18228) );
  OAI211_X1 U21293 ( .C1(n18250), .C2(n18604), .A(n18229), .B(n18228), .ZN(
        P3_U2883) );
  INV_X1 U21294 ( .A(n18293), .ZN(n18287) );
  NAND2_X1 U21295 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18253), .ZN(
        n18254) );
  NOR2_X2 U21296 ( .A1(n18254), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18315) );
  INV_X1 U21297 ( .A(n18315), .ZN(n18311) );
  AOI21_X1 U21298 ( .B1(n18287), .B2(n18311), .A(n18509), .ZN(n18246) );
  AOI22_X1 U21299 ( .A1(n18548), .A2(n18267), .B1(n18547), .B2(n18246), .ZN(
        n18233) );
  AOI221_X1 U21300 ( .B1(n18230), .B2(n18287), .C1(n18512), .C2(n18287), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18231) );
  OAI21_X1 U21301 ( .B1(n18315), .B2(n18231), .A(n18463), .ZN(n18247) );
  AOI22_X1 U21302 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18247), .B1(
        n18553), .B2(n18315), .ZN(n18232) );
  OAI211_X1 U21303 ( .C1(n18250), .C2(n18556), .A(n18233), .B(n18232), .ZN(
        P3_U2884) );
  AOI22_X1 U21304 ( .A1(n18267), .A2(n18441), .B1(n18557), .B2(n18246), .ZN(
        n18235) );
  AOI22_X1 U21305 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18247), .B1(
        n18559), .B2(n18315), .ZN(n18234) );
  OAI211_X1 U21306 ( .C1(n18250), .C2(n18444), .A(n18235), .B(n18234), .ZN(
        P3_U2885) );
  AOI22_X1 U21307 ( .A1(n18267), .A2(n18520), .B1(n18563), .B2(n18246), .ZN(
        n18237) );
  AOI22_X1 U21308 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18247), .B1(
        n18565), .B2(n18315), .ZN(n18236) );
  OAI211_X1 U21309 ( .C1(n18250), .C2(n18523), .A(n18237), .B(n18236), .ZN(
        P3_U2886) );
  AOI22_X1 U21310 ( .A1(n18267), .A2(n18570), .B1(n18569), .B2(n18246), .ZN(
        n18239) );
  AOI22_X1 U21311 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18247), .B1(
        n18571), .B2(n18315), .ZN(n18238) );
  OAI211_X1 U21312 ( .C1(n18250), .C2(n18574), .A(n18239), .B(n18238), .ZN(
        P3_U2887) );
  INV_X1 U21313 ( .A(n18267), .ZN(n18274) );
  AOI22_X1 U21314 ( .A1(n18600), .A2(n18449), .B1(n18575), .B2(n18246), .ZN(
        n18241) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18247), .B1(
        n18577), .B2(n18315), .ZN(n18240) );
  OAI211_X1 U21316 ( .C1(n18274), .C2(n18452), .A(n18241), .B(n18240), .ZN(
        P3_U2888) );
  AOI22_X1 U21317 ( .A1(n18267), .A2(n18582), .B1(n18581), .B2(n18246), .ZN(
        n18243) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18247), .B1(
        n18583), .B2(n18315), .ZN(n18242) );
  OAI211_X1 U21319 ( .C1(n18250), .C2(n18586), .A(n18243), .B(n18242), .ZN(
        P3_U2889) );
  AOI22_X1 U21320 ( .A1(n18267), .A2(n18588), .B1(n18587), .B2(n18246), .ZN(
        n18245) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18247), .B1(
        n18590), .B2(n18315), .ZN(n18244) );
  OAI211_X1 U21322 ( .C1(n18250), .C2(n18594), .A(n18245), .B(n18244), .ZN(
        P3_U2890) );
  AOI22_X1 U21323 ( .A1(n18267), .A2(n18540), .B1(n18596), .B2(n18246), .ZN(
        n18249) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18247), .B1(
        n18599), .B2(n18315), .ZN(n18248) );
  OAI211_X1 U21325 ( .C1(n18250), .C2(n18546), .A(n18249), .B(n18248), .ZN(
        P3_U2891) );
  AOI211_X1 U21326 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(n18644), .A(n18252), 
        .B(n18251), .ZN(n18342) );
  NAND2_X1 U21327 ( .A1(n18253), .A2(n18342), .ZN(n18271) );
  NOR2_X1 U21328 ( .A1(n18509), .A2(n18254), .ZN(n18270) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18271), .B1(
        n18547), .B2(n18270), .ZN(n18256) );
  INV_X1 U21330 ( .A(n18254), .ZN(n18298) );
  NAND2_X1 U21331 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18298), .ZN(
        n18335) );
  INV_X1 U21332 ( .A(n18335), .ZN(n18337) );
  AOI22_X1 U21333 ( .A1(n18548), .A2(n18293), .B1(n18553), .B2(n18337), .ZN(
        n18255) );
  OAI211_X1 U21334 ( .C1(n18274), .C2(n18556), .A(n18256), .B(n18255), .ZN(
        P3_U2892) );
  AOI22_X1 U21335 ( .A1(n18557), .A2(n18270), .B1(n18441), .B2(n18293), .ZN(
        n18258) );
  AOI22_X1 U21336 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18271), .B1(
        n18559), .B2(n18337), .ZN(n18257) );
  OAI211_X1 U21337 ( .C1(n18274), .C2(n18444), .A(n18258), .B(n18257), .ZN(
        P3_U2893) );
  AOI22_X1 U21338 ( .A1(n18267), .A2(n18564), .B1(n18563), .B2(n18270), .ZN(
        n18260) );
  AOI22_X1 U21339 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18271), .B1(
        n18565), .B2(n18337), .ZN(n18259) );
  OAI211_X1 U21340 ( .C1(n18568), .C2(n18287), .A(n18260), .B(n18259), .ZN(
        P3_U2894) );
  AOI22_X1 U21341 ( .A1(n18569), .A2(n18270), .B1(n18570), .B2(n18293), .ZN(
        n18262) );
  AOI22_X1 U21342 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18271), .B1(
        n18571), .B2(n18337), .ZN(n18261) );
  OAI211_X1 U21343 ( .C1(n18274), .C2(n18574), .A(n18262), .B(n18261), .ZN(
        P3_U2895) );
  AOI22_X1 U21344 ( .A1(n18576), .A2(n18293), .B1(n18575), .B2(n18270), .ZN(
        n18264) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18271), .B1(
        n18577), .B2(n18337), .ZN(n18263) );
  OAI211_X1 U21346 ( .C1(n18274), .C2(n18580), .A(n18264), .B(n18263), .ZN(
        P3_U2896) );
  AOI22_X1 U21347 ( .A1(n18267), .A2(n18530), .B1(n18581), .B2(n18270), .ZN(
        n18266) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18271), .B1(
        n18583), .B2(n18337), .ZN(n18265) );
  OAI211_X1 U21349 ( .C1(n18533), .C2(n18287), .A(n18266), .B(n18265), .ZN(
        P3_U2897) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18271), .B1(
        n18587), .B2(n18270), .ZN(n18269) );
  AOI22_X1 U21351 ( .A1(n18267), .A2(n18535), .B1(n18590), .B2(n18337), .ZN(
        n18268) );
  OAI211_X1 U21352 ( .C1(n18538), .C2(n18287), .A(n18269), .B(n18268), .ZN(
        P3_U2898) );
  AOI22_X1 U21353 ( .A1(n18540), .A2(n18293), .B1(n18596), .B2(n18270), .ZN(
        n18273) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18271), .B1(
        n18599), .B2(n18337), .ZN(n18272) );
  OAI211_X1 U21355 ( .C1(n18274), .C2(n18546), .A(n18273), .B(n18272), .ZN(
        P3_U2899) );
  NOR2_X2 U21356 ( .A1(n18646), .A2(n18343), .ZN(n18361) );
  NOR2_X1 U21357 ( .A1(n18337), .A2(n18361), .ZN(n18319) );
  NOR2_X1 U21358 ( .A1(n18509), .A2(n18319), .ZN(n18292) );
  AOI22_X1 U21359 ( .A1(n18413), .A2(n18293), .B1(n18547), .B2(n18292), .ZN(
        n18278) );
  NOR2_X1 U21360 ( .A1(n18293), .A2(n18315), .ZN(n18275) );
  OAI21_X1 U21361 ( .B1(n18275), .B2(n18512), .A(n18319), .ZN(n18276) );
  OAI211_X1 U21362 ( .C1(n18361), .C2(n18515), .A(n18463), .B(n18276), .ZN(
        n18294) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18294), .B1(
        n18553), .B2(n18361), .ZN(n18277) );
  OAI211_X1 U21364 ( .C1(n18418), .C2(n18311), .A(n18278), .B(n18277), .ZN(
        P3_U2900) );
  AOI22_X1 U21365 ( .A1(n18557), .A2(n18292), .B1(n18441), .B2(n18315), .ZN(
        n18280) );
  AOI22_X1 U21366 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18294), .B1(
        n18559), .B2(n18361), .ZN(n18279) );
  OAI211_X1 U21367 ( .C1(n18444), .C2(n18287), .A(n18280), .B(n18279), .ZN(
        P3_U2901) );
  AOI22_X1 U21368 ( .A1(n18564), .A2(n18293), .B1(n18563), .B2(n18292), .ZN(
        n18282) );
  AOI22_X1 U21369 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18294), .B1(
        n18565), .B2(n18361), .ZN(n18281) );
  OAI211_X1 U21370 ( .C1(n18568), .C2(n18311), .A(n18282), .B(n18281), .ZN(
        P3_U2902) );
  AOI22_X1 U21371 ( .A1(n18524), .A2(n18293), .B1(n18569), .B2(n18292), .ZN(
        n18284) );
  AOI22_X1 U21372 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18294), .B1(
        n18571), .B2(n18361), .ZN(n18283) );
  OAI211_X1 U21373 ( .C1(n18527), .C2(n18311), .A(n18284), .B(n18283), .ZN(
        P3_U2903) );
  AOI22_X1 U21374 ( .A1(n18576), .A2(n18315), .B1(n18575), .B2(n18292), .ZN(
        n18286) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18294), .B1(
        n18577), .B2(n18361), .ZN(n18285) );
  OAI211_X1 U21376 ( .C1(n18580), .C2(n18287), .A(n18286), .B(n18285), .ZN(
        P3_U2904) );
  AOI22_X1 U21377 ( .A1(n18581), .A2(n18292), .B1(n18530), .B2(n18293), .ZN(
        n18289) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18294), .B1(
        n18583), .B2(n18361), .ZN(n18288) );
  OAI211_X1 U21379 ( .C1(n18533), .C2(n18311), .A(n18289), .B(n18288), .ZN(
        P3_U2905) );
  AOI22_X1 U21380 ( .A1(n18535), .A2(n18293), .B1(n18587), .B2(n18292), .ZN(
        n18291) );
  AOI22_X1 U21381 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18294), .B1(
        n18590), .B2(n18361), .ZN(n18290) );
  OAI211_X1 U21382 ( .C1(n18538), .C2(n18311), .A(n18291), .B(n18290), .ZN(
        P3_U2906) );
  AOI22_X1 U21383 ( .A1(n18598), .A2(n18293), .B1(n18596), .B2(n18292), .ZN(
        n18296) );
  AOI22_X1 U21384 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18294), .B1(
        n18599), .B2(n18361), .ZN(n18295) );
  OAI211_X1 U21385 ( .C1(n18604), .C2(n18311), .A(n18296), .B(n18295), .ZN(
        P3_U2907) );
  NOR2_X1 U21386 ( .A1(n18386), .A2(n18343), .ZN(n18314) );
  AOI22_X1 U21387 ( .A1(n18548), .A2(n18337), .B1(n18547), .B2(n18314), .ZN(
        n18300) );
  AOI22_X1 U21388 ( .A1(n18552), .A2(n18298), .B1(n18297), .B2(n18341), .ZN(
        n18316) );
  NOR2_X2 U21389 ( .A1(n18390), .A2(n18343), .ZN(n18376) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18316), .B1(
        n18553), .B2(n18376), .ZN(n18299) );
  OAI211_X1 U21391 ( .C1(n18556), .C2(n18311), .A(n18300), .B(n18299), .ZN(
        P3_U2908) );
  AOI22_X1 U21392 ( .A1(n18558), .A2(n18315), .B1(n18557), .B2(n18314), .ZN(
        n18302) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18316), .B1(
        n18559), .B2(n18376), .ZN(n18301) );
  OAI211_X1 U21394 ( .C1(n18562), .C2(n18335), .A(n18302), .B(n18301), .ZN(
        P3_U2909) );
  AOI22_X1 U21395 ( .A1(n18520), .A2(n18337), .B1(n18563), .B2(n18314), .ZN(
        n18304) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18316), .B1(
        n18565), .B2(n18376), .ZN(n18303) );
  OAI211_X1 U21397 ( .C1(n18523), .C2(n18311), .A(n18304), .B(n18303), .ZN(
        P3_U2910) );
  AOI22_X1 U21398 ( .A1(n18569), .A2(n18314), .B1(n18570), .B2(n18337), .ZN(
        n18306) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18316), .B1(
        n18571), .B2(n18376), .ZN(n18305) );
  OAI211_X1 U21400 ( .C1(n18574), .C2(n18311), .A(n18306), .B(n18305), .ZN(
        P3_U2911) );
  AOI22_X1 U21401 ( .A1(n18576), .A2(n18337), .B1(n18575), .B2(n18314), .ZN(
        n18308) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18316), .B1(
        n18577), .B2(n18376), .ZN(n18307) );
  OAI211_X1 U21403 ( .C1(n18580), .C2(n18311), .A(n18308), .B(n18307), .ZN(
        P3_U2912) );
  AOI22_X1 U21404 ( .A1(n18582), .A2(n18337), .B1(n18581), .B2(n18314), .ZN(
        n18310) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18316), .B1(
        n18583), .B2(n18376), .ZN(n18309) );
  OAI211_X1 U21406 ( .C1(n18586), .C2(n18311), .A(n18310), .B(n18309), .ZN(
        P3_U2913) );
  AOI22_X1 U21407 ( .A1(n18535), .A2(n18315), .B1(n18587), .B2(n18314), .ZN(
        n18313) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18316), .B1(
        n18590), .B2(n18376), .ZN(n18312) );
  OAI211_X1 U21409 ( .C1(n18538), .C2(n18335), .A(n18313), .B(n18312), .ZN(
        P3_U2914) );
  AOI22_X1 U21410 ( .A1(n18598), .A2(n18315), .B1(n18596), .B2(n18314), .ZN(
        n18318) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18316), .B1(
        n18599), .B2(n18376), .ZN(n18317) );
  OAI211_X1 U21412 ( .C1(n18604), .C2(n18335), .A(n18318), .B(n18317), .ZN(
        P3_U2915) );
  NOR3_X1 U21413 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n18387), .ZN(n18393) );
  INV_X1 U21414 ( .A(n18393), .ZN(n18402) );
  INV_X1 U21415 ( .A(n18402), .ZN(n18403) );
  NOR2_X1 U21416 ( .A1(n18376), .A2(n18403), .ZN(n18364) );
  NOR2_X1 U21417 ( .A1(n18509), .A2(n18364), .ZN(n18336) );
  AOI22_X1 U21418 ( .A1(n18548), .A2(n18361), .B1(n18547), .B2(n18336), .ZN(
        n18322) );
  OAI21_X1 U21419 ( .B1(n18319), .B2(n18512), .A(n18364), .ZN(n18320) );
  OAI211_X1 U21420 ( .C1(n18403), .C2(n18515), .A(n18463), .B(n18320), .ZN(
        n18338) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18338), .B1(
        n18553), .B2(n18393), .ZN(n18321) );
  OAI211_X1 U21422 ( .C1(n18556), .C2(n18335), .A(n18322), .B(n18321), .ZN(
        P3_U2916) );
  AOI22_X1 U21423 ( .A1(n18557), .A2(n18336), .B1(n18441), .B2(n18361), .ZN(
        n18324) );
  AOI22_X1 U21424 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18338), .B1(
        n18559), .B2(n18393), .ZN(n18323) );
  OAI211_X1 U21425 ( .C1(n18444), .C2(n18335), .A(n18324), .B(n18323), .ZN(
        P3_U2917) );
  INV_X1 U21426 ( .A(n18361), .ZN(n18358) );
  AOI22_X1 U21427 ( .A1(n18564), .A2(n18337), .B1(n18563), .B2(n18336), .ZN(
        n18326) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18338), .B1(
        n18565), .B2(n18403), .ZN(n18325) );
  OAI211_X1 U21429 ( .C1(n18568), .C2(n18358), .A(n18326), .B(n18325), .ZN(
        P3_U2918) );
  AOI22_X1 U21430 ( .A1(n18524), .A2(n18337), .B1(n18569), .B2(n18336), .ZN(
        n18328) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18338), .B1(
        n18571), .B2(n18393), .ZN(n18327) );
  OAI211_X1 U21432 ( .C1(n18527), .C2(n18358), .A(n18328), .B(n18327), .ZN(
        P3_U2919) );
  AOI22_X1 U21433 ( .A1(n18449), .A2(n18337), .B1(n18575), .B2(n18336), .ZN(
        n18330) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18338), .B1(
        n18577), .B2(n18403), .ZN(n18329) );
  OAI211_X1 U21435 ( .C1(n18452), .C2(n18358), .A(n18330), .B(n18329), .ZN(
        P3_U2920) );
  AOI22_X1 U21436 ( .A1(n18581), .A2(n18336), .B1(n18530), .B2(n18337), .ZN(
        n18332) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18338), .B1(
        n18583), .B2(n18403), .ZN(n18331) );
  OAI211_X1 U21438 ( .C1(n18533), .C2(n18358), .A(n18332), .B(n18331), .ZN(
        P3_U2921) );
  AOI22_X1 U21439 ( .A1(n18588), .A2(n18361), .B1(n18587), .B2(n18336), .ZN(
        n18334) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18338), .B1(
        n18590), .B2(n18403), .ZN(n18333) );
  OAI211_X1 U21441 ( .C1(n18594), .C2(n18335), .A(n18334), .B(n18333), .ZN(
        P3_U2922) );
  AOI22_X1 U21442 ( .A1(n18598), .A2(n18337), .B1(n18596), .B2(n18336), .ZN(
        n18340) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18338), .B1(
        n18599), .B2(n18403), .ZN(n18339) );
  OAI211_X1 U21444 ( .C1(n18604), .C2(n18358), .A(n18340), .B(n18339), .ZN(
        P3_U2923) );
  NAND2_X1 U21445 ( .A1(n18342), .A2(n18341), .ZN(n18360) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18360), .B1(
        n18547), .B2(n18359), .ZN(n18345) );
  NOR2_X2 U21447 ( .A1(n18644), .A2(n18343), .ZN(n18425) );
  AOI22_X1 U21448 ( .A1(n18548), .A2(n18376), .B1(n18553), .B2(n18425), .ZN(
        n18344) );
  OAI211_X1 U21449 ( .C1(n18556), .C2(n18358), .A(n18345), .B(n18344), .ZN(
        P3_U2924) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18360), .B1(
        n18557), .B2(n18359), .ZN(n18347) );
  AOI22_X1 U21451 ( .A1(n18559), .A2(n18425), .B1(n18441), .B2(n18376), .ZN(
        n18346) );
  OAI211_X1 U21452 ( .C1(n18444), .C2(n18358), .A(n18347), .B(n18346), .ZN(
        P3_U2925) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18360), .B1(
        n18563), .B2(n18359), .ZN(n18349) );
  AOI22_X1 U21454 ( .A1(n18520), .A2(n18376), .B1(n18565), .B2(n18425), .ZN(
        n18348) );
  OAI211_X1 U21455 ( .C1(n18523), .C2(n18358), .A(n18349), .B(n18348), .ZN(
        P3_U2926) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18360), .B1(
        n18569), .B2(n18359), .ZN(n18351) );
  AOI22_X1 U21457 ( .A1(n18571), .A2(n18425), .B1(n18570), .B2(n18376), .ZN(
        n18350) );
  OAI211_X1 U21458 ( .C1(n18574), .C2(n18358), .A(n18351), .B(n18350), .ZN(
        P3_U2927) );
  INV_X1 U21459 ( .A(n18376), .ZN(n18385) );
  AOI22_X1 U21460 ( .A1(n18449), .A2(n18361), .B1(n18575), .B2(n18359), .ZN(
        n18353) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18360), .B1(
        n18577), .B2(n18425), .ZN(n18352) );
  OAI211_X1 U21462 ( .C1(n18452), .C2(n18385), .A(n18353), .B(n18352), .ZN(
        P3_U2928) );
  AOI22_X1 U21463 ( .A1(n18582), .A2(n18376), .B1(n18581), .B2(n18359), .ZN(
        n18355) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18360), .B1(
        n18583), .B2(n18425), .ZN(n18354) );
  OAI211_X1 U21465 ( .C1(n18586), .C2(n18358), .A(n18355), .B(n18354), .ZN(
        P3_U2929) );
  AOI22_X1 U21466 ( .A1(n18588), .A2(n18376), .B1(n18587), .B2(n18359), .ZN(
        n18357) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18360), .B1(
        n18590), .B2(n18425), .ZN(n18356) );
  OAI211_X1 U21468 ( .C1(n18594), .C2(n18358), .A(n18357), .B(n18356), .ZN(
        P3_U2930) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18360), .B1(
        n18596), .B2(n18359), .ZN(n18363) );
  AOI22_X1 U21470 ( .A1(n18599), .A2(n18425), .B1(n18598), .B2(n18361), .ZN(
        n18362) );
  OAI211_X1 U21471 ( .C1(n18604), .C2(n18385), .A(n18363), .B(n18362), .ZN(
        P3_U2931) );
  NOR2_X2 U21472 ( .A1(n18646), .A2(n18438), .ZN(n18455) );
  NOR2_X1 U21473 ( .A1(n18425), .A2(n18455), .ZN(n18414) );
  NOR2_X1 U21474 ( .A1(n18509), .A2(n18414), .ZN(n18381) );
  AOI22_X1 U21475 ( .A1(n18413), .A2(n18376), .B1(n18547), .B2(n18381), .ZN(
        n18367) );
  OAI21_X1 U21476 ( .B1(n18364), .B2(n18512), .A(n18414), .ZN(n18365) );
  OAI211_X1 U21477 ( .C1(n18455), .C2(n18515), .A(n18463), .B(n18365), .ZN(
        n18382) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18382), .B1(
        n18553), .B2(n18455), .ZN(n18366) );
  OAI211_X1 U21479 ( .C1(n18418), .C2(n18402), .A(n18367), .B(n18366), .ZN(
        P3_U2932) );
  AOI22_X1 U21480 ( .A1(n18558), .A2(n18376), .B1(n18557), .B2(n18381), .ZN(
        n18369) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18382), .B1(
        n18559), .B2(n18455), .ZN(n18368) );
  OAI211_X1 U21482 ( .C1(n18562), .C2(n18402), .A(n18369), .B(n18368), .ZN(
        P3_U2933) );
  AOI22_X1 U21483 ( .A1(n18520), .A2(n18393), .B1(n18563), .B2(n18381), .ZN(
        n18371) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18382), .B1(
        n18565), .B2(n18455), .ZN(n18370) );
  OAI211_X1 U21485 ( .C1(n18523), .C2(n18385), .A(n18371), .B(n18370), .ZN(
        P3_U2934) );
  AOI22_X1 U21486 ( .A1(n18524), .A2(n18376), .B1(n18569), .B2(n18381), .ZN(
        n18373) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18382), .B1(
        n18571), .B2(n18455), .ZN(n18372) );
  OAI211_X1 U21488 ( .C1(n18527), .C2(n18402), .A(n18373), .B(n18372), .ZN(
        P3_U2935) );
  AOI22_X1 U21489 ( .A1(n18576), .A2(n18403), .B1(n18575), .B2(n18381), .ZN(
        n18375) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18382), .B1(
        n18577), .B2(n18455), .ZN(n18374) );
  OAI211_X1 U21491 ( .C1(n18580), .C2(n18385), .A(n18375), .B(n18374), .ZN(
        P3_U2936) );
  AOI22_X1 U21492 ( .A1(n18581), .A2(n18381), .B1(n18530), .B2(n18376), .ZN(
        n18378) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18382), .B1(
        n18583), .B2(n18455), .ZN(n18377) );
  OAI211_X1 U21494 ( .C1(n18533), .C2(n18402), .A(n18378), .B(n18377), .ZN(
        P3_U2937) );
  AOI22_X1 U21495 ( .A1(n18588), .A2(n18403), .B1(n18587), .B2(n18381), .ZN(
        n18380) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18382), .B1(
        n18590), .B2(n18455), .ZN(n18379) );
  OAI211_X1 U21497 ( .C1(n18594), .C2(n18385), .A(n18380), .B(n18379), .ZN(
        P3_U2938) );
  AOI22_X1 U21498 ( .A1(n18540), .A2(n18403), .B1(n18596), .B2(n18381), .ZN(
        n18384) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18382), .B1(
        n18599), .B2(n18455), .ZN(n18383) );
  OAI211_X1 U21500 ( .C1(n18546), .C2(n18385), .A(n18384), .B(n18383), .ZN(
        P3_U2939) );
  INV_X1 U21501 ( .A(n18425), .ZN(n18436) );
  NOR2_X1 U21502 ( .A1(n18386), .A2(n18438), .ZN(n18408) );
  AOI22_X1 U21503 ( .A1(n18413), .A2(n18393), .B1(n18547), .B2(n18408), .ZN(
        n18392) );
  NOR2_X1 U21504 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18387), .ZN(
        n18389) );
  INV_X1 U21505 ( .A(n18388), .ZN(n18549) );
  NOR2_X1 U21506 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18438), .ZN(
        n18437) );
  AOI22_X1 U21507 ( .A1(n18552), .A2(n18389), .B1(n18549), .B2(n18437), .ZN(
        n18409) );
  NOR2_X2 U21508 ( .A1(n18390), .A2(n18438), .ZN(n18477) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18409), .B1(
        n18553), .B2(n18477), .ZN(n18391) );
  OAI211_X1 U21510 ( .C1(n18418), .C2(n18436), .A(n18392), .B(n18391), .ZN(
        P3_U2940) );
  AOI22_X1 U21511 ( .A1(n18558), .A2(n18393), .B1(n18557), .B2(n18408), .ZN(
        n18395) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18409), .B1(
        n18559), .B2(n18477), .ZN(n18394) );
  OAI211_X1 U21513 ( .C1(n18562), .C2(n18436), .A(n18395), .B(n18394), .ZN(
        P3_U2941) );
  AOI22_X1 U21514 ( .A1(n18564), .A2(n18403), .B1(n18563), .B2(n18408), .ZN(
        n18397) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18409), .B1(
        n18565), .B2(n18477), .ZN(n18396) );
  OAI211_X1 U21516 ( .C1(n18568), .C2(n18436), .A(n18397), .B(n18396), .ZN(
        P3_U2942) );
  AOI22_X1 U21517 ( .A1(n18569), .A2(n18408), .B1(n18570), .B2(n18425), .ZN(
        n18399) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18409), .B1(
        n18571), .B2(n18477), .ZN(n18398) );
  OAI211_X1 U21519 ( .C1(n18574), .C2(n18402), .A(n18399), .B(n18398), .ZN(
        P3_U2943) );
  AOI22_X1 U21520 ( .A1(n18576), .A2(n18425), .B1(n18575), .B2(n18408), .ZN(
        n18401) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18409), .B1(
        n18577), .B2(n18477), .ZN(n18400) );
  OAI211_X1 U21522 ( .C1(n18580), .C2(n18402), .A(n18401), .B(n18400), .ZN(
        P3_U2944) );
  AOI22_X1 U21523 ( .A1(n18581), .A2(n18408), .B1(n18530), .B2(n18403), .ZN(
        n18405) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18409), .B1(
        n18583), .B2(n18477), .ZN(n18404) );
  OAI211_X1 U21525 ( .C1(n18533), .C2(n18436), .A(n18405), .B(n18404), .ZN(
        P3_U2945) );
  AOI22_X1 U21526 ( .A1(n18535), .A2(n18403), .B1(n18587), .B2(n18408), .ZN(
        n18407) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18409), .B1(
        n18590), .B2(n18477), .ZN(n18406) );
  OAI211_X1 U21528 ( .C1(n18538), .C2(n18436), .A(n18407), .B(n18406), .ZN(
        P3_U2946) );
  AOI22_X1 U21529 ( .A1(n18598), .A2(n18403), .B1(n18596), .B2(n18408), .ZN(
        n18411) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18409), .B1(
        n18599), .B2(n18477), .ZN(n18410) );
  OAI211_X1 U21531 ( .C1(n18604), .C2(n18436), .A(n18411), .B(n18410), .ZN(
        P3_U2947) );
  INV_X1 U21532 ( .A(n18455), .ZN(n18462) );
  NOR2_X1 U21533 ( .A1(n18645), .A2(n18438), .ZN(n18488) );
  NAND2_X1 U21534 ( .A1(n18412), .A2(n18488), .ZN(n18501) );
  NOR2_X1 U21535 ( .A1(n18477), .A2(n18505), .ZN(n18465) );
  NOR2_X1 U21536 ( .A1(n18509), .A2(n18465), .ZN(n18432) );
  AOI22_X1 U21537 ( .A1(n18413), .A2(n18425), .B1(n18547), .B2(n18432), .ZN(
        n18417) );
  OAI21_X1 U21538 ( .B1(n18414), .B2(n18512), .A(n18465), .ZN(n18415) );
  OAI211_X1 U21539 ( .C1(n18505), .C2(n18515), .A(n18463), .B(n18415), .ZN(
        n18433) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18433), .B1(
        n18553), .B2(n18505), .ZN(n18416) );
  OAI211_X1 U21541 ( .C1(n18418), .C2(n18462), .A(n18417), .B(n18416), .ZN(
        P3_U2948) );
  AOI22_X1 U21542 ( .A1(n18557), .A2(n18432), .B1(n18441), .B2(n18455), .ZN(
        n18420) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18433), .B1(
        n18559), .B2(n18505), .ZN(n18419) );
  OAI211_X1 U21544 ( .C1(n18444), .C2(n18436), .A(n18420), .B(n18419), .ZN(
        P3_U2949) );
  AOI22_X1 U21545 ( .A1(n18564), .A2(n18425), .B1(n18563), .B2(n18432), .ZN(
        n18422) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18433), .B1(
        n18565), .B2(n18505), .ZN(n18421) );
  OAI211_X1 U21547 ( .C1(n18568), .C2(n18462), .A(n18422), .B(n18421), .ZN(
        P3_U2950) );
  AOI22_X1 U21548 ( .A1(n18524), .A2(n18425), .B1(n18569), .B2(n18432), .ZN(
        n18424) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18433), .B1(
        n18571), .B2(n18505), .ZN(n18423) );
  OAI211_X1 U21550 ( .C1(n18527), .C2(n18462), .A(n18424), .B(n18423), .ZN(
        P3_U2951) );
  AOI22_X1 U21551 ( .A1(n18449), .A2(n18425), .B1(n18575), .B2(n18432), .ZN(
        n18427) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18433), .B1(
        n18577), .B2(n18505), .ZN(n18426) );
  OAI211_X1 U21553 ( .C1(n18452), .C2(n18462), .A(n18427), .B(n18426), .ZN(
        P3_U2952) );
  AOI22_X1 U21554 ( .A1(n18582), .A2(n18455), .B1(n18581), .B2(n18432), .ZN(
        n18429) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18433), .B1(
        n18583), .B2(n18505), .ZN(n18428) );
  OAI211_X1 U21556 ( .C1(n18586), .C2(n18436), .A(n18429), .B(n18428), .ZN(
        P3_U2953) );
  AOI22_X1 U21557 ( .A1(n18588), .A2(n18455), .B1(n18587), .B2(n18432), .ZN(
        n18431) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18433), .B1(
        n18590), .B2(n18505), .ZN(n18430) );
  OAI211_X1 U21559 ( .C1(n18594), .C2(n18436), .A(n18431), .B(n18430), .ZN(
        P3_U2954) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18433), .B1(
        n18596), .B2(n18432), .ZN(n18435) );
  AOI22_X1 U21561 ( .A1(n18540), .A2(n18455), .B1(n18599), .B2(n18505), .ZN(
        n18434) );
  OAI211_X1 U21562 ( .C1(n18546), .C2(n18436), .A(n18435), .B(n18434), .ZN(
        P3_U2955) );
  AND2_X1 U21563 ( .A1(n18674), .A2(n18488), .ZN(n18458) );
  AOI22_X1 U21564 ( .A1(n18548), .A2(n18477), .B1(n18547), .B2(n18458), .ZN(
        n18440) );
  AOI22_X1 U21565 ( .A1(n18552), .A2(n18437), .B1(n18549), .B2(n18488), .ZN(
        n18459) );
  NOR2_X2 U21566 ( .A1(n18644), .A2(n18438), .ZN(n18534) );
  AOI22_X1 U21567 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18459), .B1(
        n18553), .B2(n18534), .ZN(n18439) );
  OAI211_X1 U21568 ( .C1(n18556), .C2(n18462), .A(n18440), .B(n18439), .ZN(
        P3_U2956) );
  AOI22_X1 U21569 ( .A1(n18557), .A2(n18458), .B1(n18441), .B2(n18477), .ZN(
        n18443) );
  AOI22_X1 U21570 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18459), .B1(
        n18559), .B2(n18534), .ZN(n18442) );
  OAI211_X1 U21571 ( .C1(n18444), .C2(n18462), .A(n18443), .B(n18442), .ZN(
        P3_U2957) );
  AOI22_X1 U21572 ( .A1(n18520), .A2(n18477), .B1(n18563), .B2(n18458), .ZN(
        n18446) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18459), .B1(
        n18565), .B2(n18534), .ZN(n18445) );
  OAI211_X1 U21574 ( .C1(n18523), .C2(n18462), .A(n18446), .B(n18445), .ZN(
        P3_U2958) );
  AOI22_X1 U21575 ( .A1(n18569), .A2(n18458), .B1(n18570), .B2(n18477), .ZN(
        n18448) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18459), .B1(
        n18571), .B2(n18534), .ZN(n18447) );
  OAI211_X1 U21577 ( .C1(n18574), .C2(n18462), .A(n18448), .B(n18447), .ZN(
        P3_U2959) );
  INV_X1 U21578 ( .A(n18477), .ZN(n18486) );
  AOI22_X1 U21579 ( .A1(n18449), .A2(n18455), .B1(n18575), .B2(n18458), .ZN(
        n18451) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18459), .B1(
        n18577), .B2(n18534), .ZN(n18450) );
  OAI211_X1 U21581 ( .C1(n18452), .C2(n18486), .A(n18451), .B(n18450), .ZN(
        P3_U2960) );
  AOI22_X1 U21582 ( .A1(n18582), .A2(n18477), .B1(n18581), .B2(n18458), .ZN(
        n18454) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18459), .B1(
        n18583), .B2(n18534), .ZN(n18453) );
  OAI211_X1 U21584 ( .C1(n18586), .C2(n18462), .A(n18454), .B(n18453), .ZN(
        P3_U2961) );
  AOI22_X1 U21585 ( .A1(n18535), .A2(n18455), .B1(n18587), .B2(n18458), .ZN(
        n18457) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18459), .B1(
        n18590), .B2(n18534), .ZN(n18456) );
  OAI211_X1 U21587 ( .C1(n18538), .C2(n18486), .A(n18457), .B(n18456), .ZN(
        P3_U2962) );
  AOI22_X1 U21588 ( .A1(n18540), .A2(n18477), .B1(n18596), .B2(n18458), .ZN(
        n18461) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18459), .B1(
        n18599), .B2(n18534), .ZN(n18460) );
  OAI211_X1 U21590 ( .C1(n18546), .C2(n18462), .A(n18461), .B(n18460), .ZN(
        P3_U2963) );
  INV_X1 U21591 ( .A(n18534), .ZN(n18545) );
  INV_X1 U21592 ( .A(n18551), .ZN(n18487) );
  NOR2_X2 U21593 ( .A1(n18487), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18597) );
  INV_X1 U21594 ( .A(n18597), .ZN(n18593) );
  AOI21_X1 U21595 ( .B1(n18545), .B2(n18593), .A(n18509), .ZN(n18482) );
  AOI22_X1 U21596 ( .A1(n18548), .A2(n18505), .B1(n18547), .B2(n18482), .ZN(
        n18468) );
  OAI21_X1 U21597 ( .B1(n18534), .B2(n18597), .A(n18463), .ZN(n18511) );
  OAI21_X1 U21598 ( .B1(n18465), .B2(n18464), .A(n18511), .ZN(n18466) );
  OAI21_X1 U21599 ( .B1(n18597), .B2(n18515), .A(n18466), .ZN(n18483) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18483), .B1(
        n18553), .B2(n18597), .ZN(n18467) );
  OAI211_X1 U21601 ( .C1(n18556), .C2(n18486), .A(n18468), .B(n18467), .ZN(
        P3_U2964) );
  AOI22_X1 U21602 ( .A1(n18558), .A2(n18477), .B1(n18557), .B2(n18482), .ZN(
        n18470) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18483), .B1(
        n18559), .B2(n18597), .ZN(n18469) );
  OAI211_X1 U21604 ( .C1(n18562), .C2(n18501), .A(n18470), .B(n18469), .ZN(
        P3_U2965) );
  AOI22_X1 U21605 ( .A1(n18520), .A2(n18505), .B1(n18563), .B2(n18482), .ZN(
        n18472) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18483), .B1(
        n18565), .B2(n18597), .ZN(n18471) );
  OAI211_X1 U21607 ( .C1(n18523), .C2(n18486), .A(n18472), .B(n18471), .ZN(
        P3_U2966) );
  AOI22_X1 U21608 ( .A1(n18524), .A2(n18477), .B1(n18569), .B2(n18482), .ZN(
        n18474) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18483), .B1(
        n18571), .B2(n18597), .ZN(n18473) );
  OAI211_X1 U21610 ( .C1(n18527), .C2(n18501), .A(n18474), .B(n18473), .ZN(
        P3_U2967) );
  AOI22_X1 U21611 ( .A1(n18576), .A2(n18505), .B1(n18575), .B2(n18482), .ZN(
        n18476) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18483), .B1(
        n18577), .B2(n18597), .ZN(n18475) );
  OAI211_X1 U21613 ( .C1(n18580), .C2(n18486), .A(n18476), .B(n18475), .ZN(
        P3_U2968) );
  AOI22_X1 U21614 ( .A1(n18581), .A2(n18482), .B1(n18530), .B2(n18477), .ZN(
        n18479) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18483), .B1(
        n18583), .B2(n18597), .ZN(n18478) );
  OAI211_X1 U21616 ( .C1(n18533), .C2(n18501), .A(n18479), .B(n18478), .ZN(
        P3_U2969) );
  AOI22_X1 U21617 ( .A1(n18588), .A2(n18505), .B1(n18587), .B2(n18482), .ZN(
        n18481) );
  AOI22_X1 U21618 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18483), .B1(
        n18590), .B2(n18597), .ZN(n18480) );
  OAI211_X1 U21619 ( .C1(n18594), .C2(n18486), .A(n18481), .B(n18480), .ZN(
        P3_U2970) );
  AOI22_X1 U21620 ( .A1(n18540), .A2(n18505), .B1(n18596), .B2(n18482), .ZN(
        n18485) );
  AOI22_X1 U21621 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18483), .B1(
        n18599), .B2(n18597), .ZN(n18484) );
  OAI211_X1 U21622 ( .C1(n18546), .C2(n18486), .A(n18485), .B(n18484), .ZN(
        P3_U2971) );
  NOR2_X1 U21623 ( .A1(n18509), .A2(n18487), .ZN(n18504) );
  AOI22_X1 U21624 ( .A1(n18548), .A2(n18534), .B1(n18547), .B2(n18504), .ZN(
        n18490) );
  AOI22_X1 U21625 ( .A1(n18552), .A2(n18488), .B1(n18551), .B2(n18549), .ZN(
        n18506) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18506), .B1(
        n18589), .B2(n18553), .ZN(n18489) );
  OAI211_X1 U21627 ( .C1(n18556), .C2(n18501), .A(n18490), .B(n18489), .ZN(
        P3_U2972) );
  AOI22_X1 U21628 ( .A1(n18558), .A2(n18505), .B1(n18557), .B2(n18504), .ZN(
        n18492) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18506), .B1(
        n18589), .B2(n18559), .ZN(n18491) );
  OAI211_X1 U21630 ( .C1(n18562), .C2(n18545), .A(n18492), .B(n18491), .ZN(
        P3_U2973) );
  AOI22_X1 U21631 ( .A1(n18520), .A2(n18534), .B1(n18563), .B2(n18504), .ZN(
        n18494) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18506), .B1(
        n18589), .B2(n18565), .ZN(n18493) );
  OAI211_X1 U21633 ( .C1(n18523), .C2(n18501), .A(n18494), .B(n18493), .ZN(
        P3_U2974) );
  AOI22_X1 U21634 ( .A1(n18524), .A2(n18505), .B1(n18569), .B2(n18504), .ZN(
        n18496) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18506), .B1(
        n18589), .B2(n18571), .ZN(n18495) );
  OAI211_X1 U21636 ( .C1(n18527), .C2(n18545), .A(n18496), .B(n18495), .ZN(
        P3_U2975) );
  AOI22_X1 U21637 ( .A1(n18576), .A2(n18534), .B1(n18575), .B2(n18504), .ZN(
        n18498) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18506), .B1(
        n18589), .B2(n18577), .ZN(n18497) );
  OAI211_X1 U21639 ( .C1(n18580), .C2(n18501), .A(n18498), .B(n18497), .ZN(
        P3_U2976) );
  AOI22_X1 U21640 ( .A1(n18582), .A2(n18534), .B1(n18581), .B2(n18504), .ZN(
        n18500) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18506), .B1(
        n18589), .B2(n18583), .ZN(n18499) );
  OAI211_X1 U21642 ( .C1(n18586), .C2(n18501), .A(n18500), .B(n18499), .ZN(
        P3_U2977) );
  AOI22_X1 U21643 ( .A1(n18535), .A2(n18505), .B1(n18587), .B2(n18504), .ZN(
        n18503) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18506), .B1(
        n18589), .B2(n18590), .ZN(n18502) );
  OAI211_X1 U21645 ( .C1(n18538), .C2(n18545), .A(n18503), .B(n18502), .ZN(
        P3_U2978) );
  AOI22_X1 U21646 ( .A1(n18598), .A2(n18505), .B1(n18596), .B2(n18504), .ZN(
        n18508) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18506), .B1(
        n18589), .B2(n18599), .ZN(n18507) );
  OAI211_X1 U21648 ( .C1(n18604), .C2(n18545), .A(n18508), .B(n18507), .ZN(
        P3_U2979) );
  AOI21_X1 U21649 ( .B1(n18510), .B2(n18605), .A(n18509), .ZN(n18539) );
  AOI22_X1 U21650 ( .A1(n18548), .A2(n18597), .B1(n18547), .B2(n18539), .ZN(
        n18517) );
  NOR2_X1 U21651 ( .A1(n18512), .A2(n18511), .ZN(n18513) );
  OAI22_X1 U21652 ( .A1(n18541), .A2(n18515), .B1(n18514), .B2(n18513), .ZN(
        n18542) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18553), .ZN(n18516) );
  OAI211_X1 U21654 ( .C1(n18556), .C2(n18545), .A(n18517), .B(n18516), .ZN(
        P3_U2980) );
  AOI22_X1 U21655 ( .A1(n18558), .A2(n18534), .B1(n18557), .B2(n18539), .ZN(
        n18519) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18559), .ZN(n18518) );
  OAI211_X1 U21657 ( .C1(n18562), .C2(n18593), .A(n18519), .B(n18518), .ZN(
        P3_U2981) );
  AOI22_X1 U21658 ( .A1(n18520), .A2(n18597), .B1(n18563), .B2(n18539), .ZN(
        n18522) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18565), .ZN(n18521) );
  OAI211_X1 U21660 ( .C1(n18523), .C2(n18545), .A(n18522), .B(n18521), .ZN(
        P3_U2982) );
  AOI22_X1 U21661 ( .A1(n18524), .A2(n18534), .B1(n18569), .B2(n18539), .ZN(
        n18526) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18571), .ZN(n18525) );
  OAI211_X1 U21663 ( .C1(n18527), .C2(n18593), .A(n18526), .B(n18525), .ZN(
        P3_U2983) );
  AOI22_X1 U21664 ( .A1(n18576), .A2(n18597), .B1(n18575), .B2(n18539), .ZN(
        n18529) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18577), .ZN(n18528) );
  OAI211_X1 U21666 ( .C1(n18580), .C2(n18545), .A(n18529), .B(n18528), .ZN(
        P3_U2984) );
  AOI22_X1 U21667 ( .A1(n18581), .A2(n18539), .B1(n18530), .B2(n18534), .ZN(
        n18532) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18583), .ZN(n18531) );
  OAI211_X1 U21669 ( .C1(n18533), .C2(n18593), .A(n18532), .B(n18531), .ZN(
        P3_U2985) );
  AOI22_X1 U21670 ( .A1(n18535), .A2(n18534), .B1(n18587), .B2(n18539), .ZN(
        n18537) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18590), .ZN(n18536) );
  OAI211_X1 U21672 ( .C1(n18538), .C2(n18593), .A(n18537), .B(n18536), .ZN(
        P3_U2986) );
  AOI22_X1 U21673 ( .A1(n18540), .A2(n18597), .B1(n18596), .B2(n18539), .ZN(
        n18544) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18542), .B1(
        n18541), .B2(n18599), .ZN(n18543) );
  OAI211_X1 U21675 ( .C1(n18546), .C2(n18545), .A(n18544), .B(n18543), .ZN(
        P3_U2987) );
  AND2_X1 U21676 ( .A1(n18674), .A2(n18550), .ZN(n18595) );
  AOI22_X1 U21677 ( .A1(n18548), .A2(n18589), .B1(n18547), .B2(n18595), .ZN(
        n18555) );
  AOI22_X1 U21678 ( .A1(n18552), .A2(n18551), .B1(n18550), .B2(n18549), .ZN(
        n18601) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18601), .B1(
        n18600), .B2(n18553), .ZN(n18554) );
  OAI211_X1 U21680 ( .C1(n18556), .C2(n18593), .A(n18555), .B(n18554), .ZN(
        P3_U2988) );
  AOI22_X1 U21681 ( .A1(n18558), .A2(n18597), .B1(n18557), .B2(n18595), .ZN(
        n18561) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18601), .B1(
        n18600), .B2(n18559), .ZN(n18560) );
  OAI211_X1 U21683 ( .C1(n18605), .C2(n18562), .A(n18561), .B(n18560), .ZN(
        P3_U2989) );
  AOI22_X1 U21684 ( .A1(n18564), .A2(n18597), .B1(n18563), .B2(n18595), .ZN(
        n18567) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18601), .B1(
        n18600), .B2(n18565), .ZN(n18566) );
  OAI211_X1 U21686 ( .C1(n18605), .C2(n18568), .A(n18567), .B(n18566), .ZN(
        P3_U2990) );
  AOI22_X1 U21687 ( .A1(n18589), .A2(n18570), .B1(n18569), .B2(n18595), .ZN(
        n18573) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18601), .B1(
        n18600), .B2(n18571), .ZN(n18572) );
  OAI211_X1 U21689 ( .C1(n18574), .C2(n18593), .A(n18573), .B(n18572), .ZN(
        P3_U2991) );
  AOI22_X1 U21690 ( .A1(n18589), .A2(n18576), .B1(n18575), .B2(n18595), .ZN(
        n18579) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18601), .B1(
        n18600), .B2(n18577), .ZN(n18578) );
  OAI211_X1 U21692 ( .C1(n18580), .C2(n18593), .A(n18579), .B(n18578), .ZN(
        P3_U2992) );
  AOI22_X1 U21693 ( .A1(n18589), .A2(n18582), .B1(n18581), .B2(n18595), .ZN(
        n18585) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18601), .B1(
        n18600), .B2(n18583), .ZN(n18584) );
  OAI211_X1 U21695 ( .C1(n18586), .C2(n18593), .A(n18585), .B(n18584), .ZN(
        P3_U2993) );
  AOI22_X1 U21696 ( .A1(n18589), .A2(n18588), .B1(n18587), .B2(n18595), .ZN(
        n18592) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18601), .B1(
        n18600), .B2(n18590), .ZN(n18591) );
  OAI211_X1 U21698 ( .C1(n18594), .C2(n18593), .A(n18592), .B(n18591), .ZN(
        P3_U2994) );
  AOI22_X1 U21699 ( .A1(n18598), .A2(n18597), .B1(n18596), .B2(n18595), .ZN(
        n18603) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18601), .B1(
        n18600), .B2(n18599), .ZN(n18602) );
  OAI211_X1 U21701 ( .C1(n18605), .C2(n18604), .A(n18603), .B(n18602), .ZN(
        P3_U2995) );
  AOI22_X1 U21702 ( .A1(n18609), .A2(n18608), .B1(n18607), .B2(n18606), .ZN(
        n18610) );
  OAI221_X1 U21703 ( .B1(n18613), .B2(n18612), .C1(n18613), .C2(n18611), .A(
        n18610), .ZN(n18807) );
  OAI21_X1 U21704 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18614), .ZN(n18616) );
  OAI211_X1 U21705 ( .C1(n18636), .C2(n18617), .A(n18616), .B(n18615), .ZN(
        n18659) );
  INV_X1 U21706 ( .A(n18636), .ZN(n18648) );
  AOI21_X1 U21707 ( .B1(n18637), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n18623), .ZN(n18640) );
  INV_X1 U21708 ( .A(n18640), .ZN(n18618) );
  AOI22_X1 U21709 ( .A1(n18619), .A2(n18618), .B1(n18635), .B2(n18624), .ZN(
        n18771) );
  OR2_X1 U21710 ( .A1(n18648), .A2(n18771), .ZN(n18628) );
  OAI21_X1 U21711 ( .B1(n18622), .B2(n18621), .A(n18620), .ZN(n18629) );
  AOI21_X1 U21712 ( .B1(n13971), .B2(n18623), .A(n18629), .ZN(n18625) );
  OAI21_X1 U21713 ( .B1(n18626), .B2(n18625), .A(n18624), .ZN(n18774) );
  NOR2_X1 U21714 ( .A1(n18648), .A2(n18774), .ZN(n18627) );
  MUX2_X1 U21715 ( .A(n18628), .B(n18627), .S(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n18657) );
  NAND3_X1 U21716 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18630), .A3(
        n18629), .ZN(n18631) );
  OAI221_X1 U21717 ( .B1(n18640), .B2(n18633), .C1(n18640), .C2(n18632), .A(
        n18631), .ZN(n18634) );
  AOI21_X1 U21718 ( .B1(n18635), .B2(n18780), .A(n18634), .ZN(n18782) );
  AOI22_X1 U21719 ( .A1(n18648), .A2(n10497), .B1(n18782), .B2(n18636), .ZN(
        n18652) );
  NOR2_X1 U21720 ( .A1(n18638), .A2(n18637), .ZN(n18643) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18639), .B1(
        n18643), .B2(n18796), .ZN(n18792) );
  OAI22_X1 U21722 ( .A1(n18643), .A2(n18642), .B1(n18641), .B2(n18640), .ZN(
        n18789) );
  AOI222_X1 U21723 ( .A1(n18792), .A2(n18789), .B1(n18792), .B2(n18645), .C1(
        n18789), .C2(n18644), .ZN(n18647) );
  OAI21_X1 U21724 ( .B1(n18648), .B2(n18647), .A(n18646), .ZN(n18651) );
  AND2_X1 U21725 ( .A1(n18652), .A2(n18651), .ZN(n18649) );
  OAI221_X1 U21726 ( .B1(n18652), .B2(n18651), .C1(n18650), .C2(n18649), .A(
        n18654), .ZN(n18656) );
  AOI21_X1 U21727 ( .B1(n18654), .B2(n18653), .A(n18652), .ZN(n18655) );
  AOI222_X1 U21728 ( .A1(n18657), .A2(n18656), .B1(n18657), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18656), .C2(n18655), .ZN(
        n18658) );
  NOR4_X1 U21729 ( .A1(n18660), .A2(n18807), .A3(n18659), .A4(n18658), .ZN(
        n18670) );
  INV_X1 U21730 ( .A(n18781), .ZN(n18791) );
  NOR2_X1 U21731 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18816) );
  AOI22_X1 U21732 ( .A1(n18791), .A2(n18816), .B1(n18693), .B2(n17412), .ZN(
        n18667) );
  NAND2_X1 U21733 ( .A1(n18693), .A2(n18661), .ZN(n18672) );
  OAI211_X1 U21734 ( .C1(P3_STATE2_REG_1__SCAN_IN), .C2(n18674), .A(n18672), 
        .B(n18662), .ZN(n18666) );
  OAI211_X1 U21735 ( .C1(n18665), .C2(n18664), .A(n18663), .B(n18670), .ZN(
        n18673) );
  NAND2_X1 U21736 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18673), .ZN(n18769) );
  OAI22_X1 U21737 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18667), .B1(n18666), 
        .B2(n18769), .ZN(n18668) );
  OAI21_X1 U21738 ( .B1(n18670), .B2(n18669), .A(n18668), .ZN(P3_U2996) );
  NAND2_X1 U21739 ( .A1(n18693), .A2(n17412), .ZN(n18678) );
  NOR3_X1 U21740 ( .A1(n18779), .A2(n18671), .A3(n18672), .ZN(n18681) );
  INV_X1 U21741 ( .A(n18681), .ZN(n18677) );
  NAND4_X1 U21742 ( .A1(n18675), .A2(n18674), .A3(n18673), .A4(n18672), .ZN(
        n18676) );
  NAND4_X1 U21743 ( .A1(n18679), .A2(n18678), .A3(n18677), .A4(n18676), .ZN(
        P3_U2997) );
  INV_X1 U21744 ( .A(n18680), .ZN(n18768) );
  NOR4_X1 U21745 ( .A1(n18816), .A2(n18682), .A3(n18768), .A4(n18681), .ZN(
        P3_U2998) );
  INV_X1 U21746 ( .A(n18767), .ZN(n18764) );
  AND2_X1 U21747 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18764), .ZN(
        P3_U2999) );
  AND2_X1 U21748 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18764), .ZN(
        P3_U3000) );
  AND2_X1 U21749 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18764), .ZN(
        P3_U3001) );
  AND2_X1 U21750 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18764), .ZN(
        P3_U3002) );
  AND2_X1 U21751 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18764), .ZN(
        P3_U3003) );
  AND2_X1 U21752 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18764), .ZN(
        P3_U3004) );
  AND2_X1 U21753 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18764), .ZN(
        P3_U3005) );
  AND2_X1 U21754 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18764), .ZN(
        P3_U3006) );
  AND2_X1 U21755 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18764), .ZN(
        P3_U3007) );
  AND2_X1 U21756 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18764), .ZN(
        P3_U3008) );
  AND2_X1 U21757 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18764), .ZN(
        P3_U3009) );
  AND2_X1 U21758 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18764), .ZN(
        P3_U3010) );
  AND2_X1 U21759 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18764), .ZN(
        P3_U3011) );
  AND2_X1 U21760 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18764), .ZN(
        P3_U3012) );
  AND2_X1 U21761 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18764), .ZN(
        P3_U3013) );
  AND2_X1 U21762 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18764), .ZN(
        P3_U3014) );
  AND2_X1 U21763 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18764), .ZN(
        P3_U3015) );
  AND2_X1 U21764 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18764), .ZN(
        P3_U3016) );
  AND2_X1 U21765 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18764), .ZN(
        P3_U3017) );
  AND2_X1 U21766 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18764), .ZN(
        P3_U3018) );
  AND2_X1 U21767 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18764), .ZN(
        P3_U3019) );
  AND2_X1 U21768 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18764), .ZN(
        P3_U3020) );
  INV_X1 U21769 ( .A(P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n21158) );
  NOR2_X1 U21770 ( .A1(n21158), .A2(n18767), .ZN(P3_U3021) );
  AND2_X1 U21771 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18764), .ZN(P3_U3022) );
  AND2_X1 U21772 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18764), .ZN(P3_U3023) );
  AND2_X1 U21773 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18764), .ZN(P3_U3024) );
  AND2_X1 U21774 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18764), .ZN(P3_U3025) );
  AND2_X1 U21775 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18764), .ZN(P3_U3026) );
  AND2_X1 U21776 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18764), .ZN(P3_U3027) );
  AND2_X1 U21777 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18764), .ZN(P3_U3028) );
  INV_X1 U21778 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18687) );
  AOI21_X1 U21779 ( .B1(HOLD), .B2(n18683), .A(n18687), .ZN(n18686) );
  AOI21_X1 U21780 ( .B1(n18693), .B2(P3_STATE_REG_1__SCAN_IN), .A(n18684), 
        .ZN(n18698) );
  AOI21_X1 U21781 ( .B1(NA), .B2(n18685), .A(n18699), .ZN(n18692) );
  OAI22_X1 U21782 ( .A1(n18754), .A2(n18686), .B1(n18698), .B2(n18692), .ZN(
        P3_U3029) );
  AOI21_X1 U21783 ( .B1(HOLD), .B2(n18688), .A(n18687), .ZN(n18690) );
  OAI21_X1 U21784 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n20740), .A(n18814), 
        .ZN(n18689) );
  OAI221_X1 U21785 ( .B1(n18690), .B2(P3_STATE_REG_1__SCAN_IN), .C1(n18690), 
        .C2(n18689), .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18691) );
  OAI211_X1 U21786 ( .C1(n18822), .C2(n18814), .A(n18811), .B(n18691), .ZN(
        P3_U3030) );
  INV_X1 U21787 ( .A(n18692), .ZN(n18697) );
  NAND2_X1 U21788 ( .A1(n18693), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18694) );
  OAI222_X1 U21789 ( .A1(n20740), .A2(n18699), .B1(P3_STATE_REG_1__SCAN_IN), 
        .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(n18694), .C2(NA), .ZN(n18695)
         );
  OAI211_X1 U21790 ( .C1(P3_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .B(n18695), .ZN(n18696) );
  OAI21_X1 U21791 ( .B1(n18698), .B2(n18697), .A(n18696), .ZN(P3_U3031) );
  INV_X1 U21792 ( .A(n18822), .ZN(n18821) );
  OAI222_X1 U21793 ( .A1(n18798), .A2(n18757), .B1(n18700), .B2(n18821), .C1(
        n18701), .C2(n18752), .ZN(P3_U3032) );
  OAI222_X1 U21794 ( .A1(n18752), .A2(n18703), .B1(n18702), .B2(n18754), .C1(
        n18701), .C2(n18757), .ZN(P3_U3033) );
  OAI222_X1 U21795 ( .A1(n18752), .A2(n18705), .B1(n18704), .B2(n18821), .C1(
        n18703), .C2(n18757), .ZN(P3_U3034) );
  INV_X1 U21796 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18707) );
  OAI222_X1 U21797 ( .A1(n18752), .A2(n18707), .B1(n18706), .B2(n18754), .C1(
        n18705), .C2(n18757), .ZN(P3_U3035) );
  OAI222_X1 U21798 ( .A1(n18752), .A2(n18709), .B1(n18708), .B2(n18821), .C1(
        n18707), .C2(n18757), .ZN(P3_U3036) );
  OAI222_X1 U21799 ( .A1(n18752), .A2(n18711), .B1(n18710), .B2(n18821), .C1(
        n18709), .C2(n18757), .ZN(P3_U3037) );
  OAI222_X1 U21800 ( .A1(n18752), .A2(n18713), .B1(n18712), .B2(n18754), .C1(
        n18711), .C2(n18757), .ZN(P3_U3038) );
  OAI222_X1 U21801 ( .A1(n18752), .A2(n21076), .B1(n18714), .B2(n18821), .C1(
        n18713), .C2(n18757), .ZN(P3_U3039) );
  OAI222_X1 U21802 ( .A1(n18752), .A2(n18716), .B1(n18715), .B2(n18821), .C1(
        n21076), .C2(n18757), .ZN(P3_U3040) );
  INV_X1 U21803 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18718) );
  OAI222_X1 U21804 ( .A1(n18752), .A2(n18718), .B1(n18717), .B2(n18821), .C1(
        n18716), .C2(n18757), .ZN(P3_U3041) );
  OAI222_X1 U21805 ( .A1(n18752), .A2(n18721), .B1(n18719), .B2(n18821), .C1(
        n18718), .C2(n18757), .ZN(P3_U3042) );
  OAI222_X1 U21806 ( .A1(n18721), .A2(n18757), .B1(n18720), .B2(n18821), .C1(
        n18722), .C2(n18752), .ZN(P3_U3043) );
  OAI222_X1 U21807 ( .A1(n18752), .A2(n18725), .B1(n18723), .B2(n18821), .C1(
        n18722), .C2(n18757), .ZN(P3_U3044) );
  OAI222_X1 U21808 ( .A1(n18725), .A2(n18757), .B1(n18724), .B2(n18821), .C1(
        n18726), .C2(n18752), .ZN(P3_U3045) );
  OAI222_X1 U21809 ( .A1(n18752), .A2(n18728), .B1(n18727), .B2(n18821), .C1(
        n18726), .C2(n18757), .ZN(P3_U3046) );
  OAI222_X1 U21810 ( .A1(n18752), .A2(n18731), .B1(n18729), .B2(n18821), .C1(
        n18728), .C2(n18757), .ZN(P3_U3047) );
  OAI222_X1 U21811 ( .A1(n18731), .A2(n18757), .B1(n18730), .B2(n18821), .C1(
        n21167), .C2(n18752), .ZN(P3_U3048) );
  INV_X1 U21812 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18733) );
  OAI222_X1 U21813 ( .A1(n21167), .A2(n18757), .B1(n18732), .B2(n18821), .C1(
        n18733), .C2(n18752), .ZN(P3_U3049) );
  OAI222_X1 U21814 ( .A1(n18752), .A2(n18736), .B1(n18734), .B2(n18821), .C1(
        n18733), .C2(n18757), .ZN(P3_U3050) );
  OAI222_X1 U21815 ( .A1(n18736), .A2(n18757), .B1(n18735), .B2(n18821), .C1(
        n18737), .C2(n18752), .ZN(P3_U3051) );
  OAI222_X1 U21816 ( .A1(n18752), .A2(n18739), .B1(n18738), .B2(n18821), .C1(
        n18737), .C2(n18757), .ZN(P3_U3052) );
  OAI222_X1 U21817 ( .A1(n18752), .A2(n21127), .B1(n18740), .B2(n18821), .C1(
        n18739), .C2(n18757), .ZN(P3_U3053) );
  OAI222_X1 U21818 ( .A1(n18752), .A2(n18743), .B1(n18741), .B2(n18754), .C1(
        n21127), .C2(n18757), .ZN(P3_U3054) );
  OAI222_X1 U21819 ( .A1(n18743), .A2(n18757), .B1(n18742), .B2(n18754), .C1(
        n18744), .C2(n18752), .ZN(P3_U3055) );
  INV_X1 U21820 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18746) );
  OAI222_X1 U21821 ( .A1(n18752), .A2(n18746), .B1(n18745), .B2(n18754), .C1(
        n18744), .C2(n18757), .ZN(P3_U3056) );
  OAI222_X1 U21822 ( .A1(n18752), .A2(n21068), .B1(n18747), .B2(n18754), .C1(
        n18746), .C2(n18757), .ZN(P3_U3057) );
  OAI222_X1 U21823 ( .A1(n18752), .A2(n18749), .B1(n18748), .B2(n18754), .C1(
        n21068), .C2(n18757), .ZN(P3_U3058) );
  OAI222_X1 U21824 ( .A1(n18749), .A2(n18757), .B1(n21151), .B2(n18754), .C1(
        n18750), .C2(n18752), .ZN(P3_U3059) );
  INV_X1 U21825 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18756) );
  OAI222_X1 U21826 ( .A1(n18752), .A2(n18756), .B1(n18751), .B2(n18754), .C1(
        n18750), .C2(n18757), .ZN(P3_U3060) );
  OAI222_X1 U21827 ( .A1(n18757), .A2(n18756), .B1(n18755), .B2(n18754), .C1(
        n18753), .C2(n18752), .ZN(P3_U3061) );
  INV_X1 U21828 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n21110) );
  AOI22_X1 U21829 ( .A1(n18754), .A2(n18758), .B1(n21110), .B2(n18822), .ZN(
        P3_U3274) );
  OAI22_X1 U21830 ( .A1(n18822), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18821), .ZN(n18759) );
  INV_X1 U21831 ( .A(n18759), .ZN(P3_U3275) );
  OAI22_X1 U21832 ( .A1(n18822), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18821), .ZN(n18760) );
  INV_X1 U21833 ( .A(n18760), .ZN(P3_U3276) );
  OAI22_X1 U21834 ( .A1(n18822), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18821), .ZN(n18761) );
  INV_X1 U21835 ( .A(n18761), .ZN(P3_U3277) );
  INV_X1 U21836 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18763) );
  INV_X1 U21837 ( .A(n18765), .ZN(n18762) );
  AOI21_X1 U21838 ( .B1(n18764), .B2(n18763), .A(n18762), .ZN(P3_U3280) );
  OAI21_X1 U21839 ( .B1(n18767), .B2(n18766), .A(n18765), .ZN(P3_U3281) );
  AOI21_X1 U21840 ( .B1(n18769), .B2(P3_STATE2_REG_3__SCAN_IN), .A(n18768), 
        .ZN(n18770) );
  INV_X1 U21841 ( .A(n18770), .ZN(P3_U3282) );
  NOR2_X1 U21842 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18771), .ZN(
        n18773) );
  AOI22_X1 U21843 ( .A1(n18793), .A2(n18773), .B1(n18791), .B2(n18772), .ZN(
        n18777) );
  AOI21_X1 U21844 ( .B1(n18793), .B2(n18774), .A(n18797), .ZN(n18776) );
  OAI22_X1 U21845 ( .A1(n18797), .A2(n18777), .B1(n18776), .B2(n18775), .ZN(
        P3_U3285) );
  OAI22_X1 U21846 ( .A1(n18778), .A2(n10446), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18787) );
  INV_X1 U21847 ( .A(n18787), .ZN(n18784) );
  NOR2_X1 U21848 ( .A1(n18779), .A2(n21150), .ZN(n18786) );
  OAI22_X1 U21849 ( .A1(n18782), .A2(n18824), .B1(n18781), .B2(n18780), .ZN(
        n18783) );
  AOI21_X1 U21850 ( .B1(n18784), .B2(n18786), .A(n18783), .ZN(n18785) );
  INV_X1 U21851 ( .A(n18797), .ZN(n18794) );
  AOI22_X1 U21852 ( .A1(n18797), .A2(n10497), .B1(n18785), .B2(n18794), .ZN(
        P3_U3288) );
  AOI222_X1 U21853 ( .A1(n18789), .A2(n18793), .B1(n18791), .B2(n18788), .C1(
        n18787), .C2(n18786), .ZN(n18790) );
  AOI22_X1 U21854 ( .A1(n18797), .A2(n10495), .B1(n18790), .B2(n18794), .ZN(
        P3_U3289) );
  AOI222_X1 U21855 ( .A1(n21150), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18793), 
        .B2(n18792), .C1(n18796), .C2(n18791), .ZN(n18795) );
  AOI22_X1 U21856 ( .A1(n18797), .A2(n18796), .B1(n18795), .B2(n18794), .ZN(
        P3_U3290) );
  AOI21_X1 U21857 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18799) );
  AOI22_X1 U21858 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18799), .B2(n18798), .ZN(n18802) );
  INV_X1 U21859 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18801) );
  AOI22_X1 U21860 ( .A1(n18804), .A2(n18802), .B1(n18801), .B2(n18800), .ZN(
        P3_U3292) );
  INV_X1 U21861 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21020) );
  OAI21_X1 U21862 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18804), .ZN(n18803) );
  OAI21_X1 U21863 ( .B1(n18804), .B2(n21020), .A(n18803), .ZN(P3_U3293) );
  INV_X1 U21864 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18805) );
  AOI22_X1 U21865 ( .A1(n18821), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18805), 
        .B2(n18822), .ZN(P3_U3294) );
  MUX2_X1 U21866 ( .A(P3_MORE_REG_SCAN_IN), .B(n18807), .S(n18806), .Z(
        P3_U3295) );
  OAI21_X1 U21867 ( .B1(n18809), .B2(n18808), .A(n18826), .ZN(n18810) );
  AOI21_X1 U21868 ( .B1(n17412), .B2(n18814), .A(n18810), .ZN(n18820) );
  AOI21_X1 U21869 ( .B1(n18813), .B2(n18812), .A(n18811), .ZN(n18815) );
  OAI211_X1 U21870 ( .C1(n18825), .C2(n18815), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18814), .ZN(n18817) );
  AOI21_X1 U21871 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18817), .A(n18816), 
        .ZN(n18819) );
  NAND2_X1 U21872 ( .A1(n18820), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18818) );
  OAI21_X1 U21873 ( .B1(n18820), .B2(n18819), .A(n18818), .ZN(P3_U3296) );
  OAI22_X1 U21874 ( .A1(n18822), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18821), .ZN(n18823) );
  INV_X1 U21875 ( .A(n18823), .ZN(P3_U3297) );
  OAI21_X1 U21876 ( .B1(n18824), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n18826), 
        .ZN(n18829) );
  OAI22_X1 U21877 ( .A1(n18829), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18826), 
        .B2(n18825), .ZN(n18827) );
  INV_X1 U21878 ( .A(n18827), .ZN(P3_U3298) );
  OAI21_X1 U21879 ( .B1(n18829), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18828), 
        .ZN(n18830) );
  INV_X1 U21880 ( .A(n18830), .ZN(P3_U3299) );
  INV_X1 U21881 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19769) );
  INV_X1 U21882 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19786) );
  NAND2_X1 U21883 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19786), .ZN(n19776) );
  INV_X1 U21884 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19779) );
  NAND2_X1 U21885 ( .A1(n19769), .A2(n19779), .ZN(n19773) );
  OAI21_X1 U21886 ( .B1(n19769), .B2(n19776), .A(n19773), .ZN(n19845) );
  AOI21_X1 U21887 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19845), .ZN(n18831) );
  INV_X1 U21888 ( .A(n18831), .ZN(P2_U2815) );
  INV_X1 U21889 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18833) );
  OAI22_X1 U21890 ( .A1(n19895), .A2(n18833), .B1(n19904), .B2(n18832), .ZN(
        P2_U2816) );
  OR2_X1 U21891 ( .A1(n19779), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n19913) );
  INV_X1 U21892 ( .A(n19913), .ZN(n19912) );
  AOI22_X1 U21893 ( .A1(n19912), .A2(n18833), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n19913), .ZN(n18834) );
  OAI21_X1 U21894 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n19773), .A(n18834), 
        .ZN(P2_U2817) );
  OAI21_X1 U21895 ( .B1(n19778), .B2(BS16), .A(n19845), .ZN(n19843) );
  OAI21_X1 U21896 ( .B1(n19845), .B2(n19902), .A(n19843), .ZN(P2_U2818) );
  NOR4_X1 U21897 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n18844) );
  NOR4_X1 U21898 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n18843) );
  NOR4_X1 U21899 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18835) );
  INV_X1 U21900 ( .A(P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20950) );
  INV_X1 U21901 ( .A(P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20971) );
  NAND3_X1 U21902 ( .A1(n18835), .A2(n20950), .A3(n20971), .ZN(n18841) );
  NOR4_X1 U21903 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18839) );
  NOR4_X1 U21904 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(P2_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n18838) );
  NOR4_X1 U21905 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18837) );
  NOR4_X1 U21906 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18836) );
  NAND4_X1 U21907 ( .A1(n18839), .A2(n18838), .A3(n18837), .A4(n18836), .ZN(
        n18840) );
  AOI211_X1 U21908 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n18841), .B(n18840), .ZN(n18842) );
  NAND3_X1 U21909 ( .A1(n18844), .A2(n18843), .A3(n18842), .ZN(n18852) );
  NOR2_X1 U21910 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18852), .ZN(n18847) );
  INV_X1 U21911 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19068) );
  INV_X1 U21912 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18845) );
  AOI22_X1 U21913 ( .A1(n18847), .A2(n19068), .B1(n18852), .B2(n18845), .ZN(
        P2_U2820) );
  OR3_X1 U21914 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18851) );
  INV_X1 U21915 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18846) );
  AOI22_X1 U21916 ( .A1(n18847), .A2(n18851), .B1(n18852), .B2(n18846), .ZN(
        P2_U2821) );
  INV_X1 U21917 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19844) );
  NAND2_X1 U21918 ( .A1(n18847), .A2(n19844), .ZN(n18850) );
  INV_X1 U21919 ( .A(n18852), .ZN(n18854) );
  OAI21_X1 U21920 ( .B1(n10793), .B2(n19068), .A(n18854), .ZN(n18848) );
  OAI21_X1 U21921 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18854), .A(n18848), 
        .ZN(n18849) );
  OAI221_X1 U21922 ( .B1(n18850), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18850), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18849), .ZN(P2_U2822) );
  INV_X1 U21923 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18853) );
  OAI221_X1 U21924 ( .B1(n18854), .B2(n18853), .C1(n18852), .C2(n18851), .A(
        n18850), .ZN(P2_U2823) );
  AOI22_X1 U21925 ( .A1(n18856), .A2(n19062), .B1(n18855), .B2(n19064), .ZN(
        n18866) );
  AOI211_X1 U21926 ( .C1(n18859), .C2(n18857), .A(n18858), .B(n19061), .ZN(
        n18864) );
  INV_X1 U21927 ( .A(n18860), .ZN(n18862) );
  AOI22_X1 U21928 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19080), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19049), .ZN(n18861) );
  OAI21_X1 U21929 ( .B1(n18862), .B2(n19070), .A(n18861), .ZN(n18863) );
  AOI211_X1 U21930 ( .C1(P2_EBX_REG_20__SCAN_IN), .C2(n19063), .A(n18864), .B(
        n18863), .ZN(n18865) );
  NAND2_X1 U21931 ( .A1(n18866), .A2(n18865), .ZN(P2_U2835) );
  AOI211_X1 U21932 ( .C1(n18869), .C2(n18868), .A(n18867), .B(n19061), .ZN(
        n18875) );
  INV_X1 U21933 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19811) );
  AOI22_X1 U21934 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n19063), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19080), .ZN(n18870) );
  OAI211_X1 U21935 ( .C1(n19069), .C2(n19811), .A(n18870), .B(n19034), .ZN(
        n18871) );
  AOI21_X1 U21936 ( .B1(n18872), .B2(n18999), .A(n18871), .ZN(n18873) );
  INV_X1 U21937 ( .A(n18873), .ZN(n18874) );
  AOI211_X1 U21938 ( .C1(n19062), .C2(n18876), .A(n18875), .B(n18874), .ZN(
        n18877) );
  OAI21_X1 U21939 ( .B1(n18878), .B2(n19053), .A(n18877), .ZN(P2_U2836) );
  AOI211_X1 U21940 ( .C1(n18880), .C2(n18879), .A(n9928), .B(n19061), .ZN(
        n18886) );
  NAND2_X1 U21941 ( .A1(n18881), .A2(n18999), .ZN(n18884) );
  AOI22_X1 U21942 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n19063), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19080), .ZN(n18883) );
  NAND2_X1 U21943 ( .A1(n19049), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n18882) );
  NAND4_X1 U21944 ( .A1(n18884), .A2(n18883), .A3(n19034), .A4(n18882), .ZN(
        n18885) );
  AOI211_X1 U21945 ( .C1(n19064), .C2(n18887), .A(n18886), .B(n18885), .ZN(
        n18888) );
  OAI21_X1 U21946 ( .B1(n18889), .B2(n19047), .A(n18888), .ZN(P2_U2837) );
  AOI211_X1 U21947 ( .C1(n18892), .C2(n18891), .A(n18890), .B(n19061), .ZN(
        n18898) );
  AOI22_X1 U21948 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n19063), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19080), .ZN(n18893) );
  OAI211_X1 U21949 ( .C1(n19069), .C2(n19808), .A(n18893), .B(n19034), .ZN(
        n18894) );
  INV_X1 U21950 ( .A(n18894), .ZN(n18895) );
  OAI21_X1 U21951 ( .B1(n18896), .B2(n19070), .A(n18895), .ZN(n18897) );
  AOI211_X1 U21952 ( .C1(n19062), .C2(n18899), .A(n18898), .B(n18897), .ZN(
        n18900) );
  OAI21_X1 U21953 ( .B1(n18901), .B2(n19053), .A(n18900), .ZN(P2_U2838) );
  AOI211_X1 U21954 ( .C1(n18904), .C2(n18903), .A(n18902), .B(n19061), .ZN(
        n18908) );
  AOI22_X1 U21955 ( .A1(n18905), .A2(n18999), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19080), .ZN(n18906) );
  OAI211_X1 U21956 ( .C1(n15451), .C2(n19069), .A(n18906), .B(n19034), .ZN(
        n18907) );
  AOI211_X1 U21957 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19063), .A(n18908), .B(
        n18907), .ZN(n18912) );
  INV_X1 U21958 ( .A(n19091), .ZN(n18910) );
  AOI22_X1 U21959 ( .A1(n18910), .A2(n19064), .B1(n18909), .B2(n19062), .ZN(
        n18911) );
  NAND2_X1 U21960 ( .A1(n18912), .A2(n18911), .ZN(P2_U2839) );
  NOR2_X1 U21961 ( .A1(n19061), .A2(n9925), .ZN(n19079) );
  INV_X1 U21962 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19805) );
  OAI22_X1 U21963 ( .A1(n21083), .A2(n19035), .B1(n19805), .B2(n19069), .ZN(
        n18913) );
  AOI211_X1 U21964 ( .C1(n18920), .C2(n19079), .A(n19236), .B(n18913), .ZN(
        n18916) );
  AOI22_X1 U21965 ( .A1(n18914), .A2(n18999), .B1(P2_EBX_REG_15__SCAN_IN), 
        .B2(n19063), .ZN(n18915) );
  OAI211_X1 U21966 ( .C1(n18917), .C2(n19047), .A(n18916), .B(n18915), .ZN(
        n18922) );
  NAND2_X1 U21967 ( .A1(n19764), .A2(n9925), .ZN(n19083) );
  AOI211_X1 U21968 ( .C1(n18920), .C2(n18919), .A(n18918), .B(n19083), .ZN(
        n18921) );
  NOR2_X1 U21969 ( .A1(n18922), .A2(n18921), .ZN(n18923) );
  OAI21_X1 U21970 ( .B1(n19102), .B2(n19053), .A(n18923), .ZN(P2_U2840) );
  AOI22_X1 U21971 ( .A1(n18924), .A2(n18999), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19063), .ZN(n18925) );
  OAI211_X1 U21972 ( .C1(n11341), .C2(n19069), .A(n18925), .B(n19034), .ZN(
        n18926) );
  AOI21_X1 U21973 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19080), .A(
        n18926), .ZN(n18931) );
  NOR2_X1 U21974 ( .A1(n19041), .A2(n18933), .ZN(n18928) );
  XNOR2_X1 U21975 ( .A(n18928), .B(n18927), .ZN(n18929) );
  AOI22_X1 U21976 ( .A1(n19764), .A2(n18929), .B1(n19064), .B2(n19103), .ZN(
        n18930) );
  OAI211_X1 U21977 ( .C1(n19047), .C2(n18932), .A(n18931), .B(n18930), .ZN(
        P2_U2841) );
  AOI211_X1 U21978 ( .C1(n18941), .C2(n18934), .A(n18933), .B(n19083), .ZN(
        n18939) );
  INV_X1 U21979 ( .A(n18935), .ZN(n18937) );
  AOI22_X1 U21980 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19080), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19049), .ZN(n18936) );
  OAI211_X1 U21981 ( .C1(n18937), .C2(n19070), .A(n18936), .B(n19034), .ZN(
        n18938) );
  AOI211_X1 U21982 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n19063), .A(n18939), .B(
        n18938), .ZN(n18943) );
  AOI22_X1 U21983 ( .A1(n18941), .A2(n19079), .B1(n19062), .B2(n18940), .ZN(
        n18942) );
  OAI211_X1 U21984 ( .C1(n19053), .C2(n19107), .A(n18943), .B(n18942), .ZN(
        P2_U2842) );
  NOR2_X1 U21985 ( .A1(n19041), .A2(n18944), .ZN(n18946) );
  XOR2_X1 U21986 ( .A(n18946), .B(n18945), .Z(n18953) );
  OAI21_X1 U21987 ( .B1(n11333), .B2(n19069), .A(n19034), .ZN(n18949) );
  OAI22_X1 U21988 ( .A1(n18947), .A2(n19070), .B1(n19035), .B2(n11419), .ZN(
        n18948) );
  AOI211_X1 U21989 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n19063), .A(n18949), .B(
        n18948), .ZN(n18952) );
  AOI22_X1 U21990 ( .A1(n19064), .A2(n19108), .B1(n19062), .B2(n18950), .ZN(
        n18951) );
  OAI211_X1 U21991 ( .C1(n19061), .C2(n18953), .A(n18952), .B(n18951), .ZN(
        P2_U2843) );
  OAI21_X1 U21992 ( .B1(n19800), .B2(n19069), .A(n19034), .ZN(n18957) );
  OAI22_X1 U21993 ( .A1(n18955), .A2(n19070), .B1(n18954), .B2(n19008), .ZN(
        n18956) );
  AOI211_X1 U21994 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n19080), .A(
        n18957), .B(n18956), .ZN(n18964) );
  NAND2_X1 U21995 ( .A1(n9925), .A2(n18958), .ZN(n18959) );
  XNOR2_X1 U21996 ( .A(n18960), .B(n18959), .ZN(n18962) );
  AOI22_X1 U21997 ( .A1(n19764), .A2(n18962), .B1(n19062), .B2(n18961), .ZN(
        n18963) );
  OAI211_X1 U21998 ( .C1(n19053), .C2(n19110), .A(n18964), .B(n18963), .ZN(
        P2_U2844) );
  NOR2_X1 U21999 ( .A1(n19041), .A2(n18965), .ZN(n18966) );
  XOR2_X1 U22000 ( .A(n18967), .B(n18966), .Z(n18974) );
  AOI22_X1 U22001 ( .A1(n18968), .A2(n18999), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19080), .ZN(n18969) );
  OAI211_X1 U22002 ( .C1(n19798), .C2(n19069), .A(n18969), .B(n19034), .ZN(
        n18972) );
  OAI22_X1 U22003 ( .A1(n19053), .A2(n19113), .B1(n19047), .B2(n18970), .ZN(
        n18971) );
  AOI211_X1 U22004 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n19063), .A(n18972), .B(
        n18971), .ZN(n18973) );
  OAI21_X1 U22005 ( .B1(n19061), .B2(n18974), .A(n18973), .ZN(P2_U2845) );
  OAI21_X1 U22006 ( .B1(n11324), .B2(n19069), .A(n19034), .ZN(n18978) );
  INV_X1 U22007 ( .A(n18975), .ZN(n18976) );
  OAI22_X1 U22008 ( .A1(n18976), .A2(n19070), .B1(n20978), .B2(n19008), .ZN(
        n18977) );
  AOI211_X1 U22009 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19080), .A(
        n18978), .B(n18977), .ZN(n18985) );
  NAND2_X1 U22010 ( .A1(n9925), .A2(n18979), .ZN(n18980) );
  XNOR2_X1 U22011 ( .A(n18981), .B(n18980), .ZN(n18983) );
  AOI22_X1 U22012 ( .A1(n19764), .A2(n18983), .B1(n19062), .B2(n18982), .ZN(
        n18984) );
  OAI211_X1 U22013 ( .C1(n19053), .C2(n19114), .A(n18985), .B(n18984), .ZN(
        P2_U2846) );
  AOI22_X1 U22014 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n19063), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19080), .ZN(n18986) );
  OAI21_X1 U22015 ( .B1(n18987), .B2(n19070), .A(n18986), .ZN(n18988) );
  AOI211_X1 U22016 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19049), .A(n19236), .B(
        n18988), .ZN(n18994) );
  NOR2_X1 U22017 ( .A1(n19041), .A2(n18989), .ZN(n18991) );
  XNOR2_X1 U22018 ( .A(n18991), .B(n18990), .ZN(n18992) );
  AOI22_X1 U22019 ( .A1(n19764), .A2(n18992), .B1(n19064), .B2(n19115), .ZN(
        n18993) );
  OAI211_X1 U22020 ( .C1(n19047), .C2(n18995), .A(n18994), .B(n18993), .ZN(
        P2_U2847) );
  NAND2_X1 U22021 ( .A1(n9925), .A2(n18996), .ZN(n18998) );
  XOR2_X1 U22022 ( .A(n18998), .B(n18997), .Z(n19006) );
  AOI22_X1 U22023 ( .A1(n19000), .A2(n18999), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19080), .ZN(n19001) );
  OAI211_X1 U22024 ( .C1(n19794), .C2(n19069), .A(n19001), .B(n19034), .ZN(
        n19004) );
  OAI22_X1 U22025 ( .A1(n19053), .A2(n19119), .B1(n19047), .B2(n19002), .ZN(
        n19003) );
  AOI211_X1 U22026 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n19063), .A(n19004), .B(
        n19003), .ZN(n19005) );
  OAI21_X1 U22027 ( .B1(n19006), .B2(n19061), .A(n19005), .ZN(P2_U2848) );
  OAI21_X1 U22028 ( .B1(n11312), .B2(n19069), .A(n19034), .ZN(n19011) );
  OAI22_X1 U22029 ( .A1(n19009), .A2(n19070), .B1(n19008), .B2(n19007), .ZN(
        n19010) );
  AOI211_X1 U22030 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19080), .A(
        n19011), .B(n19010), .ZN(n19018) );
  NOR2_X1 U22031 ( .A1(n19041), .A2(n19012), .ZN(n19014) );
  XNOR2_X1 U22032 ( .A(n19014), .B(n19013), .ZN(n19016) );
  AOI22_X1 U22033 ( .A1(n19764), .A2(n19016), .B1(n19062), .B2(n19015), .ZN(
        n19017) );
  OAI211_X1 U22034 ( .C1(n19053), .C2(n19122), .A(n19018), .B(n19017), .ZN(
        P2_U2849) );
  OAI21_X1 U22035 ( .B1(n11308), .B2(n19069), .A(n19034), .ZN(n19022) );
  OAI22_X1 U22036 ( .A1(n19020), .A2(n19070), .B1(n19035), .B2(n19019), .ZN(
        n19021) );
  AOI211_X1 U22037 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n19063), .A(n19022), .B(
        n19021), .ZN(n19030) );
  NAND2_X1 U22038 ( .A1(n9925), .A2(n19023), .ZN(n19025) );
  XNOR2_X1 U22039 ( .A(n19026), .B(n19025), .ZN(n19028) );
  AOI22_X1 U22040 ( .A1(n19764), .A2(n19028), .B1(n19062), .B2(n19027), .ZN(
        n19029) );
  OAI211_X1 U22041 ( .C1(n19053), .C2(n19132), .A(n19030), .B(n19029), .ZN(
        P2_U2850) );
  INV_X1 U22042 ( .A(n19031), .ZN(n19038) );
  INV_X1 U22043 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n21097) );
  AOI22_X1 U22044 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19063), .B1(n19064), .B2(
        n19032), .ZN(n19033) );
  OAI211_X1 U22045 ( .C1(n19035), .C2(n21097), .A(n19034), .B(n19033), .ZN(
        n19036) );
  AOI21_X1 U22046 ( .B1(n19049), .B2(P2_REIP_REG_4__SCAN_IN), .A(n19036), .ZN(
        n19037) );
  OAI21_X1 U22047 ( .B1(n19038), .B2(n19070), .A(n19037), .ZN(n19039) );
  AOI21_X1 U22048 ( .B1(n19128), .B2(n19077), .A(n19039), .ZN(n19046) );
  INV_X1 U22049 ( .A(n19246), .ZN(n19044) );
  NOR2_X1 U22050 ( .A1(n19041), .A2(n19040), .ZN(n19043) );
  AOI21_X1 U22051 ( .B1(n19044), .B2(n19043), .A(n19061), .ZN(n19042) );
  OAI21_X1 U22052 ( .B1(n19044), .B2(n19043), .A(n19042), .ZN(n19045) );
  OAI211_X1 U22053 ( .C1(n19048), .C2(n19047), .A(n19046), .B(n19045), .ZN(
        P2_U2851) );
  NAND2_X1 U22054 ( .A1(n19063), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n19051) );
  AOI22_X1 U22055 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19080), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19049), .ZN(n19050) );
  OAI211_X1 U22056 ( .C1(n19070), .C2(n19052), .A(n19051), .B(n19050), .ZN(
        n19056) );
  NOR2_X1 U22057 ( .A1(n19054), .A2(n19053), .ZN(n19055) );
  AOI211_X1 U22058 ( .C1(n12489), .C2(n19062), .A(n19056), .B(n19055), .ZN(
        n19059) );
  AOI22_X1 U22059 ( .A1(n19079), .A2(n19057), .B1(n19342), .B2(n19077), .ZN(
        n19058) );
  OAI211_X1 U22060 ( .C1(n19061), .C2(n19060), .A(n19059), .B(n19058), .ZN(
        P2_U2854) );
  NAND2_X1 U22061 ( .A1(n12485), .A2(n19062), .ZN(n19075) );
  NAND2_X1 U22062 ( .A1(n19063), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n19067) );
  NAND2_X1 U22063 ( .A1(n19065), .A2(n19064), .ZN(n19066) );
  OAI211_X1 U22064 ( .C1(n19069), .C2(n19068), .A(n19067), .B(n19066), .ZN(
        n19073) );
  NOR2_X1 U22065 ( .A1(n19071), .A2(n19070), .ZN(n19072) );
  NOR2_X1 U22066 ( .A1(n19073), .A2(n19072), .ZN(n19074) );
  NAND2_X1 U22067 ( .A1(n19075), .A2(n19074), .ZN(n19076) );
  AOI21_X1 U22068 ( .B1(n19078), .B2(n19077), .A(n19076), .ZN(n19082) );
  OAI21_X1 U22069 ( .B1(n19080), .B2(n19079), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19081) );
  OAI211_X1 U22070 ( .C1(n19084), .C2(n19083), .A(n19082), .B(n19081), .ZN(
        P2_U2855) );
  AOI22_X1 U22071 ( .A1(n19085), .A2(n19099), .B1(n19090), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19087) );
  AOI22_X1 U22072 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19125), .B1(n19089), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19086) );
  NAND2_X1 U22073 ( .A1(n19087), .A2(n19086), .ZN(P2_U2888) );
  AOI22_X1 U22074 ( .A1(n19088), .A2(n19204), .B1(n19125), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19098) );
  AOI22_X1 U22075 ( .A1(n19090), .A2(BUF2_REG_16__SCAN_IN), .B1(n19089), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19097) );
  OAI22_X1 U22076 ( .A1(n19094), .A2(n19093), .B1(n19092), .B2(n19091), .ZN(
        n19095) );
  INV_X1 U22077 ( .A(n19095), .ZN(n19096) );
  NAND3_X1 U22078 ( .A1(n19098), .A2(n19097), .A3(n19096), .ZN(P2_U2903) );
  INV_X1 U22079 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19174) );
  AOI22_X1 U22080 ( .A1(n19101), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19100), .ZN(n19235) );
  OAI222_X1 U22081 ( .A1(n19102), .A2(n19133), .B1(n19174), .B2(n19121), .C1(
        n19235), .C2(n19120), .ZN(P2_U2904) );
  INV_X1 U22082 ( .A(n19103), .ZN(n19106) );
  AOI22_X1 U22083 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19125), .B1(n19104), 
        .B2(n19123), .ZN(n19105) );
  OAI21_X1 U22084 ( .B1(n19133), .B2(n19106), .A(n19105), .ZN(P2_U2905) );
  INV_X1 U22085 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19178) );
  OAI222_X1 U22086 ( .A1(n19107), .A2(n19133), .B1(n19178), .B2(n19121), .C1(
        n19120), .C2(n19230), .ZN(P2_U2906) );
  INV_X1 U22087 ( .A(n19108), .ZN(n19109) );
  INV_X1 U22088 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19180) );
  OAI222_X1 U22089 ( .A1(n19109), .A2(n19133), .B1(n19180), .B2(n19121), .C1(
        n19120), .C2(n19228), .ZN(P2_U2907) );
  INV_X1 U22090 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19182) );
  OAI222_X1 U22091 ( .A1(n19110), .A2(n19133), .B1(n19182), .B2(n19121), .C1(
        n19120), .C2(n19226), .ZN(P2_U2908) );
  AOI22_X1 U22092 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19125), .B1(n19111), 
        .B2(n19123), .ZN(n19112) );
  OAI21_X1 U22093 ( .B1(n19133), .B2(n19113), .A(n19112), .ZN(P2_U2909) );
  INV_X1 U22094 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19185) );
  OAI222_X1 U22095 ( .A1(n19114), .A2(n19133), .B1(n19185), .B2(n19121), .C1(
        n19120), .C2(n19224), .ZN(P2_U2910) );
  INV_X1 U22096 ( .A(n19115), .ZN(n19118) );
  AOI22_X1 U22097 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19125), .B1(n19116), .B2(
        n19123), .ZN(n19117) );
  OAI21_X1 U22098 ( .B1(n19133), .B2(n19118), .A(n19117), .ZN(P2_U2911) );
  OAI222_X1 U22099 ( .A1(n19119), .A2(n19133), .B1(n19188), .B2(n19121), .C1(
        n19120), .C2(n19222), .ZN(P2_U2912) );
  INV_X1 U22100 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19190) );
  OAI222_X1 U22101 ( .A1(n19122), .A2(n19133), .B1(n19190), .B2(n19121), .C1(
        n19120), .C2(n19220), .ZN(P2_U2913) );
  AOI22_X1 U22102 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19125), .B1(n19124), .B2(
        n19123), .ZN(n19131) );
  INV_X1 U22103 ( .A(n19126), .ZN(n19129) );
  NAND3_X1 U22104 ( .A1(n19129), .A2(n19128), .A3(n19127), .ZN(n19130) );
  OAI211_X1 U22105 ( .C1(n19133), .C2(n19132), .A(n19131), .B(n19130), .ZN(
        P2_U2914) );
  OR2_X1 U22106 ( .A1(n19135), .A2(n19134), .ZN(n19137) );
  OAI21_X1 U22107 ( .B1(n19138), .B2(n19137), .A(n19136), .ZN(n19139) );
  OR2_X1 U22108 ( .A1(n19140), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19898) );
  NAND2_X1 U22109 ( .A1(n19203), .A2(n19898), .ZN(n19172) );
  NOR2_X1 U22110 ( .A1(n19172), .A2(n19141), .ZN(P2_U2920) );
  INV_X1 U22111 ( .A(n19168), .ZN(n19170) );
  AOI22_X1 U22112 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n19170), .B1(n9798), .B2(
        P2_UWORD_REG_14__SCAN_IN), .ZN(n19143) );
  OAI21_X1 U22113 ( .B1(n21031), .B2(n19172), .A(n19143), .ZN(P2_U2921) );
  AOI22_X1 U22114 ( .A1(n9798), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19144) );
  OAI21_X1 U22115 ( .B1(n19145), .B2(n19168), .A(n19144), .ZN(P2_U2922) );
  INV_X1 U22116 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19147) );
  AOI22_X1 U22117 ( .A1(n9798), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19146) );
  OAI21_X1 U22118 ( .B1(n19147), .B2(n19168), .A(n19146), .ZN(P2_U2923) );
  INV_X1 U22119 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19149) );
  AOI22_X1 U22120 ( .A1(n9798), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19148) );
  OAI21_X1 U22121 ( .B1(n19149), .B2(n19168), .A(n19148), .ZN(P2_U2924) );
  AOI22_X1 U22122 ( .A1(n9798), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19150) );
  OAI21_X1 U22123 ( .B1(n19151), .B2(n19168), .A(n19150), .ZN(P2_U2925) );
  INV_X1 U22124 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n21095) );
  INV_X1 U22125 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19153) );
  OAI222_X1 U22126 ( .A1(n19898), .A2(n21095), .B1(n19168), .B2(n19153), .C1(
        n19172), .C2(n19152), .ZN(P2_U2926) );
  AOI22_X1 U22127 ( .A1(n9798), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19154) );
  OAI21_X1 U22128 ( .B1(n19155), .B2(n19168), .A(n19154), .ZN(P2_U2927) );
  AOI22_X1 U22129 ( .A1(n9798), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19156) );
  OAI21_X1 U22130 ( .B1(n19157), .B2(n19168), .A(n19156), .ZN(P2_U2928) );
  AOI22_X1 U22131 ( .A1(n9798), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19158) );
  OAI21_X1 U22132 ( .B1(n21118), .B2(n19168), .A(n19158), .ZN(P2_U2929) );
  INV_X1 U22133 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19160) );
  AOI22_X1 U22134 ( .A1(n9798), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19159) );
  OAI21_X1 U22135 ( .B1(n19160), .B2(n19168), .A(n19159), .ZN(P2_U2930) );
  AOI22_X1 U22136 ( .A1(n9798), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19161) );
  OAI21_X1 U22137 ( .B1(n19162), .B2(n19168), .A(n19161), .ZN(P2_U2931) );
  INV_X1 U22138 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19164) );
  AOI22_X1 U22139 ( .A1(n9798), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19163) );
  OAI21_X1 U22140 ( .B1(n19164), .B2(n19168), .A(n19163), .ZN(P2_U2932) );
  AOI22_X1 U22141 ( .A1(n9798), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19165) );
  OAI21_X1 U22142 ( .B1(n19166), .B2(n19168), .A(n19165), .ZN(P2_U2933) );
  AOI22_X1 U22143 ( .A1(n9798), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19167) );
  OAI21_X1 U22144 ( .B1(n19169), .B2(n19168), .A(n19167), .ZN(P2_U2934) );
  AOI22_X1 U22145 ( .A1(P2_EAX_REG_16__SCAN_IN), .A2(n19170), .B1(n9798), .B2(
        P2_UWORD_REG_0__SCAN_IN), .ZN(n19171) );
  OAI21_X1 U22146 ( .B1(n21146), .B2(n19172), .A(n19171), .ZN(P2_U2935) );
  AOI22_X1 U22147 ( .A1(n9798), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19173) );
  OAI21_X1 U22148 ( .B1(n19174), .B2(n19203), .A(n19173), .ZN(P2_U2936) );
  AOI22_X1 U22149 ( .A1(n9798), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19175) );
  OAI21_X1 U22150 ( .B1(n19176), .B2(n19203), .A(n19175), .ZN(P2_U2937) );
  AOI22_X1 U22151 ( .A1(n9798), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19177) );
  OAI21_X1 U22152 ( .B1(n19178), .B2(n19203), .A(n19177), .ZN(P2_U2938) );
  AOI22_X1 U22153 ( .A1(n9798), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19179) );
  OAI21_X1 U22154 ( .B1(n19180), .B2(n19203), .A(n19179), .ZN(P2_U2939) );
  AOI22_X1 U22155 ( .A1(n9798), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19181) );
  OAI21_X1 U22156 ( .B1(n19182), .B2(n19203), .A(n19181), .ZN(P2_U2940) );
  AOI22_X1 U22157 ( .A1(n9798), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19183) );
  OAI21_X1 U22158 ( .B1(n11579), .B2(n19203), .A(n19183), .ZN(P2_U2941) );
  AOI22_X1 U22159 ( .A1(n9798), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19184) );
  OAI21_X1 U22160 ( .B1(n19185), .B2(n19203), .A(n19184), .ZN(P2_U2942) );
  AOI22_X1 U22161 ( .A1(n9798), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19186) );
  OAI21_X1 U22162 ( .B1(n11489), .B2(n19203), .A(n19186), .ZN(P2_U2943) );
  AOI22_X1 U22163 ( .A1(n9798), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19187) );
  OAI21_X1 U22164 ( .B1(n19188), .B2(n19203), .A(n19187), .ZN(P2_U2944) );
  AOI22_X1 U22165 ( .A1(n9798), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19189) );
  OAI21_X1 U22166 ( .B1(n19190), .B2(n19203), .A(n19189), .ZN(P2_U2945) );
  INV_X1 U22167 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19192) );
  AOI22_X1 U22168 ( .A1(n9798), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19191) );
  OAI21_X1 U22169 ( .B1(n19192), .B2(n19203), .A(n19191), .ZN(P2_U2946) );
  AOI22_X1 U22170 ( .A1(n9798), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19193) );
  OAI21_X1 U22171 ( .B1(n19194), .B2(n19203), .A(n19193), .ZN(P2_U2947) );
  INV_X1 U22172 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19196) );
  AOI22_X1 U22173 ( .A1(n9798), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19195) );
  OAI21_X1 U22174 ( .B1(n19196), .B2(n19203), .A(n19195), .ZN(P2_U2948) );
  AOI22_X1 U22175 ( .A1(n9798), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19197) );
  OAI21_X1 U22176 ( .B1(n19198), .B2(n19203), .A(n19197), .ZN(P2_U2949) );
  INV_X1 U22177 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19200) );
  AOI22_X1 U22178 ( .A1(n9798), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19199) );
  OAI21_X1 U22179 ( .B1(n19200), .B2(n19203), .A(n19199), .ZN(P2_U2950) );
  AOI22_X1 U22180 ( .A1(n9798), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19201), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19202) );
  OAI21_X1 U22181 ( .B1(n11501), .B2(n19203), .A(n19202), .ZN(P2_U2951) );
  AOI22_X1 U22182 ( .A1(n19232), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19231), .ZN(n19206) );
  NAND2_X1 U22183 ( .A1(n19205), .A2(n19204), .ZN(n19211) );
  NAND2_X1 U22184 ( .A1(n19206), .A2(n19211), .ZN(P2_U2952) );
  AOI22_X1 U22185 ( .A1(n19232), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19231), .ZN(n19207) );
  OAI21_X1 U22186 ( .B1(n19224), .B2(n19234), .A(n19207), .ZN(P2_U2961) );
  AOI22_X1 U22187 ( .A1(n19232), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19231), .ZN(n19208) );
  OAI21_X1 U22188 ( .B1(n19226), .B2(n19234), .A(n19208), .ZN(P2_U2963) );
  AOI22_X1 U22189 ( .A1(n19232), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n19231), .ZN(n19209) );
  OAI21_X1 U22190 ( .B1(n19228), .B2(n19234), .A(n19209), .ZN(P2_U2964) );
  AOI22_X1 U22191 ( .A1(n19232), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19231), .ZN(n19210) );
  OAI21_X1 U22192 ( .B1(n19230), .B2(n19234), .A(n19210), .ZN(P2_U2965) );
  AOI22_X1 U22193 ( .A1(n19232), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n19231), .ZN(n19212) );
  NAND2_X1 U22194 ( .A1(n19212), .A2(n19211), .ZN(P2_U2967) );
  AOI22_X1 U22195 ( .A1(n19232), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19231), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n19213) );
  OAI21_X1 U22196 ( .B1(n19214), .B2(n19234), .A(n19213), .ZN(P2_U2968) );
  AOI22_X1 U22197 ( .A1(n19232), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19231), .ZN(n19215) );
  OAI21_X1 U22198 ( .B1(n19216), .B2(n19234), .A(n19215), .ZN(P2_U2970) );
  AOI22_X1 U22199 ( .A1(n19232), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19231), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n19217) );
  OAI21_X1 U22200 ( .B1(n19218), .B2(n19234), .A(n19217), .ZN(P2_U2972) );
  AOI22_X1 U22201 ( .A1(n19232), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19231), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n19219) );
  OAI21_X1 U22202 ( .B1(n19220), .B2(n19234), .A(n19219), .ZN(P2_U2973) );
  AOI22_X1 U22203 ( .A1(n19232), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19231), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n19221) );
  OAI21_X1 U22204 ( .B1(n19222), .B2(n19234), .A(n19221), .ZN(P2_U2974) );
  AOI22_X1 U22205 ( .A1(n19232), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n19231), .ZN(n19223) );
  OAI21_X1 U22206 ( .B1(n19224), .B2(n19234), .A(n19223), .ZN(P2_U2976) );
  AOI22_X1 U22207 ( .A1(n19232), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n19231), .ZN(n19225) );
  OAI21_X1 U22208 ( .B1(n19226), .B2(n19234), .A(n19225), .ZN(P2_U2978) );
  AOI22_X1 U22209 ( .A1(n19232), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n19231), .ZN(n19227) );
  OAI21_X1 U22210 ( .B1(n19228), .B2(n19234), .A(n19227), .ZN(P2_U2979) );
  AOI22_X1 U22211 ( .A1(n19232), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19231), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n19229) );
  OAI21_X1 U22212 ( .B1(n19230), .B2(n19234), .A(n19229), .ZN(P2_U2980) );
  AOI22_X1 U22213 ( .A1(n19232), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(
        P2_EAX_REG_15__SCAN_IN), .B2(n19231), .ZN(n19233) );
  OAI21_X1 U22214 ( .B1(n19235), .B2(n19234), .A(n19233), .ZN(P2_U2982) );
  AOI22_X1 U22215 ( .A1(n19237), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19236), .ZN(n19245) );
  AOI222_X1 U22216 ( .A1(n19243), .A2(n19242), .B1(n19241), .B2(n19240), .C1(
        n9787), .C2(n19238), .ZN(n19244) );
  OAI211_X1 U22217 ( .C1(n19247), .C2(n19246), .A(n19245), .B(n19244), .ZN(
        P2_U3010) );
  INV_X1 U22218 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n21091) );
  INV_X1 U22219 ( .A(n19665), .ZN(n19702) );
  AOI22_X1 U22220 ( .A1(n19271), .A2(n19702), .B1(n19701), .B2(n19270), .ZN(
        n19250) );
  AOI22_X1 U22221 ( .A1(n19265), .A2(n19710), .B1(n19305), .B2(n19662), .ZN(
        n19249) );
  OAI211_X1 U22222 ( .C1(n19255), .C2(n21091), .A(n19250), .B(n19249), .ZN(
        P2_U3056) );
  INV_X1 U22223 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n19254) );
  AOI22_X1 U22224 ( .A1(n19271), .A2(n19715), .B1(n19714), .B2(n19270), .ZN(
        n19253) );
  AOI22_X1 U22225 ( .A1(n19265), .A2(n19716), .B1(n19305), .B2(n19666), .ZN(
        n19252) );
  OAI211_X1 U22226 ( .C1(n19255), .C2(n19254), .A(n19253), .B(n19252), .ZN(
        P2_U3057) );
  INV_X1 U22227 ( .A(n19728), .ZN(n19632) );
  AOI22_X1 U22228 ( .A1(n19271), .A2(n19727), .B1(n19726), .B2(n19270), .ZN(
        n19258) );
  AOI22_X1 U22229 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19272), .B1(
        n19305), .B2(n19674), .ZN(n19257) );
  OAI211_X1 U22230 ( .C1(n19632), .C2(n19275), .A(n19258), .B(n19257), .ZN(
        P2_U3059) );
  INV_X1 U22231 ( .A(n19305), .ZN(n19268) );
  AOI22_X1 U22232 ( .A1(n19271), .A2(n19733), .B1(n19732), .B2(n19270), .ZN(
        n19260) );
  AOI22_X1 U22233 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19272), .B1(
        n19265), .B2(n19734), .ZN(n19259) );
  OAI211_X1 U22234 ( .C1(n19737), .C2(n19268), .A(n19260), .B(n19259), .ZN(
        P2_U3060) );
  INV_X1 U22235 ( .A(n19740), .ZN(n19638) );
  AOI22_X1 U22236 ( .A1(n19271), .A2(n19739), .B1(n19738), .B2(n19270), .ZN(
        n19263) );
  AOI22_X1 U22237 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19272), .B1(
        n19305), .B2(n19682), .ZN(n19262) );
  OAI211_X1 U22238 ( .C1(n19638), .C2(n19275), .A(n19263), .B(n19262), .ZN(
        P2_U3061) );
  INV_X1 U22239 ( .A(n19686), .ZN(n19749) );
  AOI22_X1 U22240 ( .A1(n19745), .A2(n19271), .B1(n19744), .B2(n19270), .ZN(
        n19267) );
  AOI22_X1 U22241 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19272), .B1(
        n19265), .B2(n19746), .ZN(n19266) );
  OAI211_X1 U22242 ( .C1(n19749), .C2(n19268), .A(n19267), .B(n19266), .ZN(
        P2_U3062) );
  INV_X1 U22243 ( .A(n19754), .ZN(n19647) );
  AOI22_X1 U22244 ( .A1(n19271), .A2(n19752), .B1(n19750), .B2(n19270), .ZN(
        n19274) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19272), .B1(
        n19305), .B2(n19692), .ZN(n19273) );
  OAI211_X1 U22246 ( .C1(n19647), .C2(n19275), .A(n19274), .B(n19273), .ZN(
        P2_U3063) );
  NOR2_X2 U22247 ( .A1(n19401), .A2(n19847), .ZN(n19337) );
  NOR2_X1 U22248 ( .A1(n19539), .A2(n19311), .ZN(n19276) );
  AOI221_X1 U22249 ( .B1(n19337), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19305), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19276), .ZN(n19280) );
  INV_X1 U22250 ( .A(n19281), .ZN(n19277) );
  AOI21_X1 U22251 ( .B1(n19277), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19278) );
  NOR3_X2 U22252 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19873), .A3(
        n19311), .ZN(n19303) );
  NOR2_X1 U22253 ( .A1(n19278), .A2(n19303), .ZN(n19279) );
  INV_X1 U22254 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n19285) );
  OAI21_X1 U22255 ( .B1(n19281), .B2(n19303), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19282) );
  OAI21_X1 U22256 ( .B1(n19311), .B2(n19539), .A(n19282), .ZN(n19304) );
  AOI22_X1 U22257 ( .A1(n19304), .A2(n19702), .B1(n19701), .B2(n19303), .ZN(
        n19284) );
  AOI22_X1 U22258 ( .A1(n19337), .A2(n19662), .B1(n19305), .B2(n19710), .ZN(
        n19283) );
  OAI211_X1 U22259 ( .C1(n19309), .C2(n19285), .A(n19284), .B(n19283), .ZN(
        P2_U3064) );
  INV_X1 U22260 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n19288) );
  AOI22_X1 U22261 ( .A1(n19304), .A2(n19715), .B1(n19714), .B2(n19303), .ZN(
        n19287) );
  AOI22_X1 U22262 ( .A1(n19305), .A2(n19716), .B1(n19337), .B2(n19666), .ZN(
        n19286) );
  OAI211_X1 U22263 ( .C1(n19309), .C2(n19288), .A(n19287), .B(n19286), .ZN(
        P2_U3065) );
  INV_X1 U22264 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n19291) );
  AOI22_X1 U22265 ( .A1(n19304), .A2(n19721), .B1(n19720), .B2(n19303), .ZN(
        n19290) );
  AOI22_X1 U22266 ( .A1(n19305), .A2(n19722), .B1(n19337), .B2(n19670), .ZN(
        n19289) );
  OAI211_X1 U22267 ( .C1(n19309), .C2(n19291), .A(n19290), .B(n19289), .ZN(
        P2_U3066) );
  AOI22_X1 U22268 ( .A1(n19304), .A2(n19727), .B1(n19726), .B2(n19303), .ZN(
        n19293) );
  AOI22_X1 U22269 ( .A1(n19305), .A2(n19728), .B1(n19337), .B2(n19674), .ZN(
        n19292) );
  OAI211_X1 U22270 ( .C1(n19309), .C2(n19294), .A(n19293), .B(n19292), .ZN(
        P2_U3067) );
  AOI22_X1 U22271 ( .A1(n19304), .A2(n19733), .B1(n19732), .B2(n19303), .ZN(
        n19296) );
  AOI22_X1 U22272 ( .A1(n19305), .A2(n19734), .B1(n19337), .B2(n19678), .ZN(
        n19295) );
  OAI211_X1 U22273 ( .C1(n19309), .C2(n10963), .A(n19296), .B(n19295), .ZN(
        P2_U3068) );
  INV_X1 U22274 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n19299) );
  AOI22_X1 U22275 ( .A1(n19304), .A2(n19739), .B1(n19738), .B2(n19303), .ZN(
        n19298) );
  AOI22_X1 U22276 ( .A1(n19337), .A2(n19682), .B1(n19305), .B2(n19740), .ZN(
        n19297) );
  OAI211_X1 U22277 ( .C1(n19309), .C2(n19299), .A(n19298), .B(n19297), .ZN(
        P2_U3069) );
  INV_X1 U22278 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n19302) );
  AOI22_X1 U22279 ( .A1(n19745), .A2(n19304), .B1(n19744), .B2(n19303), .ZN(
        n19301) );
  AOI22_X1 U22280 ( .A1(n19305), .A2(n19746), .B1(n19337), .B2(n19686), .ZN(
        n19300) );
  OAI211_X1 U22281 ( .C1(n19309), .C2(n19302), .A(n19301), .B(n19300), .ZN(
        P2_U3070) );
  INV_X1 U22282 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n19308) );
  AOI22_X1 U22283 ( .A1(n19304), .A2(n19752), .B1(n19750), .B2(n19303), .ZN(
        n19307) );
  AOI22_X1 U22284 ( .A1(n19337), .A2(n19692), .B1(n19305), .B2(n19754), .ZN(
        n19306) );
  OAI211_X1 U22285 ( .C1(n19309), .C2(n19308), .A(n19307), .B(n19306), .ZN(
        P2_U3071) );
  INV_X1 U22286 ( .A(n19434), .ZN(n19373) );
  INV_X1 U22287 ( .A(n19847), .ZN(n19310) );
  AOI21_X1 U22288 ( .B1(n19373), .B2(n19310), .A(n15596), .ZN(n19315) );
  NOR2_X1 U22289 ( .A1(n19873), .A2(n19311), .ZN(n19320) );
  INV_X1 U22290 ( .A(n19316), .ZN(n19313) );
  NOR2_X1 U22291 ( .A1(n19312), .A2(n19311), .ZN(n19336) );
  INV_X1 U22292 ( .A(n19336), .ZN(n19317) );
  AOI21_X1 U22293 ( .B1(n19313), .B2(n19317), .A(n19654), .ZN(n19314) );
  NOR2_X2 U22294 ( .A1(n19441), .A2(n19847), .ZN(n19367) );
  AOI22_X1 U22295 ( .A1(n19662), .A2(n19367), .B1(n19701), .B2(n19336), .ZN(
        n19323) );
  INV_X1 U22296 ( .A(n19315), .ZN(n19321) );
  OAI21_X1 U22297 ( .B1(n19316), .B2(n19654), .A(n19469), .ZN(n19318) );
  AOI21_X1 U22298 ( .B1(n19318), .B2(n19317), .A(n19536), .ZN(n19319) );
  OAI21_X1 U22299 ( .B1(n19321), .B2(n19320), .A(n19319), .ZN(n19338) );
  AOI22_X1 U22300 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19338), .B1(
        n19337), .B2(n19710), .ZN(n19322) );
  OAI211_X1 U22301 ( .C1(n19341), .C2(n19665), .A(n19323), .B(n19322), .ZN(
        P2_U3072) );
  AOI22_X1 U22302 ( .A1(n19666), .A2(n19367), .B1(n19714), .B2(n19336), .ZN(
        n19325) );
  AOI22_X1 U22303 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19338), .B1(
        n19337), .B2(n19716), .ZN(n19324) );
  OAI211_X1 U22304 ( .C1(n19341), .C2(n19669), .A(n19325), .B(n19324), .ZN(
        P2_U3073) );
  AOI22_X1 U22305 ( .A1(n19722), .A2(n19337), .B1(n19720), .B2(n19336), .ZN(
        n19327) );
  AOI22_X1 U22306 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19338), .B1(
        n19367), .B2(n19670), .ZN(n19326) );
  OAI211_X1 U22307 ( .C1(n19341), .C2(n19673), .A(n19327), .B(n19326), .ZN(
        P2_U3074) );
  AOI22_X1 U22308 ( .A1(n19674), .A2(n19367), .B1(n19726), .B2(n19336), .ZN(
        n19329) );
  AOI22_X1 U22309 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19338), .B1(
        n19337), .B2(n19728), .ZN(n19328) );
  OAI211_X1 U22310 ( .C1(n19341), .C2(n19677), .A(n19329), .B(n19328), .ZN(
        P2_U3075) );
  AOI22_X1 U22311 ( .A1(n19734), .A2(n19337), .B1(n19732), .B2(n19336), .ZN(
        n19331) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19338), .B1(
        n19367), .B2(n19678), .ZN(n19330) );
  OAI211_X1 U22313 ( .C1(n19341), .C2(n19681), .A(n19331), .B(n19330), .ZN(
        P2_U3076) );
  AOI22_X1 U22314 ( .A1(n19682), .A2(n19367), .B1(n19738), .B2(n19336), .ZN(
        n19333) );
  AOI22_X1 U22315 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19338), .B1(
        n19337), .B2(n19740), .ZN(n19332) );
  OAI211_X1 U22316 ( .C1(n19341), .C2(n19685), .A(n19333), .B(n19332), .ZN(
        P2_U3077) );
  AOI22_X1 U22317 ( .A1(n19746), .A2(n19337), .B1(n19744), .B2(n19336), .ZN(
        n19335) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19338), .B1(
        n19367), .B2(n19686), .ZN(n19334) );
  OAI211_X1 U22319 ( .C1(n19341), .C2(n19689), .A(n19335), .B(n19334), .ZN(
        P2_U3078) );
  AOI22_X1 U22320 ( .A1(n19754), .A2(n19337), .B1(n19750), .B2(n19336), .ZN(
        n19340) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19338), .B1(
        n19367), .B2(n19692), .ZN(n19339) );
  OAI211_X1 U22322 ( .C1(n19341), .C2(n19696), .A(n19340), .B(n19339), .ZN(
        P2_U3079) );
  INV_X1 U22323 ( .A(n19662), .ZN(n19713) );
  INV_X1 U22324 ( .A(n19407), .ZN(n19344) );
  NOR2_X1 U22325 ( .A1(n19344), .A2(n19343), .ZN(n19591) );
  NAND2_X1 U22326 ( .A1(n19591), .A2(n19858), .ZN(n19349) );
  AND2_X1 U22327 ( .A1(n19402), .A2(n19466), .ZN(n19365) );
  OAI21_X1 U22328 ( .B1(n19346), .B2(n19365), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19345) );
  OAI21_X1 U22329 ( .B1(n19349), .B2(n15596), .A(n19345), .ZN(n19366) );
  AOI22_X1 U22330 ( .A1(n19366), .A2(n19702), .B1(n19701), .B2(n19365), .ZN(
        n19352) );
  OAI21_X1 U22331 ( .B1(n19367), .B2(n19396), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19348) );
  AOI211_X1 U22332 ( .C1(n19346), .C2(n19469), .A(n19365), .B(n19648), .ZN(
        n19347) );
  AOI211_X1 U22333 ( .C1(n19349), .C2(n19348), .A(n19536), .B(n19347), .ZN(
        n19350) );
  AOI22_X1 U22334 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19368), .B1(
        n19367), .B2(n19710), .ZN(n19351) );
  OAI211_X1 U22335 ( .C1(n19713), .C2(n19371), .A(n19352), .B(n19351), .ZN(
        P2_U3080) );
  INV_X1 U22336 ( .A(n19666), .ZN(n19719) );
  AOI22_X1 U22337 ( .A1(n19366), .A2(n19715), .B1(n19714), .B2(n19365), .ZN(
        n19354) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19368), .B1(
        n19367), .B2(n19716), .ZN(n19353) );
  OAI211_X1 U22339 ( .C1(n19719), .C2(n19371), .A(n19354), .B(n19353), .ZN(
        P2_U3081) );
  INV_X1 U22340 ( .A(n19670), .ZN(n19725) );
  AOI22_X1 U22341 ( .A1(n19366), .A2(n19721), .B1(n19720), .B2(n19365), .ZN(
        n19356) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19368), .B1(
        n19367), .B2(n19722), .ZN(n19355) );
  OAI211_X1 U22343 ( .C1(n19725), .C2(n19371), .A(n19356), .B(n19355), .ZN(
        P2_U3082) );
  INV_X1 U22344 ( .A(n19674), .ZN(n19731) );
  AOI22_X1 U22345 ( .A1(n19366), .A2(n19727), .B1(n19726), .B2(n19365), .ZN(
        n19358) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19368), .B1(
        n19367), .B2(n19728), .ZN(n19357) );
  OAI211_X1 U22347 ( .C1(n19731), .C2(n19371), .A(n19358), .B(n19357), .ZN(
        P2_U3083) );
  AOI22_X1 U22348 ( .A1(n19366), .A2(n19733), .B1(n19732), .B2(n19365), .ZN(
        n19360) );
  AOI22_X1 U22349 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19368), .B1(
        n19367), .B2(n19734), .ZN(n19359) );
  OAI211_X1 U22350 ( .C1(n19737), .C2(n19371), .A(n19360), .B(n19359), .ZN(
        P2_U3084) );
  INV_X1 U22351 ( .A(n19682), .ZN(n19743) );
  AOI22_X1 U22352 ( .A1(n19366), .A2(n19739), .B1(n19738), .B2(n19365), .ZN(
        n19362) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19368), .B1(
        n19367), .B2(n19740), .ZN(n19361) );
  OAI211_X1 U22354 ( .C1(n19743), .C2(n19371), .A(n19362), .B(n19361), .ZN(
        P2_U3085) );
  AOI22_X1 U22355 ( .A1(n19745), .A2(n19366), .B1(n19744), .B2(n19365), .ZN(
        n19364) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19368), .B1(
        n19367), .B2(n19746), .ZN(n19363) );
  OAI211_X1 U22357 ( .C1(n19749), .C2(n19371), .A(n19364), .B(n19363), .ZN(
        P2_U3086) );
  INV_X1 U22358 ( .A(n19692), .ZN(n19760) );
  AOI22_X1 U22359 ( .A1(n19366), .A2(n19752), .B1(n19750), .B2(n19365), .ZN(
        n19370) );
  AOI22_X1 U22360 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19368), .B1(
        n19367), .B2(n19754), .ZN(n19369) );
  OAI211_X1 U22361 ( .C1(n19760), .C2(n19371), .A(n19370), .B(n19369), .ZN(
        P2_U3087) );
  INV_X1 U22362 ( .A(n19619), .ZN(n19372) );
  AOI21_X1 U22363 ( .B1(n19373), .B2(n19372), .A(n15596), .ZN(n19376) );
  AND2_X1 U22364 ( .A1(n19873), .A2(n19402), .ZN(n19379) );
  NAND2_X1 U22365 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19379), .ZN(
        n19377) );
  AOI21_X1 U22366 ( .B1(n19374), .B2(n19377), .A(n19654), .ZN(n19375) );
  NOR2_X2 U22367 ( .A1(n19441), .A2(n19619), .ZN(n19429) );
  INV_X1 U22368 ( .A(n19377), .ZN(n19395) );
  AOI22_X1 U22369 ( .A1(n19662), .A2(n19429), .B1(n19701), .B2(n19395), .ZN(
        n19382) );
  INV_X1 U22370 ( .A(n19376), .ZN(n19380) );
  OAI211_X1 U22371 ( .C1(n19374), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19377), 
        .B(n15596), .ZN(n19378) );
  OAI211_X1 U22372 ( .C1(n19380), .C2(n19379), .A(n19707), .B(n19378), .ZN(
        n19397) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19397), .B1(
        n19396), .B2(n19710), .ZN(n19381) );
  OAI211_X1 U22374 ( .C1(n19400), .C2(n19665), .A(n19382), .B(n19381), .ZN(
        P2_U3088) );
  AOI22_X1 U22375 ( .A1(n19716), .A2(n19396), .B1(n19714), .B2(n19395), .ZN(
        n19384) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19397), .B1(
        n19429), .B2(n19666), .ZN(n19383) );
  OAI211_X1 U22377 ( .C1(n19400), .C2(n19669), .A(n19384), .B(n19383), .ZN(
        P2_U3089) );
  AOI22_X1 U22378 ( .A1(n19722), .A2(n19396), .B1(n19720), .B2(n19395), .ZN(
        n19386) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19397), .B1(
        n19429), .B2(n19670), .ZN(n19385) );
  OAI211_X1 U22380 ( .C1(n19400), .C2(n19673), .A(n19386), .B(n19385), .ZN(
        P2_U3090) );
  AOI22_X1 U22381 ( .A1(n19674), .A2(n19429), .B1(n19726), .B2(n19395), .ZN(
        n19388) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19397), .B1(
        n19396), .B2(n19728), .ZN(n19387) );
  OAI211_X1 U22383 ( .C1(n19400), .C2(n19677), .A(n19388), .B(n19387), .ZN(
        P2_U3091) );
  AOI22_X1 U22384 ( .A1(n19734), .A2(n19396), .B1(n19732), .B2(n19395), .ZN(
        n19390) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19397), .B1(
        n19429), .B2(n19678), .ZN(n19389) );
  OAI211_X1 U22386 ( .C1(n19400), .C2(n19681), .A(n19390), .B(n19389), .ZN(
        P2_U3092) );
  AOI22_X1 U22387 ( .A1(n19682), .A2(n19429), .B1(n19738), .B2(n19395), .ZN(
        n19392) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19397), .B1(
        n19396), .B2(n19740), .ZN(n19391) );
  OAI211_X1 U22389 ( .C1(n19400), .C2(n19685), .A(n19392), .B(n19391), .ZN(
        P2_U3093) );
  AOI22_X1 U22390 ( .A1(n19686), .A2(n19429), .B1(n19744), .B2(n19395), .ZN(
        n19394) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19397), .B1(
        n19396), .B2(n19746), .ZN(n19393) );
  OAI211_X1 U22392 ( .C1(n19400), .C2(n19689), .A(n19394), .B(n19393), .ZN(
        P2_U3094) );
  AOI22_X1 U22393 ( .A1(n19754), .A2(n19396), .B1(n19750), .B2(n19395), .ZN(
        n19399) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19397), .B1(
        n19429), .B2(n19692), .ZN(n19398) );
  OAI211_X1 U22395 ( .C1(n19400), .C2(n19696), .A(n19399), .B(n19398), .ZN(
        P2_U3095) );
  INV_X1 U22396 ( .A(n19402), .ZN(n19406) );
  NAND2_X1 U22397 ( .A1(n19699), .A2(n19858), .ZN(n19435) );
  NOR2_X1 U22398 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19435), .ZN(
        n19427) );
  OAI21_X1 U22399 ( .B1(n19408), .B2(n19427), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19403) );
  OAI21_X1 U22400 ( .B1(n19406), .B2(n19539), .A(n19403), .ZN(n19428) );
  AOI22_X1 U22401 ( .A1(n19428), .A2(n19702), .B1(n19701), .B2(n19427), .ZN(
        n19414) );
  OAI21_X1 U22402 ( .B1(n19429), .B2(n19404), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19405) );
  OAI21_X1 U22403 ( .B1(n19407), .B2(n19406), .A(n19405), .ZN(n19412) );
  INV_X1 U22404 ( .A(n19408), .ZN(n19410) );
  INV_X1 U22405 ( .A(n19427), .ZN(n19409) );
  OAI211_X1 U22406 ( .C1(n19410), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19409), 
        .B(n15596), .ZN(n19411) );
  NAND3_X1 U22407 ( .A1(n19412), .A2(n19707), .A3(n19411), .ZN(n19430) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19710), .ZN(n19413) );
  OAI211_X1 U22409 ( .C1(n19713), .C2(n19461), .A(n19414), .B(n19413), .ZN(
        P2_U3096) );
  AOI22_X1 U22410 ( .A1(n19428), .A2(n19715), .B1(n19714), .B2(n19427), .ZN(
        n19416) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19716), .ZN(n19415) );
  OAI211_X1 U22412 ( .C1(n19719), .C2(n19461), .A(n19416), .B(n19415), .ZN(
        P2_U3097) );
  AOI22_X1 U22413 ( .A1(n19428), .A2(n19721), .B1(n19720), .B2(n19427), .ZN(
        n19418) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19722), .ZN(n19417) );
  OAI211_X1 U22415 ( .C1(n19725), .C2(n19461), .A(n19418), .B(n19417), .ZN(
        P2_U3098) );
  AOI22_X1 U22416 ( .A1(n19428), .A2(n19727), .B1(n19726), .B2(n19427), .ZN(
        n19420) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19728), .ZN(n19419) );
  OAI211_X1 U22418 ( .C1(n19731), .C2(n19461), .A(n19420), .B(n19419), .ZN(
        P2_U3099) );
  AOI22_X1 U22419 ( .A1(n19428), .A2(n19733), .B1(n19732), .B2(n19427), .ZN(
        n19422) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19734), .ZN(n19421) );
  OAI211_X1 U22421 ( .C1(n19737), .C2(n19461), .A(n19422), .B(n19421), .ZN(
        P2_U3100) );
  AOI22_X1 U22422 ( .A1(n19428), .A2(n19739), .B1(n19738), .B2(n19427), .ZN(
        n19424) );
  AOI22_X1 U22423 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19740), .ZN(n19423) );
  OAI211_X1 U22424 ( .C1(n19743), .C2(n19461), .A(n19424), .B(n19423), .ZN(
        P2_U3101) );
  AOI22_X1 U22425 ( .A1(n19745), .A2(n19428), .B1(n19744), .B2(n19427), .ZN(
        n19426) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19746), .ZN(n19425) );
  OAI211_X1 U22427 ( .C1(n19749), .C2(n19461), .A(n19426), .B(n19425), .ZN(
        P2_U3102) );
  AOI22_X1 U22428 ( .A1(n19428), .A2(n19752), .B1(n19750), .B2(n19427), .ZN(
        n19432) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19754), .ZN(n19431) );
  OAI211_X1 U22430 ( .C1(n19760), .C2(n19461), .A(n19432), .B(n19431), .ZN(
        P2_U3103) );
  INV_X1 U22431 ( .A(n19710), .ZN(n19623) );
  INV_X1 U22432 ( .A(n19471), .ZN(n19456) );
  OAI21_X1 U22433 ( .B1(n19436), .B2(n19456), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19433) );
  OAI21_X1 U22434 ( .B1(n19435), .B2(n15596), .A(n19433), .ZN(n19457) );
  AOI22_X1 U22435 ( .A1(n19457), .A2(n19702), .B1(n19456), .B2(n19701), .ZN(
        n19443) );
  OR2_X1 U22436 ( .A1(n19434), .A2(n19705), .ZN(n19855) );
  INV_X1 U22437 ( .A(n19855), .ZN(n19440) );
  INV_X1 U22438 ( .A(n19435), .ZN(n19439) );
  INV_X1 U22439 ( .A(n19436), .ZN(n19437) );
  OAI211_X1 U22440 ( .C1(n19437), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19471), 
        .B(n15596), .ZN(n19438) );
  OAI211_X1 U22441 ( .C1(n19440), .C2(n19439), .A(n19707), .B(n19438), .ZN(
        n19458) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19458), .B1(
        n19489), .B2(n19662), .ZN(n19442) );
  OAI211_X1 U22443 ( .C1(n19623), .C2(n19461), .A(n19443), .B(n19442), .ZN(
        P2_U3104) );
  INV_X1 U22444 ( .A(n19716), .ZN(n19626) );
  AOI22_X1 U22445 ( .A1(n19457), .A2(n19715), .B1(n19456), .B2(n19714), .ZN(
        n19445) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19458), .B1(
        n19489), .B2(n19666), .ZN(n19444) );
  OAI211_X1 U22447 ( .C1(n19626), .C2(n19461), .A(n19445), .B(n19444), .ZN(
        P2_U3105) );
  INV_X1 U22448 ( .A(n19722), .ZN(n19629) );
  AOI22_X1 U22449 ( .A1(n19457), .A2(n19721), .B1(n19456), .B2(n19720), .ZN(
        n19447) );
  AOI22_X1 U22450 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19458), .B1(
        n19489), .B2(n19670), .ZN(n19446) );
  OAI211_X1 U22451 ( .C1(n19629), .C2(n19461), .A(n19447), .B(n19446), .ZN(
        P2_U3106) );
  AOI22_X1 U22452 ( .A1(n19457), .A2(n19727), .B1(n19456), .B2(n19726), .ZN(
        n19449) );
  AOI22_X1 U22453 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19458), .B1(
        n19489), .B2(n19674), .ZN(n19448) );
  OAI211_X1 U22454 ( .C1(n19632), .C2(n19461), .A(n19449), .B(n19448), .ZN(
        P2_U3107) );
  INV_X1 U22455 ( .A(n19734), .ZN(n19635) );
  AOI22_X1 U22456 ( .A1(n19457), .A2(n19733), .B1(n19456), .B2(n19732), .ZN(
        n19451) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19458), .B1(
        n19489), .B2(n19678), .ZN(n19450) );
  OAI211_X1 U22458 ( .C1(n19635), .C2(n19461), .A(n19451), .B(n19450), .ZN(
        P2_U3108) );
  AOI22_X1 U22459 ( .A1(n19457), .A2(n19739), .B1(n19456), .B2(n19738), .ZN(
        n19453) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19458), .B1(
        n19489), .B2(n19682), .ZN(n19452) );
  OAI211_X1 U22461 ( .C1(n19638), .C2(n19461), .A(n19453), .B(n19452), .ZN(
        P2_U3109) );
  INV_X1 U22462 ( .A(n19746), .ZN(n19641) );
  AOI22_X1 U22463 ( .A1(n19745), .A2(n19457), .B1(n19456), .B2(n19744), .ZN(
        n19455) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19458), .B1(
        n19489), .B2(n19686), .ZN(n19454) );
  OAI211_X1 U22465 ( .C1(n19641), .C2(n19461), .A(n19455), .B(n19454), .ZN(
        P2_U3110) );
  AOI22_X1 U22466 ( .A1(n19457), .A2(n19752), .B1(n19456), .B2(n19750), .ZN(
        n19460) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19458), .B1(
        n19489), .B2(n19692), .ZN(n19459) );
  OAI211_X1 U22468 ( .C1(n19647), .C2(n19461), .A(n19460), .B(n19459), .ZN(
        P2_U3111) );
  INV_X1 U22469 ( .A(n19650), .ZN(n19462) );
  INV_X1 U22470 ( .A(n19502), .ZN(n19494) );
  NAND3_X1 U22471 ( .A1(n19528), .A2(n19648), .A3(n19463), .ZN(n19464) );
  INV_X1 U22472 ( .A(n10988), .ZN(n19465) );
  AOI22_X1 U22473 ( .A1(n19467), .A2(n19465), .B1(n19654), .B2(n19471), .ZN(
        n19468) );
  AND2_X1 U22474 ( .A1(n19466), .A2(n19497), .ZN(n19488) );
  INV_X1 U22475 ( .A(n19467), .ZN(n19472) );
  AOI22_X1 U22476 ( .A1(n19710), .A2(n19489), .B1(n19701), .B2(n19488), .ZN(
        n19475) );
  OAI21_X1 U22477 ( .B1(n10988), .B2(n19654), .A(n19469), .ZN(n19470) );
  AOI21_X1 U22478 ( .B1(n19472), .B2(n19471), .A(n19470), .ZN(n19473) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19490), .B1(
        n19519), .B2(n19662), .ZN(n19474) );
  OAI211_X1 U22480 ( .C1(n19665), .C2(n19493), .A(n19475), .B(n19474), .ZN(
        P2_U3112) );
  AOI22_X1 U22481 ( .A1(n19666), .A2(n19519), .B1(n19714), .B2(n19488), .ZN(
        n19477) );
  AOI22_X1 U22482 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19490), .B1(
        n19489), .B2(n19716), .ZN(n19476) );
  OAI211_X1 U22483 ( .C1(n19669), .C2(n19493), .A(n19477), .B(n19476), .ZN(
        P2_U3113) );
  AOI22_X1 U22484 ( .A1(n19722), .A2(n19489), .B1(n19720), .B2(n19488), .ZN(
        n19479) );
  AOI22_X1 U22485 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19490), .B1(
        n19519), .B2(n19670), .ZN(n19478) );
  OAI211_X1 U22486 ( .C1(n19673), .C2(n19493), .A(n19479), .B(n19478), .ZN(
        P2_U3114) );
  AOI22_X1 U22487 ( .A1(n19728), .A2(n19489), .B1(n19726), .B2(n19488), .ZN(
        n19481) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19490), .B1(
        n19519), .B2(n19674), .ZN(n19480) );
  OAI211_X1 U22489 ( .C1(n19677), .C2(n19493), .A(n19481), .B(n19480), .ZN(
        P2_U3115) );
  AOI22_X1 U22490 ( .A1(n19734), .A2(n19489), .B1(n19732), .B2(n19488), .ZN(
        n19483) );
  AOI22_X1 U22491 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19490), .B1(
        n19519), .B2(n19678), .ZN(n19482) );
  OAI211_X1 U22492 ( .C1(n19681), .C2(n19493), .A(n19483), .B(n19482), .ZN(
        P2_U3116) );
  AOI22_X1 U22493 ( .A1(n19682), .A2(n19519), .B1(n19738), .B2(n19488), .ZN(
        n19485) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19490), .B1(
        n19489), .B2(n19740), .ZN(n19484) );
  OAI211_X1 U22495 ( .C1(n19685), .C2(n19493), .A(n19485), .B(n19484), .ZN(
        P2_U3117) );
  AOI22_X1 U22496 ( .A1(n19686), .A2(n19519), .B1(n19744), .B2(n19488), .ZN(
        n19487) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19490), .B1(
        n19489), .B2(n19746), .ZN(n19486) );
  OAI211_X1 U22498 ( .C1(n19689), .C2(n19493), .A(n19487), .B(n19486), .ZN(
        P2_U3118) );
  AOI22_X1 U22499 ( .A1(n19692), .A2(n19519), .B1(n19750), .B2(n19488), .ZN(
        n19492) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19490), .B1(
        n19489), .B2(n19754), .ZN(n19491) );
  OAI211_X1 U22501 ( .C1(n19696), .C2(n19493), .A(n19492), .B(n19491), .ZN(
        P2_U3119) );
  INV_X1 U22502 ( .A(n19706), .ZN(n19495) );
  NAND2_X1 U22503 ( .A1(n19495), .A2(n19494), .ZN(n19496) );
  NAND2_X1 U22504 ( .A1(n19497), .A2(n19873), .ZN(n19503) );
  NAND2_X1 U22505 ( .A1(n19496), .A2(n19503), .ZN(n19500) );
  NAND2_X1 U22506 ( .A1(n10997), .A2(n19469), .ZN(n19498) );
  NAND3_X1 U22507 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19497), .A3(
        n19873), .ZN(n19529) );
  NAND2_X1 U22508 ( .A1(n19498), .A2(n19529), .ZN(n19499) );
  MUX2_X1 U22509 ( .A(n19500), .B(n19499), .S(n15596), .Z(n19501) );
  NAND2_X1 U22510 ( .A1(n19501), .A2(n19707), .ZN(n19525) );
  INV_X1 U22511 ( .A(n19525), .ZN(n19522) );
  NOR2_X2 U22512 ( .A1(n19620), .A2(n19502), .ZN(n19558) );
  INV_X1 U22513 ( .A(n19529), .ZN(n19523) );
  AOI22_X1 U22514 ( .A1(n19662), .A2(n19558), .B1(n19701), .B2(n19523), .ZN(
        n19508) );
  INV_X1 U22515 ( .A(n19503), .ZN(n19504) );
  NAND2_X1 U22516 ( .A1(n19504), .A2(n19648), .ZN(n19506) );
  OAI21_X1 U22517 ( .B1(n10997), .B2(n19523), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19505) );
  NAND2_X1 U22518 ( .A1(n19506), .A2(n19505), .ZN(n19524) );
  AOI22_X1 U22519 ( .A1(n19702), .A2(n19524), .B1(n19519), .B2(n19710), .ZN(
        n19507) );
  OAI211_X1 U22520 ( .C1(n19522), .C2(n21017), .A(n19508), .B(n19507), .ZN(
        P2_U3120) );
  INV_X1 U22521 ( .A(n19558), .ZN(n19530) );
  AOI22_X1 U22522 ( .A1(n19716), .A2(n19519), .B1(n19714), .B2(n19523), .ZN(
        n19510) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19525), .B1(
        n19715), .B2(n19524), .ZN(n19509) );
  OAI211_X1 U22524 ( .C1(n19719), .C2(n19530), .A(n19510), .B(n19509), .ZN(
        P2_U3121) );
  AOI22_X1 U22525 ( .A1(n19670), .A2(n19558), .B1(n19720), .B2(n19523), .ZN(
        n19512) );
  AOI22_X1 U22526 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19525), .B1(
        n19721), .B2(n19524), .ZN(n19511) );
  OAI211_X1 U22527 ( .C1(n19629), .C2(n19528), .A(n19512), .B(n19511), .ZN(
        P2_U3122) );
  AOI22_X1 U22528 ( .A1(n19674), .A2(n19558), .B1(n19726), .B2(n19523), .ZN(
        n19514) );
  AOI22_X1 U22529 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19525), .B1(
        n19727), .B2(n19524), .ZN(n19513) );
  OAI211_X1 U22530 ( .C1(n19632), .C2(n19528), .A(n19514), .B(n19513), .ZN(
        P2_U3123) );
  AOI22_X1 U22531 ( .A1(n19734), .A2(n19519), .B1(n19732), .B2(n19523), .ZN(
        n19516) );
  AOI22_X1 U22532 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19525), .B1(
        n19733), .B2(n19524), .ZN(n19515) );
  OAI211_X1 U22533 ( .C1(n19737), .C2(n19530), .A(n19516), .B(n19515), .ZN(
        P2_U3124) );
  AOI22_X1 U22534 ( .A1(n19682), .A2(n19558), .B1(n19738), .B2(n19523), .ZN(
        n19518) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19525), .B1(
        n19739), .B2(n19524), .ZN(n19517) );
  OAI211_X1 U22536 ( .C1(n19638), .C2(n19528), .A(n19518), .B(n19517), .ZN(
        P2_U3125) );
  AOI22_X1 U22537 ( .A1(n19686), .A2(n19558), .B1(n19744), .B2(n19523), .ZN(
        n19521) );
  AOI22_X1 U22538 ( .A1(n19745), .A2(n19524), .B1(n19519), .B2(n19746), .ZN(
        n19520) );
  OAI211_X1 U22539 ( .C1(n19522), .C2(n12623), .A(n19521), .B(n19520), .ZN(
        P2_U3126) );
  AOI22_X1 U22540 ( .A1(n19692), .A2(n19558), .B1(n19750), .B2(n19523), .ZN(
        n19527) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19525), .B1(
        n19752), .B2(n19524), .ZN(n19526) );
  OAI211_X1 U22542 ( .C1(n19647), .C2(n19528), .A(n19527), .B(n19526), .ZN(
        P2_U3127) );
  OAI221_X1 U22543 ( .B1(n19902), .B2(n19572), .C1(n19902), .C2(n19530), .A(
        n19529), .ZN(n19535) );
  NAND2_X1 U22544 ( .A1(n19469), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19532) );
  NOR3_X2 U22545 ( .A1(n19873), .A2(n19540), .A3(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19556) );
  INV_X1 U22546 ( .A(n19556), .ZN(n19531) );
  OAI21_X1 U22547 ( .B1(n19533), .B2(n19532), .A(n19531), .ZN(n19534) );
  AOI21_X1 U22548 ( .B1(n19535), .B2(n19648), .A(n19534), .ZN(n19537) );
  OAI21_X1 U22549 ( .B1(n10990), .B2(n19556), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19538) );
  OAI21_X1 U22550 ( .B1(n19540), .B2(n19539), .A(n19538), .ZN(n19557) );
  AOI22_X1 U22551 ( .A1(n19557), .A2(n19702), .B1(n19701), .B2(n19556), .ZN(
        n19542) );
  AOI22_X1 U22552 ( .A1(n19578), .A2(n19662), .B1(n19558), .B2(n19710), .ZN(
        n19541) );
  OAI211_X1 U22553 ( .C1(n19561), .C2(n19543), .A(n19542), .B(n19541), .ZN(
        P2_U3128) );
  AOI22_X1 U22554 ( .A1(n19557), .A2(n19715), .B1(n19714), .B2(n19556), .ZN(
        n19545) );
  AOI22_X1 U22555 ( .A1(n19558), .A2(n19716), .B1(n19578), .B2(n19666), .ZN(
        n19544) );
  OAI211_X1 U22556 ( .C1(n19561), .C2(n12539), .A(n19545), .B(n19544), .ZN(
        P2_U3129) );
  AOI22_X1 U22557 ( .A1(n19557), .A2(n19721), .B1(n19720), .B2(n19556), .ZN(
        n19547) );
  AOI22_X1 U22558 ( .A1(n19558), .A2(n19722), .B1(n19578), .B2(n19670), .ZN(
        n19546) );
  OAI211_X1 U22559 ( .C1(n19561), .C2(n11559), .A(n19547), .B(n19546), .ZN(
        P2_U3130) );
  AOI22_X1 U22560 ( .A1(n19557), .A2(n19727), .B1(n19726), .B2(n19556), .ZN(
        n19549) );
  AOI22_X1 U22561 ( .A1(n19558), .A2(n19728), .B1(n19578), .B2(n19674), .ZN(
        n19548) );
  OAI211_X1 U22562 ( .C1(n19561), .C2(n11582), .A(n19549), .B(n19548), .ZN(
        P2_U3131) );
  AOI22_X1 U22563 ( .A1(n19557), .A2(n19733), .B1(n19732), .B2(n19556), .ZN(
        n19551) );
  AOI22_X1 U22564 ( .A1(n19558), .A2(n19734), .B1(n19578), .B2(n19678), .ZN(
        n19550) );
  OAI211_X1 U22565 ( .C1(n19561), .C2(n12591), .A(n19551), .B(n19550), .ZN(
        P2_U3132) );
  AOI22_X1 U22566 ( .A1(n19557), .A2(n19739), .B1(n19738), .B2(n19556), .ZN(
        n19553) );
  AOI22_X1 U22567 ( .A1(n19578), .A2(n19682), .B1(n19558), .B2(n19740), .ZN(
        n19552) );
  OAI211_X1 U22568 ( .C1(n19561), .C2(n12613), .A(n19553), .B(n19552), .ZN(
        P2_U3133) );
  AOI22_X1 U22569 ( .A1(n19745), .A2(n19557), .B1(n19744), .B2(n19556), .ZN(
        n19555) );
  AOI22_X1 U22570 ( .A1(n19558), .A2(n19746), .B1(n19578), .B2(n19686), .ZN(
        n19554) );
  OAI211_X1 U22571 ( .C1(n19561), .C2(n12624), .A(n19555), .B(n19554), .ZN(
        P2_U3134) );
  AOI22_X1 U22572 ( .A1(n19557), .A2(n19752), .B1(n19750), .B2(n19556), .ZN(
        n19560) );
  AOI22_X1 U22573 ( .A1(n19578), .A2(n19692), .B1(n19558), .B2(n19754), .ZN(
        n19559) );
  OAI211_X1 U22574 ( .C1(n19561), .C2(n14309), .A(n19560), .B(n19559), .ZN(
        P2_U3135) );
  INV_X1 U22575 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n21162) );
  AOI22_X1 U22576 ( .A1(n19577), .A2(n19702), .B1(n19701), .B2(n19576), .ZN(
        n19563) );
  AOI22_X1 U22577 ( .A1(n19609), .A2(n19662), .B1(n19578), .B2(n19710), .ZN(
        n19562) );
  OAI211_X1 U22578 ( .C1(n19581), .C2(n21162), .A(n19563), .B(n19562), .ZN(
        P2_U3136) );
  AOI22_X1 U22579 ( .A1(n19577), .A2(n19715), .B1(n19714), .B2(n19576), .ZN(
        n19565) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19573), .B1(
        n19609), .B2(n19666), .ZN(n19564) );
  OAI211_X1 U22581 ( .C1(n19626), .C2(n19572), .A(n19565), .B(n19564), .ZN(
        P2_U3137) );
  AOI22_X1 U22582 ( .A1(n19577), .A2(n19721), .B1(n19720), .B2(n19576), .ZN(
        n19567) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19573), .B1(
        n19609), .B2(n19670), .ZN(n19566) );
  OAI211_X1 U22584 ( .C1(n19629), .C2(n19572), .A(n19567), .B(n19566), .ZN(
        P2_U3138) );
  AOI22_X1 U22585 ( .A1(n19577), .A2(n19727), .B1(n19726), .B2(n19576), .ZN(
        n19569) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19573), .B1(
        n19609), .B2(n19674), .ZN(n19568) );
  OAI211_X1 U22587 ( .C1(n19632), .C2(n19572), .A(n19569), .B(n19568), .ZN(
        P2_U3139) );
  AOI22_X1 U22588 ( .A1(n19577), .A2(n19739), .B1(n19738), .B2(n19576), .ZN(
        n19571) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19573), .B1(
        n19609), .B2(n19682), .ZN(n19570) );
  OAI211_X1 U22590 ( .C1(n19638), .C2(n19572), .A(n19571), .B(n19570), .ZN(
        P2_U3141) );
  INV_X1 U22591 ( .A(n19609), .ZN(n19586) );
  AOI22_X1 U22592 ( .A1(n19745), .A2(n19577), .B1(n19744), .B2(n19576), .ZN(
        n19575) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19573), .B1(
        n19578), .B2(n19746), .ZN(n19574) );
  OAI211_X1 U22594 ( .C1(n19749), .C2(n19586), .A(n19575), .B(n19574), .ZN(
        P2_U3142) );
  AOI22_X1 U22595 ( .A1(n19577), .A2(n19752), .B1(n19750), .B2(n19576), .ZN(
        n19580) );
  AOI22_X1 U22596 ( .A1(n19609), .A2(n19692), .B1(n19578), .B2(n19754), .ZN(
        n19579) );
  OAI211_X1 U22597 ( .C1(n19581), .C2(n12655), .A(n19580), .B(n19579), .ZN(
        P2_U3143) );
  INV_X1 U22598 ( .A(n19582), .ZN(n19585) );
  INV_X1 U22599 ( .A(n19591), .ZN(n19584) );
  NAND3_X1 U22600 ( .A1(n19873), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19614) );
  NOR2_X1 U22601 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19614), .ZN(
        n19607) );
  OAI21_X1 U22602 ( .B1(n10989), .B2(n19607), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19583) );
  OAI21_X1 U22603 ( .B1(n19585), .B2(n19584), .A(n19583), .ZN(n19608) );
  AOI22_X1 U22604 ( .A1(n19608), .A2(n19702), .B1(n19701), .B2(n19607), .ZN(
        n19594) );
  AOI21_X1 U22605 ( .B1(n19586), .B2(n19646), .A(n19902), .ZN(n19592) );
  INV_X1 U22606 ( .A(n10989), .ZN(n19588) );
  INV_X1 U22607 ( .A(n19607), .ZN(n19587) );
  OAI211_X1 U22608 ( .C1(n19588), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19587), 
        .B(n15596), .ZN(n19589) );
  AND2_X1 U22609 ( .A1(n19589), .A2(n19707), .ZN(n19590) );
  OAI211_X1 U22610 ( .C1(n19592), .C2(n19591), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19590), .ZN(n19610) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19610), .B1(
        n19609), .B2(n19710), .ZN(n19593) );
  OAI211_X1 U22612 ( .C1(n19713), .C2(n19646), .A(n19594), .B(n19593), .ZN(
        P2_U3144) );
  AOI22_X1 U22613 ( .A1(n19608), .A2(n19715), .B1(n19714), .B2(n19607), .ZN(
        n19596) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19610), .B1(
        n19609), .B2(n19716), .ZN(n19595) );
  OAI211_X1 U22615 ( .C1(n19719), .C2(n19646), .A(n19596), .B(n19595), .ZN(
        P2_U3145) );
  AOI22_X1 U22616 ( .A1(n19608), .A2(n19721), .B1(n19720), .B2(n19607), .ZN(
        n19598) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19610), .B1(
        n19609), .B2(n19722), .ZN(n19597) );
  OAI211_X1 U22618 ( .C1(n19725), .C2(n19646), .A(n19598), .B(n19597), .ZN(
        P2_U3146) );
  AOI22_X1 U22619 ( .A1(n19608), .A2(n19727), .B1(n19726), .B2(n19607), .ZN(
        n19600) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19610), .B1(
        n19609), .B2(n19728), .ZN(n19599) );
  OAI211_X1 U22621 ( .C1(n19731), .C2(n19646), .A(n19600), .B(n19599), .ZN(
        P2_U3147) );
  AOI22_X1 U22622 ( .A1(n19608), .A2(n19733), .B1(n19732), .B2(n19607), .ZN(
        n19602) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19610), .B1(
        n19609), .B2(n19734), .ZN(n19601) );
  OAI211_X1 U22624 ( .C1(n19737), .C2(n19646), .A(n19602), .B(n19601), .ZN(
        P2_U3148) );
  AOI22_X1 U22625 ( .A1(n19608), .A2(n19739), .B1(n19738), .B2(n19607), .ZN(
        n19604) );
  AOI22_X1 U22626 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19610), .B1(
        n19609), .B2(n19740), .ZN(n19603) );
  OAI211_X1 U22627 ( .C1(n19743), .C2(n19646), .A(n19604), .B(n19603), .ZN(
        P2_U3149) );
  AOI22_X1 U22628 ( .A1(n19745), .A2(n19608), .B1(n19744), .B2(n19607), .ZN(
        n19606) );
  AOI22_X1 U22629 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19610), .B1(
        n19609), .B2(n19746), .ZN(n19605) );
  OAI211_X1 U22630 ( .C1(n19749), .C2(n19646), .A(n19606), .B(n19605), .ZN(
        P2_U3150) );
  AOI22_X1 U22631 ( .A1(n19608), .A2(n19752), .B1(n19750), .B2(n19607), .ZN(
        n19612) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19610), .B1(
        n19609), .B2(n19754), .ZN(n19611) );
  OAI211_X1 U22633 ( .C1(n19760), .C2(n19646), .A(n19612), .B(n19611), .ZN(
        P2_U3151) );
  NOR2_X1 U22634 ( .A1(n19883), .A2(n19614), .ZN(n19653) );
  OAI21_X1 U22635 ( .B1(n10996), .B2(n19653), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19613) );
  OAI21_X1 U22636 ( .B1(n19614), .B2(n15596), .A(n19613), .ZN(n19642) );
  AOI22_X1 U22637 ( .A1(n19642), .A2(n19702), .B1(n19701), .B2(n19653), .ZN(
        n19622) );
  OAI21_X1 U22638 ( .B1(n19706), .B2(n19619), .A(n19614), .ZN(n19618) );
  INV_X1 U22639 ( .A(n10996), .ZN(n19616) );
  INV_X1 U22640 ( .A(n19653), .ZN(n19615) );
  OAI211_X1 U22641 ( .C1(n19616), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19615), 
        .B(n15596), .ZN(n19617) );
  NAND3_X1 U22642 ( .A1(n19618), .A2(n19707), .A3(n19617), .ZN(n19643) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19643), .B1(
        n19691), .B2(n19662), .ZN(n19621) );
  OAI211_X1 U22644 ( .C1(n19623), .C2(n19646), .A(n19622), .B(n19621), .ZN(
        P2_U3152) );
  AOI22_X1 U22645 ( .A1(n19642), .A2(n19715), .B1(n19714), .B2(n19653), .ZN(
        n19625) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19643), .B1(
        n19691), .B2(n19666), .ZN(n19624) );
  OAI211_X1 U22647 ( .C1(n19626), .C2(n19646), .A(n19625), .B(n19624), .ZN(
        P2_U3153) );
  AOI22_X1 U22648 ( .A1(n19642), .A2(n19721), .B1(n19720), .B2(n19653), .ZN(
        n19628) );
  AOI22_X1 U22649 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19643), .B1(
        n19691), .B2(n19670), .ZN(n19627) );
  OAI211_X1 U22650 ( .C1(n19629), .C2(n19646), .A(n19628), .B(n19627), .ZN(
        P2_U3154) );
  AOI22_X1 U22651 ( .A1(n19642), .A2(n19727), .B1(n19726), .B2(n19653), .ZN(
        n19631) );
  AOI22_X1 U22652 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19643), .B1(
        n19691), .B2(n19674), .ZN(n19630) );
  OAI211_X1 U22653 ( .C1(n19632), .C2(n19646), .A(n19631), .B(n19630), .ZN(
        P2_U3155) );
  AOI22_X1 U22654 ( .A1(n19642), .A2(n19733), .B1(n19732), .B2(n19653), .ZN(
        n19634) );
  AOI22_X1 U22655 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19643), .B1(
        n19691), .B2(n19678), .ZN(n19633) );
  OAI211_X1 U22656 ( .C1(n19635), .C2(n19646), .A(n19634), .B(n19633), .ZN(
        P2_U3156) );
  AOI22_X1 U22657 ( .A1(n19642), .A2(n19739), .B1(n19738), .B2(n19653), .ZN(
        n19637) );
  AOI22_X1 U22658 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19643), .B1(
        n19691), .B2(n19682), .ZN(n19636) );
  OAI211_X1 U22659 ( .C1(n19638), .C2(n19646), .A(n19637), .B(n19636), .ZN(
        P2_U3157) );
  AOI22_X1 U22660 ( .A1(n19745), .A2(n19642), .B1(n19744), .B2(n19653), .ZN(
        n19640) );
  AOI22_X1 U22661 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19643), .B1(
        n19691), .B2(n19686), .ZN(n19639) );
  OAI211_X1 U22662 ( .C1(n19641), .C2(n19646), .A(n19640), .B(n19639), .ZN(
        P2_U3158) );
  AOI22_X1 U22663 ( .A1(n19642), .A2(n19752), .B1(n19750), .B2(n19653), .ZN(
        n19645) );
  AOI22_X1 U22664 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19643), .B1(
        n19691), .B2(n19692), .ZN(n19644) );
  OAI211_X1 U22665 ( .C1(n19647), .C2(n19646), .A(n19645), .B(n19644), .ZN(
        P2_U3159) );
  INV_X1 U22666 ( .A(n19691), .ZN(n19649) );
  NAND2_X1 U22667 ( .A1(n19649), .A2(n19648), .ZN(n19652) );
  OAI21_X1 U22668 ( .B1(n19652), .B2(n19755), .A(n19651), .ZN(n19656) );
  NAND3_X1 U22669 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19699), .A3(
        n19883), .ZN(n19657) );
  INV_X1 U22670 ( .A(n19657), .ZN(n19690) );
  OR2_X1 U22671 ( .A1(n19690), .A2(n19653), .ZN(n19660) );
  INV_X1 U22672 ( .A(n10995), .ZN(n19658) );
  AOI21_X1 U22673 ( .B1(n19658), .B2(n19657), .A(n19654), .ZN(n19655) );
  AOI22_X1 U22674 ( .A1(n19710), .A2(n19691), .B1(n19701), .B2(n19690), .ZN(
        n19664) );
  INV_X1 U22675 ( .A(n19656), .ZN(n19661) );
  OAI211_X1 U22676 ( .C1(n19658), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19657), 
        .B(n15596), .ZN(n19659) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19693), .B1(
        n19755), .B2(n19662), .ZN(n19663) );
  OAI211_X1 U22678 ( .C1(n19697), .C2(n19665), .A(n19664), .B(n19663), .ZN(
        P2_U3160) );
  AOI22_X1 U22679 ( .A1(n19666), .A2(n19755), .B1(n19714), .B2(n19690), .ZN(
        n19668) );
  AOI22_X1 U22680 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19693), .B1(
        n19691), .B2(n19716), .ZN(n19667) );
  OAI211_X1 U22681 ( .C1(n19697), .C2(n19669), .A(n19668), .B(n19667), .ZN(
        P2_U3161) );
  AOI22_X1 U22682 ( .A1(n19670), .A2(n19755), .B1(n19720), .B2(n19690), .ZN(
        n19672) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19693), .B1(
        n19691), .B2(n19722), .ZN(n19671) );
  OAI211_X1 U22684 ( .C1(n19697), .C2(n19673), .A(n19672), .B(n19671), .ZN(
        P2_U3162) );
  AOI22_X1 U22685 ( .A1(n19728), .A2(n19691), .B1(n19726), .B2(n19690), .ZN(
        n19676) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19693), .B1(
        n19755), .B2(n19674), .ZN(n19675) );
  OAI211_X1 U22687 ( .C1(n19697), .C2(n19677), .A(n19676), .B(n19675), .ZN(
        P2_U3163) );
  AOI22_X1 U22688 ( .A1(n19734), .A2(n19691), .B1(n19732), .B2(n19690), .ZN(
        n19680) );
  AOI22_X1 U22689 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19693), .B1(
        n19755), .B2(n19678), .ZN(n19679) );
  OAI211_X1 U22690 ( .C1(n19697), .C2(n19681), .A(n19680), .B(n19679), .ZN(
        P2_U3164) );
  AOI22_X1 U22691 ( .A1(n19682), .A2(n19755), .B1(n19738), .B2(n19690), .ZN(
        n19684) );
  AOI22_X1 U22692 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19693), .B1(
        n19691), .B2(n19740), .ZN(n19683) );
  OAI211_X1 U22693 ( .C1(n19697), .C2(n19685), .A(n19684), .B(n19683), .ZN(
        P2_U3165) );
  AOI22_X1 U22694 ( .A1(n19686), .A2(n19755), .B1(n19744), .B2(n19690), .ZN(
        n19688) );
  AOI22_X1 U22695 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19693), .B1(
        n19691), .B2(n19746), .ZN(n19687) );
  OAI211_X1 U22696 ( .C1(n19697), .C2(n19689), .A(n19688), .B(n19687), .ZN(
        P2_U3166) );
  AOI22_X1 U22697 ( .A1(n19754), .A2(n19691), .B1(n19750), .B2(n19690), .ZN(
        n19695) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19693), .B1(
        n19755), .B2(n19692), .ZN(n19694) );
  OAI211_X1 U22699 ( .C1(n19697), .C2(n19696), .A(n19695), .B(n19694), .ZN(
        P2_U3167) );
  NAND2_X1 U22700 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19699), .ZN(
        n19704) );
  OAI21_X1 U22701 ( .B1(n10987), .B2(n19751), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19700) );
  OAI21_X1 U22702 ( .B1(n19704), .B2(n15596), .A(n19700), .ZN(n19753) );
  AOI22_X1 U22703 ( .A1(n19753), .A2(n19702), .B1(n19751), .B2(n19701), .ZN(
        n19712) );
  INV_X1 U22704 ( .A(n10987), .ZN(n19703) );
  AOI21_X1 U22705 ( .B1(n19703), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19709) );
  OAI21_X1 U22706 ( .B1(n19706), .B2(n19705), .A(n19704), .ZN(n19708) );
  OAI211_X1 U22707 ( .C1(n19751), .C2(n19709), .A(n19708), .B(n19707), .ZN(
        n19756) );
  AOI22_X1 U22708 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19756), .B1(
        n19755), .B2(n19710), .ZN(n19711) );
  OAI211_X1 U22709 ( .C1(n19713), .C2(n19759), .A(n19712), .B(n19711), .ZN(
        P2_U3168) );
  AOI22_X1 U22710 ( .A1(n19753), .A2(n19715), .B1(n19751), .B2(n19714), .ZN(
        n19718) );
  AOI22_X1 U22711 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19756), .B1(
        n19755), .B2(n19716), .ZN(n19717) );
  OAI211_X1 U22712 ( .C1(n19719), .C2(n19759), .A(n19718), .B(n19717), .ZN(
        P2_U3169) );
  AOI22_X1 U22713 ( .A1(n19753), .A2(n19721), .B1(n19751), .B2(n19720), .ZN(
        n19724) );
  AOI22_X1 U22714 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19756), .B1(
        n19755), .B2(n19722), .ZN(n19723) );
  OAI211_X1 U22715 ( .C1(n19725), .C2(n19759), .A(n19724), .B(n19723), .ZN(
        P2_U3170) );
  AOI22_X1 U22716 ( .A1(n19753), .A2(n19727), .B1(n19751), .B2(n19726), .ZN(
        n19730) );
  AOI22_X1 U22717 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19756), .B1(
        n19755), .B2(n19728), .ZN(n19729) );
  OAI211_X1 U22718 ( .C1(n19731), .C2(n19759), .A(n19730), .B(n19729), .ZN(
        P2_U3171) );
  AOI22_X1 U22719 ( .A1(n19753), .A2(n19733), .B1(n19751), .B2(n19732), .ZN(
        n19736) );
  AOI22_X1 U22720 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19756), .B1(
        n19755), .B2(n19734), .ZN(n19735) );
  OAI211_X1 U22721 ( .C1(n19737), .C2(n19759), .A(n19736), .B(n19735), .ZN(
        P2_U3172) );
  AOI22_X1 U22722 ( .A1(n19753), .A2(n19739), .B1(n19751), .B2(n19738), .ZN(
        n19742) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19756), .B1(
        n19755), .B2(n19740), .ZN(n19741) );
  OAI211_X1 U22724 ( .C1(n19743), .C2(n19759), .A(n19742), .B(n19741), .ZN(
        P2_U3173) );
  AOI22_X1 U22725 ( .A1(n19745), .A2(n19753), .B1(n19751), .B2(n19744), .ZN(
        n19748) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19756), .B1(
        n19755), .B2(n19746), .ZN(n19747) );
  OAI211_X1 U22727 ( .C1(n19749), .C2(n19759), .A(n19748), .B(n19747), .ZN(
        P2_U3174) );
  AOI22_X1 U22728 ( .A1(n19753), .A2(n19752), .B1(n19751), .B2(n19750), .ZN(
        n19758) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19756), .B1(
        n19755), .B2(n19754), .ZN(n19757) );
  OAI211_X1 U22730 ( .C1(n19760), .C2(n19759), .A(n19758), .B(n19757), .ZN(
        P2_U3175) );
  AOI221_X1 U22731 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19654), .C1(n19899), 
        .C2(n19654), .A(n19761), .ZN(n19765) );
  AOI211_X1 U22732 ( .C1(n19762), .C2(n19766), .A(n19901), .B(n11393), .ZN(
        n19763) );
  AOI211_X1 U22733 ( .C1(n19766), .C2(n19765), .A(n19764), .B(n19763), .ZN(
        n19767) );
  INV_X1 U22734 ( .A(n19767), .ZN(P2_U3177) );
  AND2_X1 U22735 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19768), .ZN(
        P2_U3179) );
  AND2_X1 U22736 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19768), .ZN(
        P2_U3180) );
  AND2_X1 U22737 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19768), .ZN(
        P2_U3181) );
  AND2_X1 U22738 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19768), .ZN(
        P2_U3182) );
  AND2_X1 U22739 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19768), .ZN(
        P2_U3183) );
  AND2_X1 U22740 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19768), .ZN(
        P2_U3184) );
  AND2_X1 U22741 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19768), .ZN(
        P2_U3185) );
  AND2_X1 U22742 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19768), .ZN(
        P2_U3186) );
  AND2_X1 U22743 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19768), .ZN(
        P2_U3187) );
  NOR2_X1 U22744 ( .A1(n20971), .A2(n19845), .ZN(P2_U3188) );
  AND2_X1 U22745 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19768), .ZN(
        P2_U3189) );
  AND2_X1 U22746 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19768), .ZN(
        P2_U3190) );
  AND2_X1 U22747 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19768), .ZN(
        P2_U3191) );
  NOR2_X1 U22748 ( .A1(n20950), .A2(n19845), .ZN(P2_U3192) );
  AND2_X1 U22749 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19768), .ZN(
        P2_U3193) );
  AND2_X1 U22750 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19768), .ZN(
        P2_U3194) );
  AND2_X1 U22751 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19768), .ZN(
        P2_U3195) );
  AND2_X1 U22752 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19768), .ZN(
        P2_U3196) );
  AND2_X1 U22753 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19768), .ZN(
        P2_U3197) );
  AND2_X1 U22754 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19768), .ZN(
        P2_U3198) );
  AND2_X1 U22755 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19768), .ZN(
        P2_U3199) );
  AND2_X1 U22756 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19768), .ZN(
        P2_U3200) );
  AND2_X1 U22757 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19768), .ZN(P2_U3201) );
  AND2_X1 U22758 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19768), .ZN(P2_U3202) );
  AND2_X1 U22759 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19768), .ZN(P2_U3203) );
  AND2_X1 U22760 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19768), .ZN(P2_U3204) );
  AND2_X1 U22761 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19768), .ZN(P2_U3205) );
  AND2_X1 U22762 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19768), .ZN(P2_U3206) );
  AND2_X1 U22763 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19768), .ZN(P2_U3207) );
  AND2_X1 U22764 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19768), .ZN(P2_U3208) );
  NOR2_X1 U22765 ( .A1(n19901), .A2(n19779), .ZN(n19777) );
  INV_X1 U22766 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19910) );
  OR3_X1 U22767 ( .A1(n19777), .A2(n19910), .A3(n19769), .ZN(n19771) );
  AOI211_X1 U22768 ( .C1(n20740), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19778), .B(n19840), .ZN(n19770) );
  INV_X1 U22769 ( .A(NA), .ZN(n20733) );
  NOR2_X1 U22770 ( .A1(n20733), .A2(n19773), .ZN(n19783) );
  AOI211_X1 U22771 ( .C1(n19786), .C2(n19771), .A(n19770), .B(n19783), .ZN(
        n19772) );
  INV_X1 U22772 ( .A(n19772), .ZN(P2_U3209) );
  AOI21_X1 U22773 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20740), .A(n19786), 
        .ZN(n19780) );
  NOR2_X1 U22774 ( .A1(n19780), .A2(n19910), .ZN(n19774) );
  AOI211_X1 U22775 ( .C1(n19774), .C2(n19773), .A(n19906), .B(n19777), .ZN(
        n19775) );
  OAI21_X1 U22776 ( .B1(n20740), .B2(n19776), .A(n19775), .ZN(P2_U3210) );
  AOI22_X1 U22777 ( .A1(n19778), .A2(n19910), .B1(n19777), .B2(n20733), .ZN(
        n19785) );
  OAI21_X1 U22778 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19784) );
  NOR2_X1 U22779 ( .A1(n19779), .A2(n19786), .ZN(n19781) );
  AOI21_X1 U22780 ( .B1(n19781), .B2(n19899), .A(n19780), .ZN(n19782) );
  OAI22_X1 U22781 ( .A1(n19785), .A2(n19784), .B1(n19783), .B2(n19782), .ZN(
        P2_U3211) );
  OAI222_X1 U22782 ( .A1(n19832), .A2(n10808), .B1(n19787), .B2(n19912), .C1(
        n10793), .C2(n19833), .ZN(P2_U3212) );
  OAI222_X1 U22783 ( .A1(n19832), .A2(n19789), .B1(n19788), .B2(n19912), .C1(
        n10808), .C2(n19833), .ZN(P2_U3213) );
  OAI222_X1 U22784 ( .A1(n19832), .A2(n11303), .B1(n19790), .B2(n19912), .C1(
        n19789), .C2(n19833), .ZN(P2_U3214) );
  OAI222_X1 U22785 ( .A1(n19832), .A2(n11308), .B1(n19791), .B2(n19912), .C1(
        n11303), .C2(n19833), .ZN(P2_U3215) );
  OAI222_X1 U22786 ( .A1(n19832), .A2(n11312), .B1(n19792), .B2(n19912), .C1(
        n11308), .C2(n19833), .ZN(P2_U3216) );
  OAI222_X1 U22787 ( .A1(n19832), .A2(n19794), .B1(n19793), .B2(n19912), .C1(
        n11312), .C2(n19833), .ZN(P2_U3217) );
  OAI222_X1 U22788 ( .A1(n19832), .A2(n11491), .B1(n19795), .B2(n19840), .C1(
        n19794), .C2(n19833), .ZN(P2_U3218) );
  OAI222_X1 U22789 ( .A1(n19832), .A2(n11324), .B1(n19796), .B2(n19840), .C1(
        n11491), .C2(n19833), .ZN(P2_U3219) );
  OAI222_X1 U22790 ( .A1(n19832), .A2(n19798), .B1(n19797), .B2(n19840), .C1(
        n11324), .C2(n19833), .ZN(P2_U3220) );
  OAI222_X1 U22791 ( .A1(n19832), .A2(n19800), .B1(n19799), .B2(n19840), .C1(
        n19798), .C2(n19833), .ZN(P2_U3221) );
  OAI222_X1 U22792 ( .A1(n19832), .A2(n11333), .B1(n19801), .B2(n19840), .C1(
        n19800), .C2(n19833), .ZN(P2_U3222) );
  OAI222_X1 U22793 ( .A1(n19832), .A2(n11337), .B1(n19802), .B2(n19840), .C1(
        n11333), .C2(n19833), .ZN(P2_U3223) );
  OAI222_X1 U22794 ( .A1(n19832), .A2(n11341), .B1(n19803), .B2(n19840), .C1(
        n11337), .C2(n19833), .ZN(P2_U3224) );
  OAI222_X1 U22795 ( .A1(n19832), .A2(n19805), .B1(n19804), .B2(n19840), .C1(
        n11341), .C2(n19833), .ZN(P2_U3225) );
  OAI222_X1 U22796 ( .A1(n19832), .A2(n15451), .B1(n19806), .B2(n19840), .C1(
        n19805), .C2(n19833), .ZN(P2_U3226) );
  OAI222_X1 U22797 ( .A1(n19832), .A2(n19808), .B1(n19807), .B2(n19840), .C1(
        n15451), .C2(n19833), .ZN(P2_U3227) );
  INV_X1 U22798 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19809) );
  OAI222_X1 U22799 ( .A1(n19832), .A2(n19809), .B1(n21075), .B2(n19840), .C1(
        n19808), .C2(n19833), .ZN(P2_U3228) );
  OAI222_X1 U22800 ( .A1(n19832), .A2(n19811), .B1(n19810), .B2(n19840), .C1(
        n19809), .C2(n19833), .ZN(P2_U3229) );
  OAI222_X1 U22801 ( .A1(n19832), .A2(n15201), .B1(n19812), .B2(n19912), .C1(
        n19811), .C2(n19833), .ZN(P2_U3230) );
  OAI222_X1 U22802 ( .A1(n19832), .A2(n19814), .B1(n19813), .B2(n19912), .C1(
        n15201), .C2(n19833), .ZN(P2_U3231) );
  INV_X1 U22803 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19816) );
  OAI222_X1 U22804 ( .A1(n19832), .A2(n19816), .B1(n19815), .B2(n19912), .C1(
        n19814), .C2(n19833), .ZN(P2_U3232) );
  OAI222_X1 U22805 ( .A1(n19832), .A2(n19818), .B1(n19817), .B2(n19912), .C1(
        n19816), .C2(n19833), .ZN(P2_U3233) );
  OAI222_X1 U22806 ( .A1(n19832), .A2(n19820), .B1(n19819), .B2(n19912), .C1(
        n19818), .C2(n19833), .ZN(P2_U3234) );
  OAI222_X1 U22807 ( .A1(n19832), .A2(n19822), .B1(n19821), .B2(n19912), .C1(
        n19820), .C2(n19833), .ZN(P2_U3235) );
  INV_X1 U22808 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19824) );
  OAI222_X1 U22809 ( .A1(n19832), .A2(n19824), .B1(n19823), .B2(n19912), .C1(
        n19822), .C2(n19833), .ZN(P2_U3236) );
  OAI222_X1 U22810 ( .A1(n19832), .A2(n19827), .B1(n19825), .B2(n19912), .C1(
        n19824), .C2(n19833), .ZN(P2_U3237) );
  OAI222_X1 U22811 ( .A1(n19833), .A2(n19827), .B1(n19826), .B2(n19912), .C1(
        n19828), .C2(n19832), .ZN(P2_U3238) );
  INV_X1 U22812 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19830) );
  OAI222_X1 U22813 ( .A1(n19832), .A2(n19830), .B1(n19829), .B2(n19912), .C1(
        n19828), .C2(n19833), .ZN(P2_U3239) );
  INV_X1 U22814 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19834) );
  OAI222_X1 U22815 ( .A1(n19832), .A2(n19834), .B1(n19831), .B2(n19912), .C1(
        n19830), .C2(n19833), .ZN(P2_U3240) );
  OAI222_X1 U22816 ( .A1(n19832), .A2(n19836), .B1(n19835), .B2(n19912), .C1(
        n19834), .C2(n19833), .ZN(P2_U3241) );
  OAI22_X1 U22817 ( .A1(n19913), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19912), .ZN(n19837) );
  INV_X1 U22818 ( .A(n19837), .ZN(P2_U3585) );
  OAI22_X1 U22819 ( .A1(n19913), .A2(P2_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P2_BE_N_REG_2__SCAN_IN), .B2(n19912), .ZN(n19838) );
  INV_X1 U22820 ( .A(n19838), .ZN(P2_U3586) );
  OAI22_X1 U22821 ( .A1(n19913), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19912), .ZN(n19839) );
  INV_X1 U22822 ( .A(n19839), .ZN(P2_U3587) );
  OAI22_X1 U22823 ( .A1(n19913), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19840), .ZN(n19841) );
  INV_X1 U22824 ( .A(n19841), .ZN(P2_U3588) );
  OAI21_X1 U22825 ( .B1(n19845), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19843), 
        .ZN(n19842) );
  INV_X1 U22826 ( .A(n19842), .ZN(P2_U3591) );
  OAI21_X1 U22827 ( .B1(n19845), .B2(n19844), .A(n19843), .ZN(P2_U3592) );
  INV_X1 U22828 ( .A(n19882), .ZN(n19881) );
  INV_X1 U22829 ( .A(n19846), .ZN(n19853) );
  OR2_X1 U22830 ( .A1(n19847), .A2(n19865), .ZN(n19859) );
  NAND2_X1 U22831 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATEBS16_REG_SCAN_IN), .ZN(n19848) );
  OR2_X1 U22832 ( .A1(n19868), .A2(n19848), .ZN(n19849) );
  NAND2_X1 U22833 ( .A1(n19849), .A2(n19874), .ZN(n19869) );
  NAND2_X1 U22834 ( .A1(n19859), .A2(n19869), .ZN(n19852) );
  INV_X1 U22835 ( .A(n19850), .ZN(n19851) );
  AOI22_X1 U22836 ( .A1(n19853), .A2(n19852), .B1(n19851), .B2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19854) );
  OAI21_X1 U22837 ( .B1(n19855), .B2(n15596), .A(n19854), .ZN(n19856) );
  INV_X1 U22838 ( .A(n19856), .ZN(n19857) );
  AOI22_X1 U22839 ( .A1(n19881), .A2(n19858), .B1(n19857), .B2(n19882), .ZN(
        P2_U3602) );
  OAI21_X1 U22840 ( .B1(n19860), .B2(n19869), .A(n19859), .ZN(n19861) );
  AOI21_X1 U22841 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19862), .A(n19861), 
        .ZN(n19863) );
  AOI22_X1 U22842 ( .A1(n19881), .A2(n19864), .B1(n19863), .B2(n19882), .ZN(
        P2_U3603) );
  INV_X1 U22843 ( .A(n19865), .ZN(n19866) );
  NAND2_X1 U22844 ( .A1(n19868), .A2(n19866), .ZN(n19867) );
  OAI21_X1 U22845 ( .B1(n19869), .B2(n19868), .A(n19867), .ZN(n19870) );
  AOI21_X1 U22846 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19871), .A(n19870), 
        .ZN(n19872) );
  AOI22_X1 U22847 ( .A1(n19881), .A2(n19873), .B1(n19872), .B2(n19882), .ZN(
        P2_U3604) );
  INV_X1 U22848 ( .A(n19874), .ZN(n19877) );
  NAND3_X1 U22849 ( .A1(n19875), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19876) );
  OAI21_X1 U22850 ( .B1(n19878), .B2(n19877), .A(n19876), .ZN(n19879) );
  AOI21_X1 U22851 ( .B1(n19883), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19879), 
        .ZN(n19880) );
  OAI22_X1 U22852 ( .A1(n19883), .A2(n19882), .B1(n19881), .B2(n19880), .ZN(
        P2_U3605) );
  INV_X1 U22853 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19884) );
  AOI22_X1 U22854 ( .A1(n19912), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19884), 
        .B2(n19913), .ZN(P2_U3608) );
  INV_X1 U22855 ( .A(n19885), .ZN(n19886) );
  NAND2_X1 U22856 ( .A1(n19887), .A2(n19886), .ZN(n19888) );
  OAI211_X1 U22857 ( .C1(n19891), .C2(n19890), .A(n19889), .B(n19888), .ZN(
        n19893) );
  MUX2_X1 U22858 ( .A(P2_MORE_REG_SCAN_IN), .B(n19893), .S(n19892), .Z(
        P2_U3609) );
  OAI21_X1 U22859 ( .B1(n19894), .B2(n19654), .A(n19469), .ZN(n19897) );
  INV_X1 U22860 ( .A(n19895), .ZN(n19896) );
  OAI211_X1 U22861 ( .C1(n19899), .C2(n19898), .A(n19897), .B(n19896), .ZN(
        n19911) );
  AOI22_X1 U22862 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19901), .B1(n19904), 
        .B2(n19900), .ZN(n19908) );
  NAND2_X1 U22863 ( .A1(n19903), .A2(n19902), .ZN(n19905) );
  AOI211_X1 U22864 ( .C1(n19906), .C2(n19905), .A(n19904), .B(n11731), .ZN(
        n19907) );
  OAI21_X1 U22865 ( .B1(n19908), .B2(n19907), .A(n19911), .ZN(n19909) );
  OAI21_X1 U22866 ( .B1(n19911), .B2(n19910), .A(n19909), .ZN(P2_U3610) );
  OAI22_X1 U22867 ( .A1(n19913), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19912), .ZN(n19914) );
  INV_X1 U22868 ( .A(n19914), .ZN(P2_U3611) );
  AOI21_X1 U22869 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n11841), .A(n20735), 
        .ZN(n20738) );
  INV_X1 U22870 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19915) );
  NAND2_X1 U22871 ( .A1(n20735), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20832) );
  INV_X2 U22872 ( .A(n20832), .ZN(n20795) );
  AOI21_X1 U22873 ( .B1(n20738), .B2(n19915), .A(n20795), .ZN(P1_U2802) );
  NAND2_X1 U22874 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20551), .ZN(n19919) );
  OAI21_X1 U22875 ( .B1(n19917), .B2(n19916), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19918) );
  OAI21_X1 U22876 ( .B1(n19919), .B2(n20823), .A(n19918), .ZN(P1_U2803) );
  NOR2_X1 U22877 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19921) );
  OAI21_X1 U22878 ( .B1(n19921), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20832), .ZN(
        n19920) );
  OAI21_X1 U22879 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20832), .A(n19920), 
        .ZN(P1_U2804) );
  NOR2_X1 U22880 ( .A1(n20795), .A2(n20738), .ZN(n20803) );
  OAI21_X1 U22881 ( .B1(BS16), .B2(n19921), .A(n20803), .ZN(n20801) );
  OAI21_X1 U22882 ( .B1(n20803), .B2(n20622), .A(n20801), .ZN(P1_U2805) );
  OAI21_X1 U22883 ( .B1(n19924), .B2(n19923), .A(n19922), .ZN(P1_U2806) );
  NOR4_X1 U22884 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19928) );
  NOR4_X1 U22885 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19927) );
  NOR4_X1 U22886 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19926) );
  NOR4_X1 U22887 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19925) );
  NAND4_X1 U22888 ( .A1(n19928), .A2(n19927), .A3(n19926), .A4(n19925), .ZN(
        n19934) );
  NOR4_X1 U22889 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19932) );
  AOI211_X1 U22890 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_4__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19931) );
  NOR4_X1 U22891 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19930) );
  NOR4_X1 U22892 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19929) );
  NAND4_X1 U22893 ( .A1(n19932), .A2(n19931), .A3(n19930), .A4(n19929), .ZN(
        n19933) );
  NOR2_X1 U22894 ( .A1(n19934), .A2(n19933), .ZN(n20815) );
  INV_X1 U22895 ( .A(n20815), .ZN(n19937) );
  NAND2_X1 U22896 ( .A1(n20815), .A2(n21140), .ZN(n20816) );
  NOR3_X1 U22897 ( .A1(P1_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A3(n20816), .ZN(n19936) );
  AOI21_X1 U22898 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(n19937), .A(n19936), 
        .ZN(n19935) );
  OAI21_X1 U22899 ( .B1(n13222), .B2(n19937), .A(n19935), .ZN(P1_U2807) );
  NAND2_X1 U22900 ( .A1(n20815), .A2(n13222), .ZN(n20811) );
  AOI21_X1 U22901 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(n19937), .A(n19936), 
        .ZN(n19938) );
  OAI21_X1 U22902 ( .B1(P1_DATAWIDTH_REG_1__SCAN_IN), .B2(n20811), .A(n19938), 
        .ZN(P1_U2808) );
  NOR3_X1 U22903 ( .A1(n19940), .A2(n20982), .A3(n19939), .ZN(n19944) );
  AOI22_X1 U22904 ( .A1(n20013), .A2(n19988), .B1(n19996), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n19941) );
  OAI211_X1 U22905 ( .C1(n19986), .C2(n19942), .A(n19941), .B(n20135), .ZN(
        n19943) );
  AOI221_X1 U22906 ( .B1(n19945), .B2(P1_REIP_REG_9__SCAN_IN), .C1(n19944), 
        .C2(n20755), .A(n19943), .ZN(n19950) );
  OAI22_X1 U22907 ( .A1(n20016), .A2(n19947), .B1(n20002), .B2(n19946), .ZN(
        n19948) );
  INV_X1 U22908 ( .A(n19948), .ZN(n19949) );
  NAND2_X1 U22909 ( .A1(n19950), .A2(n19949), .ZN(P1_U2831) );
  INV_X1 U22910 ( .A(n20000), .ZN(n19980) );
  NOR3_X1 U22911 ( .A1(n20747), .A2(n19981), .A3(n19980), .ZN(n19975) );
  NAND3_X1 U22912 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n19975), .ZN(n19957) );
  INV_X1 U22913 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20752) );
  NAND2_X1 U22914 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19953) );
  NAND2_X1 U22915 ( .A1(n19952), .A2(n19951), .ZN(n19971) );
  OAI21_X1 U22916 ( .B1(n19953), .B2(n19971), .A(n19972), .ZN(n19962) );
  AOI22_X1 U22917 ( .A1(n19998), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19996), .B2(P1_EBX_REG_7__SCAN_IN), .ZN(n19954) );
  INV_X1 U22918 ( .A(n19954), .ZN(n19955) );
  AOI211_X1 U22919 ( .C1(n19988), .C2(n10345), .A(n12122), .B(n19955), .ZN(
        n19956) );
  OAI221_X1 U22920 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n19957), .C1(n20752), 
        .C2(n19962), .A(n19956), .ZN(n19958) );
  AOI21_X1 U22921 ( .B1(n20020), .B2(n19965), .A(n19958), .ZN(n19959) );
  OAI21_X1 U22922 ( .B1(n19960), .B2(n20002), .A(n19959), .ZN(P1_U2833) );
  INV_X1 U22923 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20751) );
  AOI22_X1 U22924 ( .A1(n19998), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n19996), .B2(P1_EBX_REG_6__SCAN_IN), .ZN(n19961) );
  OAI21_X1 U22925 ( .B1(n20751), .B2(n19962), .A(n19961), .ZN(n19963) );
  AOI211_X1 U22926 ( .C1(n19988), .C2(n19964), .A(n12122), .B(n19963), .ZN(
        n19969) );
  INV_X1 U22927 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20749) );
  NOR2_X1 U22928 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20749), .ZN(n19967) );
  AOI22_X1 U22929 ( .A1(n19975), .A2(n19967), .B1(n19966), .B2(n19965), .ZN(
        n19968) );
  OAI211_X1 U22930 ( .C1(n19970), .C2(n20002), .A(n19969), .B(n19968), .ZN(
        P1_U2834) );
  NAND2_X1 U22931 ( .A1(n19972), .A2(n19971), .ZN(n19979) );
  AOI22_X1 U22932 ( .A1(n19998), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19996), .B2(P1_EBX_REG_5__SCAN_IN), .ZN(n19973) );
  OAI21_X1 U22933 ( .B1(n20749), .B2(n19979), .A(n19973), .ZN(n19974) );
  AOI211_X1 U22934 ( .C1(n19988), .C2(n20023), .A(n12122), .B(n19974), .ZN(
        n19977) );
  AOI22_X1 U22935 ( .A1(n19975), .A2(n20749), .B1(n20026), .B2(n19982), .ZN(
        n19976) );
  OAI211_X1 U22936 ( .C1(n19978), .C2(n20002), .A(n19977), .B(n19976), .ZN(
        P1_U2835) );
  AOI221_X1 U22937 ( .B1(n19981), .B2(n20747), .C1(n19980), .C2(n20747), .A(
        n19979), .ZN(n19994) );
  AND2_X1 U22938 ( .A1(n20095), .A2(n19982), .ZN(n19993) );
  INV_X1 U22939 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n21034) );
  OR2_X1 U22940 ( .A1(n19984), .A2(n19983), .ZN(n19985) );
  OAI211_X1 U22941 ( .C1(n19986), .C2(n21034), .A(n20135), .B(n19985), .ZN(
        n19987) );
  AOI21_X1 U22942 ( .B1(n19988), .B2(n20105), .A(n19987), .ZN(n19989) );
  OAI21_X1 U22943 ( .B1(n19991), .B2(n19990), .A(n19989), .ZN(n19992) );
  NOR3_X1 U22944 ( .A1(n19994), .A2(n19993), .A3(n19992), .ZN(n19995) );
  OAI21_X1 U22945 ( .B1(n20100), .B2(n20002), .A(n19995), .ZN(P1_U2836) );
  AOI22_X1 U22946 ( .A1(n19997), .A2(P1_REIP_REG_2__SCAN_IN), .B1(n19996), 
        .B2(P1_EBX_REG_2__SCAN_IN), .ZN(n20010) );
  INV_X1 U22947 ( .A(n13091), .ZN(n20155) );
  AOI22_X1 U22948 ( .A1(n20000), .A2(n19999), .B1(n19998), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20001) );
  OAI21_X1 U22949 ( .B1(n20003), .B2(n20002), .A(n20001), .ZN(n20007) );
  NOR2_X1 U22950 ( .A1(n20005), .A2(n20004), .ZN(n20006) );
  AOI211_X1 U22951 ( .C1(n20008), .C2(n20155), .A(n20007), .B(n20006), .ZN(
        n20009) );
  OAI211_X1 U22952 ( .C1(n20012), .C2(n20011), .A(n20010), .B(n20009), .ZN(
        P1_U2838) );
  INV_X1 U22953 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20019) );
  INV_X1 U22954 ( .A(n20013), .ZN(n20014) );
  OAI22_X1 U22955 ( .A1(n20016), .A2(n14529), .B1(n20015), .B2(n20014), .ZN(
        n20017) );
  INV_X1 U22956 ( .A(n20017), .ZN(n20018) );
  OAI21_X1 U22957 ( .B1(n20029), .B2(n20019), .A(n20018), .ZN(P1_U2863) );
  INV_X1 U22958 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20022) );
  AOI22_X1 U22959 ( .A1(n20020), .A2(n20025), .B1(n20024), .B2(n10345), .ZN(
        n20021) );
  OAI21_X1 U22960 ( .B1(n20029), .B2(n20022), .A(n20021), .ZN(P1_U2865) );
  INV_X1 U22961 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20028) );
  AOI22_X1 U22962 ( .A1(n20026), .A2(n20025), .B1(n20024), .B2(n20023), .ZN(
        n20027) );
  OAI21_X1 U22963 ( .B1(n20029), .B2(n20028), .A(n20027), .ZN(P1_U2867) );
  INV_X1 U22964 ( .A(n20030), .ZN(n20031) );
  AOI22_X1 U22965 ( .A1(n20031), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20056), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n20032) );
  OAI21_X1 U22966 ( .B1(n21113), .B2(n20046), .A(n20032), .ZN(P1_U2911) );
  INV_X1 U22967 ( .A(n20046), .ZN(n20829) );
  AOI22_X1 U22968 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20829), .B1(n20056), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20033) );
  OAI21_X1 U22969 ( .B1(n13384), .B2(n20058), .A(n20033), .ZN(P1_U2921) );
  AOI22_X1 U22970 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20034) );
  OAI21_X1 U22971 ( .B1(n13911), .B2(n20058), .A(n20034), .ZN(P1_U2922) );
  AOI22_X1 U22972 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20829), .B1(n20056), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20035) );
  OAI21_X1 U22973 ( .B1(n14601), .B2(n20058), .A(n20035), .ZN(P1_U2923) );
  AOI22_X1 U22974 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20036) );
  OAI21_X1 U22975 ( .B1(n13922), .B2(n20058), .A(n20036), .ZN(P1_U2924) );
  AOI22_X1 U22976 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20829), .B1(n20056), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20037) );
  OAI21_X1 U22977 ( .B1(n13823), .B2(n20058), .A(n20037), .ZN(P1_U2925) );
  AOI22_X1 U22978 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20038) );
  OAI21_X1 U22979 ( .B1(n13797), .B2(n20058), .A(n20038), .ZN(P1_U2926) );
  INV_X1 U22980 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20040) );
  AOI22_X1 U22981 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20829), .B1(n20056), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20039) );
  OAI21_X1 U22982 ( .B1(n20040), .B2(n20058), .A(n20039), .ZN(P1_U2927) );
  AOI22_X1 U22983 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20041) );
  OAI21_X1 U22984 ( .B1(n20999), .B2(n20058), .A(n20041), .ZN(P1_U2928) );
  AOI22_X1 U22985 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20829), .B1(n20056), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20042) );
  OAI21_X1 U22986 ( .B1(n13658), .B2(n20058), .A(n20042), .ZN(P1_U2929) );
  INV_X1 U22987 ( .A(P1_LWORD_REG_6__SCAN_IN), .ZN(n21085) );
  INV_X1 U22988 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n20043) );
  OAI222_X1 U22989 ( .A1(n20046), .A2(n21085), .B1(n20058), .B2(n13640), .C1(
        n20045), .C2(n20043), .ZN(P1_U2930) );
  INV_X1 U22990 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n21053) );
  OAI222_X1 U22991 ( .A1(n20046), .A2(n21053), .B1(n20058), .B2(n13517), .C1(
        n20045), .C2(n20044), .ZN(P1_U2931) );
  AOI22_X1 U22992 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20047) );
  OAI21_X1 U22993 ( .B1(n20048), .B2(n20058), .A(n20047), .ZN(P1_U2932) );
  AOI22_X1 U22994 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20829), .B1(n20056), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20049) );
  OAI21_X1 U22995 ( .B1(n20050), .B2(n20058), .A(n20049), .ZN(P1_U2933) );
  AOI22_X1 U22996 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20051), .B1(n20056), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20052) );
  OAI21_X1 U22997 ( .B1(n20053), .B2(n20058), .A(n20052), .ZN(P1_U2934) );
  AOI22_X1 U22998 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20829), .B1(n20056), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20054) );
  OAI21_X1 U22999 ( .B1(n20055), .B2(n20058), .A(n20054), .ZN(P1_U2935) );
  AOI22_X1 U23000 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20829), .B1(n20056), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20057) );
  OAI21_X1 U23001 ( .B1(n20059), .B2(n20058), .A(n20057), .ZN(P1_U2936) );
  AOI22_X1 U23002 ( .A1(n20087), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20086), .ZN(n20062) );
  INV_X1 U23003 ( .A(n20060), .ZN(n20061) );
  NAND2_X1 U23004 ( .A1(n20074), .A2(n20061), .ZN(n20078) );
  NAND2_X1 U23005 ( .A1(n20062), .A2(n20078), .ZN(P1_U2947) );
  AOI22_X1 U23006 ( .A1(n20087), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20086), .ZN(n20065) );
  INV_X1 U23007 ( .A(n20063), .ZN(n20064) );
  NAND2_X1 U23008 ( .A1(n20074), .A2(n20064), .ZN(n20080) );
  NAND2_X1 U23009 ( .A1(n20065), .A2(n20080), .ZN(P1_U2948) );
  AOI22_X1 U23010 ( .A1(n20087), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20086), .ZN(n20068) );
  INV_X1 U23011 ( .A(n20066), .ZN(n20067) );
  NAND2_X1 U23012 ( .A1(n20074), .A2(n20067), .ZN(n20082) );
  NAND2_X1 U23013 ( .A1(n20068), .A2(n20082), .ZN(P1_U2949) );
  AOI22_X1 U23014 ( .A1(n20087), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20086), .ZN(n20071) );
  INV_X1 U23015 ( .A(n20069), .ZN(n20070) );
  NAND2_X1 U23016 ( .A1(n20074), .A2(n20070), .ZN(n20084) );
  NAND2_X1 U23017 ( .A1(n20071), .A2(n20084), .ZN(P1_U2950) );
  AOI22_X1 U23018 ( .A1(n20087), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20086), .ZN(n20075) );
  INV_X1 U23019 ( .A(n20072), .ZN(n20073) );
  NAND2_X1 U23020 ( .A1(n20074), .A2(n20073), .ZN(n20088) );
  NAND2_X1 U23021 ( .A1(n20075), .A2(n20088), .ZN(P1_U2951) );
  AOI22_X1 U23022 ( .A1(n20087), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20086), .ZN(n20077) );
  NAND2_X1 U23023 ( .A1(n20077), .A2(n20076), .ZN(P1_U2961) );
  AOI22_X1 U23024 ( .A1(n20087), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20086), .ZN(n20079) );
  NAND2_X1 U23025 ( .A1(n20079), .A2(n20078), .ZN(P1_U2962) );
  AOI22_X1 U23026 ( .A1(n20087), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20086), .ZN(n20081) );
  NAND2_X1 U23027 ( .A1(n20081), .A2(n20080), .ZN(P1_U2963) );
  AOI22_X1 U23028 ( .A1(n20087), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20086), .ZN(n20083) );
  NAND2_X1 U23029 ( .A1(n20083), .A2(n20082), .ZN(P1_U2964) );
  AOI22_X1 U23030 ( .A1(n20087), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20086), .ZN(n20085) );
  NAND2_X1 U23031 ( .A1(n20085), .A2(n20084), .ZN(P1_U2965) );
  AOI22_X1 U23032 ( .A1(n20087), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20086), .ZN(n20089) );
  NAND2_X1 U23033 ( .A1(n20089), .A2(n20088), .ZN(P1_U2966) );
  AOI22_X1 U23034 ( .A1(n20090), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n12122), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20099) );
  OAI21_X1 U23035 ( .B1(n20093), .B2(n20092), .A(n20091), .ZN(n20094) );
  INV_X1 U23036 ( .A(n20094), .ZN(n20104) );
  AOI22_X1 U23037 ( .A1(n20104), .A2(n20097), .B1(n20096), .B2(n20095), .ZN(
        n20098) );
  OAI211_X1 U23038 ( .C1(n20101), .C2(n20100), .A(n20099), .B(n20098), .ZN(
        P1_U2995) );
  OAI21_X1 U23039 ( .B1(n20132), .B2(n20127), .A(n20102), .ZN(n20103) );
  INV_X1 U23040 ( .A(n20103), .ZN(n20119) );
  AOI222_X1 U23041 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n12122), .B1(n20126), 
        .B2(n20105), .C1(n20123), .C2(n20104), .ZN(n20108) );
  OAI211_X1 U23042 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20115), .B(n20106), .ZN(n20107) );
  OAI211_X1 U23043 ( .C1(n20119), .C2(n20109), .A(n20108), .B(n20107), .ZN(
        P1_U3027) );
  INV_X1 U23044 ( .A(n20110), .ZN(n20111) );
  AOI22_X1 U23045 ( .A1(n12122), .A2(P1_REIP_REG_3__SCAN_IN), .B1(n20126), 
        .B2(n20111), .ZN(n20117) );
  INV_X1 U23046 ( .A(n20113), .ZN(n20114) );
  AOI22_X1 U23047 ( .A1(n20115), .A2(n20118), .B1(n20114), .B2(n20123), .ZN(
        n20116) );
  OAI211_X1 U23048 ( .C1(n20119), .C2(n20118), .A(n20117), .B(n20116), .ZN(
        P1_U3028) );
  AOI21_X1 U23049 ( .B1(n20122), .B2(n20121), .A(n20120), .ZN(n20140) );
  NAND3_X1 U23050 ( .A1(n9813), .A2(n20124), .A3(n20123), .ZN(n20138) );
  NAND2_X1 U23051 ( .A1(n20126), .A2(n20125), .ZN(n20134) );
  OAI21_X1 U23052 ( .B1(n20129), .B2(n20128), .A(n20127), .ZN(n20130) );
  INV_X1 U23053 ( .A(n20130), .ZN(n20131) );
  OR2_X1 U23054 ( .A1(n20132), .A2(n20131), .ZN(n20133) );
  OAI211_X1 U23055 ( .C1(n19999), .C2(n20135), .A(n20134), .B(n20133), .ZN(
        n20136) );
  INV_X1 U23056 ( .A(n20136), .ZN(n20137) );
  AND2_X1 U23057 ( .A1(n20138), .A2(n20137), .ZN(n20139) );
  OAI221_X1 U23058 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20141), .C1(
        n21116), .C2(n20140), .A(n20139), .ZN(P1_U3029) );
  NOR2_X1 U23059 ( .A1(n20143), .A2(n20142), .ZN(P1_U3032) );
  INV_X1 U23060 ( .A(DATAI_16_), .ZN(n21115) );
  INV_X1 U23061 ( .A(n20672), .ZN(n20633) );
  NAND2_X1 U23062 ( .A1(n9821), .A2(n20147), .ZN(n20509) );
  OR2_X1 U23063 ( .A1(n20666), .A2(n20509), .ZN(n20723) );
  INV_X1 U23064 ( .A(DATAI_24_), .ZN(n20148) );
  NOR2_X2 U23065 ( .A1(n20215), .A2(n20152), .ZN(n20663) );
  NAND2_X1 U23066 ( .A1(n20618), .A2(n20420), .ZN(n20278) );
  OR2_X1 U23067 ( .A1(n20545), .A2(n20278), .ZN(n20156) );
  INV_X1 U23068 ( .A(n20156), .ZN(n20216) );
  AOI22_X1 U23069 ( .A1(n20697), .A2(n20630), .B1(n20663), .B2(n20216), .ZN(
        n20165) );
  INV_X1 U23070 ( .A(n20248), .ZN(n20153) );
  OAI21_X1 U23071 ( .B1(n20153), .B2(n20697), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20154) );
  NAND2_X1 U23072 ( .A1(n20154), .A2(n20671), .ZN(n20163) );
  OR2_X1 U23073 ( .A1(n20421), .A2(n20155), .ZN(n20281) );
  NOR2_X1 U23074 ( .A1(n20281), .A2(n20625), .ZN(n20160) );
  INV_X1 U23075 ( .A(n20619), .ZN(n20423) );
  OR2_X1 U23076 ( .A1(n20423), .A2(n20422), .ZN(n20311) );
  AOI22_X1 U23077 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20311), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20156), .ZN(n20158) );
  INV_X1 U23078 ( .A(n20161), .ZN(n20157) );
  NOR2_X1 U23079 ( .A1(n20157), .A2(n13230), .ZN(n20544) );
  NOR2_X1 U23080 ( .A1(n20544), .A2(n20315), .ZN(n20488) );
  OAI211_X1 U23081 ( .C1(n20163), .C2(n20160), .A(n20158), .B(n20488), .ZN(
        n20220) );
  NAND2_X1 U23082 ( .A1(n20218), .A2(n20159), .ZN(n20555) );
  INV_X1 U23083 ( .A(n20160), .ZN(n20162) );
  OR2_X1 U23084 ( .A1(n20161), .A2(n13230), .ZN(n20425) );
  OAI22_X1 U23085 ( .A1(n20163), .A2(n20162), .B1(n20425), .B2(n20311), .ZN(
        n20219) );
  AOI22_X1 U23086 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20220), .B1(
        n20662), .B2(n20219), .ZN(n20164) );
  OAI211_X1 U23087 ( .C1(n20633), .C2(n20248), .A(n20165), .B(n20164), .ZN(
        P1_U3033) );
  INV_X1 U23088 ( .A(DATAI_17_), .ZN(n20166) );
  OAI22_X1 U23089 ( .A1(n20166), .A2(n20210), .B1(n14584), .B2(n20212), .ZN(
        n20589) );
  INV_X1 U23090 ( .A(n20589), .ZN(n20681) );
  INV_X1 U23091 ( .A(DATAI_25_), .ZN(n20167) );
  OAI22_X2 U23092 ( .A1(n20168), .A2(n20212), .B1(n20167), .B2(n20210), .ZN(
        n20678) );
  NOR2_X2 U23093 ( .A1(n20215), .A2(n20169), .ZN(n20677) );
  AOI22_X1 U23094 ( .A1(n20697), .A2(n20678), .B1(n20677), .B2(n20216), .ZN(
        n20172) );
  NAND2_X1 U23095 ( .A1(n20218), .A2(n20170), .ZN(n20558) );
  AOI22_X1 U23096 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20220), .B1(
        n20676), .B2(n20219), .ZN(n20171) );
  OAI211_X1 U23097 ( .C1(n20681), .C2(n20248), .A(n20172), .B(n20171), .ZN(
        P1_U3034) );
  INV_X1 U23098 ( .A(DATAI_18_), .ZN(n20174) );
  OAI22_X1 U23099 ( .A1(n20174), .A2(n20210), .B1(n20173), .B2(n20212), .ZN(
        n20593) );
  INV_X1 U23100 ( .A(n20593), .ZN(n20687) );
  INV_X1 U23101 ( .A(DATAI_26_), .ZN(n20175) );
  OAI22_X2 U23102 ( .A1(n20176), .A2(n20212), .B1(n20175), .B2(n20210), .ZN(
        n20684) );
  NOR2_X2 U23103 ( .A1(n20215), .A2(n20177), .ZN(n20683) );
  AOI22_X1 U23104 ( .A1(n20697), .A2(n20684), .B1(n20683), .B2(n20216), .ZN(
        n20180) );
  NAND2_X1 U23105 ( .A1(n20218), .A2(n20178), .ZN(n20561) );
  AOI22_X1 U23106 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20220), .B1(
        n20682), .B2(n20219), .ZN(n20179) );
  OAI211_X1 U23107 ( .C1(n20687), .C2(n20248), .A(n20180), .B(n20179), .ZN(
        P1_U3035) );
  INV_X1 U23108 ( .A(DATAI_19_), .ZN(n20182) );
  INV_X1 U23109 ( .A(n20690), .ZN(n20641) );
  INV_X1 U23110 ( .A(DATAI_27_), .ZN(n20183) );
  NOR2_X2 U23111 ( .A1(n20215), .A2(n20185), .ZN(n20689) );
  AOI22_X1 U23112 ( .A1(n20697), .A2(n20638), .B1(n20689), .B2(n20216), .ZN(
        n20188) );
  NAND2_X1 U23113 ( .A1(n20218), .A2(n20186), .ZN(n20564) );
  AOI22_X1 U23114 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20220), .B1(
        n20688), .B2(n20219), .ZN(n20187) );
  OAI211_X1 U23115 ( .C1(n20641), .C2(n20248), .A(n20188), .B(n20187), .ZN(
        P1_U3036) );
  INV_X1 U23116 ( .A(DATAI_20_), .ZN(n21006) );
  INV_X1 U23117 ( .A(n20696), .ZN(n20645) );
  INV_X1 U23118 ( .A(DATAI_28_), .ZN(n20190) );
  NOR2_X2 U23119 ( .A1(n20215), .A2(n20192), .ZN(n20695) );
  AOI22_X1 U23120 ( .A1(n20697), .A2(n20642), .B1(n20695), .B2(n20216), .ZN(
        n20195) );
  NAND2_X1 U23121 ( .A1(n20218), .A2(n20193), .ZN(n20567) );
  AOI22_X1 U23122 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20220), .B1(
        n20694), .B2(n20219), .ZN(n20194) );
  OAI211_X1 U23123 ( .C1(n20645), .C2(n20248), .A(n20195), .B(n20194), .ZN(
        P1_U3037) );
  INV_X1 U23124 ( .A(DATAI_21_), .ZN(n20196) );
  OAI22_X1 U23125 ( .A1(n14571), .A2(n20212), .B1(n20196), .B2(n20210), .ZN(
        n20601) );
  INV_X1 U23126 ( .A(n20601), .ZN(n20707) );
  INV_X1 U23127 ( .A(DATAI_29_), .ZN(n20197) );
  OAI22_X2 U23128 ( .A1(n20198), .A2(n20212), .B1(n20197), .B2(n20210), .ZN(
        n20704) );
  AOI22_X1 U23129 ( .A1(n20697), .A2(n20704), .B1(n20703), .B2(n20216), .ZN(
        n20202) );
  NAND2_X1 U23130 ( .A1(n20218), .A2(n20200), .ZN(n20570) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20220), .B1(
        n20702), .B2(n20219), .ZN(n20201) );
  OAI211_X1 U23132 ( .C1(n20707), .C2(n20248), .A(n20202), .B(n20201), .ZN(
        P1_U3038) );
  INV_X1 U23133 ( .A(DATAI_22_), .ZN(n20203) );
  OAI22_X1 U23134 ( .A1(n14567), .A2(n20212), .B1(n20203), .B2(n20210), .ZN(
        n20605) );
  INV_X1 U23135 ( .A(n20605), .ZN(n20713) );
  INV_X1 U23136 ( .A(DATAI_30_), .ZN(n20204) );
  OAI22_X2 U23137 ( .A1(n20205), .A2(n20212), .B1(n20204), .B2(n20210), .ZN(
        n20710) );
  NOR2_X2 U23138 ( .A1(n20215), .A2(n11984), .ZN(n20709) );
  AOI22_X1 U23139 ( .A1(n20697), .A2(n20710), .B1(n20709), .B2(n20216), .ZN(
        n20208) );
  NAND2_X1 U23140 ( .A1(n20218), .A2(n20206), .ZN(n20573) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20220), .B1(
        n20708), .B2(n20219), .ZN(n20207) );
  OAI211_X1 U23142 ( .C1(n20713), .C2(n20248), .A(n20208), .B(n20207), .ZN(
        P1_U3039) );
  INV_X1 U23143 ( .A(DATAI_23_), .ZN(n20209) );
  OAI22_X1 U23144 ( .A1(n14562), .A2(n20212), .B1(n20209), .B2(n20210), .ZN(
        n20611) );
  INV_X1 U23145 ( .A(n20611), .ZN(n20724) );
  INV_X1 U23146 ( .A(DATAI_31_), .ZN(n20211) );
  OAI22_X2 U23147 ( .A1(n20213), .A2(n20212), .B1(n20211), .B2(n20210), .ZN(
        n20718) );
  NOR2_X2 U23148 ( .A1(n20215), .A2(n20214), .ZN(n20717) );
  AOI22_X1 U23149 ( .A1(n20697), .A2(n20718), .B1(n20717), .B2(n20216), .ZN(
        n20222) );
  NAND2_X1 U23150 ( .A1(n20218), .A2(n20217), .ZN(n20579) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20220), .B1(
        n20715), .B2(n20219), .ZN(n20221) );
  OAI211_X1 U23152 ( .C1(n20724), .C2(n20248), .A(n20222), .B(n20221), .ZN(
        P1_U3040) );
  INV_X1 U23153 ( .A(n20630), .ZN(n20675) );
  NOR2_X1 U23154 ( .A1(n20278), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20228) );
  INV_X1 U23155 ( .A(n20228), .ZN(n20225) );
  NOR2_X1 U23156 ( .A1(n20581), .A2(n20225), .ZN(n20244) );
  INV_X1 U23157 ( .A(n20281), .ZN(n20224) );
  INV_X1 U23158 ( .A(n20223), .ZN(n20582) );
  AOI21_X1 U23159 ( .B1(n20224), .B2(n20582), .A(n20244), .ZN(n20226) );
  OAI22_X1 U23160 ( .A1(n20226), .A2(n20669), .B1(n20225), .B2(n13230), .ZN(
        n20243) );
  AOI22_X1 U23161 ( .A1(n20663), .A2(n20244), .B1(n20662), .B2(n20243), .ZN(
        n20230) );
  OAI211_X1 U23162 ( .C1(n20288), .C2(n20622), .A(n20671), .B(n20226), .ZN(
        n20227) );
  OAI211_X1 U23163 ( .C1(n20671), .C2(n20228), .A(n20667), .B(n20227), .ZN(
        n20245) );
  AOI22_X1 U23164 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20245), .B1(
        n20271), .B2(n20672), .ZN(n20229) );
  OAI211_X1 U23165 ( .C1(n20675), .C2(n20248), .A(n20230), .B(n20229), .ZN(
        P1_U3041) );
  INV_X1 U23166 ( .A(n20678), .ZN(n20592) );
  AOI22_X1 U23167 ( .A1(n20677), .A2(n20244), .B1(n20676), .B2(n20243), .ZN(
        n20232) );
  AOI22_X1 U23168 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20245), .B1(
        n20271), .B2(n20589), .ZN(n20231) );
  OAI211_X1 U23169 ( .C1(n20592), .C2(n20248), .A(n20232), .B(n20231), .ZN(
        P1_U3042) );
  INV_X1 U23170 ( .A(n20684), .ZN(n20596) );
  AOI22_X1 U23171 ( .A1(n20683), .A2(n20244), .B1(n20682), .B2(n20243), .ZN(
        n20234) );
  AOI22_X1 U23172 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20245), .B1(
        n20271), .B2(n20593), .ZN(n20233) );
  OAI211_X1 U23173 ( .C1(n20596), .C2(n20248), .A(n20234), .B(n20233), .ZN(
        P1_U3043) );
  INV_X1 U23174 ( .A(n20638), .ZN(n20693) );
  AOI22_X1 U23175 ( .A1(n20689), .A2(n20244), .B1(n20688), .B2(n20243), .ZN(
        n20236) );
  AOI22_X1 U23176 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20245), .B1(
        n20271), .B2(n20690), .ZN(n20235) );
  OAI211_X1 U23177 ( .C1(n20693), .C2(n20248), .A(n20236), .B(n20235), .ZN(
        P1_U3044) );
  INV_X1 U23178 ( .A(n20642), .ZN(n20701) );
  AOI22_X1 U23179 ( .A1(n20695), .A2(n20244), .B1(n20694), .B2(n20243), .ZN(
        n20238) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20245), .B1(
        n20271), .B2(n20696), .ZN(n20237) );
  OAI211_X1 U23181 ( .C1(n20701), .C2(n20248), .A(n20238), .B(n20237), .ZN(
        P1_U3045) );
  INV_X1 U23182 ( .A(n20704), .ZN(n20604) );
  AOI22_X1 U23183 ( .A1(n20703), .A2(n20244), .B1(n20702), .B2(n20243), .ZN(
        n20240) );
  AOI22_X1 U23184 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20245), .B1(
        n20271), .B2(n20601), .ZN(n20239) );
  OAI211_X1 U23185 ( .C1(n20604), .C2(n20248), .A(n20240), .B(n20239), .ZN(
        P1_U3046) );
  INV_X1 U23186 ( .A(n20710), .ZN(n20608) );
  AOI22_X1 U23187 ( .A1(n20709), .A2(n20244), .B1(n20708), .B2(n20243), .ZN(
        n20242) );
  AOI22_X1 U23188 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20245), .B1(
        n20271), .B2(n20605), .ZN(n20241) );
  OAI211_X1 U23189 ( .C1(n20608), .C2(n20248), .A(n20242), .B(n20241), .ZN(
        P1_U3047) );
  INV_X1 U23190 ( .A(n20718), .ZN(n20616) );
  AOI22_X1 U23191 ( .A1(n20717), .A2(n20244), .B1(n20715), .B2(n20243), .ZN(
        n20247) );
  AOI22_X1 U23192 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20245), .B1(
        n20271), .B2(n20611), .ZN(n20246) );
  OAI211_X1 U23193 ( .C1(n20616), .C2(n20248), .A(n20247), .B(n20246), .ZN(
        P1_U3048) );
  INV_X1 U23194 ( .A(n20271), .ZN(n20249) );
  NAND2_X1 U23195 ( .A1(n20249), .A2(n20671), .ZN(n20250) );
  NAND2_X1 U23196 ( .A1(n20671), .A2(n20622), .ZN(n20540) );
  OAI21_X1 U23197 ( .B1(n20250), .B2(n20304), .A(n20540), .ZN(n20254) );
  NOR2_X1 U23198 ( .A1(n20281), .A2(n13725), .ZN(n20251) );
  INV_X1 U23199 ( .A(n20425), .ZN(n20481) );
  NOR2_X1 U23200 ( .A1(n20619), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20362) );
  NOR2_X1 U23201 ( .A1(n20660), .A2(n20278), .ZN(n20283) );
  NAND2_X1 U23202 ( .A1(n20581), .A2(n20283), .ZN(n20252) );
  INV_X1 U23203 ( .A(n20252), .ZN(n20270) );
  AOI22_X1 U23204 ( .A1(n20271), .A2(n20630), .B1(n20663), .B2(n20270), .ZN(
        n20257) );
  INV_X1 U23205 ( .A(n20251), .ZN(n20253) );
  AOI22_X1 U23206 ( .A1(n20254), .A2(n20253), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20252), .ZN(n20255) );
  OAI21_X1 U23207 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20619), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20368) );
  NAND3_X1 U23208 ( .A1(n20488), .A2(n20255), .A3(n20368), .ZN(n20272) );
  AOI22_X1 U23209 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20272), .B1(
        n20304), .B2(n20672), .ZN(n20256) );
  OAI211_X1 U23210 ( .C1(n20275), .C2(n20555), .A(n20257), .B(n20256), .ZN(
        P1_U3049) );
  AOI22_X1 U23211 ( .A1(n20271), .A2(n20678), .B1(n20677), .B2(n20270), .ZN(
        n20259) );
  AOI22_X1 U23212 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20272), .B1(
        n20304), .B2(n20589), .ZN(n20258) );
  OAI211_X1 U23213 ( .C1(n20275), .C2(n20558), .A(n20259), .B(n20258), .ZN(
        P1_U3050) );
  AOI22_X1 U23214 ( .A1(n20304), .A2(n20593), .B1(n20683), .B2(n20270), .ZN(
        n20261) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20272), .B1(
        n20271), .B2(n20684), .ZN(n20260) );
  OAI211_X1 U23216 ( .C1(n20275), .C2(n20561), .A(n20261), .B(n20260), .ZN(
        P1_U3051) );
  AOI22_X1 U23217 ( .A1(n20271), .A2(n20638), .B1(n20689), .B2(n20270), .ZN(
        n20263) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20272), .B1(
        n20304), .B2(n20690), .ZN(n20262) );
  OAI211_X1 U23219 ( .C1(n20275), .C2(n20564), .A(n20263), .B(n20262), .ZN(
        P1_U3052) );
  AOI22_X1 U23220 ( .A1(n20304), .A2(n20696), .B1(n20695), .B2(n20270), .ZN(
        n20265) );
  AOI22_X1 U23221 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20272), .B1(
        n20271), .B2(n20642), .ZN(n20264) );
  OAI211_X1 U23222 ( .C1(n20275), .C2(n20567), .A(n20265), .B(n20264), .ZN(
        P1_U3053) );
  AOI22_X1 U23223 ( .A1(n20304), .A2(n20601), .B1(n20703), .B2(n20270), .ZN(
        n20267) );
  AOI22_X1 U23224 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20272), .B1(
        n20271), .B2(n20704), .ZN(n20266) );
  OAI211_X1 U23225 ( .C1(n20275), .C2(n20570), .A(n20267), .B(n20266), .ZN(
        P1_U3054) );
  AOI22_X1 U23226 ( .A1(n20304), .A2(n20605), .B1(n20709), .B2(n20270), .ZN(
        n20269) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20272), .B1(
        n20271), .B2(n20710), .ZN(n20268) );
  OAI211_X1 U23228 ( .C1(n20275), .C2(n20573), .A(n20269), .B(n20268), .ZN(
        P1_U3055) );
  AOI22_X1 U23229 ( .A1(n20304), .A2(n20611), .B1(n20717), .B2(n20270), .ZN(
        n20274) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20272), .B1(
        n20271), .B2(n20718), .ZN(n20273) );
  OAI211_X1 U23231 ( .C1(n20275), .C2(n20579), .A(n20274), .B(n20273), .ZN(
        P1_U3056) );
  INV_X1 U23232 ( .A(n20665), .ZN(n20514) );
  AOI21_X1 U23233 ( .B1(n20276), .B2(n20514), .A(n20669), .ZN(n20282) );
  AND2_X1 U23234 ( .A1(n20277), .A2(n13147), .ZN(n20657) );
  INV_X1 U23235 ( .A(n20657), .ZN(n20280) );
  NOR2_X1 U23236 ( .A1(n20656), .A2(n20278), .ZN(n20303) );
  INV_X1 U23237 ( .A(n20303), .ZN(n20279) );
  OAI21_X1 U23238 ( .B1(n20281), .B2(n20280), .A(n20279), .ZN(n20286) );
  AOI22_X1 U23239 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20283), .B1(n20282), 
        .B2(n20286), .ZN(n20308) );
  AOI22_X1 U23240 ( .A1(n20304), .A2(n20630), .B1(n20663), .B2(n20303), .ZN(
        n20290) );
  INV_X1 U23241 ( .A(n20282), .ZN(n20287) );
  OAI21_X1 U23242 ( .B1(n20671), .B2(n20283), .A(n20667), .ZN(n20284) );
  INV_X1 U23243 ( .A(n20284), .ZN(n20285) );
  OAI21_X1 U23244 ( .B1(n20287), .B2(n20286), .A(n20285), .ZN(n20305) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20305), .B1(
        n20332), .B2(n20672), .ZN(n20289) );
  OAI211_X1 U23246 ( .C1(n20308), .C2(n20555), .A(n20290), .B(n20289), .ZN(
        P1_U3057) );
  AOI22_X1 U23247 ( .A1(n20332), .A2(n20589), .B1(n20677), .B2(n20303), .ZN(
        n20292) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20305), .B1(
        n20304), .B2(n20678), .ZN(n20291) );
  OAI211_X1 U23249 ( .C1(n20308), .C2(n20558), .A(n20292), .B(n20291), .ZN(
        P1_U3058) );
  AOI22_X1 U23250 ( .A1(n20304), .A2(n20684), .B1(n20683), .B2(n20303), .ZN(
        n20294) );
  AOI22_X1 U23251 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20305), .B1(
        n20332), .B2(n20593), .ZN(n20293) );
  OAI211_X1 U23252 ( .C1(n20308), .C2(n20561), .A(n20294), .B(n20293), .ZN(
        P1_U3059) );
  AOI22_X1 U23253 ( .A1(n20332), .A2(n20690), .B1(n20689), .B2(n20303), .ZN(
        n20296) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20305), .B1(
        n20304), .B2(n20638), .ZN(n20295) );
  OAI211_X1 U23255 ( .C1(n20308), .C2(n20564), .A(n20296), .B(n20295), .ZN(
        P1_U3060) );
  AOI22_X1 U23256 ( .A1(n20332), .A2(n20696), .B1(n20695), .B2(n20303), .ZN(
        n20298) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20305), .B1(
        n20304), .B2(n20642), .ZN(n20297) );
  OAI211_X1 U23258 ( .C1(n20308), .C2(n20567), .A(n20298), .B(n20297), .ZN(
        P1_U3061) );
  AOI22_X1 U23259 ( .A1(n20332), .A2(n20601), .B1(n20703), .B2(n20303), .ZN(
        n20300) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20305), .B1(
        n20304), .B2(n20704), .ZN(n20299) );
  OAI211_X1 U23261 ( .C1(n20308), .C2(n20570), .A(n20300), .B(n20299), .ZN(
        P1_U3062) );
  AOI22_X1 U23262 ( .A1(n20332), .A2(n20605), .B1(n20709), .B2(n20303), .ZN(
        n20302) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20305), .B1(
        n20304), .B2(n20710), .ZN(n20301) );
  OAI211_X1 U23264 ( .C1(n20308), .C2(n20573), .A(n20302), .B(n20301), .ZN(
        P1_U3063) );
  AOI22_X1 U23265 ( .A1(n20332), .A2(n20611), .B1(n20717), .B2(n20303), .ZN(
        n20307) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20305), .B1(
        n20304), .B2(n20718), .ZN(n20306) );
  OAI211_X1 U23267 ( .C1(n20308), .C2(n20579), .A(n20307), .B(n20306), .ZN(
        P1_U3064) );
  INV_X1 U23268 ( .A(n20544), .ZN(n20620) );
  NOR2_X1 U23269 ( .A1(n13091), .A2(n20309), .ZN(n20392) );
  NAND3_X1 U23270 ( .A1(n20392), .A2(n20671), .A3(n13725), .ZN(n20310) );
  OAI21_X1 U23271 ( .B1(n20620), .B2(n20311), .A(n20310), .ZN(n20331) );
  AOI22_X1 U23272 ( .A1(n20663), .A2(n9934), .B1(n20662), .B2(n20331), .ZN(
        n20318) );
  INV_X1 U23273 ( .A(n20332), .ZN(n20312) );
  AOI21_X1 U23274 ( .B1(n20312), .B2(n20359), .A(n20622), .ZN(n20313) );
  AOI21_X1 U23275 ( .B1(n20392), .B2(n13725), .A(n20313), .ZN(n20314) );
  NOR2_X1 U23276 ( .A1(n20314), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20316) );
  NOR2_X1 U23277 ( .A1(n20481), .A2(n20315), .ZN(n20628) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20630), .ZN(n20317) );
  OAI211_X1 U23279 ( .C1(n20633), .C2(n20359), .A(n20318), .B(n20317), .ZN(
        P1_U3065) );
  AOI22_X1 U23280 ( .A1(n20677), .A2(n9934), .B1(n20676), .B2(n20331), .ZN(
        n20320) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20678), .ZN(n20319) );
  OAI211_X1 U23282 ( .C1(n20681), .C2(n20359), .A(n20320), .B(n20319), .ZN(
        P1_U3066) );
  AOI22_X1 U23283 ( .A1(n20683), .A2(n9934), .B1(n20682), .B2(n20331), .ZN(
        n20322) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20684), .ZN(n20321) );
  OAI211_X1 U23285 ( .C1(n20687), .C2(n20359), .A(n20322), .B(n20321), .ZN(
        P1_U3067) );
  AOI22_X1 U23286 ( .A1(n20689), .A2(n9934), .B1(n20688), .B2(n20331), .ZN(
        n20324) );
  AOI22_X1 U23287 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20638), .ZN(n20323) );
  OAI211_X1 U23288 ( .C1(n20641), .C2(n20359), .A(n20324), .B(n20323), .ZN(
        P1_U3068) );
  AOI22_X1 U23289 ( .A1(n20695), .A2(n9934), .B1(n20694), .B2(n20331), .ZN(
        n20326) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20642), .ZN(n20325) );
  OAI211_X1 U23291 ( .C1(n20645), .C2(n20359), .A(n20326), .B(n20325), .ZN(
        P1_U3069) );
  AOI22_X1 U23292 ( .A1(n20703), .A2(n9934), .B1(n20702), .B2(n20331), .ZN(
        n20328) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20704), .ZN(n20327) );
  OAI211_X1 U23294 ( .C1(n20707), .C2(n20359), .A(n20328), .B(n20327), .ZN(
        P1_U3070) );
  AOI22_X1 U23295 ( .A1(n20709), .A2(n9934), .B1(n20708), .B2(n20331), .ZN(
        n20330) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20710), .ZN(n20329) );
  OAI211_X1 U23297 ( .C1(n20713), .C2(n20359), .A(n20330), .B(n20329), .ZN(
        P1_U3071) );
  AOI22_X1 U23298 ( .A1(n20717), .A2(n9934), .B1(n20715), .B2(n20331), .ZN(
        n20335) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20333), .B1(
        n20332), .B2(n20718), .ZN(n20334) );
  OAI211_X1 U23300 ( .C1(n20724), .C2(n20359), .A(n20335), .B(n20334), .ZN(
        P1_U3072) );
  NOR2_X1 U23301 ( .A1(n20363), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20339) );
  INV_X1 U23302 ( .A(n20339), .ZN(n20336) );
  NOR2_X1 U23303 ( .A1(n20581), .A2(n20336), .ZN(n20355) );
  AOI21_X1 U23304 ( .B1(n20392), .B2(n20582), .A(n20355), .ZN(n20337) );
  OAI22_X1 U23305 ( .A1(n20337), .A2(n20669), .B1(n20336), .B2(n13230), .ZN(
        n20354) );
  AOI22_X1 U23306 ( .A1(n20663), .A2(n20355), .B1(n20662), .B2(n20354), .ZN(
        n20341) );
  OAI211_X1 U23307 ( .C1(n20390), .C2(n20622), .A(n20671), .B(n20337), .ZN(
        n20338) );
  OAI211_X1 U23308 ( .C1(n20671), .C2(n20339), .A(n20667), .B(n20338), .ZN(
        n20356) );
  NOR2_X2 U23309 ( .A1(n20390), .A2(n20586), .ZN(n20385) );
  AOI22_X1 U23310 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20356), .B1(
        n20385), .B2(n20672), .ZN(n20340) );
  OAI211_X1 U23311 ( .C1(n20675), .C2(n20359), .A(n20341), .B(n20340), .ZN(
        P1_U3073) );
  AOI22_X1 U23312 ( .A1(n20677), .A2(n20355), .B1(n20676), .B2(n20354), .ZN(
        n20343) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20356), .B1(
        n20385), .B2(n20589), .ZN(n20342) );
  OAI211_X1 U23314 ( .C1(n20592), .C2(n20359), .A(n20343), .B(n20342), .ZN(
        P1_U3074) );
  AOI22_X1 U23315 ( .A1(n20683), .A2(n20355), .B1(n20682), .B2(n20354), .ZN(
        n20345) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20356), .B1(
        n20385), .B2(n20593), .ZN(n20344) );
  OAI211_X1 U23317 ( .C1(n20596), .C2(n20359), .A(n20345), .B(n20344), .ZN(
        P1_U3075) );
  AOI22_X1 U23318 ( .A1(n20689), .A2(n20355), .B1(n20688), .B2(n20354), .ZN(
        n20347) );
  AOI22_X1 U23319 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20356), .B1(
        n20385), .B2(n20690), .ZN(n20346) );
  OAI211_X1 U23320 ( .C1(n20693), .C2(n20359), .A(n20347), .B(n20346), .ZN(
        P1_U3076) );
  AOI22_X1 U23321 ( .A1(n20695), .A2(n20355), .B1(n20694), .B2(n20354), .ZN(
        n20349) );
  AOI22_X1 U23322 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20356), .B1(
        n20385), .B2(n20696), .ZN(n20348) );
  OAI211_X1 U23323 ( .C1(n20701), .C2(n20359), .A(n20349), .B(n20348), .ZN(
        P1_U3077) );
  AOI22_X1 U23324 ( .A1(n20703), .A2(n20355), .B1(n20702), .B2(n20354), .ZN(
        n20351) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20356), .B1(
        n20385), .B2(n20601), .ZN(n20350) );
  OAI211_X1 U23326 ( .C1(n20604), .C2(n20359), .A(n20351), .B(n20350), .ZN(
        P1_U3078) );
  AOI22_X1 U23327 ( .A1(n20709), .A2(n20355), .B1(n20708), .B2(n20354), .ZN(
        n20353) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20356), .B1(
        n20385), .B2(n20605), .ZN(n20352) );
  OAI211_X1 U23329 ( .C1(n20608), .C2(n20359), .A(n20353), .B(n20352), .ZN(
        P1_U3079) );
  AOI22_X1 U23330 ( .A1(n20717), .A2(n20355), .B1(n20715), .B2(n20354), .ZN(
        n20358) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20356), .B1(
        n20385), .B2(n20611), .ZN(n20357) );
  OAI211_X1 U23332 ( .C1(n20616), .C2(n20359), .A(n20358), .B(n20357), .ZN(
        P1_U3080) );
  INV_X1 U23333 ( .A(n20385), .ZN(n20360) );
  NAND2_X1 U23334 ( .A1(n20360), .A2(n20671), .ZN(n20361) );
  NOR2_X2 U23335 ( .A1(n20390), .A2(n20617), .ZN(n20415) );
  OAI21_X1 U23336 ( .B1(n20361), .B2(n20415), .A(n20540), .ZN(n20367) );
  AND2_X1 U23337 ( .A1(n20392), .A2(n20625), .ZN(n20364) );
  NOR2_X1 U23338 ( .A1(n20660), .A2(n20363), .ZN(n20398) );
  NAND2_X1 U23339 ( .A1(n20581), .A2(n20398), .ZN(n20365) );
  INV_X1 U23340 ( .A(n20365), .ZN(n20384) );
  AOI22_X1 U23341 ( .A1(n20385), .A2(n20630), .B1(n20663), .B2(n20384), .ZN(
        n20371) );
  INV_X1 U23342 ( .A(n20364), .ZN(n20366) );
  AOI22_X1 U23343 ( .A1(n20367), .A2(n20366), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20365), .ZN(n20369) );
  NAND3_X1 U23344 ( .A1(n20628), .A2(n20369), .A3(n20368), .ZN(n20386) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20386), .B1(
        n20415), .B2(n20672), .ZN(n20370) );
  OAI211_X1 U23346 ( .C1(n20389), .C2(n20555), .A(n20371), .B(n20370), .ZN(
        P1_U3081) );
  AOI22_X1 U23347 ( .A1(n20385), .A2(n20678), .B1(n20677), .B2(n20384), .ZN(
        n20373) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20386), .B1(
        n20415), .B2(n20589), .ZN(n20372) );
  OAI211_X1 U23349 ( .C1(n20389), .C2(n20558), .A(n20373), .B(n20372), .ZN(
        P1_U3082) );
  AOI22_X1 U23350 ( .A1(n20415), .A2(n20593), .B1(n20683), .B2(n20384), .ZN(
        n20375) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20386), .B1(
        n20385), .B2(n20684), .ZN(n20374) );
  OAI211_X1 U23352 ( .C1(n20389), .C2(n20561), .A(n20375), .B(n20374), .ZN(
        P1_U3083) );
  AOI22_X1 U23353 ( .A1(n20415), .A2(n20690), .B1(n20689), .B2(n20384), .ZN(
        n20377) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20386), .B1(
        n20385), .B2(n20638), .ZN(n20376) );
  OAI211_X1 U23355 ( .C1(n20389), .C2(n20564), .A(n20377), .B(n20376), .ZN(
        P1_U3084) );
  AOI22_X1 U23356 ( .A1(n20385), .A2(n20642), .B1(n20695), .B2(n20384), .ZN(
        n20379) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20386), .B1(
        n20415), .B2(n20696), .ZN(n20378) );
  OAI211_X1 U23358 ( .C1(n20389), .C2(n20567), .A(n20379), .B(n20378), .ZN(
        P1_U3085) );
  AOI22_X1 U23359 ( .A1(n20385), .A2(n20704), .B1(n20703), .B2(n20384), .ZN(
        n20381) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20386), .B1(
        n20415), .B2(n20601), .ZN(n20380) );
  OAI211_X1 U23361 ( .C1(n20389), .C2(n20570), .A(n20381), .B(n20380), .ZN(
        P1_U3086) );
  AOI22_X1 U23362 ( .A1(n20415), .A2(n20605), .B1(n20709), .B2(n20384), .ZN(
        n20383) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20386), .B1(
        n20385), .B2(n20710), .ZN(n20382) );
  OAI211_X1 U23364 ( .C1(n20389), .C2(n20573), .A(n20383), .B(n20382), .ZN(
        P1_U3087) );
  AOI22_X1 U23365 ( .A1(n20385), .A2(n20718), .B1(n20717), .B2(n20384), .ZN(
        n20388) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20386), .B1(
        n20415), .B2(n20611), .ZN(n20387) );
  OAI211_X1 U23367 ( .C1(n20389), .C2(n20579), .A(n20388), .B(n20387), .ZN(
        P1_U3088) );
  INV_X1 U23368 ( .A(n20391), .ZN(n20414) );
  AOI21_X1 U23369 ( .B1(n20392), .B2(n20657), .A(n20414), .ZN(n20395) );
  INV_X1 U23370 ( .A(n20398), .ZN(n20393) );
  OAI22_X1 U23371 ( .A1(n20395), .A2(n20669), .B1(n20393), .B2(n13230), .ZN(
        n20413) );
  AOI22_X1 U23372 ( .A1(n20663), .A2(n20414), .B1(n20662), .B2(n20413), .ZN(
        n20400) );
  INV_X1 U23373 ( .A(n20394), .ZN(n20396) );
  NAND3_X1 U23374 ( .A1(n20396), .A2(n20671), .A3(n20395), .ZN(n20397) );
  OAI211_X1 U23375 ( .C1(n20671), .C2(n20398), .A(n20667), .B(n20397), .ZN(
        n20416) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20630), .ZN(n20399) );
  OAI211_X1 U23377 ( .C1(n20633), .C2(n20426), .A(n20400), .B(n20399), .ZN(
        P1_U3089) );
  AOI22_X1 U23378 ( .A1(n20677), .A2(n20414), .B1(n20676), .B2(n20413), .ZN(
        n20402) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20678), .ZN(n20401) );
  OAI211_X1 U23380 ( .C1(n20681), .C2(n20426), .A(n20402), .B(n20401), .ZN(
        P1_U3090) );
  AOI22_X1 U23381 ( .A1(n20683), .A2(n20414), .B1(n20682), .B2(n20413), .ZN(
        n20404) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20684), .ZN(n20403) );
  OAI211_X1 U23383 ( .C1(n20687), .C2(n20426), .A(n20404), .B(n20403), .ZN(
        P1_U3091) );
  AOI22_X1 U23384 ( .A1(n20689), .A2(n20414), .B1(n20688), .B2(n20413), .ZN(
        n20406) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20638), .ZN(n20405) );
  OAI211_X1 U23386 ( .C1(n20641), .C2(n20426), .A(n20406), .B(n20405), .ZN(
        P1_U3092) );
  AOI22_X1 U23387 ( .A1(n20695), .A2(n20414), .B1(n20694), .B2(n20413), .ZN(
        n20408) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20642), .ZN(n20407) );
  OAI211_X1 U23389 ( .C1(n20645), .C2(n20426), .A(n20408), .B(n20407), .ZN(
        P1_U3093) );
  AOI22_X1 U23390 ( .A1(n20703), .A2(n20414), .B1(n20702), .B2(n20413), .ZN(
        n20410) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20704), .ZN(n20409) );
  OAI211_X1 U23392 ( .C1(n20707), .C2(n20426), .A(n20410), .B(n20409), .ZN(
        P1_U3094) );
  AOI22_X1 U23393 ( .A1(n20709), .A2(n20414), .B1(n20708), .B2(n20413), .ZN(
        n20412) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20710), .ZN(n20411) );
  OAI211_X1 U23395 ( .C1(n20713), .C2(n20426), .A(n20412), .B(n20411), .ZN(
        P1_U3095) );
  AOI22_X1 U23396 ( .A1(n20717), .A2(n20414), .B1(n20715), .B2(n20413), .ZN(
        n20418) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20718), .ZN(n20417) );
  OAI211_X1 U23398 ( .C1(n20724), .C2(n20426), .A(n20418), .B(n20417), .ZN(
        P1_U3096) );
  NAND2_X1 U23399 ( .A1(n20420), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20511) );
  AND2_X1 U23400 ( .A1(n20421), .A2(n13091), .ZN(n20512) );
  AOI21_X1 U23401 ( .B1(n20512), .B2(n13725), .A(n10346), .ZN(n20428) );
  INV_X1 U23402 ( .A(n20422), .ZN(n20424) );
  NOR2_X1 U23403 ( .A1(n20424), .A2(n20423), .ZN(n20543) );
  INV_X1 U23404 ( .A(n20543), .ZN(n20547) );
  OAI22_X1 U23405 ( .A1(n20428), .A2(n20669), .B1(n20425), .B2(n20547), .ZN(
        n20445) );
  AOI22_X1 U23406 ( .A1(n20663), .A2(n10346), .B1(n20662), .B2(n20445), .ZN(
        n20432) );
  INV_X1 U23407 ( .A(n20476), .ZN(n20427) );
  OAI21_X1 U23408 ( .B1(n20427), .B2(n20446), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20429) );
  NAND2_X1 U23409 ( .A1(n20429), .A2(n20428), .ZN(n20430) );
  OAI211_X1 U23410 ( .C1(n10346), .C2(n20551), .A(n20488), .B(n20430), .ZN(
        n20447) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20447), .B1(
        n20446), .B2(n20630), .ZN(n20431) );
  OAI211_X1 U23412 ( .C1(n20633), .C2(n20476), .A(n20432), .B(n20431), .ZN(
        P1_U3097) );
  AOI22_X1 U23413 ( .A1(n20677), .A2(n10346), .B1(n20676), .B2(n20445), .ZN(
        n20434) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20447), .B1(
        n20446), .B2(n20678), .ZN(n20433) );
  OAI211_X1 U23415 ( .C1(n20681), .C2(n20476), .A(n20434), .B(n20433), .ZN(
        P1_U3098) );
  AOI22_X1 U23416 ( .A1(n20683), .A2(n10346), .B1(n20682), .B2(n20445), .ZN(
        n20436) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20447), .B1(
        n20446), .B2(n20684), .ZN(n20435) );
  OAI211_X1 U23418 ( .C1(n20687), .C2(n20476), .A(n20436), .B(n20435), .ZN(
        P1_U3099) );
  AOI22_X1 U23419 ( .A1(n20689), .A2(n10346), .B1(n20688), .B2(n20445), .ZN(
        n20438) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20447), .B1(
        n20446), .B2(n20638), .ZN(n20437) );
  OAI211_X1 U23421 ( .C1(n20641), .C2(n20476), .A(n20438), .B(n20437), .ZN(
        P1_U3100) );
  AOI22_X1 U23422 ( .A1(n20695), .A2(n10346), .B1(n20694), .B2(n20445), .ZN(
        n20440) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20447), .B1(
        n20446), .B2(n20642), .ZN(n20439) );
  OAI211_X1 U23424 ( .C1(n20645), .C2(n20476), .A(n20440), .B(n20439), .ZN(
        P1_U3101) );
  AOI22_X1 U23425 ( .A1(n20703), .A2(n10346), .B1(n20702), .B2(n20445), .ZN(
        n20442) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20447), .B1(
        n20446), .B2(n20704), .ZN(n20441) );
  OAI211_X1 U23427 ( .C1(n20707), .C2(n20476), .A(n20442), .B(n20441), .ZN(
        P1_U3102) );
  AOI22_X1 U23428 ( .A1(n20709), .A2(n10346), .B1(n20708), .B2(n20445), .ZN(
        n20444) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20447), .B1(
        n20446), .B2(n20710), .ZN(n20443) );
  OAI211_X1 U23430 ( .C1(n20713), .C2(n20476), .A(n20444), .B(n20443), .ZN(
        P1_U3103) );
  AOI22_X1 U23431 ( .A1(n20717), .A2(n10346), .B1(n20715), .B2(n20445), .ZN(
        n20449) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20447), .B1(
        n20446), .B2(n20718), .ZN(n20448) );
  OAI211_X1 U23433 ( .C1(n20724), .C2(n20476), .A(n20449), .B(n20448), .ZN(
        P1_U3104) );
  NOR2_X1 U23434 ( .A1(n20511), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20455) );
  INV_X1 U23435 ( .A(n20455), .ZN(n20450) );
  NOR2_X1 U23436 ( .A1(n20581), .A2(n20450), .ZN(n20472) );
  AOI21_X1 U23437 ( .B1(n20512), .B2(n20582), .A(n20472), .ZN(n20451) );
  OAI22_X1 U23438 ( .A1(n20451), .A2(n20669), .B1(n20450), .B2(n13230), .ZN(
        n20471) );
  AOI22_X1 U23439 ( .A1(n20663), .A2(n20472), .B1(n20662), .B2(n20471), .ZN(
        n20458) );
  INV_X1 U23440 ( .A(n20515), .ZN(n20453) );
  INV_X1 U23441 ( .A(n20540), .ZN(n20452) );
  OAI21_X1 U23442 ( .B1(n20453), .B2(n20452), .A(n20451), .ZN(n20454) );
  OAI211_X1 U23443 ( .C1(n20671), .C2(n20455), .A(n20667), .B(n20454), .ZN(
        n20473) );
  INV_X1 U23444 ( .A(n20586), .ZN(n20456) );
  AOI22_X1 U23445 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20473), .B1(
        n20504), .B2(n20672), .ZN(n20457) );
  OAI211_X1 U23446 ( .C1(n20675), .C2(n20476), .A(n20458), .B(n20457), .ZN(
        P1_U3105) );
  AOI22_X1 U23447 ( .A1(n20677), .A2(n20472), .B1(n20676), .B2(n20471), .ZN(
        n20460) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20473), .B1(
        n20504), .B2(n20589), .ZN(n20459) );
  OAI211_X1 U23449 ( .C1(n20592), .C2(n20476), .A(n20460), .B(n20459), .ZN(
        P1_U3106) );
  AOI22_X1 U23450 ( .A1(n20683), .A2(n20472), .B1(n20682), .B2(n20471), .ZN(
        n20462) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20473), .B1(
        n20504), .B2(n20593), .ZN(n20461) );
  OAI211_X1 U23452 ( .C1(n20596), .C2(n20476), .A(n20462), .B(n20461), .ZN(
        P1_U3107) );
  AOI22_X1 U23453 ( .A1(n20689), .A2(n20472), .B1(n20688), .B2(n20471), .ZN(
        n20464) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20473), .B1(
        n20504), .B2(n20690), .ZN(n20463) );
  OAI211_X1 U23455 ( .C1(n20693), .C2(n20476), .A(n20464), .B(n20463), .ZN(
        P1_U3108) );
  AOI22_X1 U23456 ( .A1(n20695), .A2(n20472), .B1(n20694), .B2(n20471), .ZN(
        n20466) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20473), .B1(
        n20504), .B2(n20696), .ZN(n20465) );
  OAI211_X1 U23458 ( .C1(n20701), .C2(n20476), .A(n20466), .B(n20465), .ZN(
        P1_U3109) );
  AOI22_X1 U23459 ( .A1(n20703), .A2(n20472), .B1(n20702), .B2(n20471), .ZN(
        n20468) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20473), .B1(
        n20504), .B2(n20601), .ZN(n20467) );
  OAI211_X1 U23461 ( .C1(n20604), .C2(n20476), .A(n20468), .B(n20467), .ZN(
        P1_U3110) );
  AOI22_X1 U23462 ( .A1(n20709), .A2(n20472), .B1(n20708), .B2(n20471), .ZN(
        n20470) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20473), .B1(
        n20504), .B2(n20605), .ZN(n20469) );
  OAI211_X1 U23464 ( .C1(n20608), .C2(n20476), .A(n20470), .B(n20469), .ZN(
        P1_U3111) );
  AOI22_X1 U23465 ( .A1(n20717), .A2(n20472), .B1(n20715), .B2(n20471), .ZN(
        n20475) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20473), .B1(
        n20504), .B2(n20611), .ZN(n20474) );
  OAI211_X1 U23467 ( .C1(n20616), .C2(n20476), .A(n20475), .B(n20474), .ZN(
        P1_U3112) );
  INV_X1 U23468 ( .A(n20504), .ZN(n20477) );
  NAND2_X1 U23469 ( .A1(n20477), .A2(n20671), .ZN(n20479) );
  OAI21_X1 U23470 ( .B1(n20479), .B2(n20535), .A(n20540), .ZN(n20486) );
  AND2_X1 U23471 ( .A1(n20512), .A2(n20625), .ZN(n20483) );
  NOR2_X1 U23472 ( .A1(n20619), .A2(n20618), .ZN(n20480) );
  INV_X1 U23473 ( .A(n20511), .ZN(n20482) );
  NAND2_X1 U23474 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20482), .ZN(
        n20516) );
  NOR2_X1 U23475 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20516), .ZN(
        n20503) );
  AOI22_X1 U23476 ( .A1(n20504), .A2(n20630), .B1(n20503), .B2(n20663), .ZN(
        n20490) );
  INV_X1 U23477 ( .A(n20483), .ZN(n20485) );
  INV_X1 U23478 ( .A(n20503), .ZN(n20484) );
  AOI22_X1 U23479 ( .A1(n20486), .A2(n20485), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20484), .ZN(n20487) );
  OAI21_X1 U23480 ( .B1(n20618), .B2(n20619), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20627) );
  NAND3_X1 U23481 ( .A1(n20488), .A2(n20487), .A3(n20627), .ZN(n20505) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20505), .B1(
        n20535), .B2(n20672), .ZN(n20489) );
  OAI211_X1 U23483 ( .C1(n20508), .C2(n20555), .A(n20490), .B(n20489), .ZN(
        P1_U3113) );
  AOI22_X1 U23484 ( .A1(n20504), .A2(n20678), .B1(n20503), .B2(n20677), .ZN(
        n20492) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20505), .B1(
        n20535), .B2(n20589), .ZN(n20491) );
  OAI211_X1 U23486 ( .C1(n20508), .C2(n20558), .A(n20492), .B(n20491), .ZN(
        P1_U3114) );
  AOI22_X1 U23487 ( .A1(n20535), .A2(n20593), .B1(n20683), .B2(n20503), .ZN(
        n20494) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20505), .B1(
        n20504), .B2(n20684), .ZN(n20493) );
  OAI211_X1 U23489 ( .C1(n20508), .C2(n20561), .A(n20494), .B(n20493), .ZN(
        P1_U3115) );
  AOI22_X1 U23490 ( .A1(n20504), .A2(n20638), .B1(n20503), .B2(n20689), .ZN(
        n20496) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20505), .B1(
        n20535), .B2(n20690), .ZN(n20495) );
  OAI211_X1 U23492 ( .C1(n20508), .C2(n20564), .A(n20496), .B(n20495), .ZN(
        P1_U3116) );
  AOI22_X1 U23493 ( .A1(n20535), .A2(n20696), .B1(n20503), .B2(n20695), .ZN(
        n20498) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20505), .B1(
        n20504), .B2(n20642), .ZN(n20497) );
  OAI211_X1 U23495 ( .C1(n20508), .C2(n20567), .A(n20498), .B(n20497), .ZN(
        P1_U3117) );
  AOI22_X1 U23496 ( .A1(n20504), .A2(n20704), .B1(n20503), .B2(n20703), .ZN(
        n20500) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20505), .B1(
        n20535), .B2(n20601), .ZN(n20499) );
  OAI211_X1 U23498 ( .C1(n20508), .C2(n20570), .A(n20500), .B(n20499), .ZN(
        P1_U3118) );
  AOI22_X1 U23499 ( .A1(n20504), .A2(n20710), .B1(n20503), .B2(n20709), .ZN(
        n20502) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20505), .B1(
        n20535), .B2(n20605), .ZN(n20501) );
  OAI211_X1 U23501 ( .C1(n20508), .C2(n20573), .A(n20502), .B(n20501), .ZN(
        P1_U3119) );
  AOI22_X1 U23502 ( .A1(n20504), .A2(n20718), .B1(n20503), .B2(n20717), .ZN(
        n20507) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20505), .B1(
        n20535), .B2(n20611), .ZN(n20506) );
  OAI211_X1 U23504 ( .C1(n20508), .C2(n20579), .A(n20507), .B(n20506), .ZN(
        P1_U3120) );
  INV_X1 U23505 ( .A(n20509), .ZN(n20510) );
  NOR2_X1 U23506 ( .A1(n20656), .A2(n20511), .ZN(n20534) );
  AOI21_X1 U23507 ( .B1(n20512), .B2(n20657), .A(n20534), .ZN(n20513) );
  OAI22_X1 U23508 ( .A1(n20513), .A2(n20669), .B1(n20516), .B2(n13230), .ZN(
        n20533) );
  AOI22_X1 U23509 ( .A1(n20663), .A2(n20534), .B1(n20662), .B2(n20533), .ZN(
        n20520) );
  NAND3_X1 U23510 ( .A1(n20515), .A2(n20671), .A3(n20514), .ZN(n20517) );
  NAND2_X1 U23511 ( .A1(n20517), .A2(n20516), .ZN(n20518) );
  NAND2_X1 U23512 ( .A1(n20518), .A2(n20667), .ZN(n20536) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20630), .ZN(n20519) );
  OAI211_X1 U23514 ( .C1(n20633), .C2(n20552), .A(n20520), .B(n20519), .ZN(
        P1_U3121) );
  AOI22_X1 U23515 ( .A1(n20677), .A2(n20534), .B1(n20676), .B2(n20533), .ZN(
        n20522) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20678), .ZN(n20521) );
  OAI211_X1 U23517 ( .C1(n20681), .C2(n20552), .A(n20522), .B(n20521), .ZN(
        P1_U3122) );
  AOI22_X1 U23518 ( .A1(n20683), .A2(n20534), .B1(n20682), .B2(n20533), .ZN(
        n20524) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20684), .ZN(n20523) );
  OAI211_X1 U23520 ( .C1(n20687), .C2(n20552), .A(n20524), .B(n20523), .ZN(
        P1_U3123) );
  AOI22_X1 U23521 ( .A1(n20689), .A2(n20534), .B1(n20688), .B2(n20533), .ZN(
        n20526) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20638), .ZN(n20525) );
  OAI211_X1 U23523 ( .C1(n20641), .C2(n20552), .A(n20526), .B(n20525), .ZN(
        P1_U3124) );
  AOI22_X1 U23524 ( .A1(n20695), .A2(n20534), .B1(n20694), .B2(n20533), .ZN(
        n20528) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20642), .ZN(n20527) );
  OAI211_X1 U23526 ( .C1(n20645), .C2(n20552), .A(n20528), .B(n20527), .ZN(
        P1_U3125) );
  AOI22_X1 U23527 ( .A1(n20703), .A2(n20534), .B1(n20702), .B2(n20533), .ZN(
        n20530) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20704), .ZN(n20529) );
  OAI211_X1 U23529 ( .C1(n20707), .C2(n20552), .A(n20530), .B(n20529), .ZN(
        P1_U3126) );
  AOI22_X1 U23530 ( .A1(n20709), .A2(n20534), .B1(n20708), .B2(n20533), .ZN(
        n20532) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20710), .ZN(n20531) );
  OAI211_X1 U23532 ( .C1(n20713), .C2(n20552), .A(n20532), .B(n20531), .ZN(
        P1_U3127) );
  AOI22_X1 U23533 ( .A1(n20717), .A2(n20534), .B1(n20715), .B2(n20533), .ZN(
        n20538) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20718), .ZN(n20537) );
  OAI211_X1 U23535 ( .C1(n20724), .C2(n20552), .A(n20538), .B(n20537), .ZN(
        P1_U3128) );
  NAND3_X1 U23536 ( .A1(n20552), .A2(n20671), .A3(n20615), .ZN(n20541) );
  NAND2_X1 U23537 ( .A1(n20541), .A2(n20540), .ZN(n20549) );
  OR2_X1 U23538 ( .A1(n13091), .A2(n20542), .ZN(n20621) );
  NOR2_X1 U23539 ( .A1(n20621), .A2(n20625), .ZN(n20546) );
  AOI22_X1 U23540 ( .A1(n20549), .A2(n20546), .B1(n20544), .B2(n20543), .ZN(
        n20580) );
  NAND2_X1 U23541 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20659) );
  AOI22_X1 U23542 ( .A1(n20574), .A2(n20672), .B1(n20663), .B2(n9935), .ZN(
        n20554) );
  INV_X1 U23543 ( .A(n20546), .ZN(n20548) );
  AOI22_X1 U23544 ( .A1(n20549), .A2(n20548), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20547), .ZN(n20550) );
  OAI211_X1 U23545 ( .C1(n9935), .C2(n20551), .A(n20628), .B(n20550), .ZN(
        n20576) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20630), .ZN(n20553) );
  OAI211_X1 U23547 ( .C1(n20580), .C2(n20555), .A(n20554), .B(n20553), .ZN(
        P1_U3129) );
  AOI22_X1 U23548 ( .A1(n20574), .A2(n20589), .B1(n20677), .B2(n9935), .ZN(
        n20557) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20678), .ZN(n20556) );
  OAI211_X1 U23550 ( .C1(n20580), .C2(n20558), .A(n20557), .B(n20556), .ZN(
        P1_U3130) );
  AOI22_X1 U23551 ( .A1(n20574), .A2(n20593), .B1(n20683), .B2(n9935), .ZN(
        n20560) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20684), .ZN(n20559) );
  OAI211_X1 U23553 ( .C1(n20580), .C2(n20561), .A(n20560), .B(n20559), .ZN(
        P1_U3131) );
  AOI22_X1 U23554 ( .A1(n20574), .A2(n20690), .B1(n20689), .B2(n9935), .ZN(
        n20563) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20638), .ZN(n20562) );
  OAI211_X1 U23556 ( .C1(n20580), .C2(n20564), .A(n20563), .B(n20562), .ZN(
        P1_U3132) );
  AOI22_X1 U23557 ( .A1(n20574), .A2(n20696), .B1(n20695), .B2(n9935), .ZN(
        n20566) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20642), .ZN(n20565) );
  OAI211_X1 U23559 ( .C1(n20580), .C2(n20567), .A(n20566), .B(n20565), .ZN(
        P1_U3133) );
  AOI22_X1 U23560 ( .A1(n20574), .A2(n20601), .B1(n20703), .B2(n9935), .ZN(
        n20569) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20704), .ZN(n20568) );
  OAI211_X1 U23562 ( .C1(n20580), .C2(n20570), .A(n20569), .B(n20568), .ZN(
        P1_U3134) );
  AOI22_X1 U23563 ( .A1(n20574), .A2(n20605), .B1(n20709), .B2(n9935), .ZN(
        n20572) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20710), .ZN(n20571) );
  OAI211_X1 U23565 ( .C1(n20580), .C2(n20573), .A(n20572), .B(n20571), .ZN(
        P1_U3135) );
  AOI22_X1 U23566 ( .A1(n20574), .A2(n20611), .B1(n20717), .B2(n9935), .ZN(
        n20578) );
  AOI22_X1 U23567 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20718), .ZN(n20577) );
  OAI211_X1 U23568 ( .C1(n20580), .C2(n20579), .A(n20578), .B(n20577), .ZN(
        P1_U3136) );
  NOR3_X2 U23569 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20581), .A3(
        n20659), .ZN(n20610) );
  INV_X1 U23570 ( .A(n20621), .ZN(n20658) );
  AOI21_X1 U23571 ( .B1(n20658), .B2(n20582), .A(n20610), .ZN(n20584) );
  NOR2_X1 U23572 ( .A1(n20659), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20585) );
  INV_X1 U23573 ( .A(n20585), .ZN(n20583) );
  OAI22_X1 U23574 ( .A1(n20584), .A2(n20669), .B1(n20583), .B2(n13230), .ZN(
        n20609) );
  AOI22_X1 U23575 ( .A1(n20663), .A2(n20610), .B1(n20662), .B2(n20609), .ZN(
        n20588) );
  OAI21_X1 U23576 ( .B1(n10331), .B2(n20585), .A(n20667), .ZN(n20612) );
  OR2_X1 U23577 ( .A1(n20666), .A2(n20586), .ZN(n20623) );
  AOI22_X1 U23578 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20612), .B1(
        n20652), .B2(n20672), .ZN(n20587) );
  OAI211_X1 U23579 ( .C1(n20675), .C2(n20615), .A(n20588), .B(n20587), .ZN(
        P1_U3137) );
  AOI22_X1 U23580 ( .A1(n20677), .A2(n20610), .B1(n20676), .B2(n20609), .ZN(
        n20591) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20612), .B1(
        n20652), .B2(n20589), .ZN(n20590) );
  OAI211_X1 U23582 ( .C1(n20592), .C2(n20615), .A(n20591), .B(n20590), .ZN(
        P1_U3138) );
  AOI22_X1 U23583 ( .A1(n20683), .A2(n20610), .B1(n20682), .B2(n20609), .ZN(
        n20595) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20612), .B1(
        n20652), .B2(n20593), .ZN(n20594) );
  OAI211_X1 U23585 ( .C1(n20596), .C2(n20615), .A(n20595), .B(n20594), .ZN(
        P1_U3139) );
  AOI22_X1 U23586 ( .A1(n20689), .A2(n20610), .B1(n20688), .B2(n20609), .ZN(
        n20598) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20612), .B1(
        n20652), .B2(n20690), .ZN(n20597) );
  OAI211_X1 U23588 ( .C1(n20693), .C2(n20615), .A(n20598), .B(n20597), .ZN(
        P1_U3140) );
  AOI22_X1 U23589 ( .A1(n20695), .A2(n20610), .B1(n20694), .B2(n20609), .ZN(
        n20600) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20612), .B1(
        n20652), .B2(n20696), .ZN(n20599) );
  OAI211_X1 U23591 ( .C1(n20701), .C2(n20615), .A(n20600), .B(n20599), .ZN(
        P1_U3141) );
  AOI22_X1 U23592 ( .A1(n20703), .A2(n20610), .B1(n20702), .B2(n20609), .ZN(
        n20603) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20612), .B1(
        n20652), .B2(n20601), .ZN(n20602) );
  OAI211_X1 U23594 ( .C1(n20604), .C2(n20615), .A(n20603), .B(n20602), .ZN(
        P1_U3142) );
  AOI22_X1 U23595 ( .A1(n20709), .A2(n20610), .B1(n20708), .B2(n20609), .ZN(
        n20607) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20612), .B1(
        n20652), .B2(n20605), .ZN(n20606) );
  OAI211_X1 U23597 ( .C1(n20608), .C2(n20615), .A(n20607), .B(n20606), .ZN(
        P1_U3143) );
  AOI22_X1 U23598 ( .A1(n20717), .A2(n20610), .B1(n20715), .B2(n20609), .ZN(
        n20614) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20612), .B1(
        n20652), .B2(n20611), .ZN(n20613) );
  OAI211_X1 U23600 ( .C1(n20616), .C2(n20615), .A(n20614), .B(n20613), .ZN(
        P1_U3144) );
  OAI33_X1 U23601 ( .A1(n20669), .A2(n13725), .A3(n20621), .B1(n20620), .B2(
        n20619), .B3(n20618), .ZN(n20650) );
  AOI22_X1 U23602 ( .A1(n20663), .A2(n20651), .B1(n20662), .B2(n9939), .ZN(
        n20632) );
  AOI21_X1 U23603 ( .B1(n20700), .B2(n20623), .A(n20622), .ZN(n20624) );
  AOI21_X1 U23604 ( .B1(n20658), .B2(n20625), .A(n20624), .ZN(n20626) );
  NOR2_X1 U23605 ( .A1(n20626), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20629) );
  OAI211_X1 U23606 ( .C1(n20651), .C2(n20629), .A(n20628), .B(n20627), .ZN(
        n20653) );
  AOI22_X1 U23607 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20653), .B1(
        n20652), .B2(n20630), .ZN(n20631) );
  OAI211_X1 U23608 ( .C1(n20633), .C2(n20700), .A(n20632), .B(n20631), .ZN(
        P1_U3145) );
  AOI22_X1 U23609 ( .A1(n20677), .A2(n20651), .B1(n9939), .B2(n20676), .ZN(
        n20635) );
  AOI22_X1 U23610 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20653), .B1(
        n20652), .B2(n20678), .ZN(n20634) );
  OAI211_X1 U23611 ( .C1(n20681), .C2(n20700), .A(n20635), .B(n20634), .ZN(
        P1_U3146) );
  AOI22_X1 U23612 ( .A1(n20683), .A2(n20651), .B1(n9939), .B2(n20682), .ZN(
        n20637) );
  AOI22_X1 U23613 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20653), .B1(
        n20652), .B2(n20684), .ZN(n20636) );
  OAI211_X1 U23614 ( .C1(n20687), .C2(n20700), .A(n20637), .B(n20636), .ZN(
        P1_U3147) );
  AOI22_X1 U23615 ( .A1(n20689), .A2(n20651), .B1(n9939), .B2(n20688), .ZN(
        n20640) );
  AOI22_X1 U23616 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20653), .B1(
        n20652), .B2(n20638), .ZN(n20639) );
  OAI211_X1 U23617 ( .C1(n20641), .C2(n20700), .A(n20640), .B(n20639), .ZN(
        P1_U3148) );
  AOI22_X1 U23618 ( .A1(n20695), .A2(n20651), .B1(n9939), .B2(n20694), .ZN(
        n20644) );
  AOI22_X1 U23619 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20653), .B1(
        n20652), .B2(n20642), .ZN(n20643) );
  OAI211_X1 U23620 ( .C1(n20645), .C2(n20700), .A(n20644), .B(n20643), .ZN(
        P1_U3149) );
  AOI22_X1 U23621 ( .A1(n20703), .A2(n20651), .B1(n9939), .B2(n20702), .ZN(
        n20647) );
  AOI22_X1 U23622 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20653), .B1(
        n20652), .B2(n20704), .ZN(n20646) );
  OAI211_X1 U23623 ( .C1(n20707), .C2(n20700), .A(n20647), .B(n20646), .ZN(
        P1_U3150) );
  AOI22_X1 U23624 ( .A1(n20709), .A2(n20651), .B1(n9939), .B2(n20708), .ZN(
        n20649) );
  AOI22_X1 U23625 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20653), .B1(
        n20652), .B2(n20710), .ZN(n20648) );
  OAI211_X1 U23626 ( .C1(n20713), .C2(n20700), .A(n20649), .B(n20648), .ZN(
        P1_U3151) );
  AOI22_X1 U23627 ( .A1(n20717), .A2(n20651), .B1(n9939), .B2(n20715), .ZN(
        n20655) );
  AOI22_X1 U23628 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20653), .B1(
        n20652), .B2(n20718), .ZN(n20654) );
  OAI211_X1 U23629 ( .C1(n20724), .C2(n20700), .A(n20655), .B(n20654), .ZN(
        P1_U3152) );
  NOR2_X1 U23630 ( .A1(n20656), .A2(n20659), .ZN(n20716) );
  AOI21_X1 U23631 ( .B1(n20658), .B2(n20657), .A(n20716), .ZN(n20664) );
  NOR2_X1 U23632 ( .A1(n20660), .A2(n20659), .ZN(n20670) );
  INV_X1 U23633 ( .A(n20670), .ZN(n20661) );
  OAI22_X1 U23634 ( .A1(n20664), .A2(n20669), .B1(n20661), .B2(n13230), .ZN(
        n20714) );
  AOI22_X1 U23635 ( .A1(n20663), .A2(n20716), .B1(n20662), .B2(n20714), .ZN(
        n20674) );
  OAI21_X1 U23636 ( .B1(n20666), .B2(n20665), .A(n20664), .ZN(n20668) );
  OAI221_X1 U23637 ( .B1(n20671), .B2(n20670), .C1(n20669), .C2(n20668), .A(
        n20667), .ZN(n20720) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20720), .B1(
        n20697), .B2(n20672), .ZN(n20673) );
  OAI211_X1 U23639 ( .C1(n20675), .C2(n20700), .A(n20674), .B(n20673), .ZN(
        P1_U3153) );
  AOI22_X1 U23640 ( .A1(n20677), .A2(n20716), .B1(n20676), .B2(n20714), .ZN(
        n20680) );
  INV_X1 U23641 ( .A(n20700), .ZN(n20719) );
  AOI22_X1 U23642 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20720), .B1(
        n20719), .B2(n20678), .ZN(n20679) );
  OAI211_X1 U23643 ( .C1(n20681), .C2(n20723), .A(n20680), .B(n20679), .ZN(
        P1_U3154) );
  AOI22_X1 U23644 ( .A1(n20683), .A2(n20716), .B1(n20682), .B2(n20714), .ZN(
        n20686) );
  AOI22_X1 U23645 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20720), .B1(
        n20719), .B2(n20684), .ZN(n20685) );
  OAI211_X1 U23646 ( .C1(n20687), .C2(n20723), .A(n20686), .B(n20685), .ZN(
        P1_U3155) );
  AOI22_X1 U23647 ( .A1(n20689), .A2(n20716), .B1(n20688), .B2(n20714), .ZN(
        n20692) );
  AOI22_X1 U23648 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20720), .B1(
        n20697), .B2(n20690), .ZN(n20691) );
  OAI211_X1 U23649 ( .C1(n20693), .C2(n20700), .A(n20692), .B(n20691), .ZN(
        P1_U3156) );
  AOI22_X1 U23650 ( .A1(n20695), .A2(n20716), .B1(n20694), .B2(n20714), .ZN(
        n20699) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20720), .B1(
        n20697), .B2(n20696), .ZN(n20698) );
  OAI211_X1 U23652 ( .C1(n20701), .C2(n20700), .A(n20699), .B(n20698), .ZN(
        P1_U3157) );
  AOI22_X1 U23653 ( .A1(n20703), .A2(n20716), .B1(n20702), .B2(n20714), .ZN(
        n20706) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20720), .B1(
        n20719), .B2(n20704), .ZN(n20705) );
  OAI211_X1 U23655 ( .C1(n20707), .C2(n20723), .A(n20706), .B(n20705), .ZN(
        P1_U3158) );
  AOI22_X1 U23656 ( .A1(n20709), .A2(n20716), .B1(n20708), .B2(n20714), .ZN(
        n20712) );
  AOI22_X1 U23657 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20720), .B1(
        n20719), .B2(n20710), .ZN(n20711) );
  OAI211_X1 U23658 ( .C1(n20713), .C2(n20723), .A(n20712), .B(n20711), .ZN(
        P1_U3159) );
  AOI22_X1 U23659 ( .A1(n20717), .A2(n20716), .B1(n20715), .B2(n20714), .ZN(
        n20722) );
  AOI22_X1 U23660 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20720), .B1(
        n20719), .B2(n20718), .ZN(n20721) );
  OAI211_X1 U23661 ( .C1(n20724), .C2(n20723), .A(n20722), .B(n20721), .ZN(
        P1_U3160) );
  OR2_X1 U23662 ( .A1(n20726), .A2(n20725), .ZN(P1_U3163) );
  AND2_X1 U23663 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20727), .ZN(
        P1_U3164) );
  AND2_X1 U23664 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20727), .ZN(
        P1_U3165) );
  AND2_X1 U23665 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20727), .ZN(
        P1_U3166) );
  AND2_X1 U23666 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20727), .ZN(
        P1_U3167) );
  AND2_X1 U23667 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20727), .ZN(
        P1_U3168) );
  AND2_X1 U23668 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20727), .ZN(
        P1_U3169) );
  AND2_X1 U23669 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20727), .ZN(
        P1_U3170) );
  AND2_X1 U23670 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20727), .ZN(
        P1_U3171) );
  AND2_X1 U23671 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20727), .ZN(
        P1_U3172) );
  AND2_X1 U23672 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20727), .ZN(
        P1_U3173) );
  AND2_X1 U23673 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20727), .ZN(
        P1_U3174) );
  AND2_X1 U23674 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20727), .ZN(
        P1_U3175) );
  AND2_X1 U23675 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20727), .ZN(
        P1_U3176) );
  AND2_X1 U23676 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20727), .ZN(
        P1_U3177) );
  AND2_X1 U23677 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20727), .ZN(
        P1_U3178) );
  AND2_X1 U23678 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20727), .ZN(
        P1_U3179) );
  AND2_X1 U23679 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20727), .ZN(
        P1_U3180) );
  AND2_X1 U23680 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20727), .ZN(
        P1_U3181) );
  AND2_X1 U23681 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20727), .ZN(
        P1_U3182) );
  AND2_X1 U23682 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20727), .ZN(
        P1_U3183) );
  AND2_X1 U23683 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20727), .ZN(
        P1_U3184) );
  AND2_X1 U23684 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20727), .ZN(
        P1_U3185) );
  AND2_X1 U23685 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20727), .ZN(P1_U3186) );
  AND2_X1 U23686 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20727), .ZN(P1_U3187) );
  AND2_X1 U23687 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20727), .ZN(P1_U3188) );
  AND2_X1 U23688 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20727), .ZN(P1_U3189) );
  AND2_X1 U23689 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20727), .ZN(P1_U3190) );
  AND2_X1 U23690 ( .A1(n20727), .A2(P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(P1_U3191) );
  AND2_X1 U23691 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20727), .ZN(P1_U3192) );
  AND2_X1 U23692 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20727), .ZN(P1_U3193) );
  AND2_X1 U23693 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20728), .ZN(n20742) );
  OAI21_X1 U23694 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20733), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20729) );
  AOI211_X1 U23695 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n20730), .B(
        n20729), .ZN(n20731) );
  OAI22_X1 U23696 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20742), .B1(n20795), 
        .B2(n20731), .ZN(P1_U3194) );
  AND2_X1 U23697 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20734) );
  INV_X1 U23698 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20736) );
  NOR2_X1 U23699 ( .A1(n20735), .A2(n20736), .ZN(n20732) );
  OAI22_X1 U23700 ( .A1(n20734), .A2(n20733), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20732), .ZN(n20741) );
  NOR3_X1 U23701 ( .A1(NA), .A2(n20735), .A3(n20828), .ZN(n20737) );
  OAI22_X1 U23702 ( .A1(n20738), .A2(n20737), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20736), .ZN(n20739) );
  OAI22_X1 U23703 ( .A1(n20742), .A2(n20741), .B1(n20740), .B2(n20739), .ZN(
        P1_U3196) );
  NOR2_X1 U23704 ( .A1(n20832), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20768) );
  INV_X1 U23705 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20743) );
  OAI222_X1 U23706 ( .A1(n20771), .A2(n19999), .B1(n20743), .B2(n20795), .C1(
        n13222), .C2(n20798), .ZN(P1_U3197) );
  AOI22_X1 U23707 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20832), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n20768), .ZN(n20744) );
  OAI21_X1 U23708 ( .B1(n19999), .B2(n20798), .A(n20744), .ZN(P1_U3198) );
  INV_X1 U23709 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20746) );
  OAI222_X1 U23710 ( .A1(n20798), .A2(n20746), .B1(n20745), .B2(n20795), .C1(
        n20747), .C2(n20771), .ZN(P1_U3199) );
  INV_X1 U23711 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21130) );
  OAI222_X1 U23712 ( .A1(n20771), .A2(n20749), .B1(n21130), .B2(n20795), .C1(
        n20747), .C2(n20798), .ZN(P1_U3200) );
  INV_X1 U23713 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20748) );
  OAI222_X1 U23714 ( .A1(n20798), .A2(n20749), .B1(n20748), .B2(n20795), .C1(
        n20751), .C2(n20771), .ZN(P1_U3201) );
  INV_X1 U23715 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20750) );
  OAI222_X1 U23716 ( .A1(n20798), .A2(n20751), .B1(n20750), .B2(n20795), .C1(
        n20752), .C2(n20771), .ZN(P1_U3202) );
  INV_X1 U23717 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21131) );
  OAI222_X1 U23718 ( .A1(n20798), .A2(n20752), .B1(n21131), .B2(n20795), .C1(
        n20982), .C2(n20771), .ZN(P1_U3203) );
  INV_X1 U23719 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20753) );
  OAI222_X1 U23720 ( .A1(n20771), .A2(n20755), .B1(n20753), .B2(n20795), .C1(
        n20982), .C2(n20798), .ZN(P1_U3204) );
  INV_X1 U23721 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20754) );
  OAI222_X1 U23722 ( .A1(n20798), .A2(n20755), .B1(n20754), .B2(n20795), .C1(
        n20756), .C2(n20771), .ZN(P1_U3205) );
  INV_X1 U23723 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20757) );
  OAI222_X1 U23724 ( .A1(n20771), .A2(n20758), .B1(n20757), .B2(n20795), .C1(
        n20756), .C2(n20798), .ZN(P1_U3206) );
  INV_X1 U23725 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20759) );
  OAI222_X1 U23726 ( .A1(n20771), .A2(n20760), .B1(n20759), .B2(n20795), .C1(
        n20758), .C2(n20798), .ZN(P1_U3207) );
  INV_X1 U23727 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20761) );
  OAI222_X1 U23728 ( .A1(n20771), .A2(n20763), .B1(n20761), .B2(n20795), .C1(
        n20760), .C2(n20798), .ZN(P1_U3208) );
  INV_X1 U23729 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20762) );
  OAI222_X1 U23730 ( .A1(n20798), .A2(n20763), .B1(n20762), .B2(n20795), .C1(
        n20765), .C2(n20771), .ZN(P1_U3209) );
  INV_X1 U23731 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20764) );
  OAI222_X1 U23732 ( .A1(n20798), .A2(n20765), .B1(n20764), .B2(n20795), .C1(
        n20767), .C2(n20771), .ZN(P1_U3210) );
  INV_X1 U23733 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20766) );
  OAI222_X1 U23734 ( .A1(n20798), .A2(n20767), .B1(n20766), .B2(n20795), .C1(
        n14715), .C2(n20771), .ZN(P1_U3211) );
  AOI22_X1 U23735 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20832), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20768), .ZN(n20769) );
  OAI21_X1 U23736 ( .B1(n14715), .B2(n20798), .A(n20769), .ZN(P1_U3212) );
  INV_X1 U23737 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n21094) );
  INV_X1 U23738 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20770) );
  OAI222_X1 U23739 ( .A1(n20771), .A2(n20773), .B1(n21094), .B2(n20795), .C1(
        n20770), .C2(n20798), .ZN(P1_U3213) );
  INV_X1 U23740 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20772) );
  OAI222_X1 U23741 ( .A1(n20798), .A2(n20773), .B1(n20772), .B2(n20795), .C1(
        n21098), .C2(n20771), .ZN(P1_U3214) );
  INV_X1 U23742 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20774) );
  OAI222_X1 U23743 ( .A1(n20798), .A2(n21098), .B1(n20774), .B2(n20795), .C1(
        n20776), .C2(n20771), .ZN(P1_U3215) );
  INV_X1 U23744 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20775) );
  OAI222_X1 U23745 ( .A1(n20798), .A2(n20776), .B1(n20775), .B2(n20795), .C1(
        n20948), .C2(n20771), .ZN(P1_U3216) );
  INV_X1 U23746 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20777) );
  OAI222_X1 U23747 ( .A1(n20798), .A2(n20948), .B1(n20777), .B2(n20795), .C1(
        n20779), .C2(n20771), .ZN(P1_U3217) );
  INV_X1 U23748 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20778) );
  OAI222_X1 U23749 ( .A1(n20798), .A2(n20779), .B1(n20778), .B2(n20795), .C1(
        n20781), .C2(n20771), .ZN(P1_U3218) );
  INV_X1 U23750 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20780) );
  OAI222_X1 U23751 ( .A1(n20798), .A2(n20781), .B1(n20780), .B2(n20795), .C1(
        n20783), .C2(n20771), .ZN(P1_U3219) );
  INV_X1 U23752 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20782) );
  INV_X1 U23753 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20785) );
  OAI222_X1 U23754 ( .A1(n20798), .A2(n20783), .B1(n20782), .B2(n20795), .C1(
        n20785), .C2(n20771), .ZN(P1_U3220) );
  INV_X1 U23755 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20784) );
  INV_X1 U23756 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20787) );
  OAI222_X1 U23757 ( .A1(n20798), .A2(n20785), .B1(n20784), .B2(n20795), .C1(
        n20787), .C2(n20771), .ZN(P1_U3221) );
  INV_X1 U23758 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20786) );
  OAI222_X1 U23759 ( .A1(n20798), .A2(n20787), .B1(n20786), .B2(n20795), .C1(
        n20789), .C2(n20771), .ZN(P1_U3222) );
  INV_X1 U23760 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20788) );
  INV_X1 U23761 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20791) );
  OAI222_X1 U23762 ( .A1(n20798), .A2(n20789), .B1(n20788), .B2(n20795), .C1(
        n20791), .C2(n20771), .ZN(P1_U3223) );
  INV_X1 U23763 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20790) );
  OAI222_X1 U23764 ( .A1(n20798), .A2(n20791), .B1(n20790), .B2(n20795), .C1(
        n20792), .C2(n20771), .ZN(P1_U3224) );
  INV_X1 U23765 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20793) );
  OAI222_X1 U23766 ( .A1(n20771), .A2(n20797), .B1(n20793), .B2(n20795), .C1(
        n20792), .C2(n20798), .ZN(P1_U3225) );
  INV_X1 U23767 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20796) );
  OAI222_X1 U23768 ( .A1(n20798), .A2(n20797), .B1(n20796), .B2(n20795), .C1(
        n20794), .C2(n20771), .ZN(P1_U3226) );
  MUX2_X1 U23769 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(P1_BE_N_REG_3__SCAN_IN), .S(n20832), .Z(P1_U3458) );
  MUX2_X1 U23770 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .B(P1_BE_N_REG_2__SCAN_IN), .S(n20832), .Z(P1_U3459) );
  MUX2_X1 U23771 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .B(P1_BE_N_REG_1__SCAN_IN), .S(n20832), .Z(P1_U3460) );
  OAI22_X1 U23772 ( .A1(n20832), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20795), .ZN(n20799) );
  INV_X1 U23773 ( .A(n20799), .ZN(P1_U3461) );
  OAI21_X1 U23774 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20803), .A(n20801), 
        .ZN(n20800) );
  INV_X1 U23775 ( .A(n20800), .ZN(P1_U3464) );
  INV_X1 U23776 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20802) );
  OAI21_X1 U23777 ( .B1(n20803), .B2(n20802), .A(n20801), .ZN(P1_U3465) );
  INV_X1 U23778 ( .A(n20804), .ZN(n20808) );
  OAI22_X1 U23779 ( .A1(n20808), .A2(n20807), .B1(n20806), .B2(n20805), .ZN(
        n20810) );
  MUX2_X1 U23780 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20810), .S(
        n20809), .Z(P1_U3469) );
  NOR2_X1 U23781 ( .A1(P1_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20812) );
  AOI211_X1 U23782 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(n21140), .A(n20812), 
        .B(n20811), .ZN(n20814) );
  OAI22_X1 U23783 ( .A1(n20815), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(n13222), .B2(n20816), .ZN(n20813) );
  NOR2_X1 U23784 ( .A1(n20814), .A2(n20813), .ZN(P1_U3481) );
  OAI22_X1 U23785 ( .A1(n20816), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n20815), 
        .B2(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20817) );
  INV_X1 U23786 ( .A(n20817), .ZN(P1_U3482) );
  INV_X1 U23787 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20818) );
  AOI22_X1 U23788 ( .A1(n20795), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20818), 
        .B2(n20832), .ZN(P1_U3483) );
  AND2_X1 U23789 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20828), .ZN(n20819) );
  OAI211_X1 U23790 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20821), .A(n20820), 
        .B(n20819), .ZN(n20822) );
  INV_X1 U23791 ( .A(n20822), .ZN(n20825) );
  OAI21_X1 U23792 ( .B1(n20825), .B2(n20824), .A(n20823), .ZN(n20831) );
  AOI211_X1 U23793 ( .C1(n20829), .C2(n20828), .A(n20827), .B(n20826), .ZN(
        n20830) );
  MUX2_X1 U23794 ( .A(n20831), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20830), 
        .Z(P1_U3485) );
  AOI22_X1 U23795 ( .A1(n20795), .A2(n20833), .B1(n21065), .B2(n20832), .ZN(
        P1_U3486) );
  OAI22_X1 U23796 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(keyinput3), .B1(
        P2_DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput36), .ZN(n20834) );
  AOI221_X1 U23797 ( .B1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B2(keyinput3), 
        .C1(keyinput36), .C2(P2_DATAWIDTH_REG_18__SCAN_IN), .A(n20834), .ZN(
        n20841) );
  OAI22_X1 U23798 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(keyinput7), .B1(
        P3_EAX_REG_16__SCAN_IN), .B2(keyinput75), .ZN(n20835) );
  AOI221_X1 U23799 ( .B1(P1_DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput7), .C1(
        keyinput75), .C2(P3_EAX_REG_16__SCAN_IN), .A(n20835), .ZN(n20840) );
  OAI22_X1 U23800 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(keyinput41), 
        .B1(keyinput102), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n20836) );
  AOI221_X1 U23801 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(keyinput41), 
        .C1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .C2(keyinput102), .A(n20836), 
        .ZN(n20839) );
  OAI22_X1 U23802 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(keyinput23), 
        .B1(keyinput53), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n20837) );
  AOI221_X1 U23803 ( .B1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput23), 
        .C1(P1_REIP_REG_21__SCAN_IN), .C2(keyinput53), .A(n20837), .ZN(n20838)
         );
  NAND4_X1 U23804 ( .A1(n20841), .A2(n20840), .A3(n20839), .A4(n20838), .ZN(
        n20869) );
  OAI22_X1 U23805 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(keyinput101), 
        .B1(keyinput103), .B2(READY2), .ZN(n20842) );
  AOI221_X1 U23806 ( .B1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B2(keyinput101), 
        .C1(READY2), .C2(keyinput103), .A(n20842), .ZN(n20849) );
  OAI22_X1 U23807 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(keyinput127), 
        .B1(keyinput91), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20843)
         );
  AOI221_X1 U23808 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput127), 
        .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(keyinput91), .A(n20843), 
        .ZN(n20848) );
  OAI22_X1 U23809 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(keyinput71), .B1(
        keyinput31), .B2(P3_EAX_REG_22__SCAN_IN), .ZN(n20844) );
  AOI221_X1 U23810 ( .B1(P3_EBX_REG_30__SCAN_IN), .B2(keyinput71), .C1(
        P3_EAX_REG_22__SCAN_IN), .C2(keyinput31), .A(n20844), .ZN(n20847) );
  OAI22_X1 U23811 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(keyinput61), .B1(
        keyinput54), .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20845) );
  AOI221_X1 U23812 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(keyinput61), .C1(
        P1_UWORD_REG_14__SCAN_IN), .C2(keyinput54), .A(n20845), .ZN(n20846) );
  NAND4_X1 U23813 ( .A1(n20849), .A2(n20848), .A3(n20847), .A4(n20846), .ZN(
        n20868) );
  OAI22_X1 U23814 ( .A1(BUF1_REG_24__SCAN_IN), .A2(keyinput72), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(keyinput118), .ZN(n20850) );
  AOI221_X1 U23815 ( .B1(BUF1_REG_24__SCAN_IN), .B2(keyinput72), .C1(
        keyinput118), .C2(P3_LWORD_REG_15__SCAN_IN), .A(n20850), .ZN(n20857)
         );
  OAI22_X1 U23816 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(keyinput49), 
        .B1(keyinput95), .B2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n20851)
         );
  AOI221_X1 U23817 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput49), 
        .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(keyinput95), .A(n20851), 
        .ZN(n20856) );
  OAI22_X1 U23818 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(keyinput37), 
        .B1(P3_ADDRESS_REG_3__SCAN_IN), .B2(keyinput44), .ZN(n20852) );
  AOI221_X1 U23819 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput37), 
        .C1(keyinput44), .C2(P3_ADDRESS_REG_3__SCAN_IN), .A(n20852), .ZN(
        n20855) );
  OAI22_X1 U23820 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(keyinput48), 
        .B1(P3_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput50), .ZN(n20853) );
  AOI221_X1 U23821 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(keyinput48), 
        .C1(keyinput50), .C2(P3_BYTEENABLE_REG_0__SCAN_IN), .A(n20853), .ZN(
        n20854) );
  NAND4_X1 U23822 ( .A1(n20857), .A2(n20856), .A3(n20855), .A4(n20854), .ZN(
        n20867) );
  OAI22_X1 U23823 ( .A1(P2_EBX_REG_3__SCAN_IN), .A2(keyinput84), .B1(
        keyinput86), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n20858) );
  AOI221_X1 U23824 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(keyinput84), .C1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .C2(keyinput86), .A(n20858), .ZN(
        n20865) );
  OAI22_X1 U23825 ( .A1(BUF2_REG_9__SCAN_IN), .A2(keyinput2), .B1(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput39), .ZN(n20859) );
  AOI221_X1 U23826 ( .B1(BUF2_REG_9__SCAN_IN), .B2(keyinput2), .C1(keyinput39), 
        .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(n20859), .ZN(n20864) );
  OAI22_X1 U23827 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(keyinput47), .B1(
        keyinput63), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n20860) );
  AOI221_X1 U23828 ( .B1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(keyinput47), 
        .C1(P2_EAX_REG_30__SCAN_IN), .C2(keyinput63), .A(n20860), .ZN(n20863)
         );
  OAI22_X1 U23829 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(keyinput14), .B1(
        DATAI_20_), .B2(keyinput76), .ZN(n20861) );
  AOI221_X1 U23830 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(keyinput14), .C1(
        keyinput76), .C2(DATAI_20_), .A(n20861), .ZN(n20862) );
  NAND4_X1 U23831 ( .A1(n20865), .A2(n20864), .A3(n20863), .A4(n20862), .ZN(
        n20866) );
  NOR4_X1 U23832 ( .A1(n20869), .A2(n20868), .A3(n20867), .A4(n20866), .ZN(
        n21218) );
  AOI22_X1 U23833 ( .A1(BUF2_REG_24__SCAN_IN), .A2(keyinput234), .B1(
        BUF2_REG_9__SCAN_IN), .B2(keyinput130), .ZN(n20870) );
  OAI221_X1 U23834 ( .B1(BUF2_REG_24__SCAN_IN), .B2(keyinput234), .C1(
        BUF2_REG_9__SCAN_IN), .C2(keyinput130), .A(n20870), .ZN(n20877) );
  AOI22_X1 U23835 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(keyinput230), 
        .B1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput254), .ZN(n20871) );
  OAI221_X1 U23836 ( .B1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(keyinput230), 
        .C1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .C2(keyinput254), .A(n20871), 
        .ZN(n20876) );
  AOI22_X1 U23837 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(keyinput210), 
        .B1(P1_ADDRESS_REG_18__SCAN_IN), .B2(keyinput166), .ZN(n20872) );
  OAI221_X1 U23838 ( .B1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput210), 
        .C1(P1_ADDRESS_REG_18__SCAN_IN), .C2(keyinput166), .A(n20872), .ZN(
        n20875) );
  AOI22_X1 U23839 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(keyinput225), .B1(
        P3_REIP_REG_18__SCAN_IN), .B2(keyinput186), .ZN(n20873) );
  OAI221_X1 U23840 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(keyinput225), .C1(
        P3_REIP_REG_18__SCAN_IN), .C2(keyinput186), .A(n20873), .ZN(n20874) );
  NOR4_X1 U23841 ( .A1(n20877), .A2(n20876), .A3(n20875), .A4(n20874), .ZN(
        n20905) );
  AOI22_X1 U23842 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(keyinput205), .B1(
        P2_INSTQUEUE_REG_8__4__SCAN_IN), .B2(keyinput137), .ZN(n20878) );
  OAI221_X1 U23843 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(keyinput205), .C1(
        P2_INSTQUEUE_REG_8__4__SCAN_IN), .C2(keyinput137), .A(n20878), .ZN(
        n20885) );
  AOI22_X1 U23844 ( .A1(P1_EAX_REG_17__SCAN_IN), .A2(keyinput226), .B1(
        P1_INSTQUEUE_REG_12__3__SCAN_IN), .B2(keyinput131), .ZN(n20879) );
  OAI221_X1 U23845 ( .B1(P1_EAX_REG_17__SCAN_IN), .B2(keyinput226), .C1(
        P1_INSTQUEUE_REG_12__3__SCAN_IN), .C2(keyinput131), .A(n20879), .ZN(
        n20884) );
  AOI22_X1 U23846 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(keyinput214), 
        .B1(P1_REIP_REG_11__SCAN_IN), .B2(keyinput189), .ZN(n20880) );
  OAI221_X1 U23847 ( .B1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(keyinput214), 
        .C1(P1_REIP_REG_11__SCAN_IN), .C2(keyinput189), .A(n20880), .ZN(n20883) );
  AOI22_X1 U23848 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(keyinput161), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(keyinput149), .ZN(n20881) );
  OAI221_X1 U23849 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(keyinput161), .C1(
        P1_ADDRESS_REG_3__SCAN_IN), .C2(keyinput149), .A(n20881), .ZN(n20882)
         );
  NOR4_X1 U23850 ( .A1(n20885), .A2(n20884), .A3(n20883), .A4(n20882), .ZN(
        n20904) );
  AOI22_X1 U23851 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(keyinput135), .B1(
        BUF1_REG_24__SCAN_IN), .B2(keyinput200), .ZN(n20886) );
  OAI221_X1 U23852 ( .B1(P1_DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput135), .C1(
        BUF1_REG_24__SCAN_IN), .C2(keyinput200), .A(n20886), .ZN(n20893) );
  AOI22_X1 U23853 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput202), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(keyinput245), .ZN(n20887) );
  OAI221_X1 U23854 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput202), .C1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .C2(keyinput245), .A(n20887), .ZN(
        n20892) );
  AOI22_X1 U23855 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(keyinput197), 
        .B1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput239), .ZN(n20888) );
  OAI221_X1 U23856 ( .B1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B2(keyinput197), 
        .C1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .C2(keyinput239), .A(n20888), 
        .ZN(n20891) );
  AOI22_X1 U23857 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(keyinput217), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(keyinput175), .ZN(n20889) );
  OAI221_X1 U23858 ( .B1(P1_ADDRESS_REG_16__SCAN_IN), .B2(keyinput217), .C1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .C2(keyinput175), .A(n20889), .ZN(
        n20890) );
  NOR4_X1 U23859 ( .A1(n20893), .A2(n20892), .A3(n20891), .A4(n20890), .ZN(
        n20903) );
  AOI22_X1 U23860 ( .A1(P3_ADDRESS_REG_3__SCAN_IN), .A2(keyinput172), .B1(
        P2_REIP_REG_0__SCAN_IN), .B2(keyinput129), .ZN(n20894) );
  OAI221_X1 U23861 ( .B1(P3_ADDRESS_REG_3__SCAN_IN), .B2(keyinput172), .C1(
        P2_REIP_REG_0__SCAN_IN), .C2(keyinput129), .A(n20894), .ZN(n20901) );
  AOI22_X1 U23862 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(keyinput227), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(keyinput191), .ZN(n20895) );
  OAI221_X1 U23863 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(keyinput227), .C1(
        P2_EAX_REG_30__SCAN_IN), .C2(keyinput191), .A(n20895), .ZN(n20900) );
  AOI22_X1 U23864 ( .A1(READY2), .A2(keyinput231), .B1(
        P1_INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput158), .ZN(n20896) );
  OAI221_X1 U23865 ( .B1(READY2), .B2(keyinput231), .C1(
        P1_INSTQUEUE_REG_7__5__SCAN_IN), .C2(keyinput158), .A(n20896), .ZN(
        n20899) );
  AOI22_X1 U23866 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(keyinput182), .B1(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .B2(keyinput132), .ZN(n20897) );
  OAI221_X1 U23867 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(keyinput182), .C1(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .C2(keyinput132), .A(n20897), .ZN(
        n20898) );
  NOR4_X1 U23868 ( .A1(n20901), .A2(n20900), .A3(n20899), .A4(n20898), .ZN(
        n20902) );
  NAND4_X1 U23869 ( .A1(n20905), .A2(n20904), .A3(n20903), .A4(n20902), .ZN(
        n21046) );
  AOI22_X1 U23870 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(keyinput165), 
        .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput192), .ZN(n20906)
         );
  OAI221_X1 U23871 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput165), 
        .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(keyinput192), .A(n20906), 
        .ZN(n20913) );
  AOI22_X1 U23872 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(keyinput142), .B1(
        P1_EAX_REG_0__SCAN_IN), .B2(keyinput183), .ZN(n20907) );
  OAI221_X1 U23873 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(keyinput142), .C1(
        P1_EAX_REG_0__SCAN_IN), .C2(keyinput183), .A(n20907), .ZN(n20912) );
  AOI22_X1 U23874 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(keyinput255), 
        .B1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(keyinput153), .ZN(n20908) );
  OAI221_X1 U23875 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput255), 
        .C1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .C2(keyinput153), .A(n20908), 
        .ZN(n20911) );
  AOI22_X1 U23876 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(keyinput213), .B1(
        P3_INSTQUEUE_REG_12__5__SCAN_IN), .B2(keyinput146), .ZN(n20909) );
  OAI221_X1 U23877 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(keyinput213), .C1(
        P3_INSTQUEUE_REG_12__5__SCAN_IN), .C2(keyinput146), .A(n20909), .ZN(
        n20910) );
  NOR4_X1 U23878 ( .A1(n20913), .A2(n20912), .A3(n20911), .A4(n20910), .ZN(
        n20941) );
  AOI22_X1 U23879 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(keyinput159), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(keyinput140), .ZN(n20914) );
  OAI221_X1 U23880 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(keyinput159), .C1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .C2(keyinput140), .A(n20914), .ZN(
        n20921) );
  AOI22_X1 U23881 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(keyinput168), 
        .B1(P2_EAX_REG_22__SCAN_IN), .B2(keyinput252), .ZN(n20915) );
  OAI221_X1 U23882 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput168), 
        .C1(P2_EAX_REG_22__SCAN_IN), .C2(keyinput252), .A(n20915), .ZN(n20920)
         );
  AOI22_X1 U23883 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput138), .B1(
        P2_INSTQUEUE_REG_10__2__SCAN_IN), .B2(keyinput253), .ZN(n20916) );
  OAI221_X1 U23884 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput138), 
        .C1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .C2(keyinput253), .A(n20916), 
        .ZN(n20919) );
  AOI22_X1 U23885 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(keyinput194), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput237), .ZN(n20917) );
  OAI221_X1 U23886 ( .B1(P3_DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput194), .C1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(keyinput237), .A(n20917), .ZN(
        n20918) );
  NOR4_X1 U23887 ( .A1(n20921), .A2(n20920), .A3(n20919), .A4(n20918), .ZN(
        n20940) );
  AOI22_X1 U23888 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(keyinput174), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput177), .ZN(n20922) );
  OAI221_X1 U23889 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(keyinput174), .C1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(keyinput177), .A(n20922), .ZN(
        n20929) );
  AOI22_X1 U23890 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(keyinput176), 
        .B1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B2(keyinput139), .ZN(n20923) );
  OAI221_X1 U23891 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(keyinput176), 
        .C1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .C2(keyinput139), .A(n20923), 
        .ZN(n20928) );
  AOI22_X1 U23892 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(keyinput154), 
        .B1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B2(keyinput198), .ZN(n20924) );
  OAI221_X1 U23893 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput154), 
        .C1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .C2(keyinput198), .A(n20924), 
        .ZN(n20927) );
  AOI22_X1 U23894 ( .A1(P3_BE_N_REG_3__SCAN_IN), .A2(keyinput220), .B1(
        P2_INSTQUEUE_REG_10__0__SCAN_IN), .B2(keyinput241), .ZN(n20925) );
  OAI221_X1 U23895 ( .B1(P3_BE_N_REG_3__SCAN_IN), .B2(keyinput220), .C1(
        P2_INSTQUEUE_REG_10__0__SCAN_IN), .C2(keyinput241), .A(n20925), .ZN(
        n20926) );
  NOR4_X1 U23896 ( .A1(n20929), .A2(n20928), .A3(n20927), .A4(n20926), .ZN(
        n20939) );
  AOI22_X1 U23897 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(keyinput195), .B1(
        P3_INSTQUEUE_REG_2__3__SCAN_IN), .B2(keyinput145), .ZN(n20930) );
  OAI221_X1 U23898 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(keyinput195), .C1(
        P3_INSTQUEUE_REG_2__3__SCAN_IN), .C2(keyinput145), .A(n20930), .ZN(
        n20937) );
  AOI22_X1 U23899 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(keyinput228), .B1(
        P1_INSTQUEUE_REG_10__3__SCAN_IN), .B2(keyinput243), .ZN(n20931) );
  OAI221_X1 U23900 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(keyinput228), .C1(
        P1_INSTQUEUE_REG_10__3__SCAN_IN), .C2(keyinput243), .A(n20931), .ZN(
        n20936) );
  AOI22_X1 U23901 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(keyinput203), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(keyinput141), .ZN(n20932) );
  OAI221_X1 U23902 ( .B1(P3_EAX_REG_16__SCAN_IN), .B2(keyinput203), .C1(
        P1_M_IO_N_REG_SCAN_IN), .C2(keyinput141), .A(n20932), .ZN(n20935) );
  AOI22_X1 U23903 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(keyinput157), .B1(
        P1_EBX_REG_15__SCAN_IN), .B2(keyinput238), .ZN(n20933) );
  OAI221_X1 U23904 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(keyinput157), .C1(
        P1_EBX_REG_15__SCAN_IN), .C2(keyinput238), .A(n20933), .ZN(n20934) );
  NOR4_X1 U23905 ( .A1(n20937), .A2(n20936), .A3(n20935), .A4(n20934), .ZN(
        n20938) );
  NAND4_X1 U23906 ( .A1(n20941), .A2(n20940), .A3(n20939), .A4(n20938), .ZN(
        n21045) );
  AOI22_X1 U23907 ( .A1(n21075), .A2(keyinput173), .B1(keyinput242), .B2(
        n21060), .ZN(n20942) );
  OAI221_X1 U23908 ( .B1(n21075), .B2(keyinput173), .C1(n21060), .C2(
        keyinput242), .A(n20942), .ZN(n20946) );
  AOI22_X1 U23909 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(keyinput162), 
        .B1(P1_REIP_REG_19__SCAN_IN), .B2(keyinput134), .ZN(n20943) );
  OAI221_X1 U23910 ( .B1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B2(keyinput162), 
        .C1(P1_REIP_REG_19__SCAN_IN), .C2(keyinput134), .A(n20943), .ZN(n20945) );
  XOR2_X1 U23911 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B(keyinput249), .Z(
        n20944) );
  OR3_X1 U23912 ( .A1(n20946), .A2(n20945), .A3(n20944), .ZN(n20953) );
  AOI22_X1 U23913 ( .A1(n20949), .A2(keyinput155), .B1(n20948), .B2(
        keyinput181), .ZN(n20947) );
  OAI221_X1 U23914 ( .B1(n20949), .B2(keyinput155), .C1(n20948), .C2(
        keyinput181), .A(n20947), .ZN(n20952) );
  XNOR2_X1 U23915 ( .A(n20950), .B(keyinput164), .ZN(n20951) );
  NOR3_X1 U23916 ( .A1(n20953), .A2(n20952), .A3(n20951), .ZN(n20991) );
  AOI22_X1 U23917 ( .A1(n21119), .A2(keyinput170), .B1(n20955), .B2(
        keyinput212), .ZN(n20954) );
  OAI221_X1 U23918 ( .B1(n21119), .B2(keyinput170), .C1(n20955), .C2(
        keyinput212), .A(n20954), .ZN(n20963) );
  AOI22_X1 U23919 ( .A1(n21141), .A2(keyinput160), .B1(n11419), .B2(
        keyinput185), .ZN(n20956) );
  OAI221_X1 U23920 ( .B1(n21141), .B2(keyinput160), .C1(n11419), .C2(
        keyinput185), .A(n20956), .ZN(n20962) );
  AOI22_X1 U23921 ( .A1(n21159), .A2(keyinput147), .B1(keyinput246), .B2(
        n20958), .ZN(n20957) );
  OAI221_X1 U23922 ( .B1(n21159), .B2(keyinput147), .C1(n20958), .C2(
        keyinput246), .A(n20957), .ZN(n20961) );
  INV_X1 U23923 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21092) );
  AOI22_X1 U23924 ( .A1(n21092), .A2(keyinput179), .B1(n21066), .B2(
        keyinput236), .ZN(n20959) );
  OAI221_X1 U23925 ( .B1(n21092), .B2(keyinput179), .C1(n21066), .C2(
        keyinput236), .A(n20959), .ZN(n20960) );
  NOR4_X1 U23926 ( .A1(n20963), .A2(n20962), .A3(n20961), .A4(n20960), .ZN(
        n20990) );
  INV_X1 U23927 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n21100) );
  AOI22_X1 U23928 ( .A1(n21100), .A2(keyinput224), .B1(n15039), .B2(
        keyinput247), .ZN(n20964) );
  OAI221_X1 U23929 ( .B1(n21100), .B2(keyinput224), .C1(n15039), .C2(
        keyinput247), .A(n20964), .ZN(n20975) );
  AOI22_X1 U23930 ( .A1(n20966), .A2(keyinput223), .B1(n21134), .B2(
        keyinput133), .ZN(n20965) );
  OAI221_X1 U23931 ( .B1(n20966), .B2(keyinput223), .C1(n21134), .C2(
        keyinput133), .A(n20965), .ZN(n20974) );
  AOI22_X1 U23932 ( .A1(n20968), .A2(keyinput144), .B1(n21112), .B2(
        keyinput190), .ZN(n20967) );
  OAI221_X1 U23933 ( .B1(n20968), .B2(keyinput144), .C1(n21112), .C2(
        keyinput190), .A(n20967), .ZN(n20973) );
  AOI22_X1 U23934 ( .A1(n20971), .A2(keyinput248), .B1(n20970), .B2(
        keyinput187), .ZN(n20969) );
  OAI221_X1 U23935 ( .B1(n20971), .B2(keyinput248), .C1(n20970), .C2(
        keyinput187), .A(n20969), .ZN(n20972) );
  NOR4_X1 U23936 ( .A1(n20975), .A2(n20974), .A3(n20973), .A4(n20972), .ZN(
        n20989) );
  INV_X1 U23937 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n20977) );
  AOI22_X1 U23938 ( .A1(n20978), .A2(keyinput233), .B1(n20977), .B2(
        keyinput229), .ZN(n20976) );
  OAI221_X1 U23939 ( .B1(n20978), .B2(keyinput233), .C1(n20977), .C2(
        keyinput229), .A(n20976), .ZN(n20987) );
  AOI22_X1 U23940 ( .A1(n21142), .A2(keyinput222), .B1(n20980), .B2(
        keyinput188), .ZN(n20979) );
  OAI221_X1 U23941 ( .B1(n21142), .B2(keyinput222), .C1(n20980), .C2(
        keyinput188), .A(n20979), .ZN(n20986) );
  AOI22_X1 U23942 ( .A1(n20982), .A2(keyinput218), .B1(n21131), .B2(
        keyinput235), .ZN(n20981) );
  OAI221_X1 U23943 ( .B1(n20982), .B2(keyinput218), .C1(n21131), .C2(
        keyinput235), .A(n20981), .ZN(n20985) );
  AOI22_X1 U23944 ( .A1(n21095), .A2(keyinput184), .B1(keyinput209), .B2(
        n21151), .ZN(n20983) );
  OAI221_X1 U23945 ( .B1(n21095), .B2(keyinput184), .C1(n21151), .C2(
        keyinput209), .A(n20983), .ZN(n20984) );
  NOR4_X1 U23946 ( .A1(n20987), .A2(n20986), .A3(n20985), .A4(n20984), .ZN(
        n20988) );
  NAND4_X1 U23947 ( .A1(n20991), .A2(n20990), .A3(n20989), .A4(n20988), .ZN(
        n21044) );
  AOI22_X1 U23948 ( .A1(n20994), .A2(keyinput219), .B1(keyinput216), .B2(
        n20993), .ZN(n20992) );
  OAI221_X1 U23949 ( .B1(n20994), .B2(keyinput219), .C1(n20993), .C2(
        keyinput216), .A(n20992), .ZN(n21003) );
  AOI22_X1 U23950 ( .A1(n21069), .A2(keyinput171), .B1(n12448), .B2(
        keyinput151), .ZN(n20995) );
  OAI221_X1 U23951 ( .B1(n21069), .B2(keyinput171), .C1(n12448), .C2(
        keyinput151), .A(n20995), .ZN(n21002) );
  AOI22_X1 U23952 ( .A1(n20997), .A2(keyinput208), .B1(n21164), .B2(
        keyinput150), .ZN(n20996) );
  OAI221_X1 U23953 ( .B1(n20997), .B2(keyinput208), .C1(n21164), .C2(
        keyinput150), .A(n20996), .ZN(n21001) );
  AOI22_X1 U23954 ( .A1(n21068), .A2(keyinput156), .B1(n20999), .B2(
        keyinput163), .ZN(n20998) );
  OAI221_X1 U23955 ( .B1(n21068), .B2(keyinput156), .C1(n20999), .C2(
        keyinput163), .A(n20998), .ZN(n21000) );
  NOR4_X1 U23956 ( .A1(n21003), .A2(n21002), .A3(n21001), .A4(n21000), .ZN(
        n21042) );
  AOI22_X1 U23957 ( .A1(n21158), .A2(keyinput207), .B1(n21097), .B2(
        keyinput250), .ZN(n21004) );
  OAI221_X1 U23958 ( .B1(n21158), .B2(keyinput207), .C1(n21097), .C2(
        keyinput250), .A(n21004), .ZN(n21014) );
  AOI22_X1 U23959 ( .A1(n21007), .A2(keyinput167), .B1(n21006), .B2(
        keyinput204), .ZN(n21005) );
  OAI221_X1 U23960 ( .B1(n21007), .B2(keyinput167), .C1(n21006), .C2(
        keyinput204), .A(n21005), .ZN(n21013) );
  INV_X1 U23961 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n21147) );
  INV_X1 U23962 ( .A(DATAI_10_), .ZN(n21009) );
  AOI22_X1 U23963 ( .A1(n21147), .A2(keyinput136), .B1(keyinput211), .B2(
        n21009), .ZN(n21008) );
  OAI221_X1 U23964 ( .B1(n21147), .B2(keyinput136), .C1(n21009), .C2(
        keyinput211), .A(n21008), .ZN(n21012) );
  AOI22_X1 U23965 ( .A1(n12416), .A2(keyinput232), .B1(n10963), .B2(
        keyinput143), .ZN(n21010) );
  OAI221_X1 U23966 ( .B1(n12416), .B2(keyinput232), .C1(n10963), .C2(
        keyinput143), .A(n21010), .ZN(n21011) );
  NOR4_X1 U23967 ( .A1(n21014), .A2(n21013), .A3(n21012), .A4(n21011), .ZN(
        n21041) );
  AOI22_X1 U23968 ( .A1(n13015), .A2(keyinput169), .B1(keyinput128), .B2(
        n21127), .ZN(n21015) );
  OAI221_X1 U23969 ( .B1(n13015), .B2(keyinput169), .C1(n21127), .C2(
        keyinput128), .A(n21015), .ZN(n21025) );
  AOI22_X1 U23970 ( .A1(n21150), .A2(keyinput244), .B1(n21017), .B2(
        keyinput221), .ZN(n21016) );
  OAI221_X1 U23971 ( .B1(n21150), .B2(keyinput244), .C1(n21017), .C2(
        keyinput221), .A(n21016), .ZN(n21024) );
  AOI22_X1 U23972 ( .A1(n21115), .A2(keyinput180), .B1(keyinput240), .B2(
        n21085), .ZN(n21018) );
  OAI221_X1 U23973 ( .B1(n21115), .B2(keyinput180), .C1(n21085), .C2(
        keyinput240), .A(n21018), .ZN(n21023) );
  AOI22_X1 U23974 ( .A1(n21021), .A2(keyinput199), .B1(keyinput178), .B2(
        n21020), .ZN(n21019) );
  OAI221_X1 U23975 ( .B1(n21021), .B2(keyinput199), .C1(n21020), .C2(
        keyinput178), .A(n21019), .ZN(n21022) );
  NOR4_X1 U23976 ( .A1(n21025), .A2(n21024), .A3(n21023), .A4(n21022), .ZN(
        n21040) );
  AOI22_X1 U23977 ( .A1(n21077), .A2(keyinput193), .B1(keyinput148), .B2(
        n21027), .ZN(n21026) );
  OAI221_X1 U23978 ( .B1(n21077), .B2(keyinput193), .C1(n21027), .C2(
        keyinput148), .A(n21026), .ZN(n21038) );
  AOI22_X1 U23979 ( .A1(n21029), .A2(keyinput251), .B1(keyinput152), .B2(
        n21168), .ZN(n21028) );
  OAI221_X1 U23980 ( .B1(n21029), .B2(keyinput251), .C1(n21168), .C2(
        keyinput152), .A(n21028), .ZN(n21037) );
  INV_X1 U23981 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n21063) );
  AOI22_X1 U23982 ( .A1(n21063), .A2(keyinput196), .B1(keyinput215), .B2(
        n21031), .ZN(n21030) );
  OAI221_X1 U23983 ( .B1(n21063), .B2(keyinput196), .C1(n21031), .C2(
        keyinput215), .A(n21030), .ZN(n21036) );
  AOI22_X1 U23984 ( .A1(n21034), .A2(keyinput206), .B1(keyinput201), .B2(
        n21033), .ZN(n21032) );
  OAI221_X1 U23985 ( .B1(n21034), .B2(keyinput206), .C1(n21033), .C2(
        keyinput201), .A(n21032), .ZN(n21035) );
  NOR4_X1 U23986 ( .A1(n21038), .A2(n21037), .A3(n21036), .A4(n21035), .ZN(
        n21039) );
  NAND4_X1 U23987 ( .A1(n21042), .A2(n21041), .A3(n21040), .A4(n21039), .ZN(
        n21043) );
  NOR4_X1 U23988 ( .A1(n21046), .A2(n21045), .A3(n21044), .A4(n21043), .ZN(
        n21179) );
  AOI22_X1 U23989 ( .A1(P1_EAX_REG_8__SCAN_IN), .A2(keyinput35), .B1(
        P1_EAX_REG_0__SCAN_IN), .B2(keyinput55), .ZN(n21047) );
  OAI221_X1 U23990 ( .B1(P1_EAX_REG_8__SCAN_IN), .B2(keyinput35), .C1(
        P1_EAX_REG_0__SCAN_IN), .C2(keyinput55), .A(n21047), .ZN(n21057) );
  AOI22_X1 U23991 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(keyinput38), .B1(
        n21049), .B2(keyinput18), .ZN(n21048) );
  OAI221_X1 U23992 ( .B1(P1_ADDRESS_REG_18__SCAN_IN), .B2(keyinput38), .C1(
        n21049), .C2(keyinput18), .A(n21048), .ZN(n21056) );
  AOI22_X1 U23993 ( .A1(n12416), .A2(keyinput104), .B1(n15039), .B2(
        keyinput119), .ZN(n21050) );
  OAI221_X1 U23994 ( .B1(n12416), .B2(keyinput104), .C1(n15039), .C2(
        keyinput119), .A(n21050), .ZN(n21055) );
  AOI22_X1 U23995 ( .A1(n21053), .A2(keyinput77), .B1(n21052), .B2(keyinput98), 
        .ZN(n21051) );
  OAI221_X1 U23996 ( .B1(n21053), .B2(keyinput77), .C1(n21052), .C2(keyinput98), .A(n21051), .ZN(n21054) );
  NOR4_X1 U23997 ( .A1(n21057), .A2(n21056), .A3(n21055), .A4(n21054), .ZN(
        n21108) );
  INV_X1 U23998 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n21059) );
  AOI22_X1 U23999 ( .A1(n21060), .A2(keyinput114), .B1(n21059), .B2(
        keyinput117), .ZN(n21058) );
  OAI221_X1 U24000 ( .B1(n21060), .B2(keyinput114), .C1(n21059), .C2(
        keyinput117), .A(n21058), .ZN(n21073) );
  AOI22_X1 U24001 ( .A1(n21063), .A2(keyinput68), .B1(keyinput82), .B2(n21062), 
        .ZN(n21061) );
  OAI221_X1 U24002 ( .B1(n21063), .B2(keyinput68), .C1(n21062), .C2(keyinput82), .A(n21061), .ZN(n21072) );
  AOI22_X1 U24003 ( .A1(n21066), .A2(keyinput108), .B1(keyinput13), .B2(n21065), .ZN(n21064) );
  OAI221_X1 U24004 ( .B1(n21066), .B2(keyinput108), .C1(n21065), .C2(
        keyinput13), .A(n21064), .ZN(n21071) );
  AOI22_X1 U24005 ( .A1(n21069), .A2(keyinput43), .B1(n21068), .B2(keyinput28), 
        .ZN(n21067) );
  OAI221_X1 U24006 ( .B1(n21069), .B2(keyinput43), .C1(n21068), .C2(keyinput28), .A(n21067), .ZN(n21070) );
  NOR4_X1 U24007 ( .A1(n21073), .A2(n21072), .A3(n21071), .A4(n21070), .ZN(
        n21107) );
  AOI22_X1 U24008 ( .A1(n21076), .A2(keyinput46), .B1(n21075), .B2(keyinput45), 
        .ZN(n21074) );
  OAI221_X1 U24009 ( .B1(n21076), .B2(keyinput46), .C1(n21075), .C2(keyinput45), .A(n21074), .ZN(n21080) );
  XOR2_X1 U24010 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B(keyinput121), .Z(
        n21079) );
  XNOR2_X1 U24011 ( .A(n21077), .B(keyinput65), .ZN(n21078) );
  OR3_X1 U24012 ( .A1(n21080), .A2(n21079), .A3(n21078), .ZN(n21089) );
  AOI22_X1 U24013 ( .A1(n21083), .A2(keyinput64), .B1(keyinput67), .B2(n21082), 
        .ZN(n21081) );
  OAI221_X1 U24014 ( .B1(n21083), .B2(keyinput64), .C1(n21082), .C2(keyinput67), .A(n21081), .ZN(n21088) );
  AOI22_X1 U24015 ( .A1(n21086), .A2(keyinput106), .B1(keyinput112), .B2(
        n21085), .ZN(n21084) );
  OAI221_X1 U24016 ( .B1(n21086), .B2(keyinput106), .C1(n21085), .C2(
        keyinput112), .A(n21084), .ZN(n21087) );
  NOR3_X1 U24017 ( .A1(n21089), .A2(n21088), .A3(n21087), .ZN(n21106) );
  AOI22_X1 U24018 ( .A1(n21092), .A2(keyinput51), .B1(n21091), .B2(keyinput70), 
        .ZN(n21090) );
  OAI221_X1 U24019 ( .B1(n21092), .B2(keyinput51), .C1(n21091), .C2(keyinput70), .A(n21090), .ZN(n21104) );
  AOI22_X1 U24020 ( .A1(n21095), .A2(keyinput56), .B1(n21094), .B2(keyinput89), 
        .ZN(n21093) );
  OAI221_X1 U24021 ( .B1(n21095), .B2(keyinput56), .C1(n21094), .C2(keyinput89), .A(n21093), .ZN(n21103) );
  AOI22_X1 U24022 ( .A1(n21098), .A2(keyinput6), .B1(n21097), .B2(keyinput122), 
        .ZN(n21096) );
  OAI221_X1 U24023 ( .B1(n21098), .B2(keyinput6), .C1(n21097), .C2(keyinput122), .A(n21096), .ZN(n21102) );
  AOI22_X1 U24024 ( .A1(n21100), .A2(keyinput96), .B1(n11419), .B2(keyinput57), 
        .ZN(n21099) );
  OAI221_X1 U24025 ( .B1(n21100), .B2(keyinput96), .C1(n11419), .C2(keyinput57), .A(n21099), .ZN(n21101) );
  NOR4_X1 U24026 ( .A1(n21104), .A2(n21103), .A3(n21102), .A4(n21101), .ZN(
        n21105) );
  NAND4_X1 U24027 ( .A1(n21108), .A2(n21107), .A3(n21106), .A4(n21105), .ZN(
        n21178) );
  AOI22_X1 U24028 ( .A1(n21110), .A2(keyinput92), .B1(n10963), .B2(keyinput15), 
        .ZN(n21109) );
  OAI221_X1 U24029 ( .B1(n21110), .B2(keyinput92), .C1(n10963), .C2(keyinput15), .A(n21109), .ZN(n21123) );
  AOI22_X1 U24030 ( .A1(n21113), .A2(keyinput100), .B1(n21112), .B2(keyinput62), .ZN(n21111) );
  OAI221_X1 U24031 ( .B1(n21113), .B2(keyinput100), .C1(n21112), .C2(
        keyinput62), .A(n21111), .ZN(n21122) );
  AOI22_X1 U24032 ( .A1(n21116), .A2(keyinput109), .B1(keyinput52), .B2(n21115), .ZN(n21114) );
  OAI221_X1 U24033 ( .B1(n21116), .B2(keyinput109), .C1(n21115), .C2(
        keyinput52), .A(n21114), .ZN(n21121) );
  AOI22_X1 U24034 ( .A1(n21119), .A2(keyinput42), .B1(n21118), .B2(keyinput124), .ZN(n21117) );
  OAI221_X1 U24035 ( .B1(n21119), .B2(keyinput42), .C1(n21118), .C2(
        keyinput124), .A(n21117), .ZN(n21120) );
  NOR4_X1 U24036 ( .A1(n21123), .A2(n21122), .A3(n21121), .A4(n21120), .ZN(
        n21176) );
  INV_X1 U24037 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n21125) );
  AOI22_X1 U24038 ( .A1(n11134), .A2(keyinput111), .B1(keyinput126), .B2(
        n21125), .ZN(n21124) );
  OAI221_X1 U24039 ( .B1(n11134), .B2(keyinput111), .C1(n21125), .C2(
        keyinput126), .A(n21124), .ZN(n21138) );
  AOI22_X1 U24040 ( .A1(n21128), .A2(keyinput34), .B1(keyinput0), .B2(n21127), 
        .ZN(n21126) );
  OAI221_X1 U24041 ( .B1(n21128), .B2(keyinput34), .C1(n21127), .C2(keyinput0), 
        .A(n21126), .ZN(n21137) );
  AOI22_X1 U24042 ( .A1(n21131), .A2(keyinput107), .B1(keyinput21), .B2(n21130), .ZN(n21129) );
  OAI221_X1 U24043 ( .B1(n21131), .B2(keyinput107), .C1(n21130), .C2(
        keyinput21), .A(n21129), .ZN(n21136) );
  AOI22_X1 U24044 ( .A1(n21134), .A2(keyinput5), .B1(n21133), .B2(keyinput40), 
        .ZN(n21132) );
  OAI221_X1 U24045 ( .B1(n21134), .B2(keyinput5), .C1(n21133), .C2(keyinput40), 
        .A(n21132), .ZN(n21135) );
  NOR4_X1 U24046 ( .A1(n21138), .A2(n21137), .A3(n21136), .A4(n21135), .ZN(
        n21175) );
  AOI22_X1 U24047 ( .A1(n21141), .A2(keyinput32), .B1(keyinput33), .B2(n21140), 
        .ZN(n21139) );
  OAI221_X1 U24048 ( .B1(n21141), .B2(keyinput32), .C1(n21140), .C2(keyinput33), .A(n21139), .ZN(n21144) );
  XNOR2_X1 U24049 ( .A(n21142), .B(keyinput94), .ZN(n21143) );
  NOR2_X1 U24050 ( .A1(n21144), .A2(n21143), .ZN(n21156) );
  AOI22_X1 U24051 ( .A1(n21147), .A2(keyinput8), .B1(keyinput74), .B2(n21146), 
        .ZN(n21145) );
  OAI221_X1 U24052 ( .B1(n21147), .B2(keyinput8), .C1(n21146), .C2(keyinput74), 
        .A(n21145), .ZN(n21148) );
  INV_X1 U24053 ( .A(n21148), .ZN(n21155) );
  AOI22_X1 U24054 ( .A1(n21151), .A2(keyinput81), .B1(n21150), .B2(keyinput116), .ZN(n21149) );
  OAI221_X1 U24055 ( .B1(n21151), .B2(keyinput81), .C1(n21150), .C2(
        keyinput116), .A(n21149), .ZN(n21152) );
  INV_X1 U24056 ( .A(n21152), .ZN(n21154) );
  XNOR2_X1 U24057 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B(keyinput9), .ZN(
        n21153) );
  AND4_X1 U24058 ( .A1(n21156), .A2(n21155), .A3(n21154), .A4(n21153), .ZN(
        n21174) );
  AOI22_X1 U24059 ( .A1(n21159), .A2(keyinput19), .B1(keyinput79), .B2(n21158), 
        .ZN(n21157) );
  OAI221_X1 U24060 ( .B1(n21159), .B2(keyinput19), .C1(n21158), .C2(keyinput79), .A(n21157), .ZN(n21172) );
  AOI22_X1 U24061 ( .A1(n21162), .A2(keyinput11), .B1(keyinput4), .B2(n21161), 
        .ZN(n21160) );
  OAI221_X1 U24062 ( .B1(n21162), .B2(keyinput11), .C1(n21161), .C2(keyinput4), 
        .A(n21160), .ZN(n21171) );
  INV_X1 U24063 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n21165) );
  AOI22_X1 U24064 ( .A1(n21165), .A2(keyinput69), .B1(keyinput22), .B2(n21164), 
        .ZN(n21163) );
  OAI221_X1 U24065 ( .B1(n21165), .B2(keyinput69), .C1(n21164), .C2(keyinput22), .A(n21163), .ZN(n21170) );
  AOI22_X1 U24066 ( .A1(n21168), .A2(keyinput24), .B1(keyinput58), .B2(n21167), 
        .ZN(n21166) );
  OAI221_X1 U24067 ( .B1(n21168), .B2(keyinput24), .C1(n21167), .C2(keyinput58), .A(n21166), .ZN(n21169) );
  NOR4_X1 U24068 ( .A1(n21172), .A2(n21171), .A3(n21170), .A4(n21169), .ZN(
        n21173) );
  NAND4_X1 U24069 ( .A1(n21176), .A2(n21175), .A3(n21174), .A4(n21173), .ZN(
        n21177) );
  NOR3_X1 U24070 ( .A1(n21179), .A2(n21178), .A3(n21177), .ZN(n21217) );
  OAI22_X1 U24071 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(keyinput85), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(keyinput87), .ZN(n21180) );
  AOI221_X1 U24072 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(keyinput85), .C1(
        keyinput87), .C2(P2_DATAO_REG_30__SCAN_IN), .A(n21180), .ZN(n21187) );
  OAI22_X1 U24073 ( .A1(P2_EBX_REG_9__SCAN_IN), .A2(keyinput105), .B1(
        keyinput88), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n21181) );
  AOI221_X1 U24074 ( .B1(P2_EBX_REG_9__SCAN_IN), .B2(keyinput105), .C1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(keyinput88), .A(n21181), .ZN(
        n21186) );
  OAI22_X1 U24075 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(keyinput26), 
        .B1(keyinput115), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n21182) );
  AOI221_X1 U24076 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput26), 
        .C1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .C2(keyinput115), .A(n21182), 
        .ZN(n21185) );
  OAI22_X1 U24077 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(keyinput97), .B1(
        keyinput10), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21183) );
  AOI221_X1 U24078 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(keyinput97), .C1(
        P2_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput10), .A(n21183), .ZN(
        n21184) );
  NAND4_X1 U24079 ( .A1(n21187), .A2(n21186), .A3(n21185), .A4(n21184), .ZN(
        n21215) );
  OAI22_X1 U24080 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(keyinput120), .B1(
        keyinput73), .B2(P3_EAX_REG_17__SCAN_IN), .ZN(n21188) );
  AOI221_X1 U24081 ( .B1(P2_DATAWIDTH_REG_22__SCAN_IN), .B2(keyinput120), .C1(
        P3_EAX_REG_17__SCAN_IN), .C2(keyinput73), .A(n21188), .ZN(n21195) );
  OAI22_X1 U24082 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(keyinput25), 
        .B1(keyinput99), .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n21189) );
  AOI221_X1 U24083 ( .B1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(keyinput25), 
        .C1(P1_DATAO_REG_30__SCAN_IN), .C2(keyinput99), .A(n21189), .ZN(n21194) );
  OAI22_X1 U24084 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(keyinput16), 
        .B1(P3_DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput66), .ZN(n21190) );
  AOI221_X1 U24085 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(keyinput16), 
        .C1(keyinput66), .C2(P3_DATAWIDTH_REG_10__SCAN_IN), .A(n21190), .ZN(
        n21193) );
  OAI22_X1 U24086 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(keyinput125), 
        .B1(keyinput1), .B2(P2_REIP_REG_0__SCAN_IN), .ZN(n21191) );
  AOI221_X1 U24087 ( .B1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B2(keyinput125), 
        .C1(P2_REIP_REG_0__SCAN_IN), .C2(keyinput1), .A(n21191), .ZN(n21192)
         );
  NAND4_X1 U24088 ( .A1(n21195), .A2(n21194), .A3(n21193), .A4(n21192), .ZN(
        n21214) );
  OAI22_X1 U24089 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(keyinput93), .B1(
        keyinput83), .B2(DATAI_10_), .ZN(n21196) );
  AOI221_X1 U24090 ( .B1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B2(keyinput93), 
        .C1(DATAI_10_), .C2(keyinput83), .A(n21196), .ZN(n21203) );
  OAI22_X1 U24091 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(keyinput17), .B1(
        keyinput20), .B2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n21197) );
  AOI221_X1 U24092 ( .B1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B2(keyinput17), 
        .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(keyinput20), .A(n21197), 
        .ZN(n21202) );
  OAI22_X1 U24093 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(keyinput123), 
        .B1(keyinput80), .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n21198) );
  AOI221_X1 U24094 ( .B1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B2(keyinput123), 
        .C1(P1_UWORD_REG_6__SCAN_IN), .C2(keyinput80), .A(n21198), .ZN(n21201)
         );
  OAI22_X1 U24095 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(keyinput78), 
        .B1(keyinput27), .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n21199) );
  AOI221_X1 U24096 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(keyinput78), 
        .C1(P3_DATAO_REG_16__SCAN_IN), .C2(keyinput27), .A(n21199), .ZN(n21200) );
  NAND4_X1 U24097 ( .A1(n21203), .A2(n21202), .A3(n21201), .A4(n21200), .ZN(
        n21213) );
  OAI22_X1 U24098 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(keyinput113), 
        .B1(P1_EBX_REG_15__SCAN_IN), .B2(keyinput110), .ZN(n21204) );
  AOI221_X1 U24099 ( .B1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B2(keyinput113), 
        .C1(keyinput110), .C2(P1_EBX_REG_15__SCAN_IN), .A(n21204), .ZN(n21211)
         );
  OAI22_X1 U24100 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(keyinput30), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(keyinput90), .ZN(n21205) );
  AOI221_X1 U24101 ( .B1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput30), 
        .C1(keyinput90), .C2(P1_REIP_REG_8__SCAN_IN), .A(n21205), .ZN(n21210)
         );
  OAI22_X1 U24102 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(keyinput12), .B1(
        keyinput29), .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n21206) );
  AOI221_X1 U24103 ( .B1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(keyinput12), 
        .C1(P1_UWORD_REG_11__SCAN_IN), .C2(keyinput29), .A(n21206), .ZN(n21209) );
  OAI22_X1 U24104 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(keyinput60), .B1(
        P3_INSTQUEUE_REG_5__4__SCAN_IN), .B2(keyinput59), .ZN(n21207) );
  AOI221_X1 U24105 ( .B1(P2_EBX_REG_31__SCAN_IN), .B2(keyinput60), .C1(
        keyinput59), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(n21207), .ZN(
        n21208) );
  NAND4_X1 U24106 ( .A1(n21211), .A2(n21210), .A3(n21209), .A4(n21208), .ZN(
        n21212) );
  NOR4_X1 U24107 ( .A1(n21215), .A2(n21214), .A3(n21213), .A4(n21212), .ZN(
        n21216) );
  NAND3_X1 U24108 ( .A1(n21218), .A2(n21217), .A3(n21216), .ZN(n21226) );
  AOI22_X1 U24109 ( .A1(n9790), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n21220), 
        .B2(n21219), .ZN(n21223) );
  NAND3_X1 U24110 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n9796), .A3(
        n21221), .ZN(n21222) );
  OAI211_X1 U24111 ( .C1(n21224), .C2(n10104), .A(n21223), .B(n21222), .ZN(
        n21225) );
  XNOR2_X1 U24112 ( .A(n21226), .B(n21225), .ZN(P3_U2845) );
  AND2_X1 U14927 ( .A1(n11832), .A2(n13318), .ZN(n11865) );
  INV_X1 U11350 ( .A(n12256), .ZN(n20199) );
  CLKBUF_X1 U11285 ( .A(n14382), .Z(n12099) );
  CLKBUF_X1 U12123 ( .A(n10188), .Z(n9925) );
  CLKBUF_X1 U12362 ( .A(n16202), .Z(n19236) );
  CLKBUF_X1 U12482 ( .A(n16390), .Z(n16404) );
endmodule

