

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, 
        P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, 
        P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, 
        P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, 
        P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, 
        P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, 
        P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, 
        P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, 
        P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, 
        P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, 
        P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN,
         P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN,
         P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN,
         P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN,
         P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN,
         P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN,
         P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN,
         P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN,
         P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN,
         P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN,
         P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
         P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
         P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
         P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
         P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
         P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
         P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN,
         P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN,
         P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
         P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN,
         P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
         P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
         P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
         P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
         P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
         P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
         P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
         P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
         P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
         P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
         P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
         P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
         P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
         P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
         P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
         P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
         P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
         P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
         P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
         P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
         P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
         P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
         P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
         P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN,
         P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN,
         P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
         P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN,
         P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN,
         P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN,
         P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN,
         P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN,
         P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN,
         P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN,
         P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN,
         P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN,
         P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN,
         P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN,
         P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN,
         P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN,
         P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
         P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN,
         P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN,
         P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
         P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
         P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
         P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
         P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
         P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
         P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
         P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
         P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
         P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
         P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
         P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
         P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
         P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN,
         P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN,
         P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
         P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN,
         P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN,
         P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN,
         P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN,
         P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN,
         P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN,
         P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN,
         P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN,
         P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN,
         P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN,
         P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN,
         P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN,
         P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN,
         P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN,
         P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN,
         P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN,
         P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN,
         P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7198, n7199, n7201, n7202, n7203, n7204, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16168;

  AND2_X1 U7298 ( .A1(n14558), .A2(n7701), .ZN(n14487) );
  INV_X1 U7299 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n15500) );
  NAND2_X1 U7300 ( .A1(n7836), .A2(n7837), .ZN(n13931) );
  INV_X1 U7301 ( .A(n13474), .ZN(n13509) );
  INV_X1 U7302 ( .A(n11879), .ZN(n10679) );
  CLKBUF_X2 U7303 ( .A(n8370), .Z(n12960) );
  INV_X1 U7304 ( .A(n9902), .ZN(n10176) );
  INV_X1 U7305 ( .A(n7213), .ZN(n10183) );
  CLKBUF_X3 U7306 ( .A(n9798), .Z(n7404) );
  BUF_X2 U7308 ( .A(n9334), .Z(n9624) );
  BUF_X1 U7309 ( .A(n9606), .Z(n7208) );
  INV_X1 U7310 ( .A(n11419), .ZN(n8048) );
  XNOR2_X1 U7311 ( .A(n9744), .B(n9741), .ZN(n12255) );
  XNOR2_X1 U7312 ( .A(n8868), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8872) );
  AND4_X1 U7313 ( .A1(n7622), .A2(n9992), .A3(n8231), .A4(n9735), .ZN(n7621)
         );
  INV_X1 U7315 ( .A(n16168), .ZN(n7198) );
  INV_X1 U7316 ( .A(n15500), .ZN(n7199) );
  INV_X1 U7317 ( .A(n7199), .ZN(P1_U3086) );
  INV_X1 U7318 ( .A(n7199), .ZN(n7201) );
  INV_X1 U7319 ( .A(n9958), .ZN(n14905) );
  NOR2_X1 U7320 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n9730) );
  INV_X1 U7321 ( .A(n13743), .ZN(n13755) );
  INV_X1 U7322 ( .A(n14229), .ZN(n14188) );
  NAND2_X1 U7323 ( .A1(n8872), .A2(n12578), .ZN(n9606) );
  INV_X1 U7324 ( .A(n9894), .ZN(n7210) );
  INV_X1 U7325 ( .A(n7421), .ZN(n10175) );
  OR2_X1 U7326 ( .A1(n15433), .A2(n15256), .ZN(n15242) );
  AND4_X1 U7327 ( .A1(n8231), .A2(n8221), .A3(n9992), .A4(n7946), .ZN(n7930)
         );
  XNOR2_X1 U7328 ( .A(n8702), .B(n8700), .ZN(n13316) );
  AND2_X1 U7329 ( .A1(n13783), .A2(n13782), .ZN(n13791) );
  NAND2_X1 U7330 ( .A1(n13931), .A2(n13930), .ZN(n13933) );
  NOR2_X1 U7332 ( .A1(n12575), .A2(n13588), .ZN(n11264) );
  NAND2_X1 U7333 ( .A1(n8305), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8307) );
  NAND2_X2 U7334 ( .A1(n14807), .A2(n10658), .ZN(n10662) );
  CLKBUF_X3 U7335 ( .A(n8917), .Z(n9621) );
  BUF_X1 U7336 ( .A(n9606), .Z(n7209) );
  INV_X1 U7337 ( .A(n14617), .ZN(n7690) );
  CLKBUF_X2 U7338 ( .A(n10697), .Z(n14633) );
  AOI21_X1 U7339 ( .B1(n7587), .B2(n9901), .A(n7586), .ZN(n7585) );
  INV_X1 U7340 ( .A(n7210), .ZN(n7212) );
  BUF_X1 U7341 ( .A(n9870), .Z(n12829) );
  AND3_X1 U7342 ( .A1(n8355), .A2(n8354), .A3(n8353), .ZN(n11624) );
  AND4_X1 U7343 ( .A1(n8486), .A2(n8485), .A3(n8484), .A4(n8483), .ZN(n12474)
         );
  AND4_X1 U7344 ( .A1(n8442), .A2(n8441), .A3(n8440), .A4(n8439), .ZN(n12234)
         );
  AOI21_X1 U7345 ( .B1(n16059), .B2(n14019), .A(n14018), .ZN(n14093) );
  NAND2_X1 U7346 ( .A1(n9476), .A2(n9475), .ZN(n14609) );
  NAND2_X1 U7347 ( .A1(n12591), .A2(n12590), .ZN(n15425) );
  NAND2_X1 U7348 ( .A1(n12601), .A2(n12600), .ZN(n15429) );
  NAND2_X1 U7349 ( .A1(n10119), .A2(n10118), .ZN(n12755) );
  BUF_X1 U7350 ( .A(n8953), .Z(n7216) );
  NOR2_X1 U7351 ( .A1(n14743), .A2(n7678), .ZN(n14820) );
  XNOR2_X1 U7352 ( .A(n7698), .B(n8870), .ZN(n12578) );
  INV_X4 U7353 ( .A(n8315), .ZN(n10252) );
  OR2_X1 U7354 ( .A1(n8966), .A2(n8965), .ZN(n7202) );
  NAND2_X2 U7355 ( .A1(n15728), .A2(n15727), .ZN(n15730) );
  NAND2_X2 U7356 ( .A1(n15001), .A2(n7481), .ZN(n14976) );
  NAND2_X1 U7357 ( .A1(n8372), .A2(n8371), .ZN(n8378) );
  NAND4_X2 U7358 ( .A1(n8255), .A2(n8252), .A3(n10718), .A4(n7522), .ZN(n8542)
         );
  AND3_X2 U7359 ( .A1(n7420), .A2(n8254), .A3(n8253), .ZN(n8255) );
  OAI21_X2 U7360 ( .B1(n11145), .B2(n11144), .A(n11143), .ZN(n11335) );
  OR2_X1 U7361 ( .A1(n10152), .A2(n10150), .ZN(n10155) );
  NAND2_X1 U7362 ( .A1(n9755), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9757) );
  XNOR2_X2 U7363 ( .A(n7682), .B(n14524), .ZN(n14739) );
  NAND2_X1 U7364 ( .A1(n8827), .A2(n8308), .ZN(n7203) );
  NAND2_X1 U7365 ( .A1(n8827), .A2(n8308), .ZN(n7204) );
  NAND2_X2 U7366 ( .A1(n8827), .A2(n8308), .ZN(n10628) );
  NAND2_X1 U7368 ( .A1(n10231), .A2(n15508), .ZN(n10267) );
  MUX2_X2 U7370 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8265), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8267) );
  NAND4_X2 U7371 ( .A1(n8981), .A2(n8980), .A3(n8979), .A4(n8978), .ZN(n14373)
         );
  OAI21_X2 U7372 ( .B1(n9274), .B2(n8012), .A(n9280), .ZN(n9298) );
  OAI21_X2 U7373 ( .B1(n9223), .B2(n9222), .A(n9225), .ZN(n9274) );
  AOI22_X1 U7374 ( .A1(n12924), .A2(n12923), .B1(n15190), .B2(n15413), .ZN(
        n15179) );
  XNOR2_X2 U7375 ( .A(n16031), .B(n15067), .ZN(n12737) );
  NAND4_X2 U7376 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n8898), .ZN(n14377)
         );
  NAND2_X2 U7377 ( .A1(n8092), .A2(n8094), .ZN(n8659) );
  NAND3_X2 U7378 ( .A1(n9748), .A2(n10200), .A3(n9747), .ZN(n10226) );
  NAND2_X2 U7379 ( .A1(n7954), .A2(n7953), .ZN(n15274) );
  INV_X1 U7380 ( .A(n8885), .ZN(n7206) );
  INV_X1 U7381 ( .A(n8885), .ZN(n9077) );
  INV_X4 U7382 ( .A(n9636), .ZN(n9634) );
  AOI21_X2 U7383 ( .B1(n13789), .B2(n13970), .A(n13788), .ZN(n13790) );
  OAI21_X2 U7384 ( .B1(n7253), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9783) );
  XOR2_X2 U7385 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(n15671), .Z(n15672) );
  INV_X2 U7386 ( .A(n7720), .ZN(n15671) );
  XNOR2_X2 U7387 ( .A(n8307), .B(n8306), .ZN(n8308) );
  NAND2_X4 U7389 ( .A1(n7256), .A2(n9876), .ZN(n15074) );
  AND3_X1 U7390 ( .A1(n9875), .A2(n9874), .A3(n9873), .ZN(n7256) );
  XNOR2_X2 U7391 ( .A(n7796), .B(n7795), .ZN(n10811) );
  NOR2_X4 U7392 ( .A1(n10771), .A2(n11375), .ZN(n8885) );
  INV_X4 U7393 ( .A(n9077), .ZN(n9615) );
  NOR2_X2 U7394 ( .A1(n12922), .A2(n12923), .ZN(n12921) );
  NAND2_X1 U7395 ( .A1(n11673), .A2(n11624), .ZN(n13393) );
  OAI222_X1 U7396 ( .A1(P3_U3151), .A2(n8827), .B1(n14158), .B2(n14157), .C1(
        n14156), .C2(n14155), .ZN(P3_U3267) );
  OAI21_X2 U7397 ( .B1(n8465), .B2(n8464), .A(n8466), .ZN(n8487) );
  INV_X1 U7398 ( .A(n7210), .ZN(n7211) );
  INV_X4 U7399 ( .A(n7210), .ZN(n7213) );
  AOI21_X2 U7400 ( .B1(n15075), .B2(n9887), .A(n9850), .ZN(n9851) );
  BUF_X2 U7401 ( .A(n10902), .Z(n15075) );
  AND2_X4 U7402 ( .A1(n10226), .A2(n11065), .ZN(n9798) );
  OAI21_X2 U7403 ( .B1(n8378), .B2(n8377), .A(n8379), .ZN(n8406) );
  OR2_X2 U7404 ( .A1(n15498), .A2(n15501), .ZN(n9769) );
  MUX2_X1 U7405 ( .A(n10729), .B(n10240), .S(n10628), .Z(n13380) );
  XNOR2_X2 U7406 ( .A(n8314), .B(n8313), .ZN(n10729) );
  INV_X1 U7407 ( .A(n14229), .ZN(n7214) );
  INV_X1 U7408 ( .A(n8315), .ZN(n7215) );
  INV_X2 U7409 ( .A(n8926), .ZN(n8315) );
  AOI22_X2 U7410 ( .A1(n13865), .A2(n12945), .B1(n14114), .B2(n13880), .ZN(
        n13856) );
  XNOR2_X2 U7411 ( .A(n8369), .B(n8368), .ZN(n10974) );
  AOI21_X2 U7412 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(n15699), .A(n15698), .ZN(
        n15826) );
  NAND2_X1 U7413 ( .A1(n13797), .A2(n13798), .ZN(n12985) );
  NAND2_X1 U7414 ( .A1(n13392), .A2(n13384), .ZN(n13386) );
  INV_X2 U7415 ( .A(n8790), .ZN(n8711) );
  INV_X1 U7416 ( .A(n12703), .ZN(n11440) );
  INV_X1 U7417 ( .A(n11270), .ZN(n12575) );
  CLKBUF_X2 U7418 ( .A(n8887), .Z(n11375) );
  BUF_X1 U7419 ( .A(n10267), .Z(n7421) );
  NAND2_X1 U7420 ( .A1(n7929), .A2(n7930), .ZN(n9755) );
  INV_X1 U7421 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7795) );
  NAND2_X1 U7422 ( .A1(n7588), .A2(n7590), .ZN(n12920) );
  NAND2_X1 U7423 ( .A1(n14915), .A2(n14916), .ZN(n14952) );
  OR3_X1 U7424 ( .A1(n7589), .A2(n12821), .A3(n7342), .ZN(n7588) );
  OR2_X1 U7425 ( .A1(n15418), .A2(n7499), .ZN(n15483) );
  OAI21_X1 U7426 ( .B1(n12985), .B2(n7844), .A(n7841), .ZN(n13553) );
  NAND2_X1 U7427 ( .A1(n12985), .A2(n7845), .ZN(n13783) );
  NAND2_X1 U7428 ( .A1(n15002), .A2(n15003), .ZN(n15001) );
  AOI21_X1 U7429 ( .B1(n12926), .B2(n16119), .A(n12925), .ZN(n12927) );
  AOI21_X1 U7430 ( .B1(n14238), .B2(n7399), .A(n7398), .ZN(n7397) );
  AND2_X1 U7431 ( .A1(n7969), .A2(n7968), .ZN(n15188) );
  NOR2_X1 U7432 ( .A1(n10217), .A2(n10218), .ZN(n14887) );
  NAND3_X1 U7433 ( .A1(n14333), .A2(n14198), .A3(n14334), .ZN(n14345) );
  NAND2_X1 U7434 ( .A1(n7684), .A2(n7246), .ZN(n14533) );
  NAND2_X1 U7435 ( .A1(n13507), .A2(n13506), .ZN(n13771) );
  NAND2_X1 U7436 ( .A1(n7733), .A2(n15445), .ZN(n15394) );
  NAND2_X1 U7437 ( .A1(n13497), .A2(n13496), .ZN(n13785) );
  XNOR2_X1 U7438 ( .A(n15159), .B(n7734), .ZN(n7733) );
  NAND2_X1 U7439 ( .A1(n7856), .A2(n7857), .ZN(n13853) );
  INV_X1 U7440 ( .A(n12950), .ZN(n14096) );
  NAND2_X1 U7441 ( .A1(n12955), .A2(n12956), .ZN(n13210) );
  NAND2_X1 U7442 ( .A1(n7464), .A2(n7355), .ZN(n8022) );
  NAND2_X1 U7443 ( .A1(n7454), .A2(n7453), .ZN(n7464) );
  NAND2_X1 U7444 ( .A1(n13842), .A2(n13841), .ZN(n13840) );
  NAND2_X1 U7445 ( .A1(n8767), .A2(n8766), .ZN(n12950) );
  XNOR2_X1 U7446 ( .A(n9567), .B(n9566), .ZN(n14851) );
  OR2_X1 U7447 ( .A1(n8780), .A2(n8779), .ZN(n12954) );
  INV_X1 U7448 ( .A(n15240), .ZN(n7217) );
  NAND2_X1 U7449 ( .A1(n9545), .A2(n9544), .ZN(n14563) );
  NAND2_X1 U7450 ( .A1(n7674), .A2(n14581), .ZN(n7673) );
  AND2_X1 U7451 ( .A1(n7718), .A2(n7715), .ZN(n15798) );
  NAND2_X1 U7452 ( .A1(n7383), .A2(n12872), .ZN(n16120) );
  NAND2_X1 U7453 ( .A1(n10070), .A2(n10069), .ZN(n12258) );
  AND2_X1 U7454 ( .A1(n8665), .A2(n8664), .ZN(n14118) );
  NAND2_X1 U7455 ( .A1(n15354), .A2(n15353), .ZN(n7928) );
  NAND2_X1 U7456 ( .A1(n15372), .A2(n12655), .ZN(n15354) );
  NAND2_X1 U7457 ( .A1(n7850), .A2(n7283), .ZN(n12369) );
  NAND2_X1 U7458 ( .A1(n12614), .A2(n12613), .ZN(n15433) );
  NAND2_X1 U7459 ( .A1(n11692), .A2(n11691), .ZN(n12284) );
  NAND2_X1 U7460 ( .A1(n12164), .A2(n13421), .ZN(n12242) );
  NAND2_X1 U7461 ( .A1(n8613), .A2(n8612), .ZN(n14123) );
  NAND2_X1 U7462 ( .A1(n9451), .A2(n9450), .ZN(n9471) );
  XNOR2_X1 U7463 ( .A(n9449), .B(n13105), .ZN(n9752) );
  NAND2_X1 U7464 ( .A1(n15748), .A2(n15749), .ZN(n15751) );
  NAND2_X2 U7465 ( .A1(n9228), .A2(n9227), .ZN(n16111) );
  NAND2_X1 U7466 ( .A1(n9284), .A2(n9283), .ZN(n14808) );
  NAND2_X1 U7467 ( .A1(n8606), .A2(n8605), .ZN(n8626) );
  CLKBUF_X1 U7468 ( .A(n9403), .Z(n7441) );
  NAND2_X1 U7469 ( .A1(n9118), .A2(n9117), .ZN(n12157) );
  OR2_X1 U7470 ( .A1(n12056), .A2(n12057), .ZN(n7759) );
  NAND2_X1 U7471 ( .A1(n8545), .A2(n8544), .ZN(n14141) );
  NAND2_X1 U7472 ( .A1(n10056), .A2(n10055), .ZN(n12744) );
  NAND2_X1 U7473 ( .A1(n7647), .A2(n9094), .ZN(n11795) );
  NAND2_X1 U7474 ( .A1(n11757), .A2(n11762), .ZN(n11758) );
  NAND2_X1 U7475 ( .A1(n10016), .A2(n10015), .ZN(n16019) );
  NAND2_X1 U7476 ( .A1(n7433), .A2(n7300), .ZN(n7432) );
  OR2_X1 U7477 ( .A1(n8559), .A2(n8569), .ZN(n8098) );
  CLKBUF_X1 U7478 ( .A(n8557), .Z(n7498) );
  NAND2_X1 U7479 ( .A1(n14937), .A2(n14938), .ZN(n14936) );
  AND2_X1 U7480 ( .A1(n12026), .A2(n11540), .ZN(n12057) );
  NAND2_X1 U7481 ( .A1(n8539), .A2(n8538), .ZN(n8558) );
  AND2_X1 U7482 ( .A1(n10986), .A2(n9892), .ZN(n14937) );
  XNOR2_X1 U7483 ( .A(n9135), .B(n9136), .ZN(n9110) );
  OAI21_X1 U7484 ( .B1(n9135), .B2(n8007), .A(n8004), .ZN(n9171) );
  NAND2_X1 U7485 ( .A1(n9044), .A2(n9043), .ZN(n11510) );
  OR2_X1 U7486 ( .A1(n8537), .A2(n8536), .ZN(n8539) );
  NAND2_X1 U7487 ( .A1(n9021), .A2(n9020), .ZN(n11400) );
  AND3_X1 U7488 ( .A1(n8496), .A2(n8495), .A3(n8494), .ZN(n12394) );
  OAI21_X1 U7489 ( .B1(n8941), .B2(n8940), .A(n8939), .ZN(n8966) );
  NAND2_X2 U7490 ( .A1(n11641), .A2(n13983), .ZN(n13966) );
  NAND2_X1 U7491 ( .A1(n7971), .A2(n7972), .ZN(n9087) );
  XNOR2_X1 U7492 ( .A(n13582), .B(n11955), .ZN(n13533) );
  NAND2_X1 U7493 ( .A1(n7736), .A2(n11440), .ZN(n11568) );
  INV_X2 U7494 ( .A(n16001), .ZN(n7218) );
  INV_X2 U7495 ( .A(n8614), .ZN(n7238) );
  NAND2_X1 U7496 ( .A1(n8991), .A2(n8990), .ZN(n9013) );
  AND2_X1 U7497 ( .A1(n8271), .A2(n8270), .ZN(n8359) );
  INV_X1 U7499 ( .A(n14153), .ZN(n8270) );
  NOR2_X1 U7500 ( .A1(n15691), .A2(n15690), .ZN(n15697) );
  BUF_X2 U7501 ( .A(n8943), .Z(n9608) );
  BUF_X2 U7502 ( .A(n8942), .Z(n9547) );
  OAI211_X1 U7503 ( .C1(n9621), .C2(n10259), .A(n8931), .B(n8930), .ZN(n10587)
         );
  NAND2_X1 U7504 ( .A1(n7203), .A2(n10252), .ZN(n8370) );
  AOI21_X1 U7505 ( .B1(n7242), .B2(n7974), .A(n7326), .ZN(n7972) );
  INV_X2 U7506 ( .A(n9621), .ZN(n9354) );
  INV_X2 U7507 ( .A(n9958), .ZN(n7219) );
  INV_X1 U7508 ( .A(n12676), .ZN(n11065) );
  NAND2_X1 U7509 ( .A1(n7227), .A2(n15513), .ZN(n12672) );
  OAI21_X1 U7510 ( .B1(n8406), .B2(n8405), .A(n8407), .ZN(n8422) );
  INV_X2 U7511 ( .A(n9893), .ZN(n12834) );
  AND2_X1 U7512 ( .A1(n11430), .A2(n10475), .ZN(n11734) );
  AND2_X1 U7513 ( .A1(n14860), .A2(n12578), .ZN(n9095) );
  INV_X1 U7514 ( .A(n11027), .ZN(n15513) );
  BUF_X2 U7515 ( .A(n9840), .Z(n12833) );
  NAND2_X1 U7516 ( .A1(n8905), .A2(n8315), .ZN(n8917) );
  NAND2_X1 U7517 ( .A1(n8857), .A2(n8856), .ZN(n11430) );
  CLKBUF_X2 U7518 ( .A(n8905), .Z(n10428) );
  NAND2_X1 U7519 ( .A1(n8048), .A2(n12838), .ZN(n12676) );
  XNOR2_X1 U7520 ( .A(n8297), .B(n8296), .ZN(n11426) );
  NOR2_X1 U7521 ( .A1(n15680), .A2(n15681), .ZN(n15693) );
  AND2_X2 U7522 ( .A1(n8860), .A2(n8859), .ZN(n12410) );
  NAND2_X1 U7523 ( .A1(n8859), .A2(n8855), .ZN(n8856) );
  XNOR2_X1 U7524 ( .A(n9786), .B(n9785), .ZN(n11027) );
  CLKBUF_X2 U7525 ( .A(n12885), .Z(n7228) );
  OR2_X1 U7526 ( .A1(n10267), .A2(n10331), .ZN(n7912) );
  AND2_X1 U7527 ( .A1(n12936), .A2(n9771), .ZN(n9872) );
  OR2_X1 U7528 ( .A1(n8858), .A2(n8853), .ZN(n8860) );
  NAND2_X1 U7529 ( .A1(n14852), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8868) );
  XNOR2_X1 U7530 ( .A(n15678), .B(n15677), .ZN(n15679) );
  XNOR2_X1 U7531 ( .A(n8862), .B(n8861), .ZN(n8887) );
  MUX2_X1 U7532 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8847), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n8851) );
  NAND2_X1 U7533 ( .A1(n9760), .A2(n9784), .ZN(n11419) );
  OR3_X1 U7534 ( .A1(n8879), .A2(n8880), .A3(n8878), .ZN(n8051) );
  NOR2_X1 U7535 ( .A1(n15673), .A2(n15674), .ZN(n15678) );
  INV_X1 U7536 ( .A(n8919), .ZN(n8923) );
  NAND2_X1 U7537 ( .A1(n8136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8862) );
  XNOR2_X1 U7538 ( .A(n9770), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9773) );
  NAND2_X2 U7539 ( .A1(n7215), .A2(P3_U3151), .ZN(n14155) );
  NAND2_X1 U7540 ( .A1(n9758), .A2(n9736), .ZN(n9784) );
  AND2_X1 U7541 ( .A1(n8881), .A2(n8232), .ZN(n8869) );
  AND2_X1 U7542 ( .A1(n8881), .A2(n8883), .ZN(n8879) );
  OAI21_X1 U7543 ( .B1(n8926), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n7440), .ZN(
        n8919) );
  OAI21_X1 U7544 ( .B1(n9755), .B2(n8208), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9770) );
  OAI211_X1 U7545 ( .C1(n8926), .C2(P2_DATAO_REG_0__SCAN_IN), .A(n7417), .B(
        SI_0_), .ZN(n8953) );
  NAND2_X1 U7546 ( .A1(n7621), .A2(n7932), .ZN(n9763) );
  NAND2_X2 U7547 ( .A1(n7641), .A2(n7643), .ZN(n8926) );
  AND2_X1 U7548 ( .A1(n7931), .A2(n7932), .ZN(n7929) );
  AND2_X1 U7549 ( .A1(n7932), .A2(n7622), .ZN(n9738) );
  NAND2_X1 U7550 ( .A1(n7645), .A2(n7644), .ZN(n7643) );
  NOR2_X1 U7551 ( .A1(n9729), .A2(n9737), .ZN(n7931) );
  AND2_X1 U7552 ( .A1(n8251), .A2(n8250), .ZN(n8252) );
  NAND3_X1 U7553 ( .A1(n7990), .A2(n7989), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7645) );
  AND4_X1 U7554 ( .A1(n9175), .A2(n8843), .A3(n8842), .A4(n8841), .ZN(n9193)
         );
  XNOR2_X1 U7555 ( .A(n15664), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n15662) );
  NOR2_X1 U7556 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n7468) );
  NOR2_X1 U7557 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n9731) );
  INV_X1 U7558 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10136) );
  NOR2_X1 U7559 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n8253) );
  NOR2_X1 U7560 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n8221) );
  NOR2_X1 U7561 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8259) );
  NOR2_X1 U7562 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8254) );
  NOR2_X1 U7563 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n7420) );
  NOR2_X1 U7564 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n8258) );
  INV_X1 U7565 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9734) );
  INV_X1 U7566 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9785) );
  INV_X4 U7567 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7568 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9736) );
  INV_X1 U7569 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9735) );
  NOR2_X1 U7570 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8250) );
  INV_X1 U7571 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9781) );
  NOR2_X1 U7572 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9726) );
  NOR2_X1 U7573 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9725) );
  INV_X1 U7574 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9782) );
  NOR2_X1 U7575 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n9732) );
  INV_X4 U7576 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  AND2_X1 U7577 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n8855) );
  NOR2_X2 U7578 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n10718) );
  INV_X1 U7579 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9197) );
  INV_X1 U7580 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7987) );
  INV_X1 U7581 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7989) );
  INV_X1 U7582 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7990) );
  NOR2_X1 U7583 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n9175) );
  NOR2_X1 U7584 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n8839) );
  NOR2_X1 U7585 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n8838) );
  XNOR2_X1 U7586 ( .A(n13746), .B(n7220), .ZN(n13756) );
  OR2_X1 U7587 ( .A1(n13739), .A2(n13738), .ZN(n7220) );
  OR2_X2 U7588 ( .A1(n8302), .A2(n7221), .ZN(n8268) );
  OR2_X1 U7589 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_29__SCAN_IN), .ZN(
        n7221) );
  OAI21_X1 U7590 ( .B1(n13940), .B2(n7328), .A(n8188), .ZN(n7222) );
  XNOR2_X1 U7591 ( .A(n13586), .B(n13380), .ZN(n7223) );
  OAI21_X1 U7592 ( .B1(n12520), .B2(n12519), .A(n12518), .ZN(n7224) );
  BUF_X1 U7593 ( .A(n13810), .Z(n7225) );
  CLKBUF_X1 U7594 ( .A(n13856), .Z(n7226) );
  NOR2_X1 U7595 ( .A1(n8302), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n8266) );
  OAI21_X1 U7596 ( .B1(n13940), .B2(n7328), .A(n8188), .ZN(n13913) );
  XNOR2_X1 U7597 ( .A(n13586), .B(n13380), .ZN(n11271) );
  OAI21_X1 U7598 ( .B1(n12520), .B2(n12519), .A(n12518), .ZN(n13990) );
  AND2_X1 U7599 ( .A1(n8271), .A2(n14153), .ZN(n8438) );
  INV_X1 U7600 ( .A(n8271), .ZN(n13213) );
  AOI21_X2 U7601 ( .B1(n15235), .B2(n7923), .A(n7460), .ZN(n15224) );
  NAND2_X1 U7602 ( .A1(n8903), .A2(n8836), .ZN(n8959) );
  OAI222_X1 U7603 ( .A1(P3_U3151), .A2(n14153), .B1(n14158), .B2(n14152), .C1(
        n14151), .C2(n14155), .ZN(P3_U3266) );
  AND2_X1 U7604 ( .A1(n13213), .A2(n14153), .ZN(n8362) );
  AND2_X1 U7605 ( .A1(n7795), .A2(n8256), .ZN(n7522) );
  XNOR2_X1 U7607 ( .A(n9783), .B(n9782), .ZN(n12885) );
  AOI21_X2 U7608 ( .B1(n13702), .B2(n13701), .A(n13700), .ZN(n13704) );
  NAND2_X1 U7609 ( .A1(n8359), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8320) );
  NAND3_X2 U7610 ( .A1(n8051), .A2(n8050), .A3(n8049), .ZN(n9707) );
  NAND2_X2 U7611 ( .A1(n13955), .A2(n12940), .ZN(n13940) );
  AND2_X1 U7612 ( .A1(n10679), .A2(n10775), .ZN(n10499) );
  NAND2_X2 U7613 ( .A1(n13957), .A2(n13956), .ZN(n13955) );
  NAND2_X1 U7614 ( .A1(n8872), .A2(n8871), .ZN(n9334) );
  NAND2_X1 U7615 ( .A1(n10231), .A2(n15508), .ZN(n7229) );
  NAND2_X1 U7616 ( .A1(n10231), .A2(n15508), .ZN(n7230) );
  INV_X4 U7617 ( .A(n12702), .ZN(n12826) );
  AND2_X1 U7618 ( .A1(n8270), .A2(n13213), .ZN(n8361) );
  NAND2_X2 U7619 ( .A1(n8976), .A2(n8975), .ZN(n11738) );
  BUF_X4 U7620 ( .A(n8359), .Z(n7231) );
  OAI222_X1 U7621 ( .A1(n13213), .A2(P3_U3151), .B1(n14155), .B2(n13372), .C1(
        n14158), .C2(n13212), .ZN(P3_U3265) );
  BUF_X4 U7622 ( .A(n7587), .Z(n7232) );
  INV_X1 U7623 ( .A(n9846), .ZN(n7587) );
  NOR2_X2 U7624 ( .A1(n11758), .A2(n11795), .ZN(n7709) );
  AOI21_X1 U7625 ( .B1(n13769), .B2(n13770), .A(n13768), .ZN(n14014) );
  AND2_X1 U7626 ( .A1(n8270), .A2(n13213), .ZN(n7233) );
  AOI21_X1 U7627 ( .B1(n9162), .B2(n9161), .A(n9160), .ZN(n9164) );
  OAI22_X2 U7628 ( .A1(n12128), .A2(n8074), .B1(n8075), .B2(n8073), .ZN(n12422) );
  XNOR2_X1 U7629 ( .A(n14377), .B(n11879), .ZN(n10492) );
  AND2_X1 U7630 ( .A1(n13213), .A2(n14153), .ZN(n7234) );
  AND2_X1 U7631 ( .A1(n10718), .A2(n7795), .ZN(n8351) );
  AOI21_X2 U7632 ( .B1(n13799), .B2(n12983), .A(n7507), .ZN(n13786) );
  OAI22_X2 U7633 ( .A1(n13810), .A2(n13811), .B1(n13827), .B2(n14104), .ZN(
        n13799) );
  NAND2_X1 U7634 ( .A1(n7229), .A2(n10252), .ZN(n7235) );
  NAND2_X1 U7635 ( .A1(n7229), .A2(n10252), .ZN(n7236) );
  NAND2_X1 U7636 ( .A1(n7230), .A2(n7215), .ZN(n9902) );
  OAI22_X2 U7637 ( .A1(n8022), .A2(n8021), .B1(n10159), .B2(n14993), .ZN(
        n15024) );
  INV_X1 U7638 ( .A(n8614), .ZN(n7237) );
  NOR2_X2 U7639 ( .A1(n15976), .A2(n16019), .ZN(n11972) );
  OR2_X2 U7640 ( .A1(n15975), .A2(n15992), .ZN(n15976) );
  OR2_X1 U7641 ( .A1(n12674), .A2(n15878), .ZN(n11005) );
  NOR2_X1 U7642 ( .A1(n7814), .A2(n14514), .ZN(n7813) );
  AND2_X1 U7643 ( .A1(n7690), .A2(n14513), .ZN(n7814) );
  NAND2_X1 U7644 ( .A1(n7991), .A2(n7995), .ZN(n9375) );
  OR2_X1 U7645 ( .A1(n14091), .A2(n13787), .ZN(n13507) );
  NAND2_X1 U7646 ( .A1(n11268), .A2(n13565), .ZN(n13474) );
  INV_X1 U7647 ( .A(n7962), .ZN(n7961) );
  OAI22_X1 U7648 ( .A1(n12879), .A2(n7968), .B1(n15057), .B2(n15198), .ZN(
        n7962) );
  OR2_X1 U7649 ( .A1(n15460), .A2(n15299), .ZN(n7742) );
  NAND2_X1 U7650 ( .A1(n10994), .A2(n12690), .ZN(n11200) );
  AND2_X1 U7651 ( .A1(n13494), .A2(n13575), .ZN(n7507) );
  INV_X1 U7652 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8200) );
  OAI22_X1 U7653 ( .A1(n14573), .A2(n9634), .B1(n14484), .B2(n9615), .ZN(n9533) );
  NAND2_X1 U7654 ( .A1(n7809), .A2(n7810), .ZN(n7674) );
  OAI21_X1 U7655 ( .B1(n15513), .B2(n7228), .A(n12672), .ZN(n12843) );
  INV_X1 U7656 ( .A(n8964), .ZN(n7450) );
  NAND2_X1 U7657 ( .A1(n7515), .A2(n7514), .ZN(n7513) );
  INV_X1 U7658 ( .A(n9189), .ZN(n7514) );
  NAND2_X1 U7659 ( .A1(n12748), .A2(n12750), .ZN(n8210) );
  AOI21_X1 U7660 ( .B1(n14723), .B2(n9615), .A(n9314), .ZN(n9320) );
  NAND2_X1 U7661 ( .A1(n9468), .A2(n7243), .ZN(n8125) );
  AOI21_X1 U7662 ( .B1(n8126), .B2(n8125), .A(n7311), .ZN(n8124) );
  NOR2_X1 U7663 ( .A1(n13544), .A2(n7313), .ZN(n8086) );
  AND2_X1 U7664 ( .A1(n7764), .A2(n7763), .ZN(n10880) );
  NAND2_X1 U7665 ( .A1(n7754), .A2(n7780), .ZN(n7749) );
  NAND2_X1 U7666 ( .A1(n7759), .A2(n7758), .ZN(n7757) );
  INV_X1 U7667 ( .A(n15840), .ZN(n7758) );
  AND2_X1 U7668 ( .A1(n13501), .A2(n12984), .ZN(n7845) );
  OR2_X1 U7669 ( .A1(n12949), .A2(n13827), .ZN(n13493) );
  OR2_X1 U7670 ( .A1(n14054), .A2(n13899), .ZN(n13378) );
  NAND2_X1 U7671 ( .A1(n11649), .A2(n11648), .ZN(n8181) );
  AOI21_X1 U7672 ( .B1(n8106), .B2(n8108), .A(n7377), .ZN(n8103) );
  INV_X1 U7673 ( .A(n8542), .ZN(n8182) );
  NAND2_X1 U7674 ( .A1(n10262), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8407) );
  INV_X1 U7675 ( .A(n12578), .ZN(n8871) );
  NAND2_X1 U7676 ( .A1(n14860), .A2(n8871), .ZN(n9629) );
  INV_X1 U7677 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8837) );
  NOR2_X1 U7678 ( .A1(n15282), .A2(n7958), .ZN(n7957) );
  INV_X1 U7679 ( .A(n12610), .ZN(n7958) );
  NAND2_X1 U7680 ( .A1(n9579), .A2(n9559), .ZN(n9619) );
  NAND2_X1 U7681 ( .A1(n9519), .A2(n9518), .ZN(n9537) );
  OR2_X1 U7682 ( .A1(n9517), .A2(n9516), .ZN(n9519) );
  NAND2_X1 U7683 ( .A1(n9404), .A2(SI_21_), .ZN(n9424) );
  XNOR2_X1 U7684 ( .A(n9375), .B(SI_18_), .ZN(n9345) );
  NAND2_X1 U7685 ( .A1(n7330), .A2(n9278), .ZN(n8012) );
  AOI21_X1 U7686 ( .B1(n9279), .B2(n9278), .A(n9277), .ZN(n9280) );
  XNOR2_X1 U7687 ( .A(n9038), .B(SI_6_), .ZN(n9035) );
  AOI21_X1 U7688 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15738), .A(n15737), .ZN(
        n15745) );
  NOR2_X1 U7689 ( .A1(n15736), .A2(n15735), .ZN(n15737) );
  AND2_X1 U7690 ( .A1(n13248), .A2(n8149), .ZN(n8148) );
  OR2_X1 U7691 ( .A1(n13324), .A2(n8150), .ZN(n8149) );
  NAND2_X1 U7692 ( .A1(n7568), .A2(n7567), .ZN(n7566) );
  AND2_X1 U7693 ( .A1(n8335), .A2(n8333), .ZN(n7471) );
  OR2_X1 U7694 ( .A1(n8327), .A2(n10280), .ZN(n8334) );
  NAND2_X1 U7695 ( .A1(n7521), .A2(n13231), .ZN(n13341) );
  NAND2_X1 U7696 ( .A1(n13229), .A2(n13230), .ZN(n7521) );
  NAND2_X1 U7697 ( .A1(n13517), .A2(n13551), .ZN(n8084) );
  BUF_X4 U7699 ( .A(n8361), .Z(n13365) );
  NOR2_X1 U7700 ( .A1(n7779), .A2(n10977), .ZN(n7778) );
  NAND2_X1 U7701 ( .A1(n7463), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7467) );
  NAND2_X1 U7702 ( .A1(n13754), .A2(n13755), .ZN(n7555) );
  NAND2_X1 U7703 ( .A1(n13784), .A2(n8187), .ZN(n13770) );
  AND2_X1 U7704 ( .A1(n13771), .A2(n12952), .ZN(n8187) );
  NAND2_X1 U7705 ( .A1(n13786), .A2(n13785), .ZN(n13784) );
  AND2_X1 U7706 ( .A1(n12980), .A2(n13843), .ZN(n7493) );
  AOI21_X1 U7707 ( .B1(n7239), .B2(n7863), .A(n7308), .ZN(n7857) );
  AOI21_X1 U7708 ( .B1(n7864), .B2(n7862), .A(n7861), .ZN(n7860) );
  INV_X1 U7709 ( .A(n8237), .ZN(n7862) );
  INV_X1 U7710 ( .A(n13476), .ZN(n7861) );
  OR2_X1 U7711 ( .A1(n14054), .A2(n13924), .ZN(n12942) );
  NAND2_X1 U7712 ( .A1(n13938), .A2(n12941), .ZN(n13920) );
  AOI21_X1 U7713 ( .B1(n7838), .B2(n7840), .A(n7365), .ZN(n7837) );
  OR2_X1 U7714 ( .A1(n14141), .A2(n13237), .ZN(n12937) );
  INV_X1 U7715 ( .A(n8327), .ZN(n13370) );
  INV_X1 U7716 ( .A(n12960), .ZN(n8647) );
  OR2_X1 U7717 ( .A1(n8327), .A2(n10254), .ZN(n8311) );
  AND2_X1 U7718 ( .A1(n8282), .A2(n12349), .ZN(n8286) );
  AND2_X2 U7719 ( .A1(n8182), .A2(n7846), .ZN(n8262) );
  AND2_X1 U7720 ( .A1(n7259), .A2(n7847), .ZN(n7846) );
  AND2_X1 U7721 ( .A1(n7849), .A2(n8805), .ZN(n7847) );
  OAI21_X1 U7722 ( .B1(n8487), .B2(n8488), .A(n8490), .ZN(n8508) );
  OR2_X1 U7723 ( .A1(n9332), .A2(n12340), .ZN(n9359) );
  NOR2_X1 U7724 ( .A1(n7909), .A2(n7901), .ZN(n7900) );
  OR2_X1 U7725 ( .A1(n14243), .A2(n14180), .ZN(n7909) );
  OR2_X1 U7726 ( .A1(n14185), .A2(n14184), .ZN(n14186) );
  NAND2_X1 U7727 ( .A1(n7403), .A2(n7402), .ZN(n7437) );
  NAND2_X1 U7728 ( .A1(n12280), .A2(n12181), .ZN(n7402) );
  INV_X1 U7729 ( .A(n12180), .ZN(n7403) );
  INV_X1 U7730 ( .A(n9608), .ZN(n9626) );
  NOR2_X1 U7731 ( .A1(n14461), .A2(n7700), .ZN(n7699) );
  INV_X1 U7732 ( .A(n7701), .ZN(n7700) );
  INV_X1 U7733 ( .A(n14555), .ZN(n7684) );
  INV_X1 U7734 ( .A(n8063), .ZN(n8060) );
  INV_X1 U7735 ( .A(n7809), .ZN(n7394) );
  INV_X1 U7736 ( .A(n7673), .ZN(n7395) );
  NAND2_X1 U7737 ( .A1(n14593), .A2(n14573), .ZN(n14570) );
  NAND2_X1 U7738 ( .A1(n14511), .A2(n14510), .ZN(n14614) );
  NOR2_X1 U7739 ( .A1(n7655), .A2(n14508), .ZN(n7654) );
  OR2_X1 U7740 ( .A1(n14784), .A2(n14507), .ZN(n8072) );
  AOI21_X1 U7741 ( .B1(n7661), .B2(n7658), .A(n7322), .ZN(n7657) );
  INV_X1 U7742 ( .A(n14506), .ZN(n7658) );
  OAI21_X2 U7743 ( .B1(n14659), .B2(n14473), .A(n14475), .ZN(n14645) );
  AND2_X1 U7744 ( .A1(n7650), .A2(n7335), .ZN(n7648) );
  OR2_X1 U7745 ( .A1(n14711), .A2(n7653), .ZN(n7649) );
  INV_X1 U7746 ( .A(n14498), .ZN(n7653) );
  OR2_X1 U7747 ( .A1(n7705), .A2(n14723), .ZN(n7704) );
  OR2_X1 U7748 ( .A1(n11722), .A2(n7820), .ZN(n7817) );
  NAND2_X1 U7749 ( .A1(n11398), .A2(n11397), .ZN(n11512) );
  NAND2_X1 U7750 ( .A1(n10483), .A2(n12414), .ZN(n14807) );
  NAND4_X1 U7751 ( .A1(n11707), .A2(n11706), .A3(n7820), .A4(n11861), .ZN(
        n8057) );
  AND2_X1 U7752 ( .A1(n12451), .A2(n10462), .ZN(n15519) );
  NAND2_X1 U7753 ( .A1(n9697), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9705) );
  OR2_X1 U7754 ( .A1(n9696), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9697) );
  NAND2_X1 U7755 ( .A1(n9752), .A2(n9426), .ZN(n9451) );
  NAND2_X1 U7756 ( .A1(n9975), .A2(n9974), .ZN(n12725) );
  INV_X1 U7757 ( .A(n8023), .ZN(n7418) );
  OAI21_X1 U7758 ( .B1(n8026), .B2(n8024), .A(n14894), .ZN(n8023) );
  NAND2_X1 U7759 ( .A1(n9862), .A2(n9861), .ZN(n10447) );
  NAND2_X1 U7760 ( .A1(n12843), .A2(n11419), .ZN(n7619) );
  AND4_X1 U7761 ( .A1(n12647), .A2(n12646), .A3(n12645), .A4(n12644), .ZN(
        n14962) );
  NAND2_X1 U7762 ( .A1(n9871), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U7763 ( .A1(n12841), .A2(n12840), .ZN(n15153) );
  NOR2_X1 U7764 ( .A1(n12921), .A2(n7569), .ZN(n12666) );
  NOR2_X1 U7765 ( .A1(n15413), .A2(n15056), .ZN(n7569) );
  XNOR2_X1 U7766 ( .A(n15413), .B(n15056), .ZN(n12923) );
  INV_X1 U7767 ( .A(n15057), .ZN(n14918) );
  AND2_X1 U7768 ( .A1(n15433), .A2(n12615), .ZN(n7460) );
  NAND2_X1 U7769 ( .A1(n7741), .A2(n15439), .ZN(n7740) );
  INV_X1 U7770 ( .A(n7742), .ZN(n7741) );
  OAI21_X1 U7771 ( .B1(n15268), .B2(n12663), .A(n12662), .ZN(n15251) );
  OR2_X1 U7772 ( .A1(n15444), .A2(n15259), .ZN(n12662) );
  NAND2_X1 U7773 ( .A1(n15452), .A2(n15061), .ZN(n7959) );
  OAI22_X1 U7774 ( .A1(n7928), .A2(n7572), .B1(n7573), .B2(n12659), .ZN(n15308) );
  NAND2_X1 U7775 ( .A1(n7576), .A2(n12658), .ZN(n7572) );
  INV_X1 U7776 ( .A(n7574), .ZN(n7573) );
  NAND2_X1 U7777 ( .A1(n12302), .A2(n7935), .ZN(n12386) );
  AND2_X1 U7778 ( .A1(n12303), .A2(n12301), .ZN(n7935) );
  NAND2_X1 U7779 ( .A1(n11993), .A2(n12868), .ZN(n7571) );
  NAND2_X1 U7780 ( .A1(n11915), .A2(n11914), .ZN(n7934) );
  NAND2_X1 U7781 ( .A1(n11355), .A2(n11199), .ZN(n11352) );
  OAI21_X1 U7782 ( .B1(n12683), .B2(n7916), .A(n12673), .ZN(n7915) );
  INV_X1 U7783 ( .A(n10908), .ZN(n7916) );
  NAND2_X1 U7784 ( .A1(n10901), .A2(n12675), .ZN(n16119) );
  NAND2_X1 U7785 ( .A1(n15791), .A2(n7276), .ZN(n7718) );
  AND2_X1 U7786 ( .A1(n15813), .A2(n15812), .ZN(n15816) );
  NAND2_X1 U7787 ( .A1(n8804), .A2(n8803), .ZN(n9751) );
  XNOR2_X1 U7788 ( .A(n14187), .B(n8241), .ZN(n14209) );
  NAND2_X1 U7789 ( .A1(n9641), .A2(n9642), .ZN(n8130) );
  NAND2_X1 U7790 ( .A1(n14540), .A2(n14539), .ZN(n14743) );
  NAND2_X1 U7791 ( .A1(n7806), .A2(n7807), .ZN(n14536) );
  NAND2_X1 U7792 ( .A1(n14566), .A2(n14485), .ZN(n14553) );
  INV_X1 U7793 ( .A(n15058), .ZN(n15191) );
  INV_X1 U7794 ( .A(n7228), .ZN(n15150) );
  NOR2_X1 U7795 ( .A1(n15807), .A2(n15808), .ZN(n15822) );
  NAND2_X1 U7796 ( .A1(n8985), .A2(n7262), .ZN(n8134) );
  INV_X1 U7797 ( .A(n9082), .ZN(n7424) );
  NAND2_X1 U7798 ( .A1(n8220), .A2(n12738), .ZN(n8217) );
  AND2_X1 U7799 ( .A1(n8218), .A2(n12737), .ZN(n8215) );
  INV_X1 U7800 ( .A(n12738), .ZN(n8219) );
  AND2_X1 U7801 ( .A1(n9189), .A2(n9190), .ZN(n8144) );
  OAI21_X1 U7802 ( .B1(n12184), .B2(n9634), .A(n9212), .ZN(n9213) );
  INV_X1 U7803 ( .A(n9240), .ZN(n8141) );
  NAND2_X1 U7804 ( .A1(n7614), .A2(n7613), .ZN(n12760) );
  AOI21_X1 U7805 ( .B1(n7615), .B2(n7618), .A(n7327), .ZN(n7613) );
  NOR2_X1 U7806 ( .A1(n7617), .A2(n12752), .ZN(n7618) );
  AOI22_X1 U7807 ( .A1(n14808), .A2(n9615), .B1(n14463), .B2(n9634), .ZN(n9291) );
  NOR2_X1 U7808 ( .A1(n7319), .A2(n7610), .ZN(n7609) );
  NOR2_X1 U7809 ( .A1(n8223), .A2(n12767), .ZN(n7610) );
  INV_X1 U7810 ( .A(n12766), .ZN(n8223) );
  AND2_X1 U7811 ( .A1(n12769), .A2(n12771), .ZN(n7611) );
  AND2_X1 U7812 ( .A1(n7609), .A2(n8224), .ZN(n7608) );
  NOR2_X1 U7813 ( .A1(n8225), .A2(n12766), .ZN(n8224) );
  INV_X1 U7814 ( .A(n12767), .ZN(n8225) );
  NAND2_X1 U7815 ( .A1(n7476), .A2(n7475), .ZN(n7474) );
  INV_X1 U7816 ( .A(n9343), .ZN(n7475) );
  NAND2_X1 U7817 ( .A1(n7600), .A2(n7599), .ZN(n12783) );
  AOI21_X1 U7818 ( .B1(n7601), .B2(n7604), .A(n7329), .ZN(n7599) );
  NAND2_X1 U7819 ( .A1(n8201), .A2(n12789), .ZN(n12795) );
  NAND2_X1 U7820 ( .A1(n12790), .A2(n12791), .ZN(n8201) );
  INV_X1 U7821 ( .A(n12796), .ZN(n8222) );
  AOI21_X1 U7822 ( .B1(n8124), .B2(n8122), .A(n9487), .ZN(n8121) );
  INV_X1 U7823 ( .A(n8125), .ZN(n8122) );
  NOR2_X1 U7824 ( .A1(n9468), .A2(n7243), .ZN(n8126) );
  NOR2_X1 U7825 ( .A1(n9647), .A2(n7798), .ZN(n9648) );
  NAND2_X1 U7826 ( .A1(n8089), .A2(n8088), .ZN(n13502) );
  INV_X1 U7827 ( .A(n9293), .ZN(n9297) );
  AND2_X1 U7828 ( .A1(n9142), .A2(n8009), .ZN(n8008) );
  INV_X1 U7829 ( .A(n9165), .ZN(n8009) );
  INV_X1 U7830 ( .A(n9134), .ZN(n8006) );
  OAI21_X1 U7831 ( .B1(n10252), .B2(n10273), .A(n7415), .ZN(n9038) );
  NAND2_X1 U7832 ( .A1(n10252), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7415) );
  AOI21_X1 U7833 ( .B1(n10880), .B2(n7756), .A(n7278), .ZN(n7754) );
  NAND2_X1 U7834 ( .A1(n7751), .A2(n10977), .ZN(n7750) );
  INV_X1 U7835 ( .A(n7754), .ZN(n7751) );
  NAND2_X1 U7836 ( .A1(n7744), .A2(n7752), .ZN(n7745) );
  NOR2_X1 U7837 ( .A1(n7755), .A2(n7780), .ZN(n7752) );
  NAND2_X1 U7838 ( .A1(n7757), .A2(n7363), .ZN(n12060) );
  NAND2_X1 U7839 ( .A1(n12060), .A2(n15855), .ZN(n12059) );
  OR2_X1 U7840 ( .A1(n15838), .A2(n15837), .ZN(n15835) );
  NOR2_X1 U7841 ( .A1(n13597), .A2(n13617), .ZN(n13633) );
  INV_X1 U7842 ( .A(n7845), .ZN(n7843) );
  OAI21_X1 U7843 ( .B1(n12979), .B2(n7870), .A(n7868), .ZN(n12981) );
  INV_X1 U7844 ( .A(n7869), .ZN(n7868) );
  OAI21_X1 U7845 ( .B1(n7871), .B2(n7870), .A(n13499), .ZN(n7869) );
  OR2_X1 U7846 ( .A1(n12980), .A2(n13812), .ZN(n13500) );
  NOR2_X1 U7847 ( .A1(n13841), .A2(n7872), .ZN(n7871) );
  INV_X1 U7848 ( .A(n13376), .ZN(n7872) );
  AND2_X1 U7849 ( .A1(n14123), .A2(n13914), .ZN(n8193) );
  INV_X1 U7850 ( .A(n8191), .ZN(n8190) );
  NAND2_X1 U7851 ( .A1(n8181), .A2(n8179), .ZN(n11890) );
  INV_X1 U7852 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8261) );
  INV_X1 U7853 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8805) );
  INV_X1 U7854 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7849) );
  NOR2_X1 U7855 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n8260) );
  NOR2_X1 U7856 ( .A1(n8641), .A2(n8624), .ZN(n8093) );
  INV_X1 U7857 ( .A(n8627), .ZN(n8095) );
  XNOR2_X1 U7858 ( .A(n8558), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8557) );
  INV_X1 U7859 ( .A(n10937), .ZN(n7876) );
  INV_X1 U7860 ( .A(n11364), .ZN(n7881) );
  AND2_X1 U7861 ( .A1(n11592), .A2(n11311), .ZN(n7880) );
  INV_X1 U7862 ( .A(n14298), .ZN(n7910) );
  NOR2_X1 U7863 ( .A1(n7889), .A2(n14354), .ZN(n7888) );
  INV_X1 U7864 ( .A(n9095), .ZN(n8943) );
  AND2_X1 U7865 ( .A1(n14646), .A2(n7662), .ZN(n7661) );
  NAND2_X1 U7866 ( .A1(n14504), .A2(n14506), .ZN(n7662) );
  NAND2_X1 U7867 ( .A1(n10468), .A2(n10467), .ZN(n10697) );
  OAI21_X1 U7868 ( .B1(n14465), .B2(n8065), .A(n7325), .ZN(n7681) );
  INV_X1 U7869 ( .A(n14467), .ZN(n8065) );
  XNOR2_X1 U7870 ( .A(n11795), .B(n14368), .ZN(n11714) );
  NOR2_X1 U7871 ( .A1(n11403), .A2(n8071), .ZN(n8070) );
  INV_X1 U7872 ( .A(n11401), .ZN(n8071) );
  NOR2_X1 U7873 ( .A1(n8973), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9194) );
  NOR2_X1 U7874 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8903) );
  NAND2_X1 U7875 ( .A1(n12676), .A2(n10226), .ZN(n9958) );
  OR2_X1 U7876 ( .A1(n16031), .A2(n11982), .ZN(n11983) );
  INV_X1 U7877 ( .A(n11446), .ZN(n7948) );
  XNOR2_X1 U7878 ( .A(n15073), .B(n15906), .ZN(n12855) );
  NAND2_X1 U7879 ( .A1(n7738), .A2(n7737), .ZN(n15380) );
  AND2_X1 U7880 ( .A1(n11027), .A2(n12838), .ZN(n12849) );
  INV_X1 U7881 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7946) );
  OAI21_X1 U7882 ( .B1(n9471), .B2(SI_23_), .A(n9470), .ZN(n9473) );
  NAND2_X1 U7883 ( .A1(n7980), .A2(SI_20_), .ZN(n7979) );
  INV_X1 U7884 ( .A(n9402), .ZN(n7980) );
  INV_X1 U7885 ( .A(n9729), .ZN(n7622) );
  INV_X1 U7886 ( .A(n9302), .ZN(n7997) );
  OR2_X1 U7887 ( .A1(n9298), .A2(n9297), .ZN(n7998) );
  NAND2_X1 U7888 ( .A1(n9192), .A2(n9191), .ZN(n9223) );
  NAND2_X1 U7889 ( .A1(n9171), .A2(n8244), .ZN(n9192) );
  AND4_X2 U7890 ( .A1(n9730), .A2(n15634), .A3(n9879), .A4(n9845), .ZN(n8231)
         );
  XNOR2_X1 U7891 ( .A(n8970), .B(SI_3_), .ZN(n8967) );
  AND2_X1 U7892 ( .A1(n7216), .A2(SI_2_), .ZN(n7416) );
  AOI22_X1 U7893 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15707), .B1(n15706), .B2(
        n15705), .ZN(n15710) );
  OR2_X1 U7894 ( .A1(n15707), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n15706) );
  OAI22_X1 U7895 ( .A1(n15757), .A2(n15756), .B1(P3_ADDR_REG_11__SCAN_IN), 
        .B2(n15755), .ZN(n15764) );
  AND2_X1 U7896 ( .A1(n7528), .A2(n8168), .ZN(n7526) );
  NAND2_X1 U7897 ( .A1(n7534), .A2(n7529), .ZN(n7528) );
  INV_X1 U7898 ( .A(n13262), .ZN(n7529) );
  OAI21_X1 U7899 ( .B1(n8703), .B2(n13316), .A(n7532), .ZN(n7535) );
  INV_X1 U7900 ( .A(n7544), .ZN(n7543) );
  OAI21_X1 U7901 ( .B1(n7545), .B2(n8623), .A(n8147), .ZN(n7544) );
  AOI21_X1 U7902 ( .B1(n8148), .B2(n8150), .A(n7307), .ZN(n8147) );
  OR2_X1 U7903 ( .A1(n8499), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8522) );
  NOR2_X1 U7904 ( .A1(n8184), .A2(n7539), .ZN(n7538) );
  INV_X1 U7905 ( .A(n11207), .ZN(n7539) );
  INV_X1 U7906 ( .A(n8376), .ZN(n8184) );
  NOR2_X1 U7907 ( .A1(n11388), .A2(n8186), .ZN(n8185) );
  INV_X1 U7908 ( .A(n8358), .ZN(n8186) );
  OR2_X1 U7909 ( .A1(n11943), .A2(n11944), .ZN(n11941) );
  AND4_X1 U7910 ( .A1(n13369), .A2(n13368), .A3(n13367), .A4(n13366), .ZN(
        n13760) );
  NOR2_X1 U7911 ( .A1(n10880), .A2(n7762), .ZN(n10854) );
  NOR2_X1 U7912 ( .A1(n7764), .A2(n7763), .ZN(n7762) );
  INV_X1 U7913 ( .A(n7776), .ZN(n7775) );
  NAND2_X1 U7914 ( .A1(n7467), .A2(n7320), .ZN(n7761) );
  NAND2_X1 U7915 ( .A1(n7761), .A2(n7760), .ZN(n11537) );
  INV_X1 U7916 ( .A(n11500), .ZN(n7760) );
  NAND2_X1 U7917 ( .A1(n7790), .A2(n7794), .ZN(n7792) );
  INV_X1 U7918 ( .A(n7757), .ZN(n15839) );
  NAND2_X1 U7919 ( .A1(n12059), .A2(n7462), .ZN(n15859) );
  OR2_X1 U7920 ( .A1(n12060), .A2(n15855), .ZN(n7462) );
  NOR2_X1 U7921 ( .A1(n15858), .A2(n15859), .ZN(n15857) );
  AND2_X1 U7922 ( .A1(n13592), .A2(n13608), .ZN(n13624) );
  OR2_X1 U7923 ( .A1(n13648), .A2(n13657), .ZN(n7766) );
  NAND3_X1 U7924 ( .A1(n7766), .A2(P3_REG1_REG_15__SCAN_IN), .A3(n13666), .ZN(
        n7767) );
  AOI21_X1 U7925 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n13695), .A(n13691), .ZN(
        n13715) );
  NAND2_X1 U7926 ( .A1(n13725), .A2(n7523), .ZN(n13728) );
  OR2_X1 U7927 ( .A1(n13726), .A2(n13727), .ZN(n7523) );
  INV_X1 U7928 ( .A(n7781), .ZN(n13726) );
  INV_X1 U7929 ( .A(n13751), .ZN(n7455) );
  NOR2_X1 U7930 ( .A1(n13748), .A2(n7457), .ZN(n7456) );
  NAND2_X1 U7931 ( .A1(n12979), .A2(n7871), .ZN(n13839) );
  INV_X1 U7932 ( .A(n13475), .ZN(n7865) );
  NOR2_X1 U7933 ( .A1(n13930), .A2(n8192), .ZN(n8191) );
  INV_X1 U7934 ( .A(n12941), .ZN(n8192) );
  AND2_X1 U7935 ( .A1(n13379), .A2(n13906), .ZN(n13930) );
  OR2_X1 U7936 ( .A1(n14133), .A2(n13974), .ZN(n13459) );
  INV_X1 U7937 ( .A(n7839), .ZN(n7838) );
  OAI21_X1 U7938 ( .B1(n13953), .B2(n7840), .A(n13941), .ZN(n7839) );
  INV_X1 U7939 ( .A(n13459), .ZN(n7840) );
  NAND2_X1 U7940 ( .A1(n8195), .A2(n8194), .ZN(n13938) );
  NAND2_X1 U7941 ( .A1(n13980), .A2(n13454), .ZN(n13954) );
  NAND2_X1 U7942 ( .A1(n13954), .A2(n13953), .ZN(n13952) );
  AND2_X1 U7943 ( .A1(n8171), .A2(n13972), .ZN(n8170) );
  NAND2_X1 U7944 ( .A1(n13447), .A2(n12937), .ZN(n8171) );
  NAND2_X1 U7945 ( .A1(n13991), .A2(n13448), .ZN(n12517) );
  OR2_X1 U7946 ( .A1(n12524), .A2(n13447), .ZN(n12938) );
  NAND2_X1 U7947 ( .A1(n12369), .A2(n13435), .ZN(n12370) );
  NAND2_X1 U7948 ( .A1(n11961), .A2(n11960), .ZN(n12162) );
  INV_X1 U7949 ( .A(n14002), .ZN(n13970) );
  NAND2_X1 U7950 ( .A1(n13401), .A2(n13400), .ZN(n11648) );
  AND2_X1 U7951 ( .A1(n11266), .A2(n13509), .ZN(n13997) );
  NAND2_X1 U7952 ( .A1(n8783), .A2(n8782), .ZN(n14091) );
  OR2_X1 U7953 ( .A1(n12960), .A2(n14156), .ZN(n8782) );
  NAND2_X1 U7954 ( .A1(n8736), .A2(n8735), .ZN(n12949) );
  OR2_X1 U7955 ( .A1(n12960), .A2(n12348), .ZN(n8735) );
  OR2_X1 U7956 ( .A1(n12960), .A2(n13105), .ZN(n8693) );
  NAND2_X1 U7957 ( .A1(n8593), .A2(n8592), .ZN(n13468) );
  NAND2_X1 U7958 ( .A1(n13388), .A2(n11259), .ZN(n16054) );
  INV_X1 U7959 ( .A(n16054), .ZN(n15940) );
  INV_X1 U7960 ( .A(n13944), .ZN(n13996) );
  AND2_X1 U7961 ( .A1(n8306), .A2(n8263), .ZN(n7834) );
  NAND2_X1 U7962 ( .A1(n8708), .A2(n12599), .ZN(n8111) );
  NAND2_X1 U7963 ( .A1(n8692), .A2(n8691), .ZN(n8705) );
  AND2_X1 U7965 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n11428), .ZN(n8115) );
  NAND2_X1 U7966 ( .A1(n8661), .A2(n11428), .ZN(n8116) );
  NAND2_X1 U7967 ( .A1(n8117), .A2(n8116), .ZN(n8662) );
  NAND2_X1 U7968 ( .A1(n8114), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8117) );
  INV_X1 U7969 ( .A(n8661), .ZN(n8114) );
  INV_X1 U7970 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8256) );
  OR2_X1 U7971 ( .A1(n8505), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U7972 ( .A1(n8424), .A2(n8423), .ZN(n8446) );
  NAND2_X1 U7973 ( .A1(n11226), .A2(n11225), .ZN(n11309) );
  AND2_X1 U7974 ( .A1(n14178), .A2(n14172), .ZN(n14216) );
  NOR2_X1 U7975 ( .A1(n14202), .A2(n7884), .ZN(n7883) );
  INV_X1 U7976 ( .A(n7885), .ZN(n7884) );
  INV_X1 U7977 ( .A(n9310), .ZN(n9308) );
  XNOR2_X1 U7978 ( .A(n11795), .B(n14188), .ZN(n11588) );
  NAND2_X1 U7979 ( .A1(n9151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9204) );
  INV_X1 U7980 ( .A(n9152), .ZN(n9151) );
  INV_X1 U7981 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n12288) );
  AOI21_X1 U7982 ( .B1(n7900), .B2(n7898), .A(n7289), .ZN(n7897) );
  INV_X1 U7983 ( .A(n7900), .ZN(n7899) );
  XNOR2_X1 U7984 ( .A(n9663), .B(n9662), .ZN(n10761) );
  NAND2_X1 U7985 ( .A1(n9255), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9285) );
  AOI21_X1 U7986 ( .B1(n14571), .B2(n9546), .A(n9528), .ZN(n14484) );
  CLKBUF_X1 U7987 ( .A(n9629), .Z(n7494) );
  OR2_X1 U7988 ( .A1(n8943), .A2(n8911), .ZN(n8915) );
  OR2_X1 U7989 ( .A1(n8943), .A2(n8897), .ZN(n8900) );
  NAND4_X1 U7990 ( .A1(n7388), .A2(n8874), .A3(n8875), .A4(n8873), .ZN(n9645)
         );
  NAND2_X1 U7991 ( .A1(n9095), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8875) );
  OR2_X1 U7992 ( .A1(n9334), .A2(n10443), .ZN(n8873) );
  OAI211_X1 U7993 ( .C1(n7670), .C2(n14614), .A(n14576), .B(n7671), .ZN(n14519) );
  NAND2_X1 U7994 ( .A1(n7672), .A2(n7673), .ZN(n7671) );
  INV_X1 U7995 ( .A(n7672), .ZN(n7670) );
  INV_X1 U7996 ( .A(n7813), .ZN(n7810) );
  AOI21_X1 U7997 ( .B1(n7813), .B2(n7815), .A(n7294), .ZN(n7809) );
  INV_X1 U7998 ( .A(n14513), .ZN(n7815) );
  INV_X1 U7999 ( .A(n8072), .ZN(n7695) );
  OR2_X1 U8000 ( .A1(n14645), .A2(n7275), .ZN(n7696) );
  OR2_X1 U8001 ( .A1(n14668), .A2(n7659), .ZN(n7656) );
  INV_X1 U8002 ( .A(n7661), .ZN(n7659) );
  OR2_X1 U8003 ( .A1(n9386), .A2(n14304), .ZN(n9410) );
  AND2_X1 U8004 ( .A1(n7651), .A2(n14500), .ZN(n7650) );
  NAND2_X1 U8005 ( .A1(n14498), .A2(n7652), .ZN(n7651) );
  INV_X1 U8006 ( .A(n14496), .ZN(n7652) );
  INV_X1 U8007 ( .A(n14468), .ZN(n14691) );
  AOI21_X1 U8008 ( .B1(n7666), .B2(n12423), .A(n7665), .ZN(n7664) );
  NAND2_X1 U8009 ( .A1(n14465), .A2(n8068), .ZN(n14704) );
  NAND2_X1 U8010 ( .A1(n7668), .A2(n7669), .ZN(n7667) );
  INV_X1 U8011 ( .A(n12424), .ZN(n7668) );
  NAND2_X1 U8012 ( .A1(n7667), .A2(n7666), .ZN(n14708) );
  OR2_X2 U8013 ( .A1(n12019), .A2(n12192), .ZN(n12120) );
  NAND2_X1 U8014 ( .A1(n7817), .A2(n7816), .ZN(n12011) );
  NOR2_X1 U8015 ( .A1(n7819), .A2(n11861), .ZN(n7816) );
  OR2_X1 U8016 ( .A1(n12145), .A2(n11719), .ZN(n11722) );
  NAND2_X1 U8017 ( .A1(n7709), .A2(n7708), .ZN(n12152) );
  OAI21_X1 U8018 ( .B1(n7801), .B2(n11512), .A(n7799), .ZN(n11715) );
  AOI21_X1 U8019 ( .B1(n7802), .B2(n7800), .A(n7317), .ZN(n7799) );
  OR2_X1 U8020 ( .A1(n11510), .A2(n11511), .ZN(n7803) );
  NAND2_X1 U8021 ( .A1(n10694), .A2(n10693), .ZN(n10829) );
  XNOR2_X1 U8022 ( .A(n14374), .B(n12099), .ZN(n10691) );
  NAND2_X1 U8023 ( .A1(n7409), .A2(n10683), .ZN(n10488) );
  INV_X1 U8024 ( .A(n10492), .ZN(n7409) );
  CLKBUF_X1 U8025 ( .A(n10492), .Z(n7425) );
  NAND2_X1 U8026 ( .A1(n9623), .A2(n9622), .ZN(n14736) );
  NAND2_X1 U8027 ( .A1(n9409), .A2(n9408), .ZN(n14784) );
  NAND2_X1 U8028 ( .A1(n9385), .A2(n9384), .ZN(n14789) );
  NAND2_X1 U8029 ( .A1(n8076), .A2(n12419), .ZN(n8074) );
  INV_X1 U8030 ( .A(n12419), .ZN(n8073) );
  NAND2_X1 U8031 ( .A1(n12422), .A2(n12427), .ZN(n14465) );
  AND2_X1 U8032 ( .A1(n12357), .A2(n12356), .ZN(n8075) );
  AND2_X1 U8033 ( .A1(n8058), .A2(n12007), .ZN(n7697) );
  NAND2_X1 U8034 ( .A1(n11861), .A2(n8059), .ZN(n8058) );
  INV_X1 U8035 ( .A(n11853), .ZN(n8059) );
  NAND2_X1 U8036 ( .A1(n11705), .A2(n11720), .ZN(n11707) );
  OR2_X1 U8037 ( .A1(n12143), .A2(n12157), .ZN(n11706) );
  NAND2_X1 U8038 ( .A1(n11046), .A2(n11045), .ZN(n11402) );
  NAND2_X1 U8039 ( .A1(n11402), .A2(n8070), .ZN(n11508) );
  INV_X1 U8040 ( .A(n7449), .ZN(n10494) );
  NAND2_X1 U8041 ( .A1(n12451), .A2(n9706), .ZN(n10762) );
  AND2_X1 U8042 ( .A1(n10761), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9749) );
  NOR2_X2 U8043 ( .A1(n9305), .A2(n8867), .ZN(n8881) );
  NAND2_X1 U8044 ( .A1(n9698), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9701) );
  INV_X1 U8045 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9700) );
  NAND2_X1 U8046 ( .A1(n9701), .A2(n9700), .ZN(n9703) );
  NAND2_X1 U8047 ( .A1(n8846), .A2(n7911), .ZN(n8848) );
  AND2_X1 U8048 ( .A1(n8135), .A2(n8861), .ZN(n7911) );
  OR2_X1 U8049 ( .A1(n8959), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8973) );
  INV_X1 U8050 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8876) );
  INV_X1 U8051 ( .A(n14886), .ZN(n8028) );
  AND2_X1 U8052 ( .A1(n14885), .A2(n14884), .ZN(n14886) );
  AOI21_X1 U8053 ( .B1(n7273), .B2(n8020), .A(n8017), .ZN(n8016) );
  INV_X1 U8054 ( .A(n15033), .ZN(n8017) );
  AOI21_X1 U8055 ( .B1(n14880), .B2(n14879), .A(n14951), .ZN(n14916) );
  NAND2_X1 U8056 ( .A1(n11454), .A2(n7302), .ZN(n11664) );
  AOI21_X1 U8057 ( .B1(n8041), .B2(n8040), .A(n7312), .ZN(n8039) );
  INV_X1 U8058 ( .A(n8041), .ZN(n8038) );
  INV_X1 U8059 ( .A(n12509), .ZN(n8040) );
  INV_X1 U8060 ( .A(n14986), .ZN(n7453) );
  NOR2_X1 U8061 ( .A1(n15014), .A2(n8045), .ZN(n8044) );
  OR2_X1 U8062 ( .A1(n10197), .A2(n10198), .ZN(n7511) );
  OR2_X1 U8063 ( .A1(n10183), .A2(n9914), .ZN(n9916) );
  INV_X1 U8064 ( .A(n15403), .ZN(n15167) );
  AND2_X1 U8065 ( .A1(n12643), .A2(n12638), .ZN(n14960) );
  INV_X1 U8066 ( .A(n7578), .ZN(n7577) );
  INV_X1 U8067 ( .A(n12879), .ZN(n15187) );
  NAND2_X1 U8068 ( .A1(n15433), .A2(n15257), .ZN(n7926) );
  NAND2_X1 U8069 ( .A1(n7217), .A2(n12877), .ZN(n7927) );
  OR2_X1 U8070 ( .A1(n15276), .A2(n7959), .ZN(n7953) );
  NOR2_X1 U8071 ( .A1(n15276), .A2(n7956), .ZN(n7955) );
  OR2_X1 U8072 ( .A1(n15452), .A2(n15310), .ZN(n8235) );
  NAND2_X1 U8073 ( .A1(n15302), .A2(n7957), .ZN(n7960) );
  NAND2_X1 U8074 ( .A1(n15302), .A2(n12610), .ZN(n15283) );
  NAND2_X1 U8075 ( .A1(n15308), .A2(n15307), .ZN(n15306) );
  NAND2_X1 U8076 ( .A1(n12604), .A2(n12603), .ZN(n15388) );
  NOR2_X1 U8077 ( .A1(n7265), .A2(n7951), .ZN(n7950) );
  AOI21_X1 U8078 ( .B1(n7919), .B2(n12869), .A(n8246), .ZN(n7917) );
  NOR2_X1 U8079 ( .A1(n7918), .A2(n7584), .ZN(n7583) );
  INV_X1 U8080 ( .A(n12385), .ZN(n7584) );
  INV_X1 U8081 ( .A(n7919), .ZN(n7918) );
  NAND2_X1 U8082 ( .A1(n7582), .A2(n7581), .ZN(n15372) );
  AND2_X1 U8083 ( .A1(n7917), .A2(n15387), .ZN(n7581) );
  NOR2_X1 U8084 ( .A1(n12871), .A2(n7920), .ZN(n7919) );
  INV_X1 U8085 ( .A(n12446), .ZN(n7920) );
  NAND2_X1 U8086 ( .A1(n12445), .A2(n12444), .ZN(n7921) );
  XNOR2_X1 U8087 ( .A(n12755), .B(n15374), .ZN(n12871) );
  NAND2_X1 U8088 ( .A1(n12386), .A2(n12385), .ZN(n12445) );
  NAND2_X1 U8089 ( .A1(n7944), .A2(n11930), .ZN(n15980) );
  AND2_X1 U8090 ( .A1(n15983), .A2(n11916), .ZN(n7933) );
  NAND2_X1 U8091 ( .A1(n9957), .A2(n9956), .ZN(n12716) );
  AND2_X1 U8092 ( .A1(n10231), .A2(n10265), .ZN(n15376) );
  OR2_X1 U8093 ( .A1(n11020), .A2(n15150), .ZN(n12928) );
  NAND2_X1 U8094 ( .A1(n10909), .A2(n10908), .ZN(n10993) );
  NAND2_X1 U8095 ( .A1(n12628), .A2(n12627), .ZN(n15413) );
  AND2_X1 U8096 ( .A1(n15425), .A2(n16134), .ZN(n7382) );
  INV_X1 U8097 ( .A(n12674), .ZN(n10903) );
  NAND2_X1 U8098 ( .A1(n9562), .A2(n8013), .ZN(n9598) );
  AND2_X1 U8099 ( .A1(n8014), .A2(n9561), .ZN(n8013) );
  INV_X1 U8100 ( .A(n9763), .ZN(n9758) );
  NAND2_X1 U8101 ( .A1(n7984), .A2(n7983), .ZN(n7982) );
  NAND2_X1 U8102 ( .A1(n9402), .A2(n13114), .ZN(n7983) );
  NAND2_X1 U8103 ( .A1(n7985), .A2(n7986), .ZN(n9406) );
  NAND2_X1 U8104 ( .A1(n7441), .A2(n13114), .ZN(n7986) );
  NAND2_X1 U8105 ( .A1(n7981), .A2(n9402), .ZN(n7985) );
  OR2_X1 U8106 ( .A1(n7441), .A2(n13114), .ZN(n7981) );
  NAND2_X1 U8107 ( .A1(n7441), .A2(n7979), .ZN(n7976) );
  AND2_X1 U8108 ( .A1(n10116), .A2(n10098), .ZN(n11837) );
  XNOR2_X1 U8109 ( .A(n9110), .B(SI_9_), .ZN(n10380) );
  OR2_X1 U8110 ( .A1(n9993), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9920) );
  NAND2_X1 U8111 ( .A1(n15501), .A2(n9845), .ZN(n7630) );
  AOI22_X1 U8112 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n10886), .B1(n15693), .B2(
        n15692), .ZN(n15702) );
  OR2_X1 U8113 ( .A1(n10886), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n15692) );
  OAI21_X1 U8114 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n15781), .A(n15780), .ZN(
        n15787) );
  NAND2_X1 U8115 ( .A1(n15792), .A2(n7719), .ZN(n7717) );
  NAND2_X1 U8116 ( .A1(n8175), .A2(n8173), .ZN(n11813) );
  AOI21_X1 U8117 ( .B1(n11944), .B2(n8417), .A(n8174), .ZN(n8173) );
  NAND2_X1 U8118 ( .A1(n11943), .A2(n8417), .ZN(n8175) );
  INV_X1 U8119 ( .A(n11814), .ZN(n8174) );
  AND4_X1 U8120 ( .A1(n8637), .A2(n8636), .A3(n8635), .A4(n8634), .ZN(n13899)
         );
  NAND2_X1 U8121 ( .A1(n12002), .A2(n12001), .ZN(n12000) );
  AOI21_X1 U8122 ( .B1(n7272), .B2(n8157), .A(n8155), .ZN(n8154) );
  INV_X1 U8123 ( .A(n13270), .ZN(n8155) );
  INV_X1 U8124 ( .A(n13899), .ZN(n13924) );
  OR2_X1 U8125 ( .A1(n15851), .A2(n15852), .ZN(n7410) );
  OAI21_X1 U8126 ( .B1(n13724), .B2(n7466), .A(n7465), .ZN(n13698) );
  INV_X1 U8127 ( .A(n13725), .ZN(n13724) );
  MUX2_X1 U8128 ( .A(n10639), .B(P3_U3897), .S(n12963), .Z(n13754) );
  OR2_X1 U8129 ( .A1(n10638), .A2(n13603), .ZN(n15866) );
  XNOR2_X1 U8130 ( .A(n13553), .B(n13546), .ZN(n13221) );
  NAND2_X1 U8131 ( .A1(n13783), .A2(n12986), .ZN(n13774) );
  NAND2_X1 U8132 ( .A1(n13784), .A2(n12952), .ZN(n13766) );
  INV_X1 U8133 ( .A(n13791), .ZN(n14019) );
  NAND2_X1 U8134 ( .A1(n8727), .A2(n8726), .ZN(n14035) );
  NAND2_X1 U8135 ( .A1(n8631), .A2(n8630), .ZN(n14054) );
  INV_X1 U8136 ( .A(n14091), .ZN(n14017) );
  NAND2_X1 U8137 ( .A1(n14091), .A2(n14124), .ZN(n7497) );
  AND2_X1 U8138 ( .A1(n8710), .A2(n8709), .ZN(n14108) );
  AND2_X1 U8139 ( .A1(n8792), .A2(n8791), .ZN(n11635) );
  INV_X1 U8140 ( .A(n12036), .ZN(n15855) );
  NAND2_X1 U8141 ( .A1(n14209), .A2(n8240), .ZN(n14210) );
  NAND2_X1 U8142 ( .A1(n9454), .A2(n9453), .ZN(n14769) );
  NAND2_X1 U8143 ( .A1(n14345), .A2(n7883), .ZN(n14238) );
  AND2_X1 U8144 ( .A1(n10665), .A2(n10667), .ZN(n10674) );
  OR2_X1 U8145 ( .A1(n10663), .A2(n10664), .ZN(n10665) );
  NAND2_X1 U8146 ( .A1(n14196), .A2(n14251), .ZN(n14333) );
  OAI21_X1 U8147 ( .B1(n14164), .B2(n14163), .A(n14280), .ZN(n14287) );
  NAND2_X1 U8148 ( .A1(n9307), .A2(n9306), .ZN(n14723) );
  AOI21_X1 U8149 ( .B1(n10753), .B2(n10752), .A(n8242), .ZN(n10760) );
  INV_X1 U8150 ( .A(n10840), .ZN(n10752) );
  NAND2_X1 U8151 ( .A1(n7449), .A2(n10496), .ZN(n10683) );
  INV_X1 U8152 ( .A(n7371), .ZN(n7436) );
  NAND2_X1 U8153 ( .A1(n9431), .A2(n9430), .ZN(n14778) );
  OR2_X1 U8154 ( .A1(n11872), .A2(n9599), .ZN(n9431) );
  NAND2_X1 U8155 ( .A1(n9149), .A2(n9148), .ZN(n12091) );
  INV_X1 U8156 ( .A(n14573), .ZN(n14755) );
  AND2_X1 U8157 ( .A1(n9718), .A2(n7487), .ZN(n7486) );
  NOR2_X1 U8158 ( .A1(n7489), .A2(n7488), .ZN(n7487) );
  INV_X1 U8159 ( .A(n9691), .ZN(n7488) );
  INV_X1 U8160 ( .A(n9690), .ZN(n7489) );
  NAND2_X1 U8161 ( .A1(n9552), .A2(n9551), .ZN(n14520) );
  NAND2_X1 U8162 ( .A1(n9504), .A2(n9503), .ZN(n14482) );
  NAND2_X1 U8163 ( .A1(n9441), .A2(n9440), .ZN(n14476) );
  NAND2_X1 U8164 ( .A1(n9417), .A2(n9416), .ZN(n14507) );
  CLKBUF_X1 U8165 ( .A(n9645), .Z(n7449) );
  NAND2_X1 U8166 ( .A1(n7358), .A2(n12155), .ZN(n7828) );
  NAND2_X1 U8167 ( .A1(n14533), .A2(n7683), .ZN(n7682) );
  NAND2_X1 U8168 ( .A1(n14741), .A2(n9643), .ZN(n7683) );
  NAND2_X1 U8169 ( .A1(n9496), .A2(n9495), .ZN(n14759) );
  NAND2_X1 U8170 ( .A1(n8077), .A2(n8076), .ZN(n16109) );
  AND2_X1 U8171 ( .A1(n12150), .A2(n11736), .ZN(n14728) );
  OR2_X1 U8172 ( .A1(n8905), .A2(n10520), .ZN(n8908) );
  INV_X1 U8173 ( .A(n14742), .ZN(n7679) );
  NAND2_X1 U8174 ( .A1(n14747), .A2(n7429), .ZN(n14749) );
  AND2_X1 U8175 ( .A1(n14746), .A2(n7430), .ZN(n7429) );
  NAND2_X1 U8176 ( .A1(n14563), .A2(n16112), .ZN(n7430) );
  NOR2_X1 U8177 ( .A1(n14825), .A2(n14849), .ZN(n7505) );
  NAND2_X1 U8178 ( .A1(n10472), .A2(n10471), .ZN(n15524) );
  NAND2_X1 U8179 ( .A1(n10178), .A2(n10177), .ZN(n15460) );
  NOR2_X1 U8180 ( .A1(n8032), .A2(n15042), .ZN(n8030) );
  NOR2_X1 U8181 ( .A1(n8035), .A2(n8033), .ZN(n8032) );
  INV_X1 U8182 ( .A(n8036), .ZN(n8033) );
  NAND2_X1 U8183 ( .A1(n8036), .A2(n8037), .ZN(n8034) );
  INV_X1 U8184 ( .A(n14958), .ZN(n8037) );
  NAND2_X1 U8185 ( .A1(n12634), .A2(n12633), .ZN(n15408) );
  NAND2_X1 U8186 ( .A1(n9815), .A2(n9814), .ZN(n15474) );
  OR2_X1 U8187 ( .A1(n9846), .A2(n7254), .ZN(n9883) );
  NAND2_X1 U8188 ( .A1(n10162), .A2(n10161), .ZN(n15466) );
  NAND2_X1 U8189 ( .A1(n12619), .A2(n12618), .ZN(n15420) );
  NAND2_X1 U8190 ( .A1(n8003), .A2(n12894), .ZN(n12903) );
  NAND2_X1 U8191 ( .A1(n12888), .A2(n12887), .ZN(n8003) );
  NAND2_X1 U8192 ( .A1(n8002), .A2(n8001), .ZN(n8000) );
  NAND2_X1 U8193 ( .A1(n12910), .A2(n12904), .ZN(n8002) );
  NAND2_X1 U8194 ( .A1(n7591), .A2(n12827), .ZN(n7590) );
  NAND4_X1 U8195 ( .A1(n12626), .A2(n12625), .A3(n12624), .A4(n12623), .ZN(
        n15057) );
  NAND2_X1 U8196 ( .A1(n9840), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U8197 ( .A1(n9870), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9855) );
  OAI21_X1 U8198 ( .B1(n15146), .B2(n15145), .A(n7637), .ZN(n7636) );
  AOI21_X1 U8199 ( .B1(n15148), .B2(n15149), .A(n15147), .ZN(n7637) );
  AND2_X1 U8200 ( .A1(n7579), .A2(n7240), .ZN(n15206) );
  NAND2_X1 U8201 ( .A1(n7579), .A2(n7922), .ZN(n15207) );
  AOI21_X1 U8202 ( .B1(n15203), .B2(n15202), .A(n15201), .ZN(n15205) );
  NAND2_X1 U8203 ( .A1(n15222), .A2(n7970), .ZN(n15202) );
  NAND2_X1 U8204 ( .A1(n16120), .A2(n12605), .ZN(n15352) );
  NAND2_X1 U8205 ( .A1(n10141), .A2(n10140), .ZN(n15386) );
  NAND2_X1 U8206 ( .A1(n12302), .A2(n12301), .ZN(n12304) );
  NAND2_X1 U8207 ( .A1(n7218), .A2(n11028), .ZN(n15365) );
  NAND2_X1 U8208 ( .A1(n8207), .A2(n8206), .ZN(n8205) );
  INV_X1 U8209 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8206) );
  INV_X1 U8210 ( .A(n8208), .ZN(n8207) );
  NAND2_X1 U8211 ( .A1(n15739), .A2(n15740), .ZN(n15742) );
  NAND2_X1 U8212 ( .A1(n15742), .A2(n15743), .ZN(n15748) );
  NAND2_X1 U8213 ( .A1(n15734), .A2(n7710), .ZN(n15749) );
  INV_X1 U8214 ( .A(n15740), .ZN(n7710) );
  NOR2_X1 U8215 ( .A1(n15782), .A2(n15783), .ZN(n15785) );
  NAND2_X1 U8216 ( .A1(n7730), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7729) );
  OR2_X1 U8217 ( .A1(n15822), .A2(n15821), .ZN(n7728) );
  OAI21_X1 U8218 ( .B1(n10830), .B2(n9615), .A(n8984), .ZN(n8985) );
  NAND2_X1 U8219 ( .A1(n9034), .A2(n7287), .ZN(n8142) );
  NAND2_X1 U8220 ( .A1(n7623), .A2(n12726), .ZN(n8214) );
  INV_X1 U8221 ( .A(n9081), .ZN(n7423) );
  INV_X1 U8222 ( .A(n9130), .ZN(n8138) );
  INV_X1 U8223 ( .A(n9190), .ZN(n7515) );
  NAND2_X1 U8224 ( .A1(n7598), .A2(n12745), .ZN(n7596) );
  OR2_X1 U8225 ( .A1(n7597), .A2(n7595), .ZN(n7594) );
  AND2_X1 U8226 ( .A1(n12741), .A2(n12745), .ZN(n7595) );
  NOR2_X1 U8227 ( .A1(n7315), .A2(n7616), .ZN(n7615) );
  AND2_X1 U8228 ( .A1(n7617), .A2(n12752), .ZN(n7616) );
  INV_X1 U8229 ( .A(n12769), .ZN(n7612) );
  NAND2_X1 U8230 ( .A1(n8141), .A2(n8140), .ZN(n8139) );
  INV_X1 U8231 ( .A(n9239), .ZN(n8140) );
  AND2_X1 U8232 ( .A1(n9270), .A2(n9269), .ZN(n9272) );
  OAI21_X1 U8233 ( .B1(n14495), .B2(n9634), .A(n9316), .ZN(n9317) );
  INV_X1 U8234 ( .A(n9344), .ZN(n7476) );
  NAND2_X1 U8235 ( .A1(n12772), .A2(n12774), .ZN(n8212) );
  NOR2_X1 U8236 ( .A1(n7323), .A2(n7608), .ZN(n7607) );
  AND2_X1 U8237 ( .A1(n12777), .A2(n7605), .ZN(n7604) );
  INV_X1 U8238 ( .A(n12775), .ZN(n7605) );
  AND2_X1 U8239 ( .A1(n7602), .A2(n7341), .ZN(n7601) );
  NAND2_X1 U8240 ( .A1(n12775), .A2(n7603), .ZN(n7602) );
  NOR2_X1 U8241 ( .A1(n9372), .A2(n9371), .ZN(n9400) );
  INV_X1 U8242 ( .A(n9396), .ZN(n7438) );
  OAI21_X1 U8243 ( .B1(n14505), .B2(n9615), .A(n9395), .ZN(n9396) );
  OAI22_X1 U8244 ( .A1(n12798), .A2(n7310), .B1(n12797), .B2(n8222), .ZN(
        n12801) );
  NOR2_X1 U8245 ( .A1(n12983), .A2(n8091), .ZN(n8090) );
  NAND2_X1 U8246 ( .A1(n13492), .A2(n13493), .ZN(n8091) );
  AOI22_X1 U8247 ( .A1(n8121), .A2(n8123), .B1(n7258), .B2(n8126), .ZN(n8119)
         );
  INV_X1 U8248 ( .A(n8124), .ZN(n8123) );
  INV_X1 U8249 ( .A(n7995), .ZN(n7994) );
  AOI21_X1 U8250 ( .B1(n7995), .B2(n7993), .A(n9374), .ZN(n7992) );
  INV_X1 U8251 ( .A(n7255), .ZN(n7993) );
  AOI21_X1 U8252 ( .B1(n7255), .B2(n9297), .A(n7996), .ZN(n7995) );
  INV_X1 U8253 ( .A(n9324), .ZN(n7996) );
  INV_X1 U8254 ( .A(n13487), .ZN(n7870) );
  INV_X1 U8255 ( .A(n13393), .ZN(n7470) );
  INV_X1 U8256 ( .A(n8107), .ZN(n8106) );
  OAI21_X1 U8257 ( .B1(n8704), .B2(n8108), .A(n8724), .ZN(n8107) );
  INV_X1 U8258 ( .A(n8706), .ZN(n8108) );
  NAND2_X1 U8259 ( .A1(n8069), .A2(n14467), .ZN(n8064) );
  NOR2_X1 U8260 ( .A1(n12879), .A2(n7965), .ZN(n7964) );
  INV_X1 U8261 ( .A(n7966), .ZN(n7965) );
  INV_X1 U8262 ( .A(n7932), .ZN(n9780) );
  INV_X1 U8263 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7988) );
  AND2_X1 U8264 ( .A1(n8166), .A2(n8169), .ZN(n8165) );
  NAND2_X1 U8265 ( .A1(n13222), .A2(n8167), .ZN(n8166) );
  NOR2_X1 U8266 ( .A1(n8239), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U8267 ( .A1(n8087), .A2(n8085), .ZN(n13505) );
  NAND2_X1 U8268 ( .A1(n7435), .A2(n7765), .ZN(n7764) );
  NAND2_X1 U8269 ( .A1(n10853), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7765) );
  NAND2_X1 U8270 ( .A1(n7410), .A2(n12047), .ZN(n7784) );
  NAND2_X1 U8271 ( .A1(n7784), .A2(n7783), .ZN(n13590) );
  INV_X1 U8272 ( .A(n12049), .ZN(n7783) );
  NAND2_X1 U8273 ( .A1(n13654), .A2(n7459), .ZN(n13679) );
  OR2_X1 U8274 ( .A1(n13655), .A2(n13656), .ZN(n7459) );
  OR2_X1 U8275 ( .A1(n13694), .A2(n7782), .ZN(n7781) );
  NOR2_X1 U8276 ( .A1(n13688), .A2(n13670), .ZN(n7782) );
  INV_X1 U8277 ( .A(n14108), .ZN(n12980) );
  INV_X1 U8278 ( .A(n13479), .ZN(n7858) );
  OR2_X1 U8279 ( .A1(n14051), .A2(n13881), .ZN(n13521) );
  OR2_X1 U8280 ( .A1(n14141), .A2(n13995), .ZN(n13450) );
  INV_X1 U8281 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n13062) );
  INV_X1 U8282 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8306) );
  NOR2_X1 U8283 ( .A1(n8569), .A2(n8101), .ZN(n8099) );
  INV_X1 U8284 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8489) );
  AND2_X1 U8285 ( .A1(n14216), .A2(n7910), .ZN(n7905) );
  INV_X1 U8286 ( .A(n7905), .ZN(n7898) );
  NOR2_X1 U8287 ( .A1(n14736), .A2(n14545), .ZN(n7701) );
  NAND2_X1 U8288 ( .A1(n9497), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9523) );
  INV_X1 U8289 ( .A(n7657), .ZN(n7655) );
  NOR2_X1 U8290 ( .A1(n14634), .A2(n14769), .ZN(n7707) );
  NAND2_X1 U8291 ( .A1(n9432), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9457) );
  INV_X1 U8292 ( .A(n9434), .ZN(n9432) );
  INV_X1 U8293 ( .A(n14706), .ZN(n7665) );
  OR2_X1 U8294 ( .A1(n14808), .A2(n16111), .ZN(n7705) );
  AOI21_X1 U8295 ( .B1(n7268), .B2(n7803), .A(n11751), .ZN(n7802) );
  INV_X1 U8296 ( .A(n7803), .ZN(n7800) );
  NOR2_X1 U8297 ( .A1(n7826), .A2(n7823), .ZN(n7822) );
  INV_X1 U8298 ( .A(n10693), .ZN(n7823) );
  AND2_X1 U8299 ( .A1(n14563), .A2(n14520), .ZN(n8063) );
  OR2_X1 U8300 ( .A1(n8070), .A2(n7688), .ZN(n7687) );
  INV_X1 U8301 ( .A(n11507), .ZN(n7688) );
  INV_X1 U8302 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8880) );
  INV_X1 U8303 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8845) );
  AND2_X1 U8304 ( .A1(n7250), .A2(n7343), .ZN(n8135) );
  INV_X1 U8305 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9326) );
  OR2_X1 U8306 ( .A1(n9249), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n9251) );
  OR2_X1 U8307 ( .A1(n14977), .A2(n8020), .ZN(n8019) );
  INV_X1 U8308 ( .A(n14904), .ZN(n8020) );
  INV_X1 U8309 ( .A(n10218), .ZN(n8024) );
  NAND2_X1 U8310 ( .A1(n8203), .A2(n8202), .ZN(n12820) );
  NAND2_X1 U8311 ( .A1(n12815), .A2(n12817), .ZN(n8202) );
  XNOR2_X1 U8312 ( .A(n15420), .B(n14918), .ZN(n12879) );
  NOR2_X1 U8313 ( .A1(n15203), .A2(n7967), .ZN(n7966) );
  INV_X1 U8314 ( .A(n7970), .ZN(n7967) );
  NOR2_X1 U8315 ( .A1(n9791), .A2(n10232), .ZN(n10220) );
  INV_X1 U8316 ( .A(n12593), .ZN(n12580) );
  INV_X1 U8317 ( .A(n7957), .ZN(n7956) );
  OAI21_X1 U8318 ( .B1(n7266), .B2(n7575), .A(n12660), .ZN(n7574) );
  NAND2_X1 U8319 ( .A1(n10142), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10144) );
  OR2_X1 U8320 ( .A1(n10144), .A2(n9832), .ZN(n9834) );
  INV_X1 U8321 ( .A(n12438), .ZN(n7951) );
  OR2_X1 U8322 ( .A1(n10079), .A2(n10078), .ZN(n10102) );
  INV_X1 U8323 ( .A(n11983), .ZN(n7941) );
  INV_X1 U8324 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9728) );
  INV_X1 U8325 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9727) );
  NAND2_X1 U8326 ( .A1(n8011), .A2(n9540), .ZN(n9554) );
  OR2_X1 U8327 ( .A1(n9537), .A2(n9536), .ZN(n8011) );
  INV_X1 U8328 ( .A(n7978), .ZN(n7977) );
  OAI21_X1 U8329 ( .B1(n7982), .B2(n7979), .A(n9424), .ZN(n7978) );
  INV_X1 U8330 ( .A(SI_22_), .ZN(n13105) );
  AOI21_X1 U8331 ( .B1(n8008), .B2(n8006), .A(n8005), .ZN(n8004) );
  INV_X1 U8332 ( .A(n8008), .ZN(n8007) );
  INV_X1 U8333 ( .A(n9167), .ZN(n8005) );
  NOR2_X1 U8334 ( .A1(n10038), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n10074) );
  NAND2_X1 U8335 ( .A1(n9111), .A2(SI_9_), .ZN(n7433) );
  NAND2_X1 U8336 ( .A1(n7384), .A2(n8971), .ZN(n8988) );
  INV_X1 U8337 ( .A(n8967), .ZN(n8968) );
  OAI21_X1 U8338 ( .B1(n15662), .B2(n15663), .A(n7721), .ZN(n7720) );
  NAND2_X1 U8339 ( .A1(n15664), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7721) );
  AOI21_X1 U8340 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n11465), .A(n15766), .ZN(
        n15769) );
  NOR2_X1 U8341 ( .A1(n15765), .A2(n15764), .ZN(n15766) );
  INV_X1 U8342 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7719) );
  OR2_X1 U8343 ( .A1(n15800), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n15801) );
  INV_X1 U8344 ( .A(n8640), .ZN(n8150) );
  INV_X1 U8345 ( .A(n8165), .ZN(n8163) );
  OAI21_X1 U8346 ( .B1(n7241), .B2(n8162), .A(n8161), .ZN(n8160) );
  NOR2_X1 U8347 ( .A1(n8163), .A2(n7260), .ZN(n8162) );
  NAND2_X1 U8348 ( .A1(n7241), .A2(n8165), .ZN(n8161) );
  OR2_X1 U8349 ( .A1(n8584), .A2(n8157), .ZN(n8156) );
  INV_X1 U8350 ( .A(n8586), .ZN(n8157) );
  NAND2_X1 U8351 ( .A1(n11206), .A2(n8185), .ZN(n11385) );
  NAND2_X1 U8352 ( .A1(n12000), .A2(n8177), .ZN(n12230) );
  AND2_X1 U8353 ( .A1(n8436), .A2(n13062), .ZN(n8470) );
  NAND2_X1 U8354 ( .A1(n8198), .A2(n8196), .ZN(n13229) );
  AND2_X1 U8355 ( .A1(n8556), .A2(n8197), .ZN(n8196) );
  NAND2_X1 U8356 ( .A1(n12560), .A2(n13576), .ZN(n8197) );
  NAND2_X1 U8357 ( .A1(n12562), .A2(n8199), .ZN(n8198) );
  OR2_X1 U8358 ( .A1(n12560), .A2(n13576), .ZN(n8199) );
  NOR2_X1 U8359 ( .A1(n8522), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8547) );
  OR2_X1 U8360 ( .A1(n8481), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8499) );
  XNOR2_X1 U8361 ( .A(n8711), .B(n13380), .ZN(n8321) );
  NOR2_X1 U8362 ( .A1(n8576), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U8363 ( .A1(n13518), .A2(n13519), .ZN(n8082) );
  AND4_X1 U8364 ( .A1(n8504), .A2(n8503), .A3(n8502), .A4(n8501), .ZN(n8514)
         );
  OAI21_X1 U8365 ( .B1(n10811), .B2(P3_REG1_REG_2__SCAN_IN), .A(n7502), .ZN(
        n10801) );
  NAND2_X1 U8366 ( .A1(n10849), .A2(n7559), .ZN(n7787) );
  AND2_X1 U8367 ( .A1(n10848), .A2(n10872), .ZN(n7559) );
  NAND2_X1 U8368 ( .A1(n7788), .A2(n7763), .ZN(n10876) );
  OR2_X1 U8369 ( .A1(n7786), .A2(n7785), .ZN(n10878) );
  INV_X1 U8370 ( .A(n10876), .ZN(n7785) );
  NAND2_X1 U8371 ( .A1(n7746), .A2(n7745), .ZN(n10970) );
  NAND2_X1 U8372 ( .A1(n7745), .A2(n7750), .ZN(n11145) );
  OAI21_X1 U8373 ( .B1(n11327), .B2(n11326), .A(n11328), .ZN(n11333) );
  NOR2_X1 U8374 ( .A1(n7791), .A2(n12046), .ZN(n12045) );
  AND2_X1 U8375 ( .A1(n12026), .A2(n11534), .ZN(n12046) );
  NAND2_X1 U8376 ( .A1(n7792), .A2(n7247), .ZN(n7557) );
  NAND2_X1 U8377 ( .A1(n12046), .A2(n7558), .ZN(n7556) );
  INV_X1 U8378 ( .A(n15832), .ZN(n7558) );
  NOR2_X1 U8379 ( .A1(n12061), .A2(n15857), .ZN(n12062) );
  INV_X1 U8380 ( .A(n13590), .ZN(n13589) );
  INV_X1 U8381 ( .A(n7784), .ZN(n12050) );
  NAND2_X1 U8382 ( .A1(n13590), .A2(n13605), .ZN(n13592) );
  NOR2_X1 U8383 ( .A1(n13633), .A2(n7770), .ZN(n13632) );
  AND2_X1 U8384 ( .A1(n7768), .A2(n7770), .ZN(n13636) );
  NAND2_X1 U8385 ( .A1(n7789), .A2(n7376), .ZN(n13643) );
  XNOR2_X1 U8386 ( .A(n13679), .B(n7458), .ZN(n13659) );
  OR2_X1 U8387 ( .A1(n13697), .A2(n13696), .ZN(n13725) );
  XNOR2_X1 U8388 ( .A(n7781), .B(n13710), .ZN(n13697) );
  AOI21_X1 U8389 ( .B1(n12986), .B2(n7843), .A(n7842), .ZN(n7841) );
  INV_X1 U8390 ( .A(n13507), .ZN(n7842) );
  AND2_X1 U8391 ( .A1(n12962), .A2(n12961), .ZN(n12988) );
  OR2_X1 U8392 ( .A1(n8785), .A2(n13757), .ZN(n13776) );
  INV_X1 U8393 ( .A(n13771), .ZN(n13765) );
  OR2_X1 U8394 ( .A1(n12468), .A2(n8327), .ZN(n8767) );
  AND2_X1 U8395 ( .A1(n13493), .A2(n13491), .ZN(n13811) );
  AND4_X1 U8396 ( .A1(n8755), .A2(n8754), .A3(n8753), .A4(n8752), .ZN(n13813)
         );
  NAND2_X1 U8397 ( .A1(n13839), .A2(n13487), .ZN(n13823) );
  NAND2_X1 U8398 ( .A1(n14039), .A2(n7492), .ZN(n7491) );
  OR2_X1 U8399 ( .A1(n13903), .A2(n13881), .ZN(n8236) );
  INV_X1 U8400 ( .A(n13857), .ZN(n13880) );
  AND2_X1 U8401 ( .A1(n7866), .A2(n7867), .ZN(n13877) );
  NAND2_X1 U8402 ( .A1(n12976), .A2(n8237), .ZN(n7866) );
  AND2_X1 U8403 ( .A1(n12973), .A2(n12972), .ZN(n13893) );
  NAND2_X1 U8404 ( .A1(n8190), .A2(n8189), .ZN(n8188) );
  INV_X1 U8405 ( .A(n8193), .ZN(n8189) );
  AND2_X1 U8406 ( .A1(n8535), .A2(n8534), .ZN(n12564) );
  AND2_X1 U8407 ( .A1(n13439), .A2(n13443), .ZN(n13532) );
  AOI21_X1 U8408 ( .B1(n12169), .B2(n7853), .A(n7244), .ZN(n7852) );
  NAND2_X1 U8409 ( .A1(n7851), .A2(n7853), .ZN(n7850) );
  NAND2_X1 U8410 ( .A1(n8176), .A2(n12168), .ZN(n12245) );
  NOR2_X1 U8411 ( .A1(n8427), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8436) );
  OR2_X1 U8412 ( .A1(n8399), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8427) );
  NAND2_X1 U8413 ( .A1(n11885), .A2(n13403), .ZN(n11959) );
  NAND2_X1 U8414 ( .A1(n8181), .A2(n11651), .ZN(n11652) );
  INV_X1 U8415 ( .A(n11648), .ZN(n13528) );
  NAND2_X1 U8416 ( .A1(n11901), .A2(n11625), .ZN(n11649) );
  NAND2_X1 U8417 ( .A1(n11627), .A2(n13383), .ZN(n13391) );
  INV_X1 U8418 ( .A(n13885), .ZN(n13994) );
  NAND2_X1 U8419 ( .A1(n11265), .A2(n13509), .ZN(n13944) );
  INV_X1 U8420 ( .A(n13997), .ZN(n13946) );
  OR2_X1 U8421 ( .A1(n13760), .A2(n13759), .ZN(n14084) );
  NAND2_X1 U8422 ( .A1(n8748), .A2(n8747), .ZN(n13494) );
  OR2_X1 U8423 ( .A1(n12960), .A2(n13103), .ZN(n8747) );
  NAND2_X1 U8424 ( .A1(n8677), .A2(n8676), .ZN(n12977) );
  AND2_X1 U8425 ( .A1(n13885), .A2(n16011), .ZN(n14058) );
  NAND2_X1 U8426 ( .A1(n7855), .A2(n13426), .ZN(n12202) );
  NAND2_X1 U8427 ( .A1(n12242), .A2(n13527), .ZN(n7855) );
  NAND2_X1 U8428 ( .A1(n8778), .A2(n8777), .ZN(n8780) );
  NAND2_X1 U8429 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n8113), .ZN(n8112) );
  INV_X1 U8430 ( .A(n8745), .ZN(n8110) );
  XNOR2_X1 U8431 ( .A(n8806), .B(n8805), .ZN(n10625) );
  AND2_X1 U8432 ( .A1(n7259), .A2(n7849), .ZN(n7848) );
  NOR2_X1 U8433 ( .A1(n8291), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n7563) );
  INV_X1 U8434 ( .A(n7565), .ZN(n7564) );
  NAND2_X1 U8435 ( .A1(n8292), .A2(n8298), .ZN(n7565) );
  OR2_X1 U8436 ( .A1(n8290), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8591) );
  AOI21_X1 U8437 ( .B1(n8642), .B2(n8095), .A(n7373), .ZN(n8094) );
  NAND2_X1 U8438 ( .A1(n8626), .A2(n8093), .ZN(n8092) );
  INV_X1 U8439 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8298) );
  INV_X1 U8440 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8607) );
  INV_X1 U8441 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U8442 ( .A1(n7508), .A2(n8257), .ZN(n8290) );
  INV_X1 U8443 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8257) );
  AND2_X1 U8444 ( .A1(n8533), .A2(n8510), .ZN(n8531) );
  INV_X1 U8445 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8460) );
  AND2_X1 U8446 ( .A1(n8466), .A2(n8451), .ZN(n8463) );
  NAND2_X1 U8447 ( .A1(n8118), .A2(n8450), .ZN(n8465) );
  INV_X1 U8448 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8449) );
  XNOR2_X1 U8449 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8447) );
  OR2_X1 U8450 ( .A1(n8381), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U8451 ( .A1(n8407), .A2(n8380), .ZN(n8405) );
  NAND2_X1 U8452 ( .A1(n8876), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U8453 ( .A1(n7874), .A2(n7248), .ZN(n11226) );
  NOR2_X1 U8454 ( .A1(n11215), .A2(n7876), .ZN(n7875) );
  NAND2_X1 U8455 ( .A1(n14197), .A2(n7886), .ZN(n7885) );
  INV_X1 U8456 ( .A(n14199), .ZN(n7886) );
  NAND2_X1 U8457 ( .A1(n9097), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9121) );
  INV_X1 U8458 ( .A(n9098), .ZN(n9097) );
  INV_X1 U8459 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9120) );
  OR2_X1 U8460 ( .A1(n9121), .A2(n9120), .ZN(n9152) );
  NAND2_X1 U8461 ( .A1(n7269), .A2(n11592), .ZN(n7878) );
  NAND2_X1 U8462 ( .A1(n11309), .A2(n11308), .ZN(n11310) );
  NAND2_X1 U8463 ( .A1(n7904), .A2(n7910), .ZN(n7903) );
  AOI21_X1 U8464 ( .B1(n14216), .B2(n14173), .A(n7907), .ZN(n7906) );
  INV_X1 U8465 ( .A(n14178), .ZN(n7907) );
  NAND2_X1 U8466 ( .A1(n14324), .A2(n7905), .ZN(n7902) );
  NAND2_X1 U8467 ( .A1(n10931), .A2(n10930), .ZN(n14264) );
  NAND2_X1 U8468 ( .A1(n11310), .A2(n11311), .ZN(n11365) );
  NAND2_X1 U8469 ( .A1(n14264), .A2(n14265), .ZN(n14263) );
  INV_X1 U8470 ( .A(n14453), .ZN(n14338) );
  AND2_X1 U8471 ( .A1(n7892), .A2(n7896), .ZN(n7891) );
  NAND2_X1 U8472 ( .A1(n12275), .A2(n7263), .ZN(n7892) );
  NAND2_X1 U8473 ( .A1(n12277), .A2(n12275), .ZN(n7890) );
  NOR2_X1 U8474 ( .A1(n8886), .A2(n11375), .ZN(n10655) );
  NAND2_X1 U8475 ( .A1(n9640), .A2(n8133), .ZN(n8131) );
  NOR2_X1 U8476 ( .A1(n9639), .A2(n9677), .ZN(n8132) );
  INV_X1 U8477 ( .A(n8886), .ZN(n9710) );
  OR2_X1 U8478 ( .A1(n9064), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9177) );
  OR2_X1 U8479 ( .A1(n9251), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n9281) );
  OR2_X1 U8480 ( .A1(n14545), .A2(n9643), .ZN(n14522) );
  AOI21_X1 U8481 ( .B1(n14552), .B2(n7808), .A(n7299), .ZN(n7807) );
  INV_X1 U8482 ( .A(n14518), .ZN(n7808) );
  NAND2_X1 U8483 ( .A1(n7396), .A2(n14552), .ZN(n7806) );
  INV_X1 U8484 ( .A(n14519), .ZN(n7396) );
  NAND2_X1 U8485 ( .A1(n7806), .A2(n7804), .ZN(n14538) );
  NOR2_X1 U8486 ( .A1(n14535), .A2(n7805), .ZN(n7804) );
  INV_X1 U8487 ( .A(n7807), .ZN(n7805) );
  NOR2_X1 U8488 ( .A1(n14552), .A2(n8062), .ZN(n8061) );
  INV_X1 U8489 ( .A(n14485), .ZN(n8062) );
  NOR2_X1 U8490 ( .A1(n14606), .A2(n14759), .ZN(n14593) );
  NAND2_X1 U8491 ( .A1(n9455), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9477) );
  INV_X1 U8492 ( .A(n9457), .ZN(n9455) );
  NAND2_X1 U8493 ( .A1(n7707), .A2(n7706), .ZN(n14606) );
  AND2_X1 U8494 ( .A1(n14618), .A2(n14479), .ZN(n14601) );
  INV_X1 U8495 ( .A(n7707), .ZN(n14619) );
  INV_X1 U8496 ( .A(n7693), .ZN(n7692) );
  OAI21_X1 U8497 ( .B1(n14630), .B2(n7694), .A(n14477), .ZN(n7693) );
  NAND2_X1 U8498 ( .A1(n7275), .A2(n8072), .ZN(n7694) );
  NAND2_X1 U8499 ( .A1(n14645), .A2(n7261), .ZN(n7691) );
  NAND2_X1 U8500 ( .A1(n7691), .A2(n7689), .ZN(n14618) );
  AND2_X1 U8501 ( .A1(n7692), .A2(n7690), .ZN(n7689) );
  NAND2_X1 U8502 ( .A1(n9357), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9386) );
  NOR2_X2 U8503 ( .A1(n14681), .A2(n14789), .ZN(n14660) );
  NAND2_X1 U8504 ( .A1(n12354), .A2(n12353), .ZN(n12424) );
  NAND2_X1 U8505 ( .A1(n9229), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9257) );
  OR3_X1 U8506 ( .A1(n9204), .A2(n9203), .A3(n12288), .ZN(n9230) );
  NOR2_X1 U8507 ( .A1(n12120), .A2(n16111), .ZN(n12359) );
  NAND2_X1 U8508 ( .A1(n9180), .A2(n9179), .ZN(n12179) );
  NAND2_X1 U8509 ( .A1(n11867), .A2(n12294), .ZN(n12019) );
  INV_X1 U8510 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9068) );
  OR2_X1 U8511 ( .A1(n9069), .A2(n9068), .ZN(n9098) );
  INV_X1 U8512 ( .A(n10691), .ZN(n7798) );
  NAND2_X1 U8513 ( .A1(n10590), .A2(n7798), .ZN(n10688) );
  INV_X1 U8514 ( .A(n8054), .ZN(n8053) );
  OAI22_X1 U8515 ( .A1(n9621), .A2(n8056), .B1(n10428), .B2(n8055), .ZN(n8054)
         );
  NAND2_X1 U8516 ( .A1(n10597), .A2(n10596), .ZN(n10692) );
  NAND2_X1 U8517 ( .A1(n14716), .A2(n12410), .ZN(n10652) );
  NOR2_X1 U8518 ( .A1(n7449), .A2(n10775), .ZN(n10493) );
  NAND2_X1 U8519 ( .A1(n14704), .A2(n14467), .ZN(n14690) );
  NAND2_X1 U8520 ( .A1(n8057), .A2(n7305), .ZN(n12126) );
  INV_X1 U8521 ( .A(n14807), .ZN(n14803) );
  INV_X1 U8522 ( .A(n11714), .ZN(n11713) );
  NAND2_X1 U8523 ( .A1(n9066), .A2(n9065), .ZN(n16003) );
  NAND2_X1 U8524 ( .A1(n8850), .A2(n8849), .ZN(n9696) );
  INV_X1 U8525 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8854) );
  AND2_X1 U8526 ( .A1(n9194), .A2(n9017), .ZN(n9041) );
  INV_X1 U8527 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8836) );
  NOR2_X1 U8528 ( .A1(n10102), .A2(n10101), .ZN(n10120) );
  AND2_X1 U8529 ( .A1(n10120), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10142) );
  AOI21_X1 U8530 ( .B1(n8044), .B2(n14944), .A(n8047), .ZN(n8043) );
  AND2_X1 U8531 ( .A1(n10194), .A2(n10195), .ZN(n8047) );
  NOR2_X1 U8532 ( .A1(n10018), .A2(n10017), .ZN(n10057) );
  NAND2_X1 U8533 ( .A1(n12258), .A2(n7301), .ZN(n12553) );
  XNOR2_X1 U8534 ( .A(n9886), .B(n14954), .ZN(n9889) );
  NOR2_X1 U8535 ( .A1(n9834), .A2(n9816), .ZN(n10163) );
  NAND2_X1 U8536 ( .A1(n9951), .A2(n9952), .ZN(n11294) );
  OR2_X1 U8537 ( .A1(n10387), .A2(n10386), .ZN(n7639) );
  NOR2_X1 U8538 ( .A1(n10613), .A2(n7632), .ZN(n10617) );
  AND2_X1 U8539 ( .A1(n10614), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7632) );
  NAND2_X1 U8540 ( .A1(n10617), .A2(n10616), .ZN(n11158) );
  NAND2_X1 U8541 ( .A1(n11463), .A2(n7624), .ZN(n11834) );
  OR2_X1 U8542 ( .A1(n11464), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7624) );
  OR2_X1 U8543 ( .A1(n15108), .A2(n15107), .ZN(n7629) );
  NAND2_X1 U8544 ( .A1(n7629), .A2(n7628), .ZN(n7627) );
  NAND2_X1 U8545 ( .A1(n15124), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7628) );
  AND2_X1 U8546 ( .A1(n7627), .A2(n15138), .ZN(n15134) );
  NAND2_X1 U8547 ( .A1(n15165), .A2(n15397), .ZN(n15159) );
  AOI21_X1 U8548 ( .B1(n12825), .B2(n7232), .A(n12824), .ZN(n15403) );
  NAND2_X1 U8549 ( .A1(n15211), .A2(n15198), .ZN(n15192) );
  NAND2_X1 U8550 ( .A1(n15425), .A2(n15191), .ZN(n7968) );
  AOI21_X1 U8551 ( .B1(n7925), .B2(n7923), .A(n7316), .ZN(n7922) );
  NAND2_X1 U8552 ( .A1(n15240), .A2(n7925), .ZN(n7579) );
  NAND2_X1 U8553 ( .A1(n15222), .A2(n7966), .ZN(n7969) );
  OR2_X1 U8554 ( .A1(n15429), .A2(n14929), .ZN(n7970) );
  NAND2_X1 U8555 ( .A1(n12664), .A2(n14969), .ZN(n7461) );
  NOR3_X1 U8556 ( .A1(n15326), .A2(n15444), .A3(n7742), .ZN(n15269) );
  OR2_X1 U8557 ( .A1(n10180), .A2(n10179), .ZN(n10182) );
  NOR2_X1 U8558 ( .A1(n10182), .A2(n15018), .ZN(n9804) );
  AOI21_X1 U8559 ( .B1(n15335), .B2(n15338), .A(n8249), .ZN(n15323) );
  NAND2_X1 U8560 ( .A1(n11981), .A2(n12737), .ZN(n7938) );
  NOR2_X1 U8561 ( .A1(n7264), .A2(n7948), .ZN(n7947) );
  OR2_X1 U8562 ( .A1(n9977), .A2(n9976), .ZN(n10000) );
  OR2_X1 U8563 ( .A1(n10000), .A2(n9999), .ZN(n10018) );
  INV_X1 U8564 ( .A(n12855), .ZN(n11202) );
  INV_X1 U8565 ( .A(n12683), .ZN(n10909) );
  NAND2_X1 U8566 ( .A1(n10227), .A2(n15879), .ZN(n16123) );
  NAND2_X1 U8567 ( .A1(n9767), .A2(n9756), .ZN(n8208) );
  XNOR2_X1 U8568 ( .A(n9619), .B(n9618), .ZN(n12825) );
  OAI21_X1 U8569 ( .B1(n9554), .B2(n9553), .A(n9555), .ZN(n9577) );
  AND2_X1 U8570 ( .A1(n9559), .A2(n9558), .ZN(n9576) );
  NAND2_X1 U8571 ( .A1(n9577), .A2(n9576), .ZN(n9579) );
  XNOR2_X1 U8572 ( .A(n9554), .B(n9553), .ZN(n14867) );
  XNOR2_X1 U8573 ( .A(n9742), .B(P1_IR_REG_26__SCAN_IN), .ZN(n10200) );
  XNOR2_X1 U8574 ( .A(n9517), .B(n9516), .ZN(n12588) );
  XNOR2_X1 U8575 ( .A(n9489), .B(n9474), .ZN(n12598) );
  NAND2_X1 U8576 ( .A1(n9784), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9786) );
  XNOR2_X1 U8577 ( .A(n9352), .B(n9351), .ZN(n11421) );
  NAND2_X1 U8578 ( .A1(n7998), .A2(n7255), .ZN(n9325) );
  NAND2_X1 U8579 ( .A1(n7998), .A2(n9296), .ZN(n9303) );
  XNOR2_X1 U8580 ( .A(n9248), .B(n9247), .ZN(n11012) );
  NAND2_X1 U8581 ( .A1(n8010), .A2(n9142), .ZN(n9166) );
  NAND2_X1 U8582 ( .A1(n9135), .A2(n9134), .ZN(n8010) );
  OR2_X1 U8583 ( .A1(n9944), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9972) );
  NAND2_X1 U8584 ( .A1(n9037), .A2(n9036), .ZN(n7973) );
  XNOR2_X1 U8585 ( .A(n9037), .B(n9035), .ZN(n10269) );
  NAND2_X1 U8586 ( .A1(n8926), .A2(n8876), .ZN(n7417) );
  INV_X1 U8587 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n15657) );
  INV_X1 U8588 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7722) );
  XNOR2_X1 U8589 ( .A(n15693), .B(n15682), .ZN(n15689) );
  OAI22_X1 U8590 ( .A1(n15702), .A2(n15701), .B1(P3_ADDR_REG_5__SCAN_IN), .B2(
        n15700), .ZN(n15705) );
  INV_X1 U8591 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n15700) );
  AND2_X1 U8592 ( .A1(n15716), .A2(n15717), .ZN(n15718) );
  INV_X1 U8593 ( .A(n7712), .ZN(n15715) );
  AOI21_X1 U8594 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15726), .A(n15725), .ZN(
        n15736) );
  OAI21_X1 U8595 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n15833), .A(n15746), .ZN(
        n15756) );
  NAND2_X1 U8596 ( .A1(n15762), .A2(n15763), .ZN(n15774) );
  NAND2_X1 U8597 ( .A1(n11941), .A2(n8417), .ZN(n11815) );
  OAI21_X1 U8598 ( .B1(n7535), .B2(n7525), .A(n7524), .ZN(n13223) );
  AOI21_X1 U8599 ( .B1(n7526), .B2(n7533), .A(n8167), .ZN(n7524) );
  INV_X1 U8600 ( .A(n7526), .ZN(n7525) );
  NAND2_X1 U8601 ( .A1(n12230), .A2(n7547), .ZN(n12389) );
  NAND2_X1 U8602 ( .A1(n11208), .A2(n11207), .ZN(n11206) );
  AND4_X2 U8603 ( .A1(n8366), .A2(n8365), .A3(n8364), .A4(n8363), .ZN(n11904)
         );
  CLKBUF_X1 U8604 ( .A(n11620), .Z(n11905) );
  NAND2_X1 U8605 ( .A1(n13323), .A2(n8640), .ZN(n13249) );
  OAI21_X1 U8606 ( .B1(n13325), .B2(n8150), .A(n8148), .ZN(n13247) );
  NAND2_X1 U8607 ( .A1(n7527), .A2(n7528), .ZN(n13332) );
  NAND2_X1 U8608 ( .A1(n7535), .A2(n7530), .ZN(n7527) );
  NAND2_X1 U8609 ( .A1(n8160), .A2(n8164), .ZN(n8159) );
  NAND2_X1 U8610 ( .A1(n7241), .A2(n7260), .ZN(n8164) );
  AND4_X1 U8611 ( .A1(n8717), .A2(n8716), .A3(n8715), .A4(n8714), .ZN(n13812)
         );
  NAND2_X1 U8612 ( .A1(n7535), .A2(n7267), .ZN(n13263) );
  NAND2_X1 U8613 ( .A1(n13342), .A2(n8586), .ZN(n13272) );
  NAND2_X1 U8614 ( .A1(n11385), .A2(n8376), .ZN(n11478) );
  NAND2_X1 U8615 ( .A1(n11206), .A2(n8358), .ZN(n11387) );
  NAND2_X1 U8616 ( .A1(n12000), .A2(n8456), .ZN(n12232) );
  AOI21_X1 U8617 ( .B1(n13278), .B2(n7543), .A(n7541), .ZN(n7540) );
  NAND2_X1 U8618 ( .A1(n7542), .A2(n13299), .ZN(n7541) );
  NAND2_X1 U8619 ( .A1(n7543), .A2(n7545), .ZN(n7542) );
  OAI21_X1 U8620 ( .B1(n13278), .B2(n7545), .A(n7543), .ZN(n13300) );
  NAND2_X1 U8621 ( .A1(n8198), .A2(n8197), .ZN(n13306) );
  OAI21_X1 U8622 ( .B1(n12000), .B2(n7548), .A(n7546), .ZN(n12471) );
  AOI21_X1 U8623 ( .B1(n8178), .B2(n7547), .A(n7249), .ZN(n7546) );
  NAND2_X1 U8624 ( .A1(n13278), .A2(n8623), .ZN(n13325) );
  NAND2_X1 U8625 ( .A1(n13325), .A2(n13324), .ZN(n13323) );
  OAI21_X1 U8626 ( .B1(n8185), .B2(n8184), .A(n11477), .ZN(n8183) );
  AND3_X1 U8627 ( .A1(n8414), .A2(n8413), .A3(n8412), .ZN(n13411) );
  AND4_X1 U8628 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), .ZN(n13348)
         );
  NAND2_X1 U8629 ( .A1(n13341), .A2(n8584), .ZN(n13342) );
  NAND2_X1 U8630 ( .A1(n8813), .A2(n8812), .ZN(n13343) );
  OAI211_X1 U8631 ( .C1(n8081), .C2(n11179), .A(n8080), .B(n8079), .ZN(n8078)
         );
  NAND2_X1 U8632 ( .A1(n7274), .A2(n7568), .ZN(n8079) );
  NAND2_X1 U8633 ( .A1(n8081), .A2(n11683), .ZN(n8080) );
  NAND2_X1 U8634 ( .A1(n8083), .A2(n8082), .ZN(n8081) );
  INV_X1 U8635 ( .A(n13813), .ZN(n13575) );
  AND4_X1 U8636 ( .A1(n8742), .A2(n8741), .A3(n8740), .A4(n8739), .ZN(n13827)
         );
  INV_X1 U8637 ( .A(n13812), .ZN(n13843) );
  INV_X1 U8638 ( .A(n13943), .ZN(n13914) );
  INV_X1 U8639 ( .A(n13348), .ZN(n13959) );
  INV_X1 U8640 ( .A(n8514), .ZN(n13998) );
  INV_X1 U8641 ( .A(n11904), .ZN(n13583) );
  INV_X1 U8642 ( .A(n11673), .ZN(n13584) );
  OR2_X1 U8643 ( .A1(n10711), .A2(n10710), .ZN(n10818) );
  NAND2_X1 U8644 ( .A1(n10884), .A2(n10882), .ZN(n7753) );
  NAND2_X1 U8645 ( .A1(n11138), .A2(n7777), .ZN(n10978) );
  INV_X1 U8646 ( .A(n7467), .ZN(n11496) );
  INV_X1 U8647 ( .A(n7761), .ZN(n11501) );
  INV_X1 U8648 ( .A(n11537), .ZN(n11536) );
  NAND2_X1 U8649 ( .A1(n7792), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7791) );
  INV_X1 U8650 ( .A(n12046), .ZN(n7793) );
  INV_X1 U8651 ( .A(n7759), .ZN(n15841) );
  NAND2_X1 U8652 ( .A1(n7557), .A2(n7556), .ZN(n15831) );
  NOR2_X1 U8653 ( .A1(n13594), .A2(n13593), .ZN(n13623) );
  OR2_X1 U8654 ( .A1(n13610), .A2(n13609), .ZN(n13622) );
  NAND2_X1 U8655 ( .A1(n7766), .A2(n13666), .ZN(n13649) );
  AND2_X1 U8656 ( .A1(n13666), .A2(n7767), .ZN(n13669) );
  AOI21_X1 U8657 ( .B1(n13721), .B2(n13720), .A(n13719), .ZN(n13739) );
  XNOR2_X1 U8658 ( .A(n7552), .B(n7551), .ZN(n7550) );
  INV_X1 U8659 ( .A(n13747), .ZN(n7551) );
  NAND2_X1 U8660 ( .A1(n13742), .A2(n13741), .ZN(n7552) );
  NOR2_X1 U8661 ( .A1(n13753), .A2(n7554), .ZN(n7553) );
  NAND2_X1 U8662 ( .A1(n13745), .A2(n7555), .ZN(n7554) );
  XNOR2_X1 U8663 ( .A(n7408), .B(n12987), .ZN(n12969) );
  NAND2_X1 U8664 ( .A1(n13770), .A2(n7284), .ZN(n7408) );
  INV_X1 U8665 ( .A(n12988), .ZN(n13218) );
  NAND2_X1 U8666 ( .A1(n12979), .A2(n13376), .ZN(n13837) );
  NAND2_X1 U8667 ( .A1(n7859), .A2(n7860), .ZN(n13868) );
  NAND2_X1 U8668 ( .A1(n13933), .A2(n7864), .ZN(n7859) );
  AND2_X1 U8669 ( .A1(n13938), .A2(n8191), .ZN(n13923) );
  OAI21_X1 U8670 ( .B1(n13954), .B2(n7840), .A(n7838), .ZN(n13936) );
  NAND2_X1 U8671 ( .A1(n13952), .A2(n13459), .ZN(n13937) );
  NAND2_X1 U8672 ( .A1(n12938), .A2(n12937), .ZN(n13973) );
  INV_X1 U8673 ( .A(n12564), .ZN(n16055) );
  INV_X1 U8674 ( .A(n13411), .ZN(n15939) );
  NAND2_X1 U8675 ( .A1(n13966), .A2(n11640), .ZN(n12254) );
  INV_X1 U8676 ( .A(n12254), .ZN(n14008) );
  INV_X1 U8677 ( .A(n14004), .ZN(n13983) );
  AOI21_X1 U8678 ( .B1(n12989), .B2(n16061), .A(n7370), .ZN(n7510) );
  INV_X1 U8679 ( .A(n13555), .ZN(n14086) );
  INV_X1 U8680 ( .A(n13513), .ZN(n14089) );
  INV_X1 U8681 ( .A(n13494), .ZN(n14100) );
  INV_X1 U8682 ( .A(n12949), .ZN(n14104) );
  INV_X1 U8683 ( .A(n12977), .ZN(n14114) );
  INV_X1 U8684 ( .A(n13468), .ZN(n14129) );
  NAND2_X1 U8685 ( .A1(n8575), .A2(n8574), .ZN(n14133) );
  INV_X1 U8686 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8303) );
  MUX2_X1 U8687 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8284), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8285) );
  NAND2_X1 U8688 ( .A1(n8111), .A2(n8734), .ZN(n8746) );
  NAND2_X1 U8689 ( .A1(n8283), .A2(n8281), .ZN(n12349) );
  INV_X1 U8690 ( .A(n8262), .ZN(n8276) );
  NAND2_X1 U8691 ( .A1(n8708), .A2(n8734), .ZN(n8733) );
  NAND2_X1 U8692 ( .A1(n8105), .A2(n8706), .ZN(n8725) );
  NAND2_X1 U8693 ( .A1(n8705), .A2(n8704), .ZN(n8105) );
  XNOR2_X1 U8694 ( .A(n8808), .B(P3_IR_REG_22__SCAN_IN), .ZN(n13565) );
  NAND2_X1 U8695 ( .A1(n7259), .A2(n7508), .ZN(n8807) );
  XNOR2_X1 U8696 ( .A(n8294), .B(n8293), .ZN(n13388) );
  INV_X1 U8697 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8293) );
  OAI21_X1 U8698 ( .B1(n8591), .B2(n7562), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8294) );
  NAND2_X1 U8699 ( .A1(n7564), .A2(n7563), .ZN(n7562) );
  NAND2_X1 U8700 ( .A1(n7331), .A2(n8117), .ZN(n8675) );
  INV_X1 U8701 ( .A(SI_19_), .ZN(n13092) );
  INV_X1 U8702 ( .A(SI_18_), .ZN(n13093) );
  NAND2_X1 U8703 ( .A1(n8096), .A2(n8627), .ZN(n8643) );
  NAND2_X1 U8704 ( .A1(n8626), .A2(n8625), .ZN(n8096) );
  INV_X1 U8705 ( .A(SI_15_), .ZN(n13122) );
  INV_X1 U8706 ( .A(SI_14_), .ZN(n13124) );
  NAND2_X1 U8707 ( .A1(n7498), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8100) );
  INV_X1 U8708 ( .A(SI_13_), .ZN(n13121) );
  NAND2_X1 U8709 ( .A1(n8255), .A2(n8418), .ZN(n8540) );
  INV_X1 U8710 ( .A(SI_12_), .ZN(n13019) );
  INV_X1 U8711 ( .A(SI_10_), .ZN(n13133) );
  INV_X1 U8712 ( .A(SI_9_), .ZN(n13136) );
  INV_X1 U8713 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8444) );
  OAI21_X1 U8714 ( .B1(n14324), .B2(n14173), .A(n14216), .ZN(n14299) );
  AND2_X1 U8715 ( .A1(n14236), .A2(n7400), .ZN(n7399) );
  NOR2_X1 U8716 ( .A1(n7401), .A2(n14353), .ZN(n7400) );
  INV_X1 U8717 ( .A(n14237), .ZN(n7401) );
  INV_X1 U8718 ( .A(n14239), .ZN(n7398) );
  NAND2_X1 U8719 ( .A1(n7902), .A2(n7903), .ZN(n14300) );
  INV_X1 U8720 ( .A(n7437), .ZN(n12296) );
  NAND2_X1 U8721 ( .A1(n14187), .A2(n7443), .ZN(n7442) );
  INV_X1 U8722 ( .A(n8241), .ZN(n7443) );
  NAND2_X1 U8723 ( .A1(n14290), .A2(n14289), .ZN(n14288) );
  NAND2_X1 U8724 ( .A1(n11365), .A2(n11364), .ZN(n11594) );
  NAND2_X1 U8725 ( .A1(n10380), .A2(n9620), .ZN(n7647) );
  AND2_X1 U8726 ( .A1(n10661), .A2(n10748), .ZN(n7873) );
  OR2_X1 U8727 ( .A1(n10659), .A2(n10660), .ZN(n10661) );
  INV_X1 U8728 ( .A(n14341), .ZN(n14348) );
  OR2_X1 U8729 ( .A1(n14165), .A2(n14166), .ZN(n7485) );
  NAND2_X1 U8730 ( .A1(n9331), .A2(n9330), .ZN(n14698) );
  NAND2_X1 U8731 ( .A1(n14263), .A2(n10937), .ZN(n11214) );
  NAND2_X1 U8732 ( .A1(n7890), .A2(n7891), .ZN(n14355) );
  NAND2_X1 U8733 ( .A1(n9484), .A2(n9483), .ZN(n14480) );
  OR3_X1 U8734 ( .A1(n9264), .A2(n9263), .A3(n9262), .ZN(n14362) );
  NAND4_X2 U8735 ( .A1(n8948), .A2(n8947), .A3(n8946), .A4(n8945), .ZN(n14374)
         );
  OR2_X1 U8736 ( .A1(n7207), .A2(n11880), .ZN(n8901) );
  OR2_X2 U8737 ( .A1(n10762), .A2(n9750), .ZN(n14376) );
  XNOR2_X1 U8738 ( .A(n14457), .B(n7702), .ZN(n14449) );
  NAND2_X1 U8739 ( .A1(n9601), .A2(n9600), .ZN(n14461) );
  AOI21_X1 U8740 ( .B1(n14551), .B2(n14710), .A(n14550), .ZN(n14747) );
  NAND2_X1 U8741 ( .A1(n14519), .A2(n14518), .ZN(n14549) );
  AND2_X1 U8742 ( .A1(n9521), .A2(n9520), .ZN(n14573) );
  OAI21_X1 U8743 ( .B1(n7811), .B2(n7673), .A(n7672), .ZN(n14575) );
  OAI21_X1 U8744 ( .B1(n7811), .B2(n7810), .A(n7809), .ZN(n14582) );
  INV_X1 U8745 ( .A(n7812), .ZN(n14598) );
  AOI21_X1 U8746 ( .B1(n14614), .B2(n14617), .A(n7815), .ZN(n7812) );
  NAND2_X1 U8747 ( .A1(n7696), .A2(n7261), .ZN(n14631) );
  NAND2_X1 U8748 ( .A1(n7656), .A2(n7657), .ZN(n14627) );
  NAND2_X1 U8749 ( .A1(n7660), .A2(n14506), .ZN(n14647) );
  OR2_X1 U8750 ( .A1(n14668), .A2(n14504), .ZN(n7660) );
  NAND2_X1 U8751 ( .A1(n7649), .A2(n7650), .ZN(n14677) );
  NAND2_X1 U8752 ( .A1(n14711), .A2(n14496), .ZN(n14692) );
  NOR2_X1 U8753 ( .A1(n8067), .A2(n8066), .ZN(n14705) );
  INV_X1 U8754 ( .A(n14464), .ZN(n8066) );
  INV_X1 U8755 ( .A(n14465), .ZN(n8067) );
  NAND2_X1 U8756 ( .A1(n7667), .A2(n12426), .ZN(n12428) );
  NAND2_X1 U8757 ( .A1(n9201), .A2(n9200), .ZN(n12192) );
  NAND2_X1 U8758 ( .A1(n7817), .A2(n7818), .ZN(n11862) );
  NAND2_X1 U8759 ( .A1(n11722), .A2(n11721), .ZN(n11859) );
  NAND2_X1 U8760 ( .A1(n11508), .A2(n11507), .ZN(n11750) );
  OAI21_X1 U8761 ( .B1(n11512), .B2(n7268), .A(n7803), .ZN(n11752) );
  NAND2_X1 U8762 ( .A1(n7825), .A2(n10831), .ZN(n11049) );
  OR2_X1 U8763 ( .A1(n15891), .A2(n11737), .ZN(n14661) );
  NAND2_X1 U8764 ( .A1(n10688), .A2(n7797), .ZN(n12105) );
  OR2_X1 U8765 ( .A1(n10590), .A2(n7798), .ZN(n7797) );
  INV_X1 U8766 ( .A(n14728), .ZN(n14642) );
  INV_X1 U8767 ( .A(n10683), .ZN(n10490) );
  INV_X1 U8768 ( .A(n14661), .ZN(n14722) );
  OAI211_X1 U8769 ( .C1(n14739), .C2(n16006), .A(n14738), .B(n14737), .ZN(
        n14819) );
  AOI21_X1 U8770 ( .B1(n7830), .B2(n14710), .A(n7358), .ZN(n14738) );
  NAND2_X1 U8771 ( .A1(n16109), .A2(n8075), .ZN(n12420) );
  AND2_X1 U8772 ( .A1(n16109), .A2(n12356), .ZN(n12358) );
  AND2_X1 U8773 ( .A1(n8057), .A2(n8058), .ZN(n12008) );
  NAND2_X1 U8774 ( .A1(n11854), .A2(n11853), .ZN(n11856) );
  NAND2_X1 U8775 ( .A1(n11707), .A2(n11706), .ZN(n11708) );
  NAND2_X1 U8776 ( .A1(n11402), .A2(n11401), .ZN(n11404) );
  NAND2_X1 U8777 ( .A1(n10494), .A2(n10775), .ZN(n9646) );
  AND2_X1 U8778 ( .A1(n10762), .A2(n9749), .ZN(n15525) );
  INV_X1 U8779 ( .A(n8872), .ZN(n14860) );
  OR2_X1 U8780 ( .A1(n8869), .A2(n8878), .ZN(n7698) );
  NAND2_X1 U8781 ( .A1(n8882), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8052) );
  XNOR2_X1 U8782 ( .A(n9699), .B(P2_IR_REG_26__SCAN_IN), .ZN(n12451) );
  NAND2_X1 U8783 ( .A1(n9703), .A2(n9702), .ZN(n12256) );
  XNOR2_X1 U8784 ( .A(n9705), .B(n9704), .ZN(n12199) );
  INV_X1 U8785 ( .A(n12410), .ZN(n12414) );
  INV_X1 U8786 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11040) );
  INV_X1 U8787 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10923) );
  INV_X1 U8788 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10397) );
  INV_X1 U8789 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10424) );
  INV_X1 U8790 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10301) );
  INV_X1 U8791 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10271) );
  INV_X1 U8792 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10262) );
  INV_X1 U8793 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10259) );
  AND2_X1 U8794 ( .A1(n10264), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10214) );
  INV_X1 U8795 ( .A(n12725), .ZN(n15957) );
  NAND2_X1 U8796 ( .A1(n11456), .A2(n11455), .ZN(n11454) );
  AND2_X1 U8797 ( .A1(n12508), .A2(n10115), .ZN(n16084) );
  NAND2_X1 U8798 ( .A1(n12508), .A2(n8041), .ZN(n16083) );
  NAND2_X1 U8799 ( .A1(n8025), .A2(n8027), .ZN(n14925) );
  INV_X1 U8800 ( .A(n14887), .ZN(n8025) );
  NOR2_X1 U8801 ( .A1(n7421), .A2(n10390), .ZN(n7586) );
  NAND2_X1 U8802 ( .A1(n11454), .A2(n9990), .ZN(n11666) );
  OAI21_X1 U8803 ( .B1(n10447), .B2(n14954), .A(n9866), .ZN(n10794) );
  NAND2_X1 U8804 ( .A1(n12258), .A2(n10073), .ZN(n12555) );
  NAND2_X1 U8805 ( .A1(n10077), .A2(n10076), .ZN(n12747) );
  OR2_X1 U8806 ( .A1(n14896), .A2(n14897), .ZN(n7481) );
  INV_X1 U8807 ( .A(n7464), .ZN(n14985) );
  NAND2_X1 U8808 ( .A1(n9831), .A2(n9830), .ZN(n16133) );
  INV_X1 U8809 ( .A(n8022), .ZN(n14996) );
  XNOR2_X1 U8810 ( .A(n9929), .B(n14954), .ZN(n11285) );
  INV_X1 U8811 ( .A(n11846), .ZN(n10028) );
  NAND2_X1 U8812 ( .A1(n8046), .A2(n14943), .ZN(n15013) );
  AND2_X1 U8813 ( .A1(n8046), .A2(n8044), .ZN(n15012) );
  OR2_X1 U8814 ( .A1(n14946), .A2(n14944), .ZN(n8046) );
  NAND2_X1 U8815 ( .A1(n12510), .A2(n12509), .ZN(n12508) );
  NOR2_X1 U8816 ( .A1(n14994), .A2(n10158), .ZN(n8021) );
  INV_X1 U8817 ( .A(n12716), .ZN(n15948) );
  NAND2_X1 U8818 ( .A1(n8018), .A2(n14904), .ZN(n15031) );
  NAND2_X1 U8819 ( .A1(n14976), .A2(n14977), .ZN(n8018) );
  CLKBUF_X1 U8820 ( .A(n15044), .Z(n15045) );
  NAND2_X1 U8821 ( .A1(n9797), .A2(n9796), .ZN(n15259) );
  AND2_X1 U8822 ( .A1(n10780), .A2(n7640), .ZN(n10387) );
  NAND2_X1 U8823 ( .A1(n10783), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7640) );
  INV_X1 U8824 ( .A(n7639), .ZN(n10385) );
  AND2_X1 U8825 ( .A1(n7639), .A2(n7638), .ZN(n10741) );
  NAND2_X1 U8826 ( .A1(n10354), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7638) );
  NOR2_X1 U8827 ( .A1(n10401), .A2(n7633), .ZN(n10405) );
  AND2_X1 U8828 ( .A1(n10402), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7633) );
  NOR2_X1 U8829 ( .A1(n10405), .A2(n10404), .ZN(n10613) );
  NOR2_X1 U8830 ( .A1(n11235), .A2(n7625), .ZN(n11239) );
  AND2_X1 U8831 ( .A1(n11236), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U8832 ( .A1(n11239), .A2(n11238), .ZN(n11463) );
  XNOR2_X1 U8833 ( .A(n11834), .B(n11474), .ZN(n11836) );
  INV_X1 U8834 ( .A(n7629), .ZN(n15123) );
  NOR2_X1 U8835 ( .A1(n15134), .A2(n7626), .ZN(n15127) );
  NOR2_X1 U8836 ( .A1(n7627), .A2(n15138), .ZN(n7626) );
  INV_X1 U8837 ( .A(n15153), .ZN(n15397) );
  INV_X1 U8838 ( .A(n12929), .ZN(n15416) );
  INV_X1 U8839 ( .A(n15420), .ZN(n15198) );
  NAND2_X1 U8840 ( .A1(n7927), .A2(n7925), .ZN(n15219) );
  AND2_X1 U8841 ( .A1(n7960), .A2(n7959), .ZN(n15275) );
  AND2_X1 U8842 ( .A1(n15289), .A2(n15288), .ZN(n15451) );
  NAND2_X1 U8843 ( .A1(n15306), .A2(n12661), .ZN(n15291) );
  NAND2_X1 U8844 ( .A1(n9803), .A2(n9802), .ZN(n15299) );
  NAND2_X1 U8845 ( .A1(n15336), .A2(n12658), .ZN(n15320) );
  INV_X1 U8846 ( .A(n15474), .ZN(n15345) );
  INV_X1 U8847 ( .A(n15388), .ZN(n7383) );
  AND2_X1 U8848 ( .A1(n7582), .A2(n7917), .ZN(n15373) );
  NAND2_X1 U8849 ( .A1(n7921), .A2(n12446), .ZN(n12447) );
  NAND2_X1 U8850 ( .A1(n7952), .A2(n12438), .ZN(n12602) );
  NAND2_X1 U8851 ( .A1(n10100), .A2(n10099), .ZN(n12751) );
  AND2_X1 U8852 ( .A1(n11994), .A2(n11984), .ZN(n7570) );
  NAND2_X1 U8853 ( .A1(n9998), .A2(n9997), .ZN(n15992) );
  NAND2_X1 U8854 ( .A1(n7934), .A2(n11916), .ZN(n15971) );
  NAND2_X1 U8855 ( .A1(n7949), .A2(n11446), .ZN(n11926) );
  NAND2_X1 U8856 ( .A1(n12673), .A2(n10993), .ZN(n10996) );
  INV_X1 U8857 ( .A(n7413), .ZN(n7412) );
  OAI211_X1 U8858 ( .C1(n15469), .C2(n15421), .A(n7501), .B(n7500), .ZN(n7499)
         );
  NAND2_X1 U8859 ( .A1(n15420), .A2(n16134), .ZN(n7500) );
  INV_X1 U8860 ( .A(n15419), .ZN(n7501) );
  OAI21_X1 U8861 ( .B1(n15426), .B2(n15469), .A(n7381), .ZN(n7380) );
  NOR2_X1 U8862 ( .A1(n15424), .A2(n7382), .ZN(n7381) );
  NAND2_X1 U8863 ( .A1(n9597), .A2(n9598), .ZN(n14859) );
  INV_X1 U8864 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9768) );
  NAND2_X1 U8865 ( .A1(n9579), .A2(n9578), .ZN(n14862) );
  OR2_X1 U8866 ( .A1(n9577), .A2(n9576), .ZN(n9578) );
  AND2_X1 U8867 ( .A1(n7350), .A2(n8221), .ZN(n7422) );
  NAND2_X1 U8868 ( .A1(n7431), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9745) );
  XNOR2_X1 U8869 ( .A(n9471), .B(n9452), .ZN(n12611) );
  NAND2_X1 U8870 ( .A1(n9763), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9759) );
  NAND2_X1 U8871 ( .A1(n7976), .A2(n7975), .ZN(n9425) );
  INV_X1 U8872 ( .A(n7982), .ZN(n7975) );
  NAND2_X1 U8873 ( .A1(n7932), .A2(n7282), .ZN(n9761) );
  INV_X1 U8874 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11038) );
  INV_X1 U8875 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10925) );
  INV_X1 U8876 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11015) );
  INV_X1 U8877 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10929) );
  INV_X1 U8878 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10422) );
  INV_X1 U8879 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10395) );
  INV_X1 U8880 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10426) );
  INV_X1 U8881 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10298) );
  INV_X1 U8882 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10251) );
  INV_X1 U8883 ( .A(n9901), .ZN(n10249) );
  NAND2_X1 U8884 ( .A1(n7631), .A2(n7290), .ZN(n10331) );
  NAND2_X1 U8885 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n7303), .ZN(n7631) );
  XNOR2_X1 U8886 ( .A(n7712), .B(n7711), .ZN(n15709) );
  NAND2_X1 U8887 ( .A1(n15709), .A2(n15708), .ZN(n15716) );
  NOR2_X1 U8888 ( .A1(n15751), .A2(n15752), .ZN(n15753) );
  XNOR2_X1 U8889 ( .A(n15761), .B(n7725), .ZN(n15759) );
  INV_X1 U8890 ( .A(n15760), .ZN(n7725) );
  NAND2_X1 U8891 ( .A1(n15759), .A2(n15758), .ZN(n15762) );
  XNOR2_X1 U8892 ( .A(n15774), .B(n7724), .ZN(n15768) );
  INV_X1 U8893 ( .A(n15773), .ZN(n7724) );
  NOR2_X1 U8894 ( .A1(n15795), .A2(n7716), .ZN(n7715) );
  INV_X1 U8895 ( .A(n7717), .ZN(n7716) );
  INV_X1 U8896 ( .A(n7410), .ZN(n15850) );
  AOI211_X1 U8897 ( .C1(n13754), .C2(n13727), .A(n13706), .B(n13705), .ZN(
        n13707) );
  INV_X1 U8898 ( .A(n13721), .ZN(n13714) );
  OAI21_X1 U8899 ( .B1(n14090), .B2(n12991), .A(n7389), .ZN(n14016) );
  NAND2_X1 U8900 ( .A1(n12991), .A2(n7390), .ZN(n7389) );
  INV_X1 U8901 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n7390) );
  NAND2_X1 U8902 ( .A1(n7393), .A2(n14063), .ZN(n7391) );
  NAND2_X1 U8903 ( .A1(n7406), .A2(n7405), .ZN(P3_U3456) );
  NAND2_X1 U8904 ( .A1(n16062), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7405) );
  NAND2_X1 U8905 ( .A1(n7407), .A2(n16065), .ZN(n7406) );
  NAND2_X1 U8906 ( .A1(n8152), .A2(n12990), .ZN(n7407) );
  AOI21_X1 U8907 ( .B1(n14090), .B2(n16065), .A(n7495), .ZN(n14092) );
  NAND2_X1 U8908 ( .A1(n7497), .A2(n7496), .ZN(n7495) );
  NAND2_X1 U8909 ( .A1(n16062), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7496) );
  NAND2_X1 U8910 ( .A1(n7393), .A2(n14124), .ZN(n7392) );
  INV_X1 U8911 ( .A(n7483), .ZN(n7482) );
  OAI21_X1 U8912 ( .B1(n14748), .B2(n14309), .A(n14208), .ZN(n7483) );
  OAI21_X1 U8913 ( .B1(n12277), .B2(n7263), .A(n12275), .ZN(n12533) );
  AND2_X1 U8914 ( .A1(n8234), .A2(n9720), .ZN(n9721) );
  NAND2_X1 U8915 ( .A1(P2_U3947), .A2(n7449), .ZN(n10304) );
  NOR2_X1 U8916 ( .A1(n15891), .A2(n14679), .ZN(n7829) );
  NAND2_X1 U8917 ( .A1(n7831), .A2(n7828), .ZN(n7827) );
  OAI21_X1 U8918 ( .B1(n14820), .B2(n16155), .A(n7426), .ZN(P2_U3527) );
  INV_X1 U8919 ( .A(n7427), .ZN(n7426) );
  OAI21_X1 U8920 ( .B1(n14822), .B2(n14816), .A(n7428), .ZN(n7427) );
  OR2_X1 U8921 ( .A1(n16156), .A2(n14745), .ZN(n7428) );
  INV_X1 U8922 ( .A(n7676), .ZN(n7675) );
  OR2_X1 U8923 ( .A1(n14820), .A2(n16157), .ZN(n7677) );
  NOR2_X1 U8924 ( .A1(n7505), .A2(n7504), .ZN(n7503) );
  INV_X1 U8925 ( .A(n7479), .ZN(n7478) );
  OAI21_X1 U8926 ( .B1(n14924), .B2(n16091), .A(n14923), .ZN(n7479) );
  NAND2_X1 U8927 ( .A1(n8034), .A2(n16093), .ZN(n8031) );
  AOI21_X1 U8928 ( .B1(n12920), .B2(n12917), .A(n7999), .ZN(n12918) );
  OAI21_X1 U8929 ( .B1(n12903), .B2(n8000), .A(n7292), .ZN(n7999) );
  OAI21_X1 U8930 ( .B1(n15151), .B2(n15150), .A(n7634), .ZN(P1_U3262) );
  AOI21_X1 U8931 ( .B1(n7636), .B2(n15150), .A(n7635), .ZN(n7634) );
  OAI21_X1 U8932 ( .B1(n15656), .B2(n7644), .A(n15152), .ZN(n7635) );
  AOI211_X1 U8933 ( .C1(n15409), .C2(n15347), .A(n12668), .B(n12667), .ZN(
        n12669) );
  INV_X1 U8934 ( .A(n15749), .ZN(n15741) );
  NOR2_X1 U8935 ( .A1(n15791), .A2(n15792), .ZN(n15793) );
  NAND2_X1 U8936 ( .A1(n7728), .A2(n7473), .ZN(n7472) );
  XNOR2_X1 U8937 ( .A(n15823), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n7726) );
  CLKBUF_X3 U8938 ( .A(n8308), .Z(n10630) );
  AND2_X1 U8939 ( .A1(n7860), .A2(n7858), .ZN(n7239) );
  INV_X2 U8940 ( .A(n8614), .ZN(n8472) );
  NOR2_X1 U8941 ( .A1(n8238), .A2(n7865), .ZN(n7864) );
  AND2_X1 U8942 ( .A1(n15203), .A2(n7922), .ZN(n7240) );
  XOR2_X1 U8943 ( .A(n13771), .B(n8790), .Z(n7241) );
  AND2_X1 U8944 ( .A1(n9061), .A2(n7434), .ZN(n7242) );
  AND2_X1 U8945 ( .A1(n13450), .A2(n13449), .ZN(n13447) );
  INV_X1 U8946 ( .A(n12877), .ZN(n7923) );
  AND2_X1 U8947 ( .A1(n9466), .A2(n9465), .ZN(n7243) );
  AND2_X1 U8948 ( .A1(n15220), .A2(n7926), .ZN(n7925) );
  AND2_X1 U8949 ( .A1(n13578), .A2(n16010), .ZN(n7244) );
  INV_X1 U8950 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15501) );
  AND2_X1 U8951 ( .A1(n7883), .A2(n14311), .ZN(n7245) );
  INV_X1 U8952 ( .A(n9642), .ZN(n8133) );
  AND2_X1 U8953 ( .A1(n14535), .A2(n8060), .ZN(n7246) );
  INV_X1 U8954 ( .A(n7756), .ZN(n7755) );
  INV_X1 U8955 ( .A(n10883), .ZN(n7756) );
  NOR2_X1 U8956 ( .A1(n15832), .A2(n12174), .ZN(n7247) );
  INV_X1 U8957 ( .A(n7533), .ZN(n7530) );
  NAND2_X1 U8958 ( .A1(n7267), .A2(n7534), .ZN(n7533) );
  INV_X1 U8959 ( .A(n7864), .ZN(n7863) );
  OR2_X1 U8960 ( .A1(n7875), .A2(n8233), .ZN(n7248) );
  NAND2_X1 U8961 ( .A1(n9245), .A2(SI_15_), .ZN(n9278) );
  NOR2_X1 U8962 ( .A1(n12474), .A2(n8498), .ZN(n7249) );
  AND2_X1 U8963 ( .A1(n9326), .A2(n8845), .ZN(n7250) );
  NAND2_X1 U8964 ( .A1(n8694), .A2(n8693), .ZN(n14039) );
  OR2_X1 U8965 ( .A1(n7888), .A2(n7894), .ZN(n7251) );
  INV_X1 U8966 ( .A(n12727), .ZN(n7623) );
  AND2_X1 U8967 ( .A1(n10018), .A2(n10001), .ZN(n7252) );
  INV_X1 U8968 ( .A(n12423), .ZN(n7669) );
  NAND2_X1 U8969 ( .A1(n15514), .A2(n7421), .ZN(n15439) );
  INV_X1 U8970 ( .A(n14096), .ZN(n7393) );
  NAND2_X1 U8971 ( .A1(n8289), .A2(n8288), .ZN(n11174) );
  INV_X1 U8972 ( .A(n11174), .ZN(n7567) );
  OR2_X1 U8973 ( .A1(n9827), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n7253) );
  NAND2_X2 U8974 ( .A1(n7411), .A2(n10040), .ZN(n16031) );
  XOR2_X1 U8975 ( .A(n8951), .B(n8949), .Z(n7254) );
  INV_X1 U8976 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8458) );
  INV_X1 U8977 ( .A(n9870), .ZN(n9772) );
  AND2_X1 U8978 ( .A1(n7997), .A2(n9296), .ZN(n7255) );
  INV_X1 U8979 ( .A(n11858), .ZN(n7820) );
  OR2_X1 U8980 ( .A1(n8678), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7257) );
  AND2_X1 U8981 ( .A1(n8125), .A2(n7311), .ZN(n7258) );
  AND4_X1 U8982 ( .A1(n7468), .A2(n8258), .A3(n8259), .A4(n8260), .ZN(n7259)
         );
  AND2_X1 U8983 ( .A1(n13222), .A2(n8168), .ZN(n7260) );
  INV_X1 U8984 ( .A(n13331), .ZN(n8168) );
  XNOR2_X1 U8985 ( .A(n8352), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10872) );
  INV_X1 U8986 ( .A(n10872), .ZN(n7763) );
  NAND2_X1 U8987 ( .A1(n9789), .A2(n9788), .ZN(n15444) );
  NOR2_X1 U8988 ( .A1(n14630), .A2(n7695), .ZN(n7261) );
  INV_X1 U8989 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8056) );
  AND2_X1 U8990 ( .A1(n8983), .A2(n8982), .ZN(n7262) );
  NOR2_X1 U8991 ( .A1(n12274), .A2(n12268), .ZN(n7263) );
  NOR2_X1 U8992 ( .A1(n12725), .A2(n11927), .ZN(n7264) );
  NOR2_X1 U8993 ( .A1(n12755), .A2(n15050), .ZN(n7265) );
  AND2_X1 U8994 ( .A1(n12657), .A2(n12656), .ZN(n7266) );
  AND2_X1 U8995 ( .A1(n8730), .A2(n8731), .ZN(n7267) );
  AND2_X1 U8996 ( .A1(n11510), .A2(n11511), .ZN(n7268) );
  AND2_X1 U8997 ( .A1(n8252), .A2(n8351), .ZN(n8418) );
  OR2_X1 U8998 ( .A1(n11593), .A2(n7881), .ZN(n7269) );
  OR3_X1 U8999 ( .A1(n8591), .A2(P3_IR_REG_18__SCAN_IN), .A3(n8291), .ZN(n7270) );
  AND2_X1 U9000 ( .A1(n15382), .A2(n15366), .ZN(n7271) );
  INV_X1 U9001 ( .A(n13426), .ZN(n7854) );
  INV_X1 U9002 ( .A(n13941), .ZN(n8194) );
  INV_X1 U9003 ( .A(n8027), .ZN(n8026) );
  AND2_X1 U9004 ( .A1(n14927), .A2(n8028), .ZN(n8027) );
  AND2_X1 U9005 ( .A1(n8156), .A2(n13269), .ZN(n7272) );
  AND2_X1 U9006 ( .A1(n8019), .A2(n15032), .ZN(n7273) );
  XOR2_X1 U9007 ( .A(n13548), .B(n13743), .Z(n7274) );
  AND2_X1 U9008 ( .A1(n14784), .A2(n14507), .ZN(n7275) );
  OR2_X1 U9009 ( .A1(n15792), .A2(n7719), .ZN(n7276) );
  NAND2_X1 U9010 ( .A1(n12848), .A2(n12847), .ZN(n15156) );
  INV_X1 U9011 ( .A(n15156), .ZN(n7734) );
  XOR2_X1 U9012 ( .A(n9138), .B(SI_10_), .Z(n7277) );
  INV_X1 U9013 ( .A(n12099), .ZN(n10844) );
  NAND2_X1 U9014 ( .A1(n8961), .A2(n8053), .ZN(n12099) );
  INV_X1 U9015 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8870) );
  INV_X1 U9016 ( .A(n12983), .ZN(n13798) );
  AND2_X1 U9017 ( .A1(n10974), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7278) );
  INV_X1 U9018 ( .A(n12757), .ZN(n8226) );
  NOR2_X1 U9019 ( .A1(n13633), .A2(n7769), .ZN(n7279) );
  OR2_X1 U9020 ( .A1(n9130), .A2(n9132), .ZN(n7280) );
  OR2_X1 U9021 ( .A1(n9034), .A2(n7287), .ZN(n7281) );
  INV_X1 U9022 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8883) );
  INV_X1 U9023 ( .A(n12872), .ZN(n15387) );
  AND3_X1 U9024 ( .A1(n7622), .A2(n9992), .A3(n8231), .ZN(n7282) );
  AND2_X1 U9025 ( .A1(n7852), .A2(n12205), .ZN(n7283) );
  NAND2_X1 U9026 ( .A1(n9569), .A2(n9568), .ZN(n14730) );
  INV_X1 U9027 ( .A(n14730), .ZN(n7702) );
  OR2_X1 U9028 ( .A1(n14017), .A2(n13787), .ZN(n7284) );
  OR2_X1 U9029 ( .A1(n9058), .A2(n9057), .ZN(n7285) );
  AND2_X1 U9030 ( .A1(n14759), .A2(n14516), .ZN(n7286) );
  AND2_X1 U9031 ( .A1(n9032), .A2(n9031), .ZN(n7287) );
  NOR2_X1 U9032 ( .A1(n13432), .A2(n7854), .ZN(n7853) );
  AND2_X1 U9033 ( .A1(n7687), .A2(n11751), .ZN(n7288) );
  INV_X1 U9034 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8853) );
  AND2_X1 U9035 ( .A1(n14182), .A2(n14181), .ZN(n7289) );
  AND2_X1 U9036 ( .A1(n9878), .A2(n7630), .ZN(n7290) );
  AND2_X1 U9037 ( .A1(n7553), .A2(n7549), .ZN(n7291) );
  NAND2_X1 U9038 ( .A1(n10854), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10884) );
  INV_X1 U9039 ( .A(n12777), .ZN(n7603) );
  INV_X1 U9040 ( .A(n12658), .ZN(n7575) );
  AND3_X1 U9041 ( .A1(n12916), .A2(n12915), .A3(n12914), .ZN(n7292) );
  OR2_X1 U9042 ( .A1(n8985), .A2(n7262), .ZN(n7293) );
  AND2_X1 U9043 ( .A1(n14609), .A2(n14515), .ZN(n7294) );
  INV_X1 U9044 ( .A(n14545), .ZN(n14741) );
  NAND2_X1 U9045 ( .A1(n9581), .A2(n9580), .ZN(n14545) );
  INV_X1 U9046 ( .A(n7735), .ZN(n15228) );
  NOR2_X1 U9047 ( .A1(n15242), .A2(n15429), .ZN(n7735) );
  NAND2_X1 U9048 ( .A1(n13648), .A2(n13657), .ZN(n13666) );
  AND2_X1 U9049 ( .A1(n7691), .A2(n7692), .ZN(n7295) );
  AND2_X1 U9050 ( .A1(n12169), .A2(n12168), .ZN(n7296) );
  AND2_X1 U9051 ( .A1(n16019), .A2(n12083), .ZN(n7297) );
  INV_X1 U9052 ( .A(n12779), .ZN(n8227) );
  AND2_X1 U9053 ( .A1(n7696), .A2(n8072), .ZN(n7298) );
  AND2_X1 U9054 ( .A1(n14563), .A2(n14521), .ZN(n7299) );
  NAND2_X1 U9055 ( .A1(n9135), .A2(n9136), .ZN(n7300) );
  AND2_X1 U9056 ( .A1(n10089), .A2(n10073), .ZN(n7301) );
  AND2_X1 U9057 ( .A1(n10010), .A2(n9990), .ZN(n7302) );
  INV_X1 U9058 ( .A(n7819), .ZN(n7818) );
  OAI21_X1 U9059 ( .B1(n11721), .B2(n7820), .A(n11860), .ZN(n7819) );
  AND2_X1 U9060 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n7303) );
  NAND2_X1 U9061 ( .A1(n12183), .A2(n12182), .ZN(n7304) );
  AND2_X1 U9062 ( .A1(n7697), .A2(n12012), .ZN(n7305) );
  OR2_X1 U9063 ( .A1(n7241), .A2(n8163), .ZN(n7306) );
  AND2_X1 U9064 ( .A1(n8657), .A2(n13915), .ZN(n7307) );
  AND2_X1 U9065 ( .A1(n12977), .A2(n13880), .ZN(n7308) );
  AND2_X1 U9066 ( .A1(n8261), .A2(n8200), .ZN(n7309) );
  INV_X1 U9067 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9756) );
  BUF_X4 U9068 ( .A(n10662), .Z(n14229) );
  AND2_X1 U9069 ( .A1(n8222), .A2(n12797), .ZN(n7310) );
  AND2_X1 U9070 ( .A1(n9486), .A2(n9485), .ZN(n7311) );
  AND2_X1 U9071 ( .A1(n10132), .A2(n10131), .ZN(n7312) );
  AND2_X1 U9072 ( .A1(n13490), .A2(n13489), .ZN(n7313) );
  NOR2_X1 U9073 ( .A1(n12772), .A2(n12774), .ZN(n7314) );
  NOR2_X1 U9074 ( .A1(n12756), .A2(n8226), .ZN(n7315) );
  NOR2_X1 U9075 ( .A1(n15429), .A2(n15059), .ZN(n7316) );
  AND2_X1 U9076 ( .A1(n13426), .A2(n13430), .ZN(n13527) );
  NOR2_X1 U9077 ( .A1(n16003), .A2(n11514), .ZN(n7317) );
  NOR2_X1 U9078 ( .A1(n12744), .A2(n12299), .ZN(n7318) );
  AND2_X1 U9079 ( .A1(n12770), .A2(n7612), .ZN(n7319) );
  NAND2_X1 U9080 ( .A1(n9764), .A2(n9763), .ZN(n12838) );
  NAND2_X1 U9081 ( .A1(n11497), .A2(n11498), .ZN(n7320) );
  AND2_X1 U9082 ( .A1(n7893), .A2(n12275), .ZN(n7321) );
  AND2_X1 U9083 ( .A1(n14656), .A2(n14507), .ZN(n7322) );
  INV_X1 U9084 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9740) );
  OR2_X1 U9085 ( .A1(n7314), .A2(n7611), .ZN(n7323) );
  AND2_X1 U9086 ( .A1(n8042), .A2(n8043), .ZN(n7324) );
  NOR2_X1 U9087 ( .A1(n8757), .A2(n13575), .ZN(n8167) );
  INV_X1 U9088 ( .A(n8233), .ZN(n7877) );
  AND2_X1 U9089 ( .A1(n14691), .A2(n8064), .ZN(n7325) );
  AND2_X1 U9090 ( .A1(n9063), .A2(SI_7_), .ZN(n7326) );
  AND2_X1 U9091 ( .A1(n12756), .A2(n8226), .ZN(n7327) );
  INV_X1 U9092 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10273) );
  INV_X1 U9093 ( .A(n7548), .ZN(n7547) );
  NAND2_X1 U9094 ( .A1(n12390), .A2(n8480), .ZN(n7548) );
  INV_X1 U9095 ( .A(n13933), .ZN(n12976) );
  OR2_X1 U9096 ( .A1(n13941), .A2(n8193), .ZN(n7328) );
  AND2_X1 U9097 ( .A1(n8227), .A2(n12778), .ZN(n7329) );
  INV_X1 U9098 ( .A(n8178), .ZN(n8177) );
  NAND2_X1 U9099 ( .A1(n8477), .A2(n8456), .ZN(n8178) );
  OR2_X1 U9100 ( .A1(n9273), .A2(n13124), .ZN(n7330) );
  AND2_X1 U9101 ( .A1(n8116), .A2(n11325), .ZN(n7331) );
  OR2_X1 U9102 ( .A1(n12748), .A2(n12750), .ZN(n7332) );
  INV_X1 U9103 ( .A(n12828), .ZN(n7591) );
  NAND2_X1 U9104 ( .A1(n14310), .A2(n14186), .ZN(n14187) );
  INV_X1 U9105 ( .A(n8069), .ZN(n8068) );
  NAND2_X1 U9106 ( .A1(n14707), .A2(n14464), .ZN(n8069) );
  INV_X1 U9107 ( .A(n14486), .ZN(n14535) );
  AND2_X1 U9108 ( .A1(n14522), .A2(n9644), .ZN(n14486) );
  NAND2_X1 U9109 ( .A1(n8744), .A2(n13827), .ZN(n7534) );
  INV_X1 U9110 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8292) );
  INV_X1 U9111 ( .A(n12736), .ZN(n8220) );
  OR2_X1 U9112 ( .A1(n15423), .A2(n7380), .ZN(n7333) );
  INV_X1 U9113 ( .A(n12754), .ZN(n7617) );
  AND2_X1 U9114 ( .A1(n12605), .A2(n15351), .ZN(n7334) );
  OR2_X1 U9115 ( .A1(n14686), .A2(n14501), .ZN(n7335) );
  AND2_X1 U9116 ( .A1(n8043), .A2(n14967), .ZN(n7336) );
  OR2_X1 U9117 ( .A1(n8121), .A2(n7258), .ZN(n7337) );
  AND2_X1 U9118 ( .A1(n8160), .A2(n7306), .ZN(n7338) );
  AND2_X1 U9119 ( .A1(n13435), .A2(n13428), .ZN(n12205) );
  AND2_X1 U9120 ( .A1(n15282), .A2(n12661), .ZN(n7339) );
  NOR2_X1 U9121 ( .A1(n9270), .A2(n9269), .ZN(n7340) );
  OR2_X1 U9122 ( .A1(n8227), .A2(n12778), .ZN(n7341) );
  AND2_X1 U9123 ( .A1(n12828), .A2(n7592), .ZN(n7342) );
  AND2_X1 U9124 ( .A1(n8853), .A2(n8854), .ZN(n7343) );
  AND2_X1 U9125 ( .A1(n8132), .A2(n8130), .ZN(n7344) );
  AND2_X1 U9126 ( .A1(n7877), .A2(n14265), .ZN(n7345) );
  AND2_X1 U9127 ( .A1(n7927), .A2(n7926), .ZN(n7346) );
  OR2_X1 U9128 ( .A1(n8138), .A2(n9131), .ZN(n7347) );
  OR2_X1 U9129 ( .A1(n12726), .A2(n7623), .ZN(n7348) );
  NAND2_X1 U9130 ( .A1(n9291), .A2(n9292), .ZN(n7349) );
  AND2_X1 U9131 ( .A1(n7946), .A2(n9756), .ZN(n7350) );
  NAND2_X1 U9132 ( .A1(n9239), .A2(n9240), .ZN(n7351) );
  NAND2_X1 U9133 ( .A1(n9343), .A2(n9344), .ZN(n7352) );
  AND2_X1 U9134 ( .A1(n12421), .A2(n12426), .ZN(n7666) );
  AND2_X1 U9135 ( .A1(n7332), .A2(n7596), .ZN(n7353) );
  OR2_X1 U9136 ( .A1(n9421), .A2(n9423), .ZN(n7354) );
  INV_X1 U9137 ( .A(n7925), .ZN(n7924) );
  NAND2_X1 U9138 ( .A1(n11620), .A2(n11619), .ZN(n11902) );
  NAND2_X1 U9139 ( .A1(n10156), .A2(n10157), .ZN(n7355) );
  INV_X1 U9140 ( .A(n7894), .ZN(n7893) );
  OR2_X1 U9141 ( .A1(n12538), .A2(n12545), .ZN(n7894) );
  INV_X1 U9142 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U9143 ( .A1(n12816), .A2(n8204), .ZN(n7356) );
  INV_X1 U9144 ( .A(n12746), .ZN(n7598) );
  INV_X1 U9145 ( .A(n14609), .ZN(n7706) );
  AND2_X1 U9146 ( .A1(n16085), .A2(n10115), .ZN(n8041) );
  INV_X1 U9147 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7646) );
  OR2_X1 U9148 ( .A1(n15326), .A2(n7742), .ZN(n7357) );
  NAND2_X1 U9149 ( .A1(n7928), .A2(n7266), .ZN(n15336) );
  NAND2_X1 U9150 ( .A1(n14530), .A2(n14529), .ZN(n7358) );
  INV_X1 U9151 ( .A(n12026), .ZN(n7794) );
  NAND2_X1 U9152 ( .A1(n7921), .A2(n7919), .ZN(n7359) );
  INV_X1 U9153 ( .A(n14943), .ZN(n8045) );
  OR3_X1 U9154 ( .A1(n12120), .A2(n14359), .A3(n16111), .ZN(n7360) );
  MUX2_X1 U9155 ( .A(n10440), .B(n14872), .S(n8905), .Z(n10775) );
  NAND2_X1 U9156 ( .A1(n7928), .A2(n12656), .ZN(n15337) );
  INV_X1 U9157 ( .A(n15056), .ZN(n15190) );
  NAND4_X1 U9158 ( .A1(n12632), .A2(n12631), .A3(n12630), .A4(n12629), .ZN(
        n15056) );
  AND2_X1 U9159 ( .A1(n8057), .A2(n7697), .ZN(n7361) );
  AND2_X1 U9160 ( .A1(n7902), .A2(n7900), .ZN(n7362) );
  INV_X1 U9161 ( .A(n7743), .ZN(n15309) );
  NOR2_X1 U9162 ( .A1(n15326), .A2(n15460), .ZN(n7743) );
  NAND2_X1 U9163 ( .A1(n15834), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7363) );
  NAND2_X1 U9164 ( .A1(n7890), .A2(n7888), .ZN(n7895) );
  OR2_X1 U9165 ( .A1(n8591), .A2(n8291), .ZN(n7364) );
  AND2_X1 U9166 ( .A1(n13468), .A2(n13467), .ZN(n7365) );
  INV_X1 U9167 ( .A(n7703), .ZN(n14714) );
  NOR3_X1 U9168 ( .A1(n12120), .A2(n14359), .A3(n7705), .ZN(n7703) );
  INV_X1 U9169 ( .A(n7738), .ZN(n12441) );
  NOR2_X1 U9170 ( .A1(n12381), .A2(n12751), .ZN(n7738) );
  AND2_X1 U9171 ( .A1(n14476), .A2(n14633), .ZN(n7366) );
  NAND2_X1 U9172 ( .A1(n15834), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7367) );
  OR2_X1 U9173 ( .A1(n8137), .A2(n9422), .ZN(n7368) );
  AND2_X1 U9174 ( .A1(n12230), .A2(n8480), .ZN(n7369) );
  INV_X1 U9175 ( .A(n8238), .ZN(n7867) );
  AND2_X2 U9176 ( .A1(n15169), .A2(n15377), .ZN(n16001) );
  AND2_X1 U9177 ( .A1(n11126), .A2(n11125), .ZN(n16062) );
  INV_X1 U9178 ( .A(n12755), .ZN(n7737) );
  INV_X1 U9179 ( .A(n12127), .ZN(n8076) );
  INV_X1 U9180 ( .A(n16157), .ZN(n16117) );
  INV_X1 U9181 ( .A(n12157), .ZN(n7708) );
  NAND2_X1 U9182 ( .A1(n7571), .A2(n7570), .ZN(n12302) );
  INV_X1 U9183 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11325) );
  AND4_X1 U9184 ( .A1(n8699), .A2(n8698), .A3(n8697), .A4(n8696), .ZN(n13846)
         );
  INV_X1 U9185 ( .A(n13846), .ZN(n7492) );
  AND2_X1 U9186 ( .A1(n12991), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n7370) );
  XOR2_X1 U9187 ( .A(n12274), .B(n12268), .Z(n7371) );
  NAND2_X1 U9188 ( .A1(n7937), .A2(n7379), .ZN(n12375) );
  NAND2_X1 U9189 ( .A1(n15980), .A2(n11932), .ZN(n11968) );
  NAND2_X1 U9190 ( .A1(n11983), .A2(n7938), .ZN(n12298) );
  NAND2_X1 U9191 ( .A1(n7571), .A2(n11994), .ZN(n11995) );
  AND2_X1 U9192 ( .A1(n7850), .A2(n7852), .ZN(n7372) );
  INV_X1 U9193 ( .A(n7709), .ZN(n12151) );
  INV_X1 U9194 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7711) );
  INV_X1 U9195 ( .A(SI_20_), .ZN(n13114) );
  AND2_X1 U9196 ( .A1(n11323), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7373) );
  NAND2_X1 U9197 ( .A1(n7508), .A2(n7848), .ZN(n7374) );
  AND2_X1 U9198 ( .A1(n7793), .A2(n7791), .ZN(n7375) );
  INV_X1 U9199 ( .A(n13657), .ZN(n7458) );
  INV_X1 U9200 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8113) );
  INV_X1 U9201 ( .A(n15872), .ZN(n7465) );
  NOR2_X1 U9202 ( .A1(n16062), .A2(n16054), .ZN(n14124) );
  INV_X1 U9203 ( .A(n14679), .ZN(n14710) );
  AND2_X1 U9204 ( .A1(n10477), .A2(n10476), .ZN(n14679) );
  INV_X1 U9205 ( .A(n14353), .ZN(n14311) );
  OR2_X1 U9206 ( .A1(n10657), .A2(n10656), .ZN(n14353) );
  OR2_X1 U9207 ( .A1(n13656), .A2(n13625), .ZN(n7376) );
  NAND2_X1 U9208 ( .A1(n11267), .A2(n13388), .ZN(n13549) );
  INV_X1 U9209 ( .A(n13549), .ZN(n7568) );
  NAND2_X1 U9210 ( .A1(n11426), .A2(n13755), .ZN(n13550) );
  NAND2_X1 U9211 ( .A1(n8886), .A2(n11375), .ZN(n10774) );
  INV_X1 U9212 ( .A(n10774), .ZN(n10468) );
  AND2_X1 U9213 ( .A1(n10230), .A2(n10216), .ZN(n16093) );
  INV_X1 U9214 ( .A(n16093), .ZN(n15042) );
  INV_X1 U9215 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11428) );
  AND2_X1 U9216 ( .A1(n11954), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7377) );
  NAND2_X1 U9217 ( .A1(n7230), .A2(n8315), .ZN(n9846) );
  INV_X1 U9218 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12589) );
  INV_X1 U9219 ( .A(n12913), .ZN(n8001) );
  NAND2_X1 U9220 ( .A1(n10800), .A2(n10801), .ZN(n7435) );
  NAND2_X1 U9221 ( .A1(n7753), .A2(n7756), .ZN(n7378) );
  INV_X1 U9222 ( .A(n14387), .ZN(n8055) );
  INV_X1 U9223 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n8101) );
  INV_X1 U9224 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7644) );
  NOR2_X1 U9225 ( .A1(n8286), .A2(n12401), .ZN(n10309) );
  NAND2_X1 U9226 ( .A1(n10945), .A2(n15524), .ZN(n16157) );
  NOR2_X1 U9227 ( .A1(n16117), .A2(n14824), .ZN(n7504) );
  OAI22_X1 U9228 ( .A1(n14822), .A2(n14849), .B1(n16117), .B2(n14821), .ZN(
        n7676) );
  NAND2_X1 U9229 ( .A1(n11981), .A2(n7939), .ZN(n7379) );
  NAND2_X2 U9230 ( .A1(n15304), .A2(n15303), .ZN(n15302) );
  NAND2_X1 U9231 ( .A1(n15224), .A2(n15223), .ZN(n15222) );
  AOI21_X1 U9232 ( .B1(n15273), .B2(n15259), .A(n15274), .ZN(n15255) );
  NAND2_X1 U9233 ( .A1(n7642), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7641) );
  NAND2_X1 U9234 ( .A1(n8969), .A2(n8968), .ZN(n7384) );
  OAI21_X1 U9235 ( .B1(n8954), .B2(n7216), .A(n8952), .ZN(n8955) );
  INV_X1 U9236 ( .A(n7940), .ZN(n7939) );
  NAND2_X1 U9237 ( .A1(n12377), .A2(n12376), .ZN(n12437) );
  NAND2_X1 U9238 ( .A1(n8956), .A2(n8957), .ZN(n8969) );
  NAND2_X1 U9239 ( .A1(n15253), .A2(n7461), .ZN(n15235) );
  OAI21_X1 U9240 ( .B1(n7941), .B2(n12737), .A(n12863), .ZN(n7940) );
  NOR2_X4 U9241 ( .A1(n10035), .A2(n9737), .ZN(n9739) );
  NOR2_X2 U9242 ( .A1(n15023), .A2(n10174), .ZN(n14946) );
  AND4_X2 U9243 ( .A1(n9724), .A2(n9725), .A3(n9726), .A4(n10136), .ZN(n7932)
         );
  NOR2_X2 U9244 ( .A1(n9755), .A2(n8205), .ZN(n15498) );
  XNOR2_X1 U9245 ( .A(n9849), .B(n10188), .ZN(n9852) );
  NAND2_X1 U9246 ( .A1(n11379), .A2(n11378), .ZN(n11377) );
  NAND2_X1 U9247 ( .A1(n8042), .A2(n7336), .ZN(n14966) );
  NAND4_X1 U9248 ( .A1(n9844), .A2(n9841), .A3(n9842), .A4(n9843), .ZN(n10902)
         );
  NAND2_X1 U9249 ( .A1(n10029), .A2(n10028), .ZN(n11848) );
  NAND2_X1 U9250 ( .A1(n7386), .A2(n7385), .ZN(n9853) );
  NAND2_X1 U9251 ( .A1(n9868), .A2(n9867), .ZN(n10792) );
  NAND4_X2 U9252 ( .A1(n9785), .A2(n9735), .A3(n9736), .A4(n9734), .ZN(n9737)
         );
  NAND2_X1 U9253 ( .A1(n14966), .A2(n7511), .ZN(n10217) );
  NAND2_X1 U9254 ( .A1(n11377), .A2(n9971), .ZN(n11456) );
  NAND2_X1 U9255 ( .A1(n15044), .A2(n15047), .ZN(n15046) );
  NAND2_X1 U9256 ( .A1(n7387), .A2(n11293), .ZN(n11379) );
  NAND2_X1 U9257 ( .A1(n11848), .A2(n10034), .ZN(n12080) );
  NAND2_X1 U9258 ( .A1(n7512), .A2(n7285), .ZN(n9082) );
  OAI21_X1 U9259 ( .B1(n9272), .B2(n9271), .A(n7349), .ZN(n7490) );
  OAI21_X1 U9260 ( .B1(n9108), .B2(n9107), .A(n7280), .ZN(n7446) );
  AOI21_X1 U9261 ( .B1(n9058), .B2(n9057), .A(n9056), .ZN(n9059) );
  OAI21_X1 U9262 ( .B1(n7448), .B2(n7447), .A(n7368), .ZN(n9447) );
  INV_X1 U9263 ( .A(n9851), .ZN(n7385) );
  INV_X1 U9264 ( .A(n9852), .ZN(n7386) );
  NAND2_X1 U9265 ( .A1(n11295), .A2(n11294), .ZN(n7387) );
  NAND3_X1 U9266 ( .A1(n9739), .A2(n9738), .A3(n7422), .ZN(n7732) );
  NAND2_X1 U9267 ( .A1(n11664), .A2(n10013), .ZN(n11847) );
  OAI21_X1 U9268 ( .B1(n9109), .B2(n7446), .A(n7347), .ZN(n9162) );
  NAND2_X2 U9269 ( .A1(n15775), .A2(n15776), .ZN(n15782) );
  NAND2_X1 U9270 ( .A1(n7714), .A2(n7713), .ZN(n7712) );
  NAND3_X1 U9271 ( .A1(n7519), .A2(n7202), .A3(n7293), .ZN(n7439) );
  NAND2_X1 U9272 ( .A1(n8884), .A2(n10775), .ZN(n8891) );
  OAI21_X2 U9273 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(n15798), .A(n15797), .ZN(
        n15804) );
  OAI21_X1 U9274 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n15669), .A(n15668), .ZN(
        n15683) );
  NAND2_X1 U9275 ( .A1(n15822), .A2(n15821), .ZN(n7730) );
  NAND2_X1 U9276 ( .A1(n7728), .A2(n7729), .ZN(n7727) );
  XNOR2_X1 U9277 ( .A(n7727), .B(n7726), .ZN(SUB_1596_U4) );
  NAND2_X1 U9278 ( .A1(n7452), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7388) );
  AOI21_X1 U9279 ( .B1(n9370), .B2(n9369), .A(n9368), .ZN(n9372) );
  NAND2_X1 U9280 ( .A1(n9645), .A2(n8885), .ZN(n8884) );
  NAND2_X1 U9281 ( .A1(n13840), .A2(n12947), .ZN(n13824) );
  OR2_X1 U9282 ( .A1(n9445), .A2(n9448), .ZN(n9469) );
  NAND2_X1 U9283 ( .A1(n14021), .A2(n7391), .ZN(P3_U3486) );
  NAND2_X1 U9284 ( .A1(n14095), .A2(n7392), .ZN(P3_U3454) );
  NAND2_X1 U9285 ( .A1(n11271), .A2(n11272), .ZN(n11677) );
  NAND2_X1 U9286 ( .A1(n8172), .A2(n8170), .ZN(n13971) );
  AOI21_X2 U9287 ( .B1(n7395), .B2(n7394), .A(n7286), .ZN(n7672) );
  NAND2_X1 U9288 ( .A1(n9087), .A2(n9086), .ZN(n9090) );
  NAND2_X1 U9289 ( .A1(n9382), .A2(n9381), .ZN(n9403) );
  NAND3_X1 U9290 ( .A1(n8129), .A2(n8131), .A3(n8128), .ZN(n8127) );
  NAND2_X1 U9291 ( .A1(n9298), .A2(n7255), .ZN(n7991) );
  INV_X1 U9292 ( .A(n7903), .ZN(n7901) );
  NAND2_X1 U9293 ( .A1(n14240), .A2(n7397), .ZN(P2_U3192) );
  INV_X1 U9294 ( .A(n7906), .ZN(n7904) );
  NAND2_X1 U9295 ( .A1(n15293), .A2(n8235), .ZN(n15268) );
  NAND2_X1 U9296 ( .A1(n15164), .A2(n15163), .ZN(n7914) );
  OAI22_X1 U9297 ( .A1(n15186), .A2(n15187), .B1(n14918), .B2(n15198), .ZN(
        n12922) );
  OAI21_X1 U9298 ( .B1(n15407), .B2(n15469), .A(n15406), .ZN(n7413) );
  OAI21_X2 U9299 ( .B1(n12664), .B2(n15060), .A(n15249), .ZN(n15240) );
  NAND2_X1 U9300 ( .A1(n12666), .A2(n12665), .ZN(n15164) );
  NAND2_X1 U9301 ( .A1(n9473), .A2(n9472), .ZN(n9489) );
  AOI21_X1 U9302 ( .B1(n7240), .B2(n7924), .A(n7580), .ZN(n7578) );
  OAI21_X1 U9303 ( .B1(n9298), .B2(n7994), .A(n7992), .ZN(n9382) );
  NAND2_X1 U9304 ( .A1(n7945), .A2(n7412), .ZN(n15480) );
  INV_X1 U9305 ( .A(n7891), .ZN(n7889) );
  OAI21_X1 U9306 ( .B1(n14324), .B2(n7899), .A(n7897), .ZN(n7908) );
  NAND2_X1 U9307 ( .A1(n10674), .A2(n10675), .ZN(n10673) );
  NAND2_X2 U9308 ( .A1(n8905), .A2(n10252), .ZN(n9599) );
  NAND2_X2 U9309 ( .A1(n9707), .A2(n14868), .ZN(n8905) );
  NAND2_X1 U9310 ( .A1(n10447), .A2(n10448), .ZN(n9866) );
  NAND2_X1 U9311 ( .A1(n9864), .A2(n9865), .ZN(n10448) );
  OR2_X1 U9312 ( .A1(n10698), .A2(n11738), .ZN(n10827) );
  AND2_X2 U9313 ( .A1(n11056), .A2(n11777), .ZN(n11409) );
  OR2_X2 U9314 ( .A1(n14695), .A2(n14686), .ZN(n14681) );
  OAI211_X2 U9315 ( .C1(n9599), .C2(n10246), .A(n8908), .B(n8907), .ZN(n11879)
         );
  NAND2_X1 U9316 ( .A1(n10811), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7502) );
  NOR2_X1 U9317 ( .A1(n13636), .A2(n13635), .ZN(n13647) );
  NOR2_X1 U9318 ( .A1(n11541), .A2(n16015), .ZN(n12056) );
  OAI21_X1 U9319 ( .B1(n9010), .B2(n8143), .A(n8142), .ZN(n9058) );
  OAI21_X2 U9320 ( .B1(n13896), .B2(n12943), .A(n8236), .ZN(n13879) );
  NAND2_X2 U9321 ( .A1(n13911), .A2(n12942), .ZN(n13896) );
  NAND4_X2 U9322 ( .A1(n8319), .A2(n8320), .A3(n8317), .A4(n8318), .ZN(n13586)
         );
  NAND2_X1 U9323 ( .A1(n11902), .A2(n7470), .ZN(n7469) );
  NAND2_X1 U9324 ( .A1(n11044), .A2(n11043), .ZN(n11046) );
  NAND2_X1 U9325 ( .A1(n7677), .A2(n7675), .ZN(P2_U3495) );
  NAND2_X1 U9326 ( .A1(n11704), .A2(n11703), .ZN(n12143) );
  NAND2_X1 U9327 ( .A1(n10482), .A2(n10481), .ZN(n10589) );
  NAND2_X1 U9328 ( .A1(n14604), .A2(n14481), .ZN(n14587) );
  OAI22_X1 U9329 ( .A1(n7490), .A2(n7340), .B1(n9291), .B2(n9292), .ZN(n9319)
         );
  NAND2_X1 U9330 ( .A1(n7424), .A2(n7423), .ZN(n9083) );
  NAND2_X1 U9331 ( .A1(n7550), .A2(n7465), .ZN(n7549) );
  NAND2_X1 U9332 ( .A1(n10849), .A2(n10848), .ZN(n7788) );
  NAND2_X1 U9333 ( .A1(n7777), .A2(n7773), .ZN(n11140) );
  NOR2_X1 U9334 ( .A1(n13644), .A2(n13645), .ZN(n13672) );
  OAI21_X1 U9335 ( .B1(n10976), .B2(n7780), .A(n7775), .ZN(n7774) );
  NOR2_X1 U9336 ( .A1(n13674), .A2(n13675), .ZN(n13694) );
  AOI21_X1 U9337 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n11340), .A(n11339), .ZN(
        n11488) );
  AOI21_X1 U9338 ( .B1(n11498), .B2(n11490), .A(n11489), .ZN(n11492) );
  NAND2_X1 U9339 ( .A1(n10423), .A2(n7232), .ZN(n7411) );
  NAND2_X1 U9340 ( .A1(n12437), .A2(n12869), .ZN(n7952) );
  NAND3_X1 U9341 ( .A1(n7414), .A2(n8924), .A3(n8925), .ZN(n8951) );
  NAND2_X1 U9342 ( .A1(n7416), .A2(n8952), .ZN(n7414) );
  INV_X1 U9343 ( .A(n9039), .ZN(n7974) );
  NAND2_X1 U9344 ( .A1(n15255), .A2(n15254), .ZN(n15253) );
  NAND2_X1 U9345 ( .A1(n7963), .A2(n7961), .ZN(n12924) );
  OAI21_X2 U9346 ( .B1(n12510), .B2(n8038), .A(n8039), .ZN(n10152) );
  NAND2_X1 U9347 ( .A1(n7419), .A2(n7418), .ZN(n15002) );
  AND2_X4 U9348 ( .A1(n12672), .A2(n12676), .ZN(n10188) );
  NAND2_X1 U9349 ( .A1(n10792), .A2(n9869), .ZN(n10987) );
  NAND2_X1 U9350 ( .A1(n10217), .A2(n8027), .ZN(n7419) );
  NAND2_X1 U9351 ( .A1(n10987), .A2(n10988), .ZN(n10986) );
  XNOR2_X1 U9352 ( .A(n9890), .B(n9889), .ZN(n10988) );
  NAND2_X1 U9353 ( .A1(n11622), .A2(n7469), .ZN(n11623) );
  NAND2_X1 U9354 ( .A1(n11962), .A2(n13415), .ZN(n12166) );
  OAI21_X2 U9355 ( .B1(n12969), .B2(n14002), .A(n12968), .ZN(n13214) );
  NAND2_X1 U9356 ( .A1(n13913), .A2(n13912), .ZN(n13911) );
  NAND2_X1 U9357 ( .A1(n13971), .A2(n12939), .ZN(n13957) );
  NAND2_X2 U9358 ( .A1(n8262), .A2(n7309), .ZN(n8283) );
  NOR2_X1 U9359 ( .A1(n14555), .A2(n8063), .ZN(n14534) );
  NAND2_X1 U9360 ( .A1(n7680), .A2(n7679), .ZN(n7678) );
  NAND2_X1 U9361 ( .A1(n10826), .A2(n10825), .ZN(n11042) );
  NAND2_X1 U9362 ( .A1(n9515), .A2(n9514), .ZN(n9529) );
  AOI21_X1 U9363 ( .B1(n9397), .B2(n9398), .A(n7438), .ZN(n7447) );
  INV_X8 U9364 ( .A(n10188), .ZN(n14954) );
  NOR2_X1 U9365 ( .A1(n15024), .A2(n15025), .ZN(n15023) );
  NOR2_X2 U9366 ( .A1(n10035), .A2(n9780), .ZN(n9823) );
  NAND2_X1 U9367 ( .A1(n14503), .A2(n14502), .ZN(n14668) );
  INV_X1 U9368 ( .A(n7802), .ZN(n7801) );
  NAND2_X1 U9369 ( .A1(n12015), .A2(n12014), .ZN(n12117) );
  NAND2_X1 U9370 ( .A1(n15046), .A2(n10155), .ZN(n14984) );
  NAND2_X1 U9371 ( .A1(n11715), .A2(n11714), .ZN(n11718) );
  NAND2_X1 U9372 ( .A1(n9738), .A2(n9739), .ZN(n7431) );
  NAND2_X1 U9373 ( .A1(n11609), .A2(n12858), .ZN(n7949) );
  NAND2_X1 U9374 ( .A1(n11000), .A2(n10999), .ZN(n7936) );
  OAI22_X2 U9375 ( .A1(n11358), .A2(n11357), .B1(n11356), .B2(n15906), .ZN(
        n11439) );
  XNOR2_X2 U9376 ( .A(n7432), .B(n7277), .ZN(n10423) );
  INV_X1 U9377 ( .A(n9035), .ZN(n9036) );
  NAND2_X1 U9378 ( .A1(n9039), .A2(n9035), .ZN(n7434) );
  NAND2_X1 U9379 ( .A1(n8151), .A2(n7510), .ZN(n7833) );
  INV_X1 U9380 ( .A(n11651), .ZN(n8180) );
  INV_X1 U9381 ( .A(n8283), .ZN(n7509) );
  NOR2_X1 U9382 ( .A1(n10718), .A2(n8458), .ZN(n7796) );
  NOR2_X2 U9383 ( .A1(n10970), .A2(n10971), .ZN(n11144) );
  NOR2_X2 U9384 ( .A1(n13596), .A2(n13595), .ZN(n13597) );
  NAND2_X1 U9385 ( .A1(n14312), .A2(n7366), .ZN(n14310) );
  NOR2_X2 U9386 ( .A1(n14326), .A2(n14325), .ZN(n14324) );
  AOI21_X2 U9387 ( .B1(n7437), .B2(n7304), .A(n7436), .ZN(n12277) );
  NAND2_X1 U9388 ( .A1(n14210), .A2(n7442), .ZN(n14290) );
  NAND2_X1 U9389 ( .A1(n11595), .A2(n11596), .ZN(n11692) );
  NAND2_X1 U9390 ( .A1(n14201), .A2(n14202), .ZN(n7444) );
  NAND2_X1 U9391 ( .A1(n10760), .A2(n10759), .ZN(n10931) );
  OAI21_X2 U9392 ( .B1(n13885), .B2(n13791), .A(n13790), .ZN(n14018) );
  INV_X1 U9393 ( .A(n12242), .ZN(n7851) );
  INV_X1 U9394 ( .A(n9400), .ZN(n9397) );
  NAND2_X1 U9395 ( .A1(n9084), .A2(n9083), .ZN(n9108) );
  NAND2_X1 U9396 ( .A1(n7439), .A2(n8134), .ZN(n9009) );
  NAND2_X1 U9397 ( .A1(n8926), .A2(n8906), .ZN(n7440) );
  AND2_X1 U9398 ( .A1(n10680), .A2(n10666), .ZN(n10675) );
  NAND2_X1 U9399 ( .A1(n7879), .A2(n7878), .ZN(n11595) );
  NAND3_X1 U9400 ( .A1(n7444), .A2(n14238), .A3(n14311), .ZN(n7484) );
  NAND2_X1 U9401 ( .A1(n8690), .A2(n8689), .ZN(n8692) );
  NAND2_X1 U9402 ( .A1(n7445), .A2(n8329), .ZN(n8331) );
  INV_X1 U9403 ( .A(n8328), .ZN(n7445) );
  NAND2_X1 U9404 ( .A1(n8705), .A2(n8106), .ZN(n8104) );
  NOR2_X2 U9405 ( .A1(n13520), .A2(n13516), .ZN(n13554) );
  OAI21_X2 U9406 ( .B1(n8659), .B2(n8658), .A(n8660), .ZN(n8661) );
  NOR2_X1 U9407 ( .A1(n9163), .A2(n8144), .ZN(n7518) );
  NAND3_X1 U9408 ( .A1(n11430), .A2(n8886), .A3(n12410), .ZN(n10771) );
  INV_X1 U9409 ( .A(n9305), .ZN(n8846) );
  NAND2_X1 U9410 ( .A1(n8844), .A2(n9193), .ZN(n9305) );
  NAND2_X1 U9411 ( .A1(n9401), .A2(n7354), .ZN(n7448) );
  NAND2_X1 U9412 ( .A1(n7451), .A2(n7450), .ZN(n7519) );
  NAND2_X1 U9413 ( .A1(n8966), .A2(n8965), .ZN(n7451) );
  INV_X1 U9414 ( .A(n7207), .ZN(n7452) );
  XNOR2_X2 U9415 ( .A(n7731), .B(n9767), .ZN(n10231) );
  INV_X1 U9416 ( .A(n14984), .ZN(n7454) );
  NAND2_X1 U9417 ( .A1(n12078), .A2(n10053), .ZN(n12260) );
  XNOR2_X1 U9418 ( .A(n7456), .B(n7455), .ZN(n13752) );
  AND2_X1 U9419 ( .A1(n13750), .A2(n13749), .ZN(n7457) );
  NAND2_X1 U9420 ( .A1(n15398), .A2(n16119), .ZN(n7945) );
  INV_X1 U9421 ( .A(n7969), .ZN(n15201) );
  INV_X1 U9422 ( .A(n11337), .ZN(n7463) );
  NAND2_X1 U9423 ( .A1(n7718), .A2(n7717), .ZN(n15796) );
  INV_X1 U9424 ( .A(n10884), .ZN(n7744) );
  NAND2_X1 U9425 ( .A1(n15704), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U9426 ( .A1(n7748), .A2(n7747), .ZN(n7746) );
  OAI21_X2 U9427 ( .B1(n15785), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n15784), .ZN(
        n15791) );
  NAND2_X1 U9428 ( .A1(n9847), .A2(n9848), .ZN(n9849) );
  NAND2_X1 U9429 ( .A1(n7786), .A2(n10876), .ZN(n10874) );
  AND2_X1 U9430 ( .A1(n13697), .A2(n13696), .ZN(n7466) );
  OR2_X2 U9431 ( .A1(n13692), .A2(n13693), .ZN(n13721) );
  XNOR2_X1 U9432 ( .A(n13715), .B(n13727), .ZN(n13692) );
  NAND2_X1 U9433 ( .A1(n7750), .A2(n7749), .ZN(n7748) );
  NOR2_X1 U9434 ( .A1(n13669), .A2(n13668), .ZN(n13691) );
  NAND2_X1 U9435 ( .A1(n7477), .A2(n7474), .ZN(n9370) );
  NAND2_X1 U9436 ( .A1(n13854), .A2(n7491), .ZN(n13842) );
  XNOR2_X1 U9437 ( .A(n7833), .B(n13208), .ZN(P3_U3488) );
  NAND2_X1 U9438 ( .A1(n7509), .A2(n8263), .ZN(n8305) );
  NAND2_X1 U9439 ( .A1(n11890), .A2(n11889), .ZN(n11962) );
  NAND2_X1 U9440 ( .A1(n13856), .A2(n13855), .ZN(n13854) );
  INV_X1 U9441 ( .A(n11619), .ZN(n11682) );
  NAND2_X1 U9442 ( .A1(n8334), .A2(n7471), .ZN(n11619) );
  NAND2_X1 U9443 ( .A1(n15685), .A2(n15686), .ZN(n15687) );
  NAND2_X1 U9444 ( .A1(n15676), .A2(n15675), .ZN(n15685) );
  NAND2_X1 U9445 ( .A1(n15782), .A2(n15783), .ZN(n15784) );
  XOR2_X1 U9446 ( .A(n15662), .B(n15663), .Z(n15659) );
  NOR2_X2 U9447 ( .A1(n15718), .A2(n15719), .ZN(n15720) );
  NOR2_X1 U9448 ( .A1(n15661), .A2(n15828), .ZN(n15667) );
  XNOR2_X1 U9449 ( .A(n7472), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9450 ( .A1(n15822), .A2(n15821), .ZN(n7473) );
  INV_X1 U9451 ( .A(n15683), .ZN(n7723) );
  INV_X1 U9452 ( .A(n15824), .ZN(n7714) );
  OAI21_X1 U9453 ( .B1(n9009), .B2(n9008), .A(n7281), .ZN(n8143) );
  NAND3_X1 U9454 ( .A1(n9323), .A2(n9322), .A3(n7352), .ZN(n7477) );
  NAND2_X1 U9455 ( .A1(n8120), .A2(n8119), .ZN(n9510) );
  NAND2_X1 U9456 ( .A1(n7732), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U9457 ( .A1(n14936), .A2(n9926), .ZN(n11283) );
  NAND2_X1 U9458 ( .A1(n7480), .A2(n7478), .ZN(P1_U3214) );
  NAND2_X1 U9459 ( .A1(n14917), .A2(n16093), .ZN(n7480) );
  NAND3_X1 U9460 ( .A1(n8111), .A2(n8734), .A3(n8110), .ZN(n8109) );
  NAND2_X1 U9461 ( .A1(n8102), .A2(n8533), .ZN(n8537) );
  NAND2_X1 U9462 ( .A1(n8448), .A2(n8447), .ZN(n8118) );
  INV_X1 U9463 ( .A(n12986), .ZN(n7844) );
  NAND2_X1 U9464 ( .A1(n7484), .A2(n7482), .ZN(P2_U3186) );
  NAND2_X1 U9465 ( .A1(n7873), .A2(n10668), .ZN(n10749) );
  NAND2_X1 U9466 ( .A1(n14287), .A2(n7485), .ZN(n14326) );
  NAND2_X1 U9467 ( .A1(n9692), .A2(n7486), .ZN(n9722) );
  NAND2_X1 U9468 ( .A1(n7520), .A2(n8139), .ZN(n9270) );
  NAND2_X1 U9469 ( .A1(n7516), .A2(n7513), .ZN(n9215) );
  NAND2_X1 U9470 ( .A1(n8896), .A2(n8895), .ZN(n8936) );
  AOI21_X2 U9471 ( .B1(n13824), .B2(n12948), .A(n7493), .ZN(n13810) );
  NAND2_X1 U9472 ( .A1(n8869), .A2(n8870), .ZN(n14852) );
  NAND2_X1 U9473 ( .A1(n7835), .A2(n7834), .ZN(n8302) );
  NAND2_X1 U9474 ( .A1(n7518), .A2(n7517), .ZN(n7516) );
  XNOR2_X1 U9475 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8329) );
  MUX2_X1 U9476 ( .A(n13511), .B(n13510), .S(n13509), .Z(n13517) );
  NAND2_X2 U9477 ( .A1(n12553), .A2(n10094), .ZN(n12510) );
  NAND2_X1 U9478 ( .A1(n8104), .A2(n8103), .ZN(n8707) );
  NAND2_X1 U9479 ( .A1(n8084), .A2(n13554), .ZN(n8083) );
  NAND2_X1 U9480 ( .A1(n8109), .A2(n8112), .ZN(n8759) );
  INV_X1 U9481 ( .A(n8086), .ZN(n8085) );
  NAND2_X1 U9482 ( .A1(n8604), .A2(n8603), .ZN(n8606) );
  NAND2_X1 U9483 ( .A1(n8532), .A2(n8531), .ZN(n8102) );
  NOR2_X1 U9484 ( .A1(n13562), .A2(n8078), .ZN(n13569) );
  NAND2_X1 U9485 ( .A1(n7288), .A2(n7688), .ZN(n7685) );
  NAND2_X1 U9486 ( .A1(n7973), .A2(n9039), .ZN(n9062) );
  NAND2_X1 U9487 ( .A1(n7681), .A2(n14469), .ZN(n14675) );
  NAND2_X1 U9488 ( .A1(n14675), .A2(n14674), .ZN(n14472) );
  NAND2_X1 U9489 ( .A1(n14744), .A2(n14803), .ZN(n7680) );
  NAND2_X1 U9490 ( .A1(n12375), .A2(n12866), .ZN(n12377) );
  NAND2_X1 U9491 ( .A1(n16120), .A2(n7334), .ZN(n12607) );
  AND2_X2 U9492 ( .A1(n9732), .A2(n9731), .ZN(n9992) );
  NAND2_X2 U9493 ( .A1(n8231), .A2(n9992), .ZN(n10035) );
  INV_X1 U9494 ( .A(n9059), .ZN(n7512) );
  INV_X1 U9495 ( .A(n9164), .ZN(n7517) );
  NAND2_X1 U9496 ( .A1(n7506), .A2(n7503), .ZN(P2_U3494) );
  OR2_X1 U9497 ( .A1(n14823), .A2(n16157), .ZN(n7506) );
  NAND2_X2 U9498 ( .A1(n9016), .A2(n9015), .ZN(n9037) );
  OAI21_X2 U9499 ( .B1(n9403), .B2(n7982), .A(n7977), .ZN(n9449) );
  AOI21_X1 U9500 ( .B1(n9108), .B2(n9107), .A(n9106), .ZN(n9109) );
  XNOR2_X1 U9501 ( .A(n10152), .B(n10151), .ZN(n15044) );
  NAND3_X1 U9502 ( .A1(n9220), .A2(n9219), .A3(n7351), .ZN(n7520) );
  NAND3_X1 U9503 ( .A1(n9739), .A2(n9740), .A3(n9738), .ZN(n9743) );
  INV_X1 U9504 ( .A(n8703), .ZN(n7536) );
  NAND2_X1 U9505 ( .A1(n13316), .A2(n13846), .ZN(n7531) );
  AND2_X1 U9506 ( .A1(n7531), .A2(n7536), .ZN(n13287) );
  AOI21_X1 U9507 ( .B1(n7536), .B2(n7492), .A(n8732), .ZN(n7532) );
  AND2_X1 U9508 ( .A1(n7538), .A2(n11208), .ZN(n7537) );
  OAI21_X1 U9509 ( .B1(n8183), .B2(n7537), .A(n8398), .ZN(n11943) );
  INV_X1 U9510 ( .A(n7540), .ZN(n13298) );
  INV_X1 U9511 ( .A(n8148), .ZN(n7545) );
  NAND3_X1 U9512 ( .A1(n7557), .A2(n7556), .A3(n7367), .ZN(n12048) );
  INV_X1 U9513 ( .A(n7561), .ZN(n13627) );
  NAND2_X1 U9514 ( .A1(n7561), .A2(n7560), .ZN(n7789) );
  INV_X1 U9515 ( .A(n13626), .ZN(n7560) );
  OR2_X1 U9516 ( .A1(n13623), .A2(n13624), .ZN(n7561) );
  OR3_X1 U9517 ( .A1(n8591), .A2(n8291), .A3(n7565), .ZN(n8295) );
  NAND2_X4 U9518 ( .A1(n8301), .A2(n7566), .ZN(n8790) );
  INV_X1 U9519 ( .A(n12659), .ZN(n7576) );
  AOI21_X2 U9520 ( .B1(n7217), .B2(n7240), .A(n7577), .ZN(n15186) );
  AND2_X1 U9521 ( .A1(n15425), .A2(n15058), .ZN(n7580) );
  NAND2_X1 U9522 ( .A1(n12386), .A2(n7583), .ZN(n7582) );
  NAND2_X2 U9523 ( .A1(n9903), .A2(n7585), .ZN(n15906) );
  AND2_X1 U9524 ( .A1(n12822), .A2(n12823), .ZN(n7589) );
  INV_X1 U9525 ( .A(n12827), .ZN(n7592) );
  NAND2_X1 U9526 ( .A1(n12742), .A2(n7594), .ZN(n7593) );
  NAND2_X1 U9527 ( .A1(n7593), .A2(n7353), .ZN(n8209) );
  AND2_X1 U9528 ( .A1(n12741), .A2(n7598), .ZN(n7597) );
  NAND2_X1 U9529 ( .A1(n12776), .A2(n7601), .ZN(n7600) );
  NAND2_X1 U9530 ( .A1(n7606), .A2(n7607), .ZN(n8211) );
  NAND2_X1 U9531 ( .A1(n12768), .A2(n7609), .ZN(n7606) );
  NAND2_X1 U9532 ( .A1(n12753), .A2(n7615), .ZN(n7614) );
  OAI21_X2 U9533 ( .B1(n12843), .B2(n12838), .A(n7619), .ZN(n12702) );
  INV_X1 U9534 ( .A(n12838), .ZN(n7620) );
  MUX2_X1 U9535 ( .A(n12725), .B(n15069), .S(n12743), .Z(n12727) );
  MUX2_X1 U9536 ( .A(n10921), .B(P1_REG1_REG_1__SCAN_IN), .S(n10331), .Z(
        n10324) );
  NAND3_X1 U9537 ( .A1(n7988), .A2(n7987), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7642) );
  NAND2_X1 U9538 ( .A1(n7649), .A2(n7648), .ZN(n14503) );
  NAND2_X1 U9539 ( .A1(n7656), .A2(n7654), .ZN(n14511) );
  NAND2_X1 U9540 ( .A1(n12424), .A2(n7666), .ZN(n7663) );
  NAND2_X1 U9541 ( .A1(n7663), .A2(n7664), .ZN(n14494) );
  AND2_X2 U9542 ( .A1(n14566), .A2(n8061), .ZN(n14555) );
  NAND2_X1 U9543 ( .A1(n7288), .A2(n11402), .ZN(n7686) );
  NAND3_X1 U9544 ( .A1(n7686), .A2(n7685), .A3(n11509), .ZN(n11702) );
  NAND3_X1 U9545 ( .A1(n14330), .A2(n7449), .A3(n10683), .ZN(n10684) );
  NAND2_X1 U9546 ( .A1(n12126), .A2(n12125), .ZN(n12128) );
  NAND2_X1 U9547 ( .A1(n14558), .A2(n7699), .ZN(n14457) );
  NAND2_X1 U9548 ( .A1(n14558), .A2(n14741), .ZN(n14541) );
  NOR3_X4 U9549 ( .A1(n12120), .A2(n14359), .A3(n7704), .ZN(n14715) );
  NOR2_X2 U9550 ( .A1(n12152), .A2(n12091), .ZN(n11867) );
  XNOR2_X1 U9551 ( .A(n7723), .B(n15684), .ZN(n15676) );
  XNOR2_X1 U9552 ( .A(n15679), .B(n7722), .ZN(n15684) );
  NOR2_X2 U9553 ( .A1(n15166), .A2(n15167), .ZN(n15165) );
  NOR2_X2 U9554 ( .A1(n15192), .A2(n15413), .ZN(n12930) );
  NOR2_X2 U9555 ( .A1(n15228), .A2(n15425), .ZN(n15211) );
  NOR2_X2 U9556 ( .A1(n11568), .A2(n12709), .ZN(n11604) );
  INV_X1 U9557 ( .A(n11352), .ZN(n7736) );
  NOR2_X2 U9558 ( .A1(n11005), .A2(n12690), .ZN(n11199) );
  NOR2_X2 U9559 ( .A1(n15380), .A2(n15386), .ZN(n15382) );
  INV_X1 U9560 ( .A(n7739), .ZN(n15256) );
  NOR3_X2 U9561 ( .A1(n15326), .A2(n15444), .A3(n7740), .ZN(n7739) );
  NAND3_X1 U9562 ( .A1(n7744), .A2(n7754), .A3(n7756), .ZN(n7747) );
  INV_X1 U9563 ( .A(n7767), .ZN(n13667) );
  INV_X1 U9564 ( .A(n13633), .ZN(n7768) );
  INV_X1 U9565 ( .A(n7771), .ZN(n7769) );
  NAND2_X1 U9566 ( .A1(n7771), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U9567 ( .A1(n13597), .A2(n13617), .ZN(n7771) );
  INV_X1 U9568 ( .A(n7772), .ZN(n11138) );
  AOI21_X1 U9569 ( .B1(n10976), .B2(n10975), .A(n7780), .ZN(n7772) );
  NAND2_X1 U9570 ( .A1(n10976), .A2(n7778), .ZN(n7777) );
  INV_X1 U9571 ( .A(n7774), .ZN(n7773) );
  OAI21_X1 U9572 ( .B1(n7780), .B2(n10975), .A(P3_REG2_REG_5__SCAN_IN), .ZN(
        n7776) );
  INV_X1 U9573 ( .A(n10975), .ZN(n7779) );
  INV_X1 U9574 ( .A(n10977), .ZN(n7780) );
  NAND2_X1 U9575 ( .A1(n10876), .A2(n7787), .ZN(n10851) );
  NAND2_X1 U9576 ( .A1(n7787), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7786) );
  INV_X1 U9577 ( .A(n7789), .ZN(n13642) );
  NAND2_X1 U9578 ( .A1(n13643), .A2(n13657), .ZN(n13671) );
  INV_X1 U9579 ( .A(n11534), .ZN(n7790) );
  NAND2_X1 U9580 ( .A1(n7793), .A2(n7792), .ZN(n11535) );
  INV_X1 U9581 ( .A(n14614), .ZN(n7811) );
  NAND2_X1 U9582 ( .A1(n10694), .A2(n7822), .ZN(n7821) );
  NAND3_X1 U9583 ( .A1(n7821), .A2(n7824), .A3(n11048), .ZN(n11052) );
  OR2_X1 U9584 ( .A1(n7826), .A2(n10828), .ZN(n7824) );
  NAND2_X1 U9585 ( .A1(n10829), .A2(n10828), .ZN(n7825) );
  INV_X1 U9586 ( .A(n10831), .ZN(n7826) );
  XNOR2_X1 U9587 ( .A(n14523), .B(n7832), .ZN(n7830) );
  AOI21_X1 U9588 ( .B1(n7830), .B2(n7829), .A(n7827), .ZN(n14532) );
  AOI21_X1 U9589 ( .B1(n14735), .B2(n14667), .A(n14531), .ZN(n7831) );
  INV_X1 U9590 ( .A(n14524), .ZN(n7832) );
  INV_X1 U9591 ( .A(n8283), .ZN(n7835) );
  NAND2_X1 U9592 ( .A1(n13954), .A2(n7838), .ZN(n7836) );
  NAND2_X1 U9593 ( .A1(n12985), .A2(n12984), .ZN(n13781) );
  NAND2_X1 U9594 ( .A1(n12976), .A2(n7239), .ZN(n7856) );
  NAND2_X1 U9595 ( .A1(n12517), .A2(n13447), .ZN(n12970) );
  NAND2_X1 U9596 ( .A1(n12370), .A2(n13532), .ZN(n12516) );
  INV_X1 U9597 ( .A(n12989), .ZN(n12990) );
  NAND2_X1 U9598 ( .A1(n12981), .A2(n13500), .ZN(n13809) );
  NAND2_X1 U9599 ( .A1(n11263), .A2(n11264), .ZN(n11627) );
  NAND2_X1 U9600 ( .A1(n12982), .A2(n13493), .ZN(n13797) );
  NAND2_X1 U9601 ( .A1(n11628), .A2(n13528), .ZN(n11653) );
  NAND2_X1 U9602 ( .A1(n12516), .A2(n13439), .ZN(n13993) );
  INV_X1 U9603 ( .A(n7223), .ZN(n11263) );
  OAI21_X1 U9604 ( .B1(n13221), .B2(n14058), .A(n8228), .ZN(n12989) );
  OR2_X2 U9605 ( .A1(n14650), .A2(n14778), .ZN(n14634) );
  NOR2_X2 U9606 ( .A1(n10827), .A2(n14269), .ZN(n11056) );
  AND2_X2 U9607 ( .A1(n11409), .A2(n11807), .ZN(n11757) );
  NOR2_X2 U9608 ( .A1(n14563), .A2(n14570), .ZN(n14558) );
  NAND2_X1 U9609 ( .A1(n7233), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8319) );
  NAND2_X1 U9610 ( .A1(n7234), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8317) );
  AOI21_X2 U9611 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(n15754), .A(n15753), .ZN(
        n15761) );
  NAND2_X1 U9612 ( .A1(n11900), .A2(n13393), .ZN(n11628) );
  OAI21_X1 U9613 ( .B1(n7873), .B2(n10668), .A(n10749), .ZN(n10669) );
  NAND2_X1 U9614 ( .A1(n14264), .A2(n7345), .ZN(n7874) );
  NAND2_X1 U9615 ( .A1(n11310), .A2(n7880), .ZN(n7879) );
  NAND2_X1 U9616 ( .A1(n7882), .A2(n14228), .ZN(n14231) );
  NAND2_X1 U9617 ( .A1(n14345), .A2(n7245), .ZN(n7882) );
  NAND2_X1 U9618 ( .A1(n14345), .A2(n7885), .ZN(n14201) );
  NAND2_X1 U9619 ( .A1(n12277), .A2(n7321), .ZN(n7887) );
  NAND2_X1 U9620 ( .A1(n7887), .A2(n7251), .ZN(n14164) );
  INV_X1 U9621 ( .A(n7895), .ZN(n14352) );
  OR2_X1 U9622 ( .A1(n12534), .A2(n12535), .ZN(n7896) );
  INV_X1 U9623 ( .A(n7908), .ZN(n14183) );
  NAND2_X1 U9624 ( .A1(n8846), .A2(n8135), .ZN(n8136) );
  NAND2_X1 U9625 ( .A1(n8848), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8847) );
  OAI211_X2 U9626 ( .C1(n9846), .C2(n10246), .A(n7913), .B(n7912), .ZN(n12674)
         );
  OR2_X1 U9627 ( .A1(n7235), .A2(n7646), .ZN(n7913) );
  XNOR2_X2 U9628 ( .A(n7914), .B(n15182), .ZN(n15407) );
  NAND2_X1 U9629 ( .A1(n7915), .A2(n11001), .ZN(n11197) );
  INV_X1 U9630 ( .A(n7927), .ZN(n15239) );
  NAND2_X1 U9631 ( .A1(n15306), .A2(n7339), .ZN(n15293) );
  NAND2_X1 U9632 ( .A1(n7934), .A2(n7933), .ZN(n15973) );
  NAND2_X1 U9633 ( .A1(n7936), .A2(n12854), .ZN(n11201) );
  XNOR2_X1 U9634 ( .A(n7936), .B(n12854), .ZN(n11004) );
  XNOR2_X2 U9635 ( .A(n9757), .B(n9756), .ZN(n15508) );
  AOI21_X1 U9636 ( .B1(n7939), .B2(n7941), .A(n7318), .ZN(n7937) );
  INV_X1 U9637 ( .A(n15982), .ZN(n7944) );
  NAND2_X1 U9638 ( .A1(n7942), .A2(n7943), .ZN(n11970) );
  NAND2_X1 U9639 ( .A1(n15982), .A2(n11932), .ZN(n7942) );
  AOI21_X1 U9640 ( .B1(n15983), .B2(n11932), .A(n7297), .ZN(n7943) );
  XNOR2_X1 U9641 ( .A(n15183), .B(n15182), .ZN(n15398) );
  NAND3_X1 U9642 ( .A1(n9739), .A2(n9738), .A3(n8221), .ZN(n9754) );
  NAND2_X1 U9643 ( .A1(n7949), .A2(n7947), .ZN(n11929) );
  NAND2_X1 U9644 ( .A1(n7952), .A2(n7950), .ZN(n12604) );
  NAND2_X1 U9645 ( .A1(n15302), .A2(n7955), .ZN(n7954) );
  INV_X1 U9646 ( .A(n7960), .ZN(n15286) );
  NAND2_X1 U9647 ( .A1(n15222), .A2(n7964), .ZN(n7963) );
  NAND2_X2 U9648 ( .A1(n12673), .A2(n10905), .ZN(n12683) );
  NAND2_X2 U9649 ( .A1(n10903), .A2(n10904), .ZN(n12673) );
  NAND2_X1 U9650 ( .A1(n9037), .A2(n7242), .ZN(n7971) );
  INV_X1 U9651 ( .A(n9405), .ZN(n7984) );
  MUX2_X1 U9652 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n8315), .Z(n8970) );
  NAND2_X1 U9653 ( .A1(n9562), .A2(n9561), .ZN(n9596) );
  NAND3_X1 U9654 ( .A1(n9597), .A2(n9598), .A3(n7232), .ZN(n12841) );
  INV_X1 U9655 ( .A(n9595), .ZN(n8014) );
  NAND2_X1 U9656 ( .A1(n14976), .A2(n7273), .ZN(n8015) );
  NAND2_X1 U9657 ( .A1(n8015), .A2(n8016), .ZN(n14915) );
  NOR2_X1 U9658 ( .A1(n14887), .A2(n14886), .ZN(n14926) );
  NAND2_X1 U9659 ( .A1(n14952), .A2(n8030), .ZN(n8029) );
  OAI211_X1 U9660 ( .C1(n14952), .C2(n8031), .A(n8029), .B(n14965), .ZN(
        P1_U3220) );
  NOR2_X1 U9661 ( .A1(n14958), .A2(n14951), .ZN(n8035) );
  NAND2_X1 U9662 ( .A1(n14958), .A2(n14951), .ZN(n8036) );
  NAND2_X1 U9663 ( .A1(n14946), .A2(n8044), .ZN(n8042) );
  NAND2_X1 U9664 ( .A1(n8878), .A2(n8880), .ZN(n8049) );
  NAND2_X1 U9665 ( .A1(n8879), .A2(n8880), .ZN(n8050) );
  XNOR2_X2 U9666 ( .A(n8052), .B(n8883), .ZN(n14868) );
  INV_X2 U9667 ( .A(n10428), .ZN(n9353) );
  NAND3_X1 U9668 ( .A1(n11707), .A2(n7820), .A3(n11706), .ZN(n11854) );
  INV_X1 U9669 ( .A(n12128), .ZN(n8077) );
  OAI21_X1 U9670 ( .B1(n13502), .B2(n13509), .A(n13544), .ZN(n8087) );
  NAND2_X1 U9671 ( .A1(n13498), .A2(n13497), .ZN(n8088) );
  NAND2_X1 U9672 ( .A1(n13501), .A2(n8090), .ZN(n8089) );
  NAND3_X1 U9673 ( .A1(n8097), .A2(n8098), .A3(n8571), .ZN(n8588) );
  NAND2_X1 U9674 ( .A1(n8557), .A2(n8099), .ZN(n8097) );
  NAND2_X1 U9675 ( .A1(n8100), .A2(n8559), .ZN(n8570) );
  OAI21_X2 U9676 ( .B1(n8508), .B2(n8507), .A(n8509), .ZN(n8532) );
  OAI22_X2 U9677 ( .A1(n8661), .A2(n8115), .B1(n11428), .B2(
        P2_DATAO_REG_20__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U9678 ( .A1(n9469), .A2(n7337), .ZN(n8120) );
  NAND2_X1 U9679 ( .A1(n8127), .A2(n7344), .ZN(n9692) );
  NAND2_X1 U9680 ( .A1(n9532), .A2(n9531), .ZN(n8128) );
  NAND2_X1 U9681 ( .A1(n9534), .A2(n9533), .ZN(n8129) );
  INV_X1 U9682 ( .A(n9692), .ZN(n9668) );
  NAND2_X1 U9683 ( .A1(n8846), .A2(n7250), .ZN(n8852) );
  INV_X1 U9684 ( .A(n9421), .ZN(n8137) );
  NAND2_X1 U9685 ( .A1(n9215), .A2(n9216), .ZN(n9214) );
  NAND2_X1 U9686 ( .A1(n9319), .A2(n9315), .ZN(n9318) );
  AOI21_X1 U9687 ( .B1(n8146), .B2(n11189), .A(n8338), .ZN(n11208) );
  XNOR2_X1 U9688 ( .A(n8146), .B(n8145), .ZN(n11194) );
  INV_X1 U9689 ( .A(n11189), .ZN(n8145) );
  NAND2_X1 U9690 ( .A1(n11071), .A2(n8322), .ZN(n8146) );
  INV_X1 U9691 ( .A(n13214), .ZN(n8152) );
  NAND2_X1 U9692 ( .A1(n13214), .A2(n16061), .ZN(n8151) );
  NAND2_X1 U9693 ( .A1(n13341), .A2(n7272), .ZN(n8153) );
  NAND2_X1 U9694 ( .A1(n8153), .A2(n8154), .ZN(n13280) );
  NAND2_X1 U9695 ( .A1(n13332), .A2(n7338), .ZN(n8158) );
  OAI211_X1 U9696 ( .C1(n13332), .C2(n8159), .A(n13343), .B(n8158), .ZN(n8835)
         );
  NAND2_X1 U9697 ( .A1(n8776), .A2(n12951), .ZN(n8169) );
  NAND2_X1 U9698 ( .A1(n12524), .A2(n12937), .ZN(n8172) );
  NAND2_X1 U9699 ( .A1(n8176), .A2(n7296), .ZN(n12243) );
  NAND2_X1 U9700 ( .A1(n12166), .A2(n13529), .ZN(n8176) );
  NOR2_X1 U9701 ( .A1(n13533), .A2(n8180), .ZN(n8179) );
  INV_X1 U9702 ( .A(n13940), .ZN(n8195) );
  NAND2_X1 U9703 ( .A1(n8262), .A2(n8261), .ZN(n8278) );
  OAI21_X1 U9704 ( .B1(n12785), .B2(n12784), .A(n12788), .ZN(n12790) );
  NAND3_X1 U9705 ( .A1(n12814), .A2(n12813), .A3(n7356), .ZN(n8203) );
  INV_X1 U9706 ( .A(n12815), .ZN(n8204) );
  NAND2_X1 U9707 ( .A1(n8209), .A2(n8210), .ZN(n12753) );
  NAND2_X1 U9708 ( .A1(n8211), .A2(n8212), .ZN(n12776) );
  NAND2_X1 U9709 ( .A1(n8213), .A2(n8214), .ZN(n12730) );
  NAND3_X1 U9710 ( .A1(n12724), .A2(n12723), .A3(n7348), .ZN(n8213) );
  NAND2_X1 U9711 ( .A1(n8216), .A2(n8215), .ZN(n12742) );
  NAND3_X1 U9712 ( .A1(n12735), .A2(n8217), .A3(n12734), .ZN(n8216) );
  NAND2_X1 U9713 ( .A1(n12736), .A2(n8219), .ZN(n8218) );
  NAND2_X1 U9714 ( .A1(n12801), .A2(n12802), .ZN(n12800) );
  OAI21_X1 U9715 ( .B1(n15417), .B2(n12928), .A(n12927), .ZN(n12929) );
  NOR2_X1 U9716 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n8251) );
  NAND4_X2 U9717 ( .A1(n8275), .A2(n8274), .A3(n8273), .A4(n8272), .ZN(n13588)
         );
  AND2_X1 U9718 ( .A1(n11854), .A2(n11709), .ZN(n12096) );
  NAND2_X1 U9719 ( .A1(n8590), .A2(n8589), .ZN(n8604) );
  NAND2_X1 U9720 ( .A1(n8588), .A2(n8587), .ZN(n8590) );
  XNOR2_X2 U9721 ( .A(n15072), .B(n11440), .ZN(n12856) );
  NAND4_X4 U9722 ( .A1(n9918), .A2(n9917), .A3(n9916), .A4(n9915), .ZN(n15072)
         );
  INV_X1 U9723 ( .A(n8687), .ZN(n8690) );
  INV_X1 U9724 ( .A(n9629), .ZN(n8942) );
  NAND2_X1 U9725 ( .A1(n9509), .A2(n9508), .ZN(n9515) );
  INV_X1 U9726 ( .A(n8848), .ZN(n8850) );
  INV_X1 U9727 ( .A(n8446), .ZN(n8448) );
  NAND2_X1 U9728 ( .A1(n8761), .A2(n8760), .ZN(n8764) );
  NAND2_X1 U9729 ( .A1(n14096), .A2(n12951), .ZN(n12952) );
  NAND2_X1 U9730 ( .A1(n8302), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8304) );
  OR2_X1 U9731 ( .A1(n9629), .A2(n10438), .ZN(n8874) );
  NAND2_X1 U9732 ( .A1(n12812), .A2(n12811), .ZN(n12813) );
  NOR2_X1 U9733 ( .A1(n10309), .A2(n10308), .ZN(n10547) );
  NAND2_X1 U9734 ( .A1(n8852), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U9735 ( .A1(n8305), .A2(n8285), .ZN(n12401) );
  INV_X1 U9736 ( .A(n8887), .ZN(n10475) );
  NAND4_X2 U9737 ( .A1(n9857), .A2(n9856), .A3(n9855), .A4(n9854), .ZN(n10907)
         );
  NOR2_X1 U9738 ( .A1(n13553), .A2(n13552), .ZN(n13558) );
  AOI21_X2 U9739 ( .B1(n12243), .B2(n12212), .A(n8230), .ZN(n12367) );
  OR2_X1 U9740 ( .A1(n12988), .A2(n16054), .ZN(n8228) );
  INV_X1 U9741 ( .A(n8438), .ZN(n8614) );
  NAND2_X1 U9742 ( .A1(n14051), .A2(n13881), .ZN(n8229) );
  INV_X1 U9743 ( .A(n9872), .ZN(n9893) );
  INV_X1 U9744 ( .A(n15075), .ZN(n10904) );
  NOR2_X1 U9745 ( .A1(n12211), .A2(n12210), .ZN(n8230) );
  AND2_X1 U9746 ( .A1(n8880), .A2(n8883), .ZN(n8232) );
  AND2_X1 U9747 ( .A1(n11219), .A2(n11218), .ZN(n8233) );
  AND3_X1 U9748 ( .A1(n9716), .A2(n9715), .A3(n9714), .ZN(n8234) );
  NOR2_X1 U9749 ( .A1(n13892), .A2(n12975), .ZN(n8237) );
  NOR2_X1 U9750 ( .A1(n12975), .A2(n12974), .ZN(n8238) );
  OR2_X1 U9751 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(n7257), .ZN(n8239) );
  AND2_X1 U9752 ( .A1(n14478), .A2(n14633), .ZN(n8240) );
  INV_X1 U9753 ( .A(n15074), .ZN(n10994) );
  INV_X1 U9754 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8469) );
  XOR2_X1 U9755 ( .A(n14769), .B(n10662), .Z(n8241) );
  AND2_X1 U9756 ( .A1(n10751), .A2(n10750), .ZN(n8242) );
  AND2_X1 U9757 ( .A1(n13393), .A2(n13395), .ZN(n8243) );
  INV_X1 U9758 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14853) );
  AND2_X1 U9759 ( .A1(n9191), .A2(n9170), .ZN(n8244) );
  INV_X1 U9760 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9741) );
  INV_X1 U9761 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8391) );
  OR2_X1 U9762 ( .A1(n7206), .A2(n10775), .ZN(n8245) );
  AND2_X1 U9763 ( .A1(n12755), .A2(n15374), .ZN(n8246) );
  INV_X1 U9764 ( .A(n15983), .ZN(n11930) );
  INV_X1 U9765 ( .A(n15408), .ZN(n15176) );
  NAND2_X1 U9766 ( .A1(n9717), .A2(n9693), .ZN(n8247) );
  INV_X1 U9767 ( .A(n10630), .ZN(n13603) );
  AND2_X1 U9768 ( .A1(n14814), .A2(n14813), .ZN(n8248) );
  AND2_X1 U9769 ( .A1(n15474), .A2(n15360), .ZN(n8249) );
  AND2_X2 U9770 ( .A1(n11638), .A2(n11186), .ZN(n16061) );
  AOI22_X1 U9771 ( .A1(n14375), .A2(n8885), .B1(n7206), .B2(n10587), .ZN(n8938) );
  OAI21_X1 U9772 ( .B1(n15073), .B2(n12826), .A(n15906), .ZN(n12697) );
  AOI21_X1 U9773 ( .B1(n9009), .B2(n9008), .A(n9007), .ZN(n9010) );
  INV_X1 U9774 ( .A(n13826), .ZN(n12946) );
  NAND2_X1 U9775 ( .A1(n14035), .A2(n12946), .ZN(n12947) );
  NAND2_X1 U9776 ( .A1(n9513), .A2(n9512), .ZN(n9514) );
  OR4_X1 U9777 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10457) );
  OR4_X1 U9778 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10206) );
  INV_X1 U9779 ( .A(n13527), .ZN(n12169) );
  INV_X1 U9780 ( .A(n15401), .ZN(n15177) );
  INV_X1 U9781 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n15670) );
  INV_X1 U9782 ( .A(n13574), .ZN(n12951) );
  INV_X1 U9783 ( .A(n9359), .ZN(n9357) );
  INV_X1 U9784 ( .A(n14367), .ZN(n11720) );
  INV_X1 U9785 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8849) );
  INV_X1 U9786 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9935) );
  INV_X1 U9787 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9832) );
  INV_X1 U9788 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9999) );
  INV_X1 U9789 ( .A(n11062), .ZN(n10998) );
  NAND2_X1 U9790 ( .A1(n9299), .A2(n13119), .ZN(n9324) );
  INV_X1 U9791 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12995) );
  NOR2_X1 U9792 ( .A1(n8737), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8750) );
  OR2_X1 U9793 ( .A1(n14152), .A2(n8327), .ZN(n12962) );
  AND2_X1 U9794 ( .A1(n13500), .A2(n13499), .ZN(n13825) );
  INV_X1 U9795 ( .A(n13540), .ZN(n13878) );
  INV_X1 U9796 ( .A(n11430), .ZN(n10646) );
  OR2_X1 U9797 ( .A1(n9523), .A2(n9522), .ZN(n9583) );
  OR2_X1 U9798 ( .A1(n9477), .A2(n14291), .ZN(n9498) );
  OR2_X1 U9799 ( .A1(n9410), .A2(n14244), .ZN(n9434) );
  NAND2_X1 U9800 ( .A1(n9308), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9332) );
  AND2_X1 U9801 ( .A1(n15624), .A2(n11083), .ZN(n15605) );
  INV_X1 U9802 ( .A(n10646), .ZN(n10467) );
  NAND2_X1 U9803 ( .A1(n14528), .A2(n14527), .ZN(n14529) );
  AND2_X1 U9804 ( .A1(n10655), .A2(n9708), .ZN(n14525) );
  INV_X1 U9805 ( .A(n14364), .ZN(n12184) );
  INV_X1 U9806 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9662) );
  INV_X1 U9807 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10101) );
  INV_X1 U9808 ( .A(n11667), .ZN(n10010) );
  OR2_X1 U9809 ( .A1(n14893), .A2(n14892), .ZN(n14894) );
  INV_X1 U9810 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10017) );
  INV_X1 U9811 ( .A(n12556), .ZN(n10089) );
  INV_X1 U9812 ( .A(n12582), .ZN(n12592) );
  NAND2_X1 U9813 ( .A1(n9804), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U9814 ( .A1(n15176), .A2(n15401), .ZN(n15180) );
  INV_X1 U9815 ( .A(n15338), .ZN(n12657) );
  INV_X1 U9816 ( .A(n12864), .ZN(n11918) );
  NAND2_X1 U9817 ( .A1(n11200), .A2(n10995), .ZN(n11001) );
  NOR2_X1 U9818 ( .A1(n15405), .A2(n15404), .ZN(n15406) );
  OR2_X1 U9819 ( .A1(n12747), .A2(n15065), .ZN(n12385) );
  OR2_X1 U9820 ( .A1(n15974), .A2(n7228), .ZN(n11018) );
  INV_X1 U9821 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9767) );
  NAND2_X1 U9822 ( .A1(n9449), .A2(SI_22_), .ZN(n9450) );
  INV_X1 U9823 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n15677) );
  NOR2_X1 U9824 ( .A1(n15724), .A2(n15723), .ZN(n15725) );
  OR2_X1 U9825 ( .A1(n8563), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8576) );
  NOR2_X1 U9826 ( .A1(n8650), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8666) );
  AND2_X1 U9827 ( .A1(n8594), .A2(n12995), .ZN(n8615) );
  NAND2_X1 U9828 ( .A1(n8615), .A2(n13182), .ZN(n8632) );
  INV_X1 U9829 ( .A(n13915), .ZN(n13881) );
  OR2_X1 U9830 ( .A1(n8632), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8650) );
  AND2_X1 U9831 ( .A1(n9751), .A2(n14143), .ZN(n11176) );
  NOR2_X1 U9832 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(n8784), .ZN(n13757) );
  INV_X1 U9833 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15707) );
  INV_X1 U9834 ( .A(n15521), .ZN(n15853) );
  OR2_X1 U9835 ( .A1(n12960), .A2(n11785), .ZN(n8726) );
  OR2_X1 U9836 ( .A1(n7308), .A2(n13479), .ZN(n13867) );
  INV_X1 U9837 ( .A(n13956), .ZN(n13953) );
  INV_X1 U9838 ( .A(n13576), .ZN(n13309) );
  INV_X1 U9839 ( .A(n16061), .ZN(n12991) );
  INV_X1 U9840 ( .A(n11635), .ZN(n11184) );
  OR2_X1 U9841 ( .A1(n12960), .A2(n13112), .ZN(n8676) );
  INV_X1 U9842 ( .A(n10628), .ZN(n8646) );
  AND2_X1 U9843 ( .A1(n13448), .A2(n13445), .ZN(n13992) );
  AND2_X1 U9844 ( .A1(n11262), .A2(n11261), .ZN(n13885) );
  INV_X1 U9845 ( .A(n13386), .ZN(n13523) );
  AND2_X1 U9846 ( .A1(n13560), .A2(n11269), .ZN(n14002) );
  INV_X1 U9847 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n14304) );
  OR2_X1 U9848 ( .A1(n10657), .A2(n10649), .ZN(n14341) );
  INV_X1 U9849 ( .A(n14339), .ZN(n14351) );
  AND2_X1 U9850 ( .A1(n9583), .A2(n9524), .ZN(n14571) );
  INV_X1 U9851 ( .A(n9624), .ZN(n9546) );
  OR2_X1 U9852 ( .A1(n9285), .A2(n15589), .ZN(n9310) );
  OR2_X1 U9853 ( .A1(n15621), .A2(n15620), .ZN(n15624) );
  INV_X1 U9854 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n15589) );
  AND2_X1 U9855 ( .A1(n15530), .A2(n10432), .ZN(n10435) );
  INV_X1 U9856 ( .A(n14480), .ZN(n14515) );
  INV_X1 U9857 ( .A(n11855), .ZN(n11861) );
  INV_X1 U9858 ( .A(n14525), .ZN(n14313) );
  INV_X1 U9859 ( .A(n14493), .ZN(n14707) );
  NOR2_X1 U9860 ( .A1(n10645), .A2(n10651), .ZN(n11733) );
  NOR2_X1 U9861 ( .A1(n12256), .A2(n12199), .ZN(n9706) );
  NAND2_X1 U9862 ( .A1(n9703), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9699) );
  NAND2_X1 U9863 ( .A1(n12620), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n12637) );
  XOR2_X1 U9864 ( .A(n14957), .B(n14956), .Z(n14958) );
  NAND2_X1 U9865 ( .A1(n14911), .A2(n14912), .ZN(n15032) );
  AND2_X1 U9866 ( .A1(n12637), .A2(n12622), .ZN(n15195) );
  INV_X1 U9867 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n15664) );
  AND2_X1 U9868 ( .A1(n8048), .A2(n15513), .ZN(n10265) );
  INV_X1 U9869 ( .A(n16030), .ZN(n15357) );
  INV_X1 U9870 ( .A(n16123), .ZN(n16134) );
  INV_X1 U9871 ( .A(n15351), .ZN(n15353) );
  INV_X1 U9872 ( .A(n12869), .ZN(n12444) );
  INV_X1 U9873 ( .A(n12737), .ZN(n12868) );
  INV_X1 U9874 ( .A(n15376), .ZN(n15359) );
  INV_X1 U9875 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9879) );
  OAI21_X1 U9876 ( .B1(P3_ADDR_REG_13__SCAN_IN), .B2(n15772), .A(n15771), .ZN(
        n15778) );
  OAI21_X1 U9877 ( .B1(n14017), .B2(n13354), .A(n8832), .ZN(n8833) );
  INV_X1 U9878 ( .A(n13354), .ZN(n12565) );
  AND2_X1 U9879 ( .A1(n11176), .A2(n15940), .ZN(n11639) );
  AND4_X1 U9880 ( .A1(n8789), .A2(n8788), .A3(n8787), .A4(n8786), .ZN(n13787)
         );
  AND4_X1 U9881 ( .A1(n8723), .A2(n8722), .A3(n8721), .A4(n8720), .ZN(n13826)
         );
  AND4_X1 U9882 ( .A1(n8620), .A2(n8619), .A3(n8618), .A4(n8617), .ZN(n13943)
         );
  INV_X1 U9883 ( .A(n15843), .ZN(n15863) );
  INV_X1 U9884 ( .A(n15866), .ZN(n13722) );
  AND2_X1 U9885 ( .A1(n11639), .A2(n11683), .ZN(n14004) );
  NAND2_X1 U9886 ( .A1(n11638), .A2(n11637), .ZN(n11641) );
  OR2_X1 U9887 ( .A1(n12960), .A2(n13101), .ZN(n8766) );
  AND2_X1 U9888 ( .A1(n14075), .A2(n14074), .ZN(n14134) );
  INV_X1 U9889 ( .A(n16011), .ZN(n16059) );
  INV_X1 U9890 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8296) );
  AND2_X1 U9891 ( .A1(n10764), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14339) );
  NAND2_X1 U9892 ( .A1(n10648), .A2(n14718), .ZN(n14358) );
  OR2_X1 U9893 ( .A1(n14543), .A2(n9624), .ZN(n9591) );
  INV_X1 U9894 ( .A(n15543), .ZN(n15627) );
  INV_X1 U9895 ( .A(n15622), .ZN(n15602) );
  AND2_X1 U9896 ( .A1(n10435), .A2(n10434), .ZN(n15611) );
  INV_X1 U9897 ( .A(n11513), .ZN(n11751) );
  INV_X1 U9898 ( .A(n14725), .ZN(n14667) );
  NAND2_X1 U9899 ( .A1(n15525), .A2(n10647), .ZN(n14718) );
  INV_X1 U9900 ( .A(n14816), .ZN(n12464) );
  INV_X1 U9901 ( .A(n16112), .ZN(n16149) );
  INV_X1 U9902 ( .A(n14461), .ZN(n14734) );
  AND2_X1 U9903 ( .A1(n14807), .A2(n10771), .ZN(n16006) );
  INV_X1 U9904 ( .A(n12421), .ZN(n12427) );
  AND2_X1 U9905 ( .A1(n12008), .A2(n11857), .ZN(n12113) );
  INV_X1 U9906 ( .A(n10771), .ZN(n16041) );
  OR2_X1 U9907 ( .A1(n12451), .A2(n10470), .ZN(n10471) );
  INV_X1 U9908 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9704) );
  AND2_X1 U9909 ( .A1(n9146), .A2(n9116), .ZN(n14428) );
  AND2_X1 U9910 ( .A1(n10449), .A2(n15495), .ZN(n11300) );
  INV_X1 U9911 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10232) );
  INV_X1 U9912 ( .A(n16098), .ZN(n14987) );
  AND2_X1 U9913 ( .A1(n9779), .A2(n9778), .ZN(n14969) );
  OR2_X1 U9914 ( .A1(n10183), .A2(n9938), .ZN(n9940) );
  INV_X1 U9915 ( .A(n15147), .ZN(n15647) );
  NOR2_X1 U9916 ( .A1(n15641), .A2(n10332), .ZN(n15147) );
  INV_X1 U9917 ( .A(n15974), .ZN(n15445) );
  NAND2_X1 U9918 ( .A1(n12649), .A2(n12648), .ZN(n12650) );
  INV_X1 U9919 ( .A(n15377), .ZN(n15990) );
  NAND2_X1 U9920 ( .A1(n11019), .A2(n15495), .ZN(n15377) );
  AND2_X1 U9921 ( .A1(n10213), .A2(n15497), .ZN(n10917) );
  AND2_X1 U9922 ( .A1(n12928), .A2(n16021), .ZN(n15469) );
  INV_X1 U9923 ( .A(n16119), .ZN(n16136) );
  AND2_X1 U9924 ( .A1(n15973), .A2(n15972), .ZN(n15997) );
  INV_X1 U9925 ( .A(n15469), .ZN(n16139) );
  INV_X1 U9926 ( .A(n10917), .ZN(n11016) );
  AND2_X1 U9927 ( .A1(n9945), .A2(n9972), .ZN(n10368) );
  INV_X1 U9928 ( .A(n15512), .ZN(n15503) );
  INV_X1 U9929 ( .A(n14143), .ZN(n10308) );
  AND2_X1 U9930 ( .A1(n10637), .A2(n10636), .ZN(n15521) );
  INV_X1 U9931 ( .A(n8833), .ZN(n8834) );
  INV_X1 U9932 ( .A(n13343), .ZN(n13314) );
  INV_X1 U9933 ( .A(n13754), .ZN(n15856) );
  OR2_X1 U9934 ( .A1(n10638), .A2(n10629), .ZN(n15872) );
  OR2_X1 U9935 ( .A1(n11641), .A2(n11786), .ZN(n14006) );
  AND2_X1 U9936 ( .A1(n13926), .A2(n13925), .ZN(n14061) );
  AND2_X1 U9937 ( .A1(n12254), .A2(n11790), .ZN(n13968) );
  NAND2_X1 U9938 ( .A1(n16061), .A2(n15940), .ZN(n14083) );
  INV_X1 U9939 ( .A(n14124), .ZN(n14142) );
  INV_X2 U9940 ( .A(n16062), .ZN(n16065) );
  AND2_X1 U9941 ( .A1(n10625), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14143) );
  INV_X1 U9942 ( .A(SI_27_), .ZN(n13101) );
  INV_X1 U9943 ( .A(SI_11_), .ZN(n13130) );
  INV_X1 U9944 ( .A(n11342), .ZN(n11498) );
  INV_X1 U9945 ( .A(n14358), .ZN(n14309) );
  NAND2_X1 U9946 ( .A1(n9591), .A2(n9590), .ZN(n14526) );
  NAND2_X1 U9947 ( .A1(n9392), .A2(n9391), .ZN(n14474) );
  AND2_X1 U9948 ( .A1(n11090), .A2(n11089), .ZN(n11557) );
  OR2_X1 U9949 ( .A1(n15530), .A2(P2_U3088), .ZN(n15616) );
  OR2_X1 U9950 ( .A1(n11741), .A2(n12410), .ZN(n14725) );
  AND2_X1 U9951 ( .A1(n12149), .A2(n12148), .ZN(n16044) );
  OR2_X1 U9952 ( .A1(n15891), .A2(n11735), .ZN(n12150) );
  AND2_X1 U9953 ( .A1(n11741), .A2(n14718), .ZN(n14697) );
  INV_X1 U9954 ( .A(n12155), .ZN(n15891) );
  INV_X1 U9955 ( .A(n16156), .ZN(n16155) );
  AND2_X2 U9956 ( .A1(n10945), .A2(n10473), .ZN(n16156) );
  INV_X1 U9957 ( .A(n14766), .ZN(n14831) );
  AND3_X1 U9958 ( .A1(n16115), .A2(n16114), .A3(n16113), .ZN(n16116) );
  INV_X1 U9959 ( .A(n16157), .ZN(n16160) );
  OR2_X1 U9960 ( .A1(n15522), .A2(n15519), .ZN(n15520) );
  INV_X1 U9961 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10420) );
  INV_X1 U9962 ( .A(n10258), .ZN(n14871) );
  NAND2_X1 U9963 ( .A1(n10234), .A2(P1_STATE_REG_SCAN_IN), .ZN(n16098) );
  INV_X1 U9964 ( .A(n15444), .ZN(n15273) );
  INV_X1 U9965 ( .A(n15299), .ZN(n15452) );
  INV_X1 U9966 ( .A(n15020), .ZN(n15026) );
  INV_X1 U9967 ( .A(n12889), .ZN(n15155) );
  INV_X1 U9968 ( .A(n14969), .ZN(n15060) );
  INV_X1 U9969 ( .A(n15143), .ZN(n15649) );
  INV_X1 U9970 ( .A(n15639), .ZN(n15656) );
  NAND2_X1 U9971 ( .A1(n7218), .A2(n11021), .ZN(n15392) );
  INV_X1 U9972 ( .A(n16143), .ZN(n16141) );
  INV_X1 U9973 ( .A(n16147), .ZN(n16144) );
  AND2_X2 U9974 ( .A1(n10918), .A2(n11016), .ZN(n16147) );
  INV_X1 U9975 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15507) );
  INV_X1 U9976 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11323) );
  INV_X1 U9977 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10605) );
  INV_X1 U9978 ( .A(n15503), .ZN(n11951) );
  INV_X1 U9979 ( .A(n14376), .ZN(P2_U3947) );
  AND2_X1 U9980 ( .A1(n10214), .A2(n9863), .ZN(P1_U4016) );
  INV_X1 U9981 ( .A(n8266), .ZN(n8264) );
  NAND2_X1 U9982 ( .A1(n8264), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8265) );
  NAND2_X2 U9983 ( .A1(n8268), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8269) );
  XNOR2_X2 U9984 ( .A(n8269), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8271) );
  NAND2_X1 U9985 ( .A1(n7231), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8275) );
  NAND2_X1 U9986 ( .A1(n8361), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U9987 ( .A1(n8362), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8273) );
  NAND2_X1 U9988 ( .A1(n8438), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U9989 ( .A1(n8276), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8277) );
  MUX2_X1 U9990 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8277), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8279) );
  NAND2_X1 U9991 ( .A1(n8279), .A2(n8278), .ZN(n12197) );
  XNOR2_X1 U9992 ( .A(n12197), .B(P3_B_REG_SCAN_IN), .ZN(n8282) );
  NAND2_X1 U9993 ( .A1(n8278), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8280) );
  MUX2_X1 U9994 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8280), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8281) );
  NAND2_X1 U9995 ( .A1(n8283), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8284) );
  INV_X1 U9996 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U9997 ( .A1(n10309), .A2(n8287), .ZN(n8289) );
  NAND2_X1 U9998 ( .A1(n12401), .A2(n12197), .ZN(n8288) );
  NAND2_X1 U9999 ( .A1(n8607), .A2(n8610), .ZN(n8291) );
  NAND2_X1 U10000 ( .A1(n8295), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8297) );
  INV_X1 U10001 ( .A(n11426), .ZN(n11267) );
  NAND2_X1 U10002 ( .A1(n7270), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8299) );
  XNOR2_X2 U10003 ( .A(n8299), .B(n8298), .ZN(n13743) );
  NAND2_X1 U10004 ( .A1(n13388), .A2(n13755), .ZN(n8300) );
  NAND2_X1 U10005 ( .A1(n8300), .A2(n11426), .ZN(n8301) );
  INV_X1 U10006 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10717) );
  XNOR2_X2 U10007 ( .A(n8304), .B(n8303), .ZN(n8827) );
  NAND2_X2 U10008 ( .A1(n10628), .A2(n8315), .ZN(n8327) );
  INV_X1 U10009 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U10010 ( .A1(n9858), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8309) );
  AND2_X1 U10011 ( .A1(n8328), .A2(n8309), .ZN(n10254) );
  INV_X1 U10012 ( .A(SI_0_), .ZN(n10253) );
  OR2_X1 U10013 ( .A1(n8370), .A2(n10253), .ZN(n8310) );
  OAI211_X1 U10014 ( .C1(n10717), .C2(n10628), .A(n8311), .B(n8310), .ZN(
        n11270) );
  MUX2_X1 U10015 ( .A(n13588), .B(n8790), .S(n12575), .Z(n8312) );
  INV_X1 U10016 ( .A(n8312), .ZN(n11073) );
  INV_X1 U10017 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U10018 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8313) );
  XNOR2_X1 U10019 ( .A(n8329), .B(n8328), .ZN(n8316) );
  INV_X1 U10020 ( .A(SI_1_), .ZN(n8918) );
  MUX2_X1 U10021 ( .A(n8316), .B(n8918), .S(n10252), .Z(n10240) );
  NAND2_X1 U10022 ( .A1(n8438), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8318) );
  XNOR2_X1 U10023 ( .A(n8321), .B(n13586), .ZN(n11072) );
  NAND2_X1 U10024 ( .A1(n11073), .A2(n11072), .ZN(n11071) );
  INV_X1 U10025 ( .A(n13586), .ZN(n11674) );
  NAND2_X1 U10026 ( .A1(n11674), .A2(n8321), .ZN(n8322) );
  NAND2_X1 U10027 ( .A1(n7231), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8326) );
  NAND2_X1 U10028 ( .A1(n8361), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8325) );
  NAND2_X1 U10029 ( .A1(n8438), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U10030 ( .A1(n8362), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8323) );
  AND4_X2 U10031 ( .A1(n8325), .A2(n8326), .A3(n8324), .A4(n8323), .ZN(n11620)
         );
  OR2_X1 U10032 ( .A1(n8370), .A2(SI_2_), .ZN(n8335) );
  INV_X1 U10033 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U10034 ( .A1(n8906), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U10035 ( .A1(n8331), .A2(n8330), .ZN(n8344) );
  NAND2_X1 U10036 ( .A1(n10259), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8345) );
  INV_X1 U10037 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10243) );
  NAND2_X1 U10038 ( .A1(n10243), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8332) );
  AND2_X1 U10039 ( .A1(n8345), .A2(n8332), .ZN(n8343) );
  XNOR2_X1 U10040 ( .A(n8344), .B(n8343), .ZN(n10280) );
  OR2_X1 U10041 ( .A1(n7204), .A2(n10811), .ZN(n8333) );
  XNOR2_X1 U10042 ( .A(n11682), .B(n8711), .ZN(n8336) );
  XNOR2_X1 U10043 ( .A(n11905), .B(n8336), .ZN(n11189) );
  INV_X1 U10044 ( .A(n8336), .ZN(n8337) );
  AND2_X1 U10045 ( .A1(n11905), .A2(n8337), .ZN(n8338) );
  INV_X1 U10046 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10856) );
  NAND2_X1 U10047 ( .A1(n7231), .A2(n10856), .ZN(n8342) );
  NAND2_X1 U10048 ( .A1(n8361), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U10049 ( .A1(n8438), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U10050 ( .A1(n8362), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8339) );
  AND4_X2 U10051 ( .A1(n8341), .A2(n8342), .A3(n8340), .A4(n8339), .ZN(n11673)
         );
  OR2_X1 U10052 ( .A1(n8370), .A2(SI_3_), .ZN(n8355) );
  NAND2_X1 U10053 ( .A1(n8344), .A2(n8343), .ZN(n8346) );
  NAND2_X1 U10054 ( .A1(n8346), .A2(n8345), .ZN(n8349) );
  NAND2_X1 U10055 ( .A1(n8056), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8371) );
  INV_X1 U10056 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10244) );
  NAND2_X1 U10057 ( .A1(n10244), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8347) );
  AND2_X1 U10058 ( .A1(n8371), .A2(n8347), .ZN(n8348) );
  NAND2_X1 U10059 ( .A1(n8349), .A2(n8348), .ZN(n8372) );
  OR2_X1 U10060 ( .A1(n8349), .A2(n8348), .ZN(n8350) );
  NAND2_X1 U10061 ( .A1(n8372), .A2(n8350), .ZN(n10294) );
  OR2_X1 U10062 ( .A1(n8327), .A2(n10294), .ZN(n8354) );
  OR2_X1 U10063 ( .A1(n8351), .A2(n8458), .ZN(n8352) );
  OR2_X1 U10064 ( .A1(n7203), .A2(n10872), .ZN(n8353) );
  XNOR2_X1 U10065 ( .A(n11624), .B(n8711), .ZN(n8356) );
  XNOR2_X1 U10066 ( .A(n11673), .B(n8356), .ZN(n11207) );
  INV_X1 U10067 ( .A(n8356), .ZN(n8357) );
  OR2_X1 U10068 ( .A1(n11673), .A2(n8357), .ZN(n8358) );
  AND2_X1 U10069 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8360) );
  NOR2_X1 U10070 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8390) );
  OR2_X1 U10071 ( .A1(n8360), .A2(n8390), .ZN(n11642) );
  NAND2_X1 U10072 ( .A1(n7231), .A2(n11642), .ZN(n8366) );
  NAND2_X1 U10073 ( .A1(n13365), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8365) );
  BUF_X4 U10074 ( .A(n8362), .Z(n13364) );
  NAND2_X1 U10075 ( .A1(n13364), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8364) );
  NAND2_X1 U10076 ( .A1(n7238), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8363) );
  INV_X1 U10077 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8367) );
  NAND2_X1 U10078 ( .A1(n8351), .A2(n8367), .ZN(n8381) );
  NAND2_X1 U10079 ( .A1(n8381), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8369) );
  INV_X1 U10080 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8368) );
  INV_X1 U10081 ( .A(SI_4_), .ZN(n10292) );
  OR2_X1 U10082 ( .A1(n12960), .A2(n10292), .ZN(n8374) );
  INV_X1 U10083 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10242) );
  XNOR2_X1 U10084 ( .A(n10242), .B(P1_DATAO_REG_4__SCAN_IN), .ZN(n8377) );
  XNOR2_X1 U10085 ( .A(n8378), .B(n8377), .ZN(n10293) );
  OR2_X1 U10086 ( .A1(n8327), .A2(n10293), .ZN(n8373) );
  OAI211_X1 U10087 ( .C1(n10628), .C2(n10974), .A(n8374), .B(n8373), .ZN(
        n11650) );
  XNOR2_X1 U10088 ( .A(n11650), .B(n8790), .ZN(n8375) );
  XNOR2_X1 U10089 ( .A(n11904), .B(n8375), .ZN(n11388) );
  NAND2_X1 U10090 ( .A1(n11904), .A2(n8375), .ZN(n8376) );
  OR2_X1 U10091 ( .A1(n12960), .A2(SI_5_), .ZN(n8389) );
  NAND2_X1 U10092 ( .A1(n10242), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8379) );
  NAND2_X1 U10093 ( .A1(n10251), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8380) );
  XNOR2_X1 U10094 ( .A(n8406), .B(n8405), .ZN(n10286) );
  OR2_X1 U10095 ( .A1(n8327), .A2(n10286), .ZN(n8388) );
  NAND2_X1 U10096 ( .A1(n8383), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8382) );
  MUX2_X1 U10097 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8382), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8386) );
  INV_X1 U10098 ( .A(n8383), .ZN(n8385) );
  INV_X1 U10099 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8384) );
  NAND2_X1 U10100 ( .A1(n8385), .A2(n8384), .ZN(n8409) );
  NAND2_X1 U10101 ( .A1(n8386), .A2(n8409), .ZN(n10977) );
  OR2_X1 U10102 ( .A1(n7203), .A2(n7780), .ZN(n8387) );
  AND3_X2 U10103 ( .A1(n8389), .A2(n8388), .A3(n8387), .ZN(n11955) );
  XNOR2_X1 U10104 ( .A(n11955), .B(n8790), .ZN(n8397) );
  NAND2_X1 U10105 ( .A1(n8390), .A2(n8391), .ZN(n8399) );
  OR2_X1 U10106 ( .A1(n8391), .A2(n8390), .ZN(n8392) );
  NAND2_X1 U10107 ( .A1(n8399), .A2(n8392), .ZN(n11658) );
  NAND2_X1 U10108 ( .A1(n7231), .A2(n11658), .ZN(n8396) );
  NAND2_X1 U10109 ( .A1(n8361), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10110 ( .A1(n8362), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10111 ( .A1(n7237), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8393) );
  NAND4_X1 U10112 ( .A1(n8396), .A2(n8395), .A3(n8394), .A4(n8393), .ZN(n13582) );
  XNOR2_X1 U10113 ( .A(n8397), .B(n13582), .ZN(n11477) );
  INV_X1 U10114 ( .A(n13582), .ZN(n11886) );
  NAND2_X1 U10115 ( .A1(n11886), .A2(n8397), .ZN(n8398) );
  NAND2_X1 U10116 ( .A1(n8399), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U10117 ( .A1(n8427), .A2(n8400), .ZN(n11947) );
  NAND2_X1 U10118 ( .A1(n7231), .A2(n11947), .ZN(n8404) );
  NAND2_X1 U10119 ( .A1(n13365), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U10120 ( .A1(n13364), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10121 ( .A1(n8472), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8401) );
  AND4_X2 U10122 ( .A1(n8404), .A2(n8403), .A3(n8402), .A4(n8401), .ZN(n13412)
         );
  INV_X1 U10123 ( .A(SI_6_), .ZN(n10278) );
  OR2_X1 U10124 ( .A1(n12960), .A2(n10278), .ZN(n8414) );
  NAND2_X1 U10125 ( .A1(n10271), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U10126 ( .A1(n10273), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U10127 ( .A1(n8423), .A2(n8408), .ZN(n8420) );
  XNOR2_X1 U10128 ( .A(n8422), .B(n8420), .ZN(n10279) );
  OR2_X1 U10129 ( .A1(n8327), .A2(n10279), .ZN(n8413) );
  NAND2_X1 U10130 ( .A1(n8409), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8411) );
  INV_X1 U10131 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8410) );
  XNOR2_X1 U10132 ( .A(n8411), .B(n8410), .ZN(n11340) );
  OR2_X1 U10133 ( .A1(n7203), .A2(n11340), .ZN(n8412) );
  XNOR2_X1 U10134 ( .A(n13411), .B(n8711), .ZN(n8415) );
  XNOR2_X1 U10135 ( .A(n13412), .B(n8415), .ZN(n11944) );
  INV_X2 U10136 ( .A(n13412), .ZN(n13581) );
  INV_X1 U10137 ( .A(n8415), .ZN(n8416) );
  NAND2_X1 U10138 ( .A1(n13581), .A2(n8416), .ZN(n8417) );
  OR2_X1 U10139 ( .A1(n8418), .A2(n8458), .ZN(n8419) );
  XNOR2_X1 U10140 ( .A(n8419), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11342) );
  INV_X1 U10141 ( .A(n8420), .ZN(n8421) );
  NAND2_X1 U10142 ( .A1(n8422), .A2(n8421), .ZN(n8424) );
  XNOR2_X1 U10143 ( .A(n8446), .B(n8447), .ZN(n10289) );
  OR2_X1 U10144 ( .A1(n8327), .A2(n10289), .ZN(n8426) );
  OR2_X1 U10145 ( .A1(n12960), .A2(SI_7_), .ZN(n8425) );
  OAI211_X1 U10146 ( .C1(n11342), .C2(n10628), .A(n8426), .B(n8425), .ZN(
        n13420) );
  XNOR2_X1 U10147 ( .A(n13420), .B(n8711), .ZN(n8433) );
  AND2_X1 U10148 ( .A1(n8427), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8428) );
  OR2_X1 U10149 ( .A1(n8428), .A2(n8436), .ZN(n12072) );
  NAND2_X1 U10150 ( .A1(n7231), .A2(n12072), .ZN(n8432) );
  NAND2_X1 U10151 ( .A1(n13365), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U10152 ( .A1(n13364), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8430) );
  NAND2_X1 U10153 ( .A1(n7238), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8429) );
  NAND4_X1 U10154 ( .A1(n8432), .A2(n8431), .A3(n8430), .A4(n8429), .ZN(n13580) );
  XNOR2_X1 U10155 ( .A(n8433), .B(n13580), .ZN(n11814) );
  INV_X1 U10156 ( .A(n8433), .ZN(n8434) );
  NAND2_X1 U10157 ( .A1(n13580), .A2(n8434), .ZN(n8435) );
  NAND2_X1 U10158 ( .A1(n11813), .A2(n8435), .ZN(n12002) );
  NOR2_X1 U10159 ( .A1(n8436), .A2(n13062), .ZN(n8437) );
  OR2_X1 U10160 ( .A1(n8470), .A2(n8437), .ZN(n11999) );
  NAND2_X1 U10161 ( .A1(n7231), .A2(n11999), .ZN(n8442) );
  NAND2_X1 U10162 ( .A1(n13365), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U10163 ( .A1(n13364), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8440) );
  NAND2_X1 U10164 ( .A1(n8472), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8439) );
  INV_X1 U10165 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U10166 ( .A1(n8418), .A2(n8443), .ZN(n8457) );
  NAND2_X1 U10167 ( .A1(n8457), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8445) );
  XNOR2_X1 U10168 ( .A(n8445), .B(n8444), .ZN(n11499) );
  NAND2_X1 U10169 ( .A1(n8449), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8450) );
  NAND2_X1 U10170 ( .A1(n10301), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U10171 ( .A1(n10298), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8451) );
  XNOR2_X1 U10172 ( .A(n8465), .B(n8463), .ZN(n10256) );
  OR2_X1 U10173 ( .A1(n8327), .A2(n10256), .ZN(n8453) );
  INV_X1 U10174 ( .A(SI_8_), .ZN(n10255) );
  OR2_X1 U10175 ( .A1(n12960), .A2(n10255), .ZN(n8452) );
  OAI211_X1 U10176 ( .C1(n7203), .C2(n11499), .A(n8453), .B(n8452), .ZN(n12165) );
  XNOR2_X1 U10177 ( .A(n12165), .B(n8711), .ZN(n8454) );
  XNOR2_X1 U10178 ( .A(n12234), .B(n8454), .ZN(n12001) );
  INV_X1 U10179 ( .A(n8454), .ZN(n8455) );
  OR2_X1 U10180 ( .A1(n12234), .A2(n8455), .ZN(n8456) );
  NOR2_X1 U10181 ( .A1(n8457), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8461) );
  OR2_X1 U10182 ( .A1(n8461), .A2(n8458), .ZN(n8459) );
  MUX2_X1 U10183 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8459), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n8462) );
  NAND2_X1 U10184 ( .A1(n8461), .A2(n8460), .ZN(n8505) );
  NAND2_X1 U10185 ( .A1(n8462), .A2(n8505), .ZN(n12026) );
  INV_X1 U10186 ( .A(n8463), .ZN(n8464) );
  XNOR2_X1 U10187 ( .A(n8489), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n8488) );
  XNOR2_X1 U10188 ( .A(n8487), .B(n8488), .ZN(n10257) );
  OR2_X1 U10189 ( .A1(n8327), .A2(n10257), .ZN(n8468) );
  OR2_X1 U10190 ( .A1(n12960), .A2(n13136), .ZN(n8467) );
  OAI211_X1 U10191 ( .C1(n7204), .C2(n12026), .A(n8468), .B(n8467), .ZN(n12237) );
  XNOR2_X1 U10192 ( .A(n12237), .B(n8711), .ZN(n8478) );
  NAND2_X1 U10193 ( .A1(n8470), .A2(n8469), .ZN(n8481) );
  OR2_X1 U10194 ( .A1(n8470), .A2(n8469), .ZN(n8471) );
  NAND2_X1 U10195 ( .A1(n8481), .A2(n8471), .ZN(n12238) );
  NAND2_X1 U10196 ( .A1(n7231), .A2(n12238), .ZN(n8476) );
  NAND2_X1 U10197 ( .A1(n13365), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10198 ( .A1(n13364), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8474) );
  NAND2_X1 U10199 ( .A1(n7238), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8473) );
  NAND4_X1 U10200 ( .A1(n8476), .A2(n8475), .A3(n8474), .A4(n8473), .ZN(n13578) );
  XNOR2_X1 U10201 ( .A(n8478), .B(n13578), .ZN(n12233) );
  INV_X1 U10202 ( .A(n12233), .ZN(n8477) );
  INV_X1 U10203 ( .A(n13578), .ZN(n12392) );
  INV_X1 U10204 ( .A(n8478), .ZN(n8479) );
  NAND2_X1 U10205 ( .A1(n12392), .A2(n8479), .ZN(n8480) );
  NAND2_X1 U10206 ( .A1(n8481), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U10207 ( .A1(n8499), .A2(n8482), .ZN(n12217) );
  NAND2_X1 U10208 ( .A1(n7231), .A2(n12217), .ZN(n8486) );
  NAND2_X1 U10209 ( .A1(n13365), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8485) );
  NAND2_X1 U10210 ( .A1(n13364), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8484) );
  NAND2_X1 U10211 ( .A1(n8472), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U10212 ( .A1(n8489), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U10213 ( .A1(n10424), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U10214 ( .A1(n10426), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8491) );
  NAND2_X1 U10215 ( .A1(n8509), .A2(n8491), .ZN(n8507) );
  XNOR2_X1 U10216 ( .A(n8508), .B(n8507), .ZN(n10274) );
  OR2_X1 U10217 ( .A1(n8327), .A2(n10274), .ZN(n8496) );
  OR2_X1 U10218 ( .A1(n12960), .A2(SI_10_), .ZN(n8495) );
  NAND2_X1 U10219 ( .A1(n8505), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8493) );
  INV_X1 U10220 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8492) );
  XNOR2_X1 U10221 ( .A(n8493), .B(n8492), .ZN(n15834) );
  INV_X1 U10222 ( .A(n15834), .ZN(n12058) );
  OR2_X1 U10223 ( .A1(n10628), .A2(n12058), .ZN(n8494) );
  XNOR2_X1 U10224 ( .A(n12394), .B(n8711), .ZN(n8497) );
  XNOR2_X1 U10225 ( .A(n12474), .B(n8497), .ZN(n12390) );
  INV_X1 U10226 ( .A(n8497), .ZN(n8498) );
  NAND2_X1 U10227 ( .A1(n8499), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8500) );
  NAND2_X1 U10228 ( .A1(n8522), .A2(n8500), .ZN(n12477) );
  NAND2_X1 U10229 ( .A1(n7231), .A2(n12477), .ZN(n8504) );
  NAND2_X1 U10230 ( .A1(n13365), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8503) );
  NAND2_X1 U10231 ( .A1(n13364), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8502) );
  NAND2_X1 U10232 ( .A1(n7238), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8501) );
  NAND2_X1 U10233 ( .A1(n8528), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8506) );
  XNOR2_X1 U10234 ( .A(n8506), .B(P3_IR_REG_11__SCAN_IN), .ZN(n12036) );
  NAND2_X1 U10235 ( .A1(n10397), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U10236 ( .A1(n10395), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8510) );
  XNOR2_X1 U10237 ( .A(n8532), .B(n8531), .ZN(n10305) );
  OR2_X1 U10238 ( .A1(n10305), .A2(n8327), .ZN(n8512) );
  OR2_X1 U10239 ( .A1(n12960), .A2(SI_11_), .ZN(n8511) );
  OAI211_X1 U10240 ( .C1(n12036), .C2(n7203), .A(n8512), .B(n8511), .ZN(n12507) );
  INV_X1 U10241 ( .A(n12507), .ZN(n8513) );
  AND2_X1 U10242 ( .A1(n13998), .A2(n8513), .ZN(n12519) );
  NOR2_X1 U10243 ( .A1(n12519), .A2(n8790), .ZN(n8517) );
  NAND2_X1 U10244 ( .A1(n8514), .A2(n12507), .ZN(n12518) );
  NAND2_X1 U10245 ( .A1(n8517), .A2(n12518), .ZN(n8516) );
  NAND2_X1 U10246 ( .A1(n13998), .A2(n12507), .ZN(n13443) );
  AND2_X1 U10247 ( .A1(n13443), .A2(n8790), .ZN(n8518) );
  NAND2_X1 U10248 ( .A1(n8514), .A2(n8513), .ZN(n13439) );
  NAND2_X1 U10249 ( .A1(n8518), .A2(n13439), .ZN(n8515) );
  NAND2_X1 U10250 ( .A1(n8516), .A2(n8515), .ZN(n12470) );
  NAND2_X1 U10251 ( .A1(n12471), .A2(n12470), .ZN(n12469) );
  INV_X1 U10252 ( .A(n8517), .ZN(n8520) );
  INV_X1 U10253 ( .A(n8518), .ZN(n8519) );
  NAND2_X1 U10254 ( .A1(n8520), .A2(n8519), .ZN(n8521) );
  NAND2_X1 U10255 ( .A1(n12469), .A2(n8521), .ZN(n12562) );
  AND2_X1 U10256 ( .A1(n8522), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8523) );
  OR2_X1 U10257 ( .A1(n8523), .A2(n8547), .ZN(n14003) );
  NAND2_X1 U10258 ( .A1(n8823), .A2(n14003), .ZN(n8527) );
  NAND2_X1 U10259 ( .A1(n13365), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8526) );
  NAND2_X1 U10260 ( .A1(n13364), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U10261 ( .A1(n7238), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8524) );
  NAND4_X1 U10262 ( .A1(n8527), .A2(n8526), .A3(n8525), .A4(n8524), .ZN(n13576) );
  OAI21_X1 U10263 ( .B1(n8528), .B2(P3_IR_REG_11__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8530) );
  INV_X1 U10264 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8529) );
  XNOR2_X1 U10265 ( .A(n8530), .B(n8529), .ZN(n12051) );
  AOI22_X1 U10266 ( .A1(n8647), .A2(n13019), .B1(n8646), .B2(n12051), .ZN(
        n8535) );
  XNOR2_X1 U10267 ( .A(n10422), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n8536) );
  XNOR2_X1 U10268 ( .A(n8537), .B(n8536), .ZN(n10307) );
  NAND2_X1 U10269 ( .A1(n10307), .A2(n13370), .ZN(n8534) );
  XNOR2_X1 U10270 ( .A(n12564), .B(n8711), .ZN(n12560) );
  NAND2_X1 U10271 ( .A1(n10422), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8538) );
  XNOR2_X1 U10272 ( .A(n7498), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10400) );
  NAND2_X1 U10273 ( .A1(n10400), .A2(n13370), .ZN(n8545) );
  NAND2_X1 U10274 ( .A1(n8540), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8541) );
  MUX2_X1 U10275 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8541), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8543) );
  NAND2_X1 U10276 ( .A1(n8543), .A2(n8542), .ZN(n13608) );
  AOI22_X1 U10277 ( .A1(n8647), .A2(n13121), .B1(n8646), .B2(n13608), .ZN(
        n8544) );
  XNOR2_X1 U10278 ( .A(n14141), .B(n8711), .ZN(n8553) );
  INV_X1 U10279 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U10280 ( .A1(n8547), .A2(n8546), .ZN(n8563) );
  OR2_X1 U10281 ( .A1(n8547), .A2(n8546), .ZN(n8548) );
  NAND2_X1 U10282 ( .A1(n8563), .A2(n8548), .ZN(n13312) );
  NAND2_X1 U10283 ( .A1(n8823), .A2(n13312), .ZN(n8552) );
  NAND2_X1 U10284 ( .A1(n13365), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U10285 ( .A1(n13364), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U10286 ( .A1(n8472), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8549) );
  NAND4_X1 U10287 ( .A1(n8552), .A2(n8551), .A3(n8550), .A4(n8549), .ZN(n13995) );
  INV_X1 U10288 ( .A(n13995), .ZN(n13237) );
  NAND2_X1 U10289 ( .A1(n8553), .A2(n13237), .ZN(n13230) );
  INV_X1 U10290 ( .A(n8553), .ZN(n8554) );
  NAND2_X1 U10291 ( .A1(n8554), .A2(n13995), .ZN(n8555) );
  NAND2_X1 U10292 ( .A1(n13230), .A2(n8555), .ZN(n13307) );
  INV_X1 U10293 ( .A(n13307), .ZN(n8556) );
  NAND2_X1 U10294 ( .A1(n8558), .A2(n10605), .ZN(n8559) );
  XNOR2_X1 U10295 ( .A(n10929), .B(P1_DATAO_REG_14__SCAN_IN), .ZN(n8569) );
  XNOR2_X1 U10296 ( .A(n8570), .B(n8569), .ZN(n10606) );
  NAND2_X1 U10297 ( .A1(n10606), .A2(n13370), .ZN(n8562) );
  NAND2_X1 U10298 ( .A1(n8542), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8560) );
  XNOR2_X1 U10299 ( .A(n8560), .B(P3_IR_REG_14__SCAN_IN), .ZN(n13656) );
  AOI22_X1 U10300 ( .A1(n8647), .A2(SI_14_), .B1(n8646), .B2(n13656), .ZN(
        n8561) );
  NAND2_X1 U10301 ( .A1(n8562), .A2(n8561), .ZN(n13987) );
  XNOR2_X1 U10302 ( .A(n13987), .B(n8790), .ZN(n8583) );
  NAND2_X1 U10303 ( .A1(n8563), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U10304 ( .A1(n8576), .A2(n8564), .ZN(n13982) );
  NAND2_X1 U10305 ( .A1(n8823), .A2(n13982), .ZN(n8568) );
  NAND2_X1 U10306 ( .A1(n13365), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U10307 ( .A1(n13364), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U10308 ( .A1(n8472), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8565) );
  XNOR2_X1 U10309 ( .A(n8583), .B(n13959), .ZN(n13231) );
  NAND2_X1 U10310 ( .A1(n10929), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8571) );
  XNOR2_X1 U10311 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8587) );
  XNOR2_X1 U10312 ( .A(n8588), .B(n8587), .ZN(n10608) );
  NAND2_X1 U10313 ( .A1(n10608), .A2(n13370), .ZN(n8575) );
  NAND2_X1 U10314 ( .A1(n8290), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8573) );
  INV_X1 U10315 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8572) );
  XNOR2_X1 U10316 ( .A(n8573), .B(n8572), .ZN(n13657) );
  AOI22_X1 U10317 ( .A1(n8647), .A2(n13122), .B1(n8646), .B2(n13657), .ZN(
        n8574) );
  XNOR2_X1 U10318 ( .A(n14133), .B(n8790), .ZN(n8585) );
  INV_X1 U10319 ( .A(n8594), .ZN(n8578) );
  NAND2_X1 U10320 ( .A1(n8576), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U10321 ( .A1(n8578), .A2(n8577), .ZN(n13962) );
  NAND2_X1 U10322 ( .A1(n8823), .A2(n13962), .ZN(n8582) );
  NAND2_X1 U10323 ( .A1(n13365), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U10324 ( .A1(n13364), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U10325 ( .A1(n8472), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8579) );
  NAND4_X1 U10326 ( .A1(n8582), .A2(n8581), .A3(n8580), .A4(n8579), .ZN(n13974) );
  INV_X1 U10327 ( .A(n13974), .ZN(n13945) );
  XNOR2_X1 U10328 ( .A(n8585), .B(n13945), .ZN(n13344) );
  NAND2_X1 U10329 ( .A1(n8583), .A2(n13348), .ZN(n13340) );
  AND2_X1 U10330 ( .A1(n13344), .A2(n13340), .ZN(n8584) );
  NAND2_X1 U10331 ( .A1(n8585), .A2(n13974), .ZN(n8586) );
  NAND2_X1 U10332 ( .A1(n11015), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8589) );
  XNOR2_X1 U10333 ( .A(n10925), .B(P1_DATAO_REG_16__SCAN_IN), .ZN(n8602) );
  XNOR2_X1 U10334 ( .A(n8604), .B(n8602), .ZN(n10837) );
  NAND2_X1 U10335 ( .A1(n10837), .A2(n13370), .ZN(n8593) );
  NAND2_X1 U10336 ( .A1(n8591), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8608) );
  XNOR2_X1 U10337 ( .A(n8608), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13688) );
  AOI22_X1 U10338 ( .A1(n8647), .A2(SI_16_), .B1(n8646), .B2(n13688), .ZN(
        n8592) );
  XNOR2_X1 U10339 ( .A(n13468), .B(n8790), .ZN(n8600) );
  NOR2_X1 U10340 ( .A1(n8594), .A2(n12995), .ZN(n8595) );
  OR2_X1 U10341 ( .A1(n8615), .A2(n8595), .ZN(n13947) );
  NAND2_X1 U10342 ( .A1(n8823), .A2(n13947), .ZN(n8599) );
  NAND2_X1 U10343 ( .A1(n13365), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U10344 ( .A1(n13364), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U10345 ( .A1(n7238), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8596) );
  NAND4_X1 U10346 ( .A1(n8599), .A2(n8598), .A3(n8597), .A4(n8596), .ZN(n13958) );
  INV_X1 U10347 ( .A(n13958), .ZN(n13467) );
  NAND2_X1 U10348 ( .A1(n8600), .A2(n13467), .ZN(n13269) );
  INV_X1 U10349 ( .A(n8600), .ZN(n8601) );
  NAND2_X1 U10350 ( .A1(n8601), .A2(n13958), .ZN(n13270) );
  INV_X1 U10351 ( .A(n8602), .ZN(n8603) );
  NAND2_X1 U10352 ( .A1(n10925), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8605) );
  XNOR2_X1 U10353 ( .A(n11038), .B(P1_DATAO_REG_17__SCAN_IN), .ZN(n8624) );
  XNOR2_X1 U10354 ( .A(n8626), .B(n8624), .ZN(n10960) );
  NAND2_X1 U10355 ( .A1(n10960), .A2(n13370), .ZN(n8613) );
  NAND2_X1 U10356 ( .A1(n8608), .A2(n8607), .ZN(n8609) );
  NAND2_X1 U10357 ( .A1(n8609), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8611) );
  XNOR2_X1 U10358 ( .A(n8611), .B(n8610), .ZN(n13710) );
  INV_X1 U10359 ( .A(n13710), .ZN(n13727) );
  AOI22_X1 U10360 ( .A1(n8647), .A2(SI_17_), .B1(n8646), .B2(n13727), .ZN(
        n8612) );
  XNOR2_X1 U10361 ( .A(n14123), .B(n8790), .ZN(n8621) );
  NAND2_X1 U10362 ( .A1(n7238), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U10363 ( .A1(n13365), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8619) );
  INV_X1 U10364 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n13182) );
  OR2_X1 U10365 ( .A1(n8615), .A2(n13182), .ZN(n8616) );
  NAND2_X1 U10366 ( .A1(n8632), .A2(n8616), .ZN(n13927) );
  NAND2_X1 U10367 ( .A1(n8823), .A2(n13927), .ZN(n8618) );
  NAND2_X1 U10368 ( .A1(n13364), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8617) );
  XNOR2_X1 U10369 ( .A(n8621), .B(n13914), .ZN(n13279) );
  NAND2_X1 U10370 ( .A1(n13280), .A2(n13279), .ZN(n13278) );
  INV_X1 U10371 ( .A(n8621), .ZN(n8622) );
  NAND2_X1 U10372 ( .A1(n8622), .A2(n13914), .ZN(n8623) );
  INV_X1 U10373 ( .A(n8624), .ZN(n8625) );
  NAND2_X1 U10374 ( .A1(n11038), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8627) );
  XNOR2_X1 U10375 ( .A(n11323), .B(P1_DATAO_REG_18__SCAN_IN), .ZN(n8641) );
  XNOR2_X1 U10376 ( .A(n8643), .B(n8641), .ZN(n11108) );
  NAND2_X1 U10377 ( .A1(n11108), .A2(n13370), .ZN(n8631) );
  NAND2_X1 U10378 ( .A1(n7364), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8628) );
  MUX2_X1 U10379 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8628), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8629) );
  AND2_X1 U10380 ( .A1(n8629), .A2(n7270), .ZN(n13749) );
  AOI22_X1 U10381 ( .A1(n8647), .A2(SI_18_), .B1(n8646), .B2(n13749), .ZN(
        n8630) );
  XNOR2_X1 U10382 ( .A(n14054), .B(n8790), .ZN(n8638) );
  NAND2_X1 U10383 ( .A1(n8632), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8633) );
  NAND2_X1 U10384 ( .A1(n8650), .A2(n8633), .ZN(n13908) );
  NAND2_X1 U10385 ( .A1(n8823), .A2(n13908), .ZN(n8637) );
  NAND2_X1 U10386 ( .A1(n13365), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U10387 ( .A1(n7238), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U10388 ( .A1(n13364), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8634) );
  XNOR2_X1 U10389 ( .A(n8638), .B(n13924), .ZN(n13324) );
  INV_X1 U10390 ( .A(n8638), .ZN(n8639) );
  NAND2_X1 U10391 ( .A1(n8639), .A2(n13924), .ZN(n8640) );
  INV_X1 U10392 ( .A(n8641), .ZN(n8642) );
  INV_X1 U10393 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11422) );
  INV_X1 U10394 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U10395 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n11422), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n11424), .ZN(n8644) );
  INV_X1 U10396 ( .A(n8644), .ZN(n8645) );
  XNOR2_X1 U10397 ( .A(n8659), .B(n8645), .ZN(n11195) );
  NAND2_X1 U10398 ( .A1(n11195), .A2(n13370), .ZN(n8649) );
  AOI22_X1 U10399 ( .A1(n8647), .A2(SI_19_), .B1(n13755), .B2(n8646), .ZN(
        n8648) );
  NAND2_X1 U10400 ( .A1(n8649), .A2(n8648), .ZN(n14051) );
  XNOR2_X1 U10401 ( .A(n14051), .B(n8790), .ZN(n8656) );
  AND2_X1 U10402 ( .A1(n8650), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8651) );
  OR2_X1 U10403 ( .A1(n8651), .A2(n8666), .ZN(n13901) );
  NAND2_X1 U10404 ( .A1(n8823), .A2(n13901), .ZN(n8655) );
  NAND2_X1 U10405 ( .A1(n13365), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U10406 ( .A1(n13364), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U10407 ( .A1(n8472), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8652) );
  NAND4_X1 U10408 ( .A1(n8655), .A2(n8654), .A3(n8653), .A4(n8652), .ZN(n13915) );
  XNOR2_X1 U10409 ( .A(n8656), .B(n13915), .ZN(n13248) );
  INV_X1 U10410 ( .A(n8656), .ZN(n8657) );
  NOR2_X1 U10411 ( .A1(n11422), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U10412 ( .A1(n11422), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U10413 ( .A1(n8662), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8663) );
  AND2_X1 U10414 ( .A1(n8675), .A2(n8663), .ZN(n11425) );
  NAND2_X1 U10415 ( .A1(n11425), .A2(n13370), .ZN(n8665) );
  OR2_X1 U10416 ( .A1(n12960), .A2(n13114), .ZN(n8664) );
  XNOR2_X1 U10417 ( .A(n14118), .B(n8790), .ZN(n8673) );
  INV_X1 U10418 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n8667) );
  OR2_X1 U10419 ( .A1(n8666), .A2(n8667), .ZN(n8668) );
  NAND2_X1 U10420 ( .A1(n8667), .A2(n8666), .ZN(n8678) );
  NAND2_X1 U10421 ( .A1(n8668), .A2(n8678), .ZN(n13887) );
  NAND2_X1 U10422 ( .A1(n8823), .A2(n13887), .ZN(n8672) );
  NAND2_X1 U10423 ( .A1(n13365), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U10424 ( .A1(n13364), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U10425 ( .A1(n7238), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8669) );
  NAND4_X1 U10426 ( .A1(n8672), .A2(n8671), .A3(n8670), .A4(n8669), .ZN(n13866) );
  INV_X1 U10427 ( .A(n13866), .ZN(n13900) );
  XNOR2_X1 U10428 ( .A(n8673), .B(n13900), .ZN(n13299) );
  NAND2_X1 U10429 ( .A1(n8673), .A2(n13866), .ZN(n8674) );
  NAND2_X1 U10430 ( .A1(n13298), .A2(n8674), .ZN(n13257) );
  INV_X1 U10431 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11376) );
  XNOR2_X1 U10432 ( .A(n11376), .B(P2_DATAO_REG_21__SCAN_IN), .ZN(n8688) );
  XNOR2_X1 U10433 ( .A(n8687), .B(n8688), .ZN(n11550) );
  NAND2_X1 U10434 ( .A1(n11550), .A2(n13370), .ZN(n8677) );
  INV_X1 U10435 ( .A(SI_21_), .ZN(n13112) );
  XNOR2_X1 U10436 ( .A(n12977), .B(n8790), .ZN(n8684) );
  NAND2_X1 U10437 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(n8678), .ZN(n8679) );
  NAND2_X1 U10438 ( .A1(n8679), .A2(n7257), .ZN(n13872) );
  NAND2_X1 U10439 ( .A1(n8823), .A2(n13872), .ZN(n8683) );
  NAND2_X1 U10440 ( .A1(n13365), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U10441 ( .A1(n13364), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U10442 ( .A1(n7238), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8680) );
  NAND4_X1 U10443 ( .A1(n8683), .A2(n8682), .A3(n8681), .A4(n8680), .ZN(n13857) );
  XNOR2_X1 U10444 ( .A(n8684), .B(n13857), .ZN(n13256) );
  NAND2_X1 U10445 ( .A1(n13257), .A2(n13256), .ZN(n13255) );
  INV_X1 U10446 ( .A(n8684), .ZN(n8685) );
  NAND2_X1 U10447 ( .A1(n8685), .A2(n13857), .ZN(n8686) );
  NAND2_X1 U10448 ( .A1(n13255), .A2(n8686), .ZN(n8702) );
  INV_X1 U10449 ( .A(n8688), .ZN(n8689) );
  NAND2_X1 U10450 ( .A1(n11376), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8691) );
  XNOR2_X1 U10451 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .ZN(n8704) );
  XNOR2_X1 U10452 ( .A(n8705), .B(n8704), .ZN(n11580) );
  NAND2_X1 U10453 ( .A1(n11580), .A2(n13370), .ZN(n8694) );
  XNOR2_X1 U10454 ( .A(n14039), .B(n8790), .ZN(n8700) );
  NAND2_X1 U10455 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(n7257), .ZN(n8695) );
  NAND2_X1 U10456 ( .A1(n8695), .A2(n8239), .ZN(n13860) );
  NAND2_X1 U10457 ( .A1(n8823), .A2(n13860), .ZN(n8699) );
  NAND2_X1 U10458 ( .A1(n13365), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8698) );
  NAND2_X1 U10459 ( .A1(n7238), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8697) );
  NAND2_X1 U10460 ( .A1(n13364), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8696) );
  INV_X1 U10461 ( .A(n8700), .ZN(n8701) );
  NOR2_X1 U10462 ( .A1(n8702), .A2(n8701), .ZN(n8703) );
  INV_X1 U10463 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11873) );
  NAND2_X1 U10464 ( .A1(n11873), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8706) );
  XNOR2_X1 U10465 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8724) );
  INV_X1 U10466 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11954) );
  INV_X1 U10467 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12201) );
  OR2_X2 U10468 ( .A1(n8707), .A2(n12201), .ZN(n8734) );
  NAND2_X1 U10469 ( .A1(n8707), .A2(n12201), .ZN(n8708) );
  INV_X1 U10470 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12599) );
  XNOR2_X1 U10471 ( .A(n8733), .B(n12599), .ZN(n12195) );
  NAND2_X1 U10472 ( .A1(n12195), .A2(n13370), .ZN(n8710) );
  INV_X1 U10473 ( .A(SI_24_), .ZN(n13005) );
  OR2_X1 U10474 ( .A1(n12960), .A2(n13005), .ZN(n8709) );
  XNOR2_X1 U10475 ( .A(n14108), .B(n8711), .ZN(n13289) );
  NAND2_X1 U10476 ( .A1(n13364), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8717) );
  INV_X1 U10477 ( .A(n8712), .ZN(n8718) );
  NAND2_X1 U10478 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n8718), .ZN(n8713) );
  INV_X1 U10479 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n13293) );
  NAND2_X1 U10480 ( .A1(n13293), .A2(n8712), .ZN(n8737) );
  NAND2_X1 U10481 ( .A1(n8713), .A2(n8737), .ZN(n13832) );
  NAND2_X1 U10482 ( .A1(n8823), .A2(n13832), .ZN(n8716) );
  NAND2_X1 U10483 ( .A1(n13365), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U10484 ( .A1(n7238), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U10485 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(n8239), .ZN(n8719) );
  NAND2_X1 U10486 ( .A1(n8719), .A2(n8718), .ZN(n13847) );
  NAND2_X1 U10487 ( .A1(n8823), .A2(n13847), .ZN(n8723) );
  NAND2_X1 U10488 ( .A1(n13365), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U10489 ( .A1(n13364), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U10490 ( .A1(n7238), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8720) );
  XNOR2_X1 U10491 ( .A(n8725), .B(n8724), .ZN(n11783) );
  NAND2_X1 U10492 ( .A1(n11783), .A2(n13370), .ZN(n8727) );
  INV_X1 U10493 ( .A(SI_23_), .ZN(n11785) );
  XNOR2_X1 U10494 ( .A(n14035), .B(n8790), .ZN(n8728) );
  OAI22_X1 U10495 ( .A1(n13289), .A2(n13812), .B1(n13826), .B2(n8728), .ZN(
        n8732) );
  NAND3_X1 U10496 ( .A1(n8728), .A2(n13826), .A3(n13812), .ZN(n8731) );
  INV_X1 U10497 ( .A(n8728), .ZN(n13286) );
  OAI21_X1 U10498 ( .B1(n13286), .B2(n12946), .A(n13843), .ZN(n8729) );
  NAND2_X1 U10499 ( .A1(n13289), .A2(n8729), .ZN(n8730) );
  XNOR2_X1 U10500 ( .A(n8113), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8745) );
  XNOR2_X1 U10501 ( .A(n8746), .B(n8745), .ZN(n12346) );
  NAND2_X1 U10502 ( .A1(n12346), .A2(n13370), .ZN(n8736) );
  INV_X1 U10503 ( .A(SI_25_), .ZN(n12348) );
  XNOR2_X1 U10504 ( .A(n14104), .B(n8790), .ZN(n8743) );
  NAND2_X1 U10505 ( .A1(n13364), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U10506 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(n8737), .ZN(n8738) );
  INV_X1 U10507 ( .A(n8750), .ZN(n8749) );
  NAND2_X1 U10508 ( .A1(n8738), .A2(n8749), .ZN(n13818) );
  NAND2_X1 U10509 ( .A1(n8823), .A2(n13818), .ZN(n8741) );
  NAND2_X1 U10510 ( .A1(n13365), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U10511 ( .A1(n8472), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8739) );
  XNOR2_X1 U10512 ( .A(n8743), .B(n13827), .ZN(n13262) );
  INV_X1 U10513 ( .A(n8743), .ZN(n8744) );
  XNOR2_X1 U10514 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n8758) );
  XNOR2_X1 U10515 ( .A(n8759), .B(n8758), .ZN(n12399) );
  NAND2_X1 U10516 ( .A1(n12399), .A2(n13370), .ZN(n8748) );
  INV_X1 U10517 ( .A(SI_26_), .ZN(n13103) );
  XNOR2_X1 U10518 ( .A(n13494), .B(n8790), .ZN(n8756) );
  NAND2_X1 U10519 ( .A1(n13364), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U10520 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(n8749), .ZN(n8751) );
  INV_X1 U10521 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n13334) );
  NAND2_X1 U10522 ( .A1(n13334), .A2(n8750), .ZN(n8768) );
  NAND2_X1 U10523 ( .A1(n8751), .A2(n8768), .ZN(n13804) );
  NAND2_X1 U10524 ( .A1(n8823), .A2(n13804), .ZN(n8754) );
  NAND2_X1 U10525 ( .A1(n13365), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U10526 ( .A1(n8472), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8752) );
  XNOR2_X1 U10527 ( .A(n8756), .B(n13813), .ZN(n13331) );
  INV_X1 U10528 ( .A(n8756), .ZN(n8757) );
  NAND2_X1 U10529 ( .A1(n8759), .A2(n8758), .ZN(n8761) );
  INV_X1 U10530 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12452) );
  NAND2_X1 U10531 ( .A1(n12452), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8760) );
  INV_X1 U10532 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15511) );
  NAND2_X1 U10533 ( .A1(n15511), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8777) );
  INV_X1 U10534 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14870) );
  NAND2_X1 U10535 ( .A1(n14870), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U10536 ( .A1(n8777), .A2(n8762), .ZN(n8763) );
  OR2_X2 U10537 ( .A1(n8764), .A2(n8763), .ZN(n8778) );
  NAND2_X1 U10538 ( .A1(n8764), .A2(n8763), .ZN(n8765) );
  NAND2_X1 U10539 ( .A1(n8778), .A2(n8765), .ZN(n12468) );
  XNOR2_X1 U10540 ( .A(n14096), .B(n8790), .ZN(n8775) );
  NAND2_X1 U10541 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(n8768), .ZN(n8770) );
  INV_X1 U10542 ( .A(n8768), .ZN(n8769) );
  INV_X1 U10543 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n13052) );
  NAND2_X1 U10544 ( .A1(n8769), .A2(n13052), .ZN(n8784) );
  NAND2_X1 U10545 ( .A1(n8770), .A2(n8784), .ZN(n13792) );
  NAND2_X1 U10546 ( .A1(n8823), .A2(n13792), .ZN(n8774) );
  NAND2_X1 U10547 ( .A1(n13365), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U10548 ( .A1(n13364), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U10549 ( .A1(n8472), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8771) );
  NAND4_X1 U10550 ( .A1(n8774), .A2(n8773), .A3(n8772), .A4(n8771), .ZN(n13574) );
  XNOR2_X1 U10551 ( .A(n8775), .B(n12951), .ZN(n13222) );
  INV_X1 U10552 ( .A(n8775), .ZN(n8776) );
  INV_X1 U10553 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14865) );
  XNOR2_X1 U10554 ( .A(n14865), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8779) );
  NAND2_X1 U10555 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  NAND2_X1 U10556 ( .A1(n12954), .A2(n8781), .ZN(n14154) );
  NAND2_X1 U10557 ( .A1(n14154), .A2(n13370), .ZN(n8783) );
  INV_X1 U10558 ( .A(SI_28_), .ZN(n14156) );
  AND2_X1 U10559 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(n8784), .ZN(n8785) );
  NAND2_X1 U10560 ( .A1(n8823), .A2(n13776), .ZN(n8789) );
  NAND2_X1 U10561 ( .A1(n13365), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8788) );
  NAND2_X1 U10562 ( .A1(n13364), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U10563 ( .A1(n7238), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8786) );
  NAND2_X1 U10564 ( .A1(n14091), .A2(n13787), .ZN(n13506) );
  INV_X1 U10565 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U10566 ( .A1(n10309), .A2(n10303), .ZN(n8792) );
  NAND2_X1 U10567 ( .A1(n12401), .A2(n12349), .ZN(n8791) );
  NOR2_X1 U10568 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n8796) );
  NOR4_X1 U10569 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n8795) );
  NOR4_X1 U10570 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8794) );
  NOR4_X1 U10571 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8793) );
  NAND4_X1 U10572 ( .A1(n8796), .A2(n8795), .A3(n8794), .A4(n8793), .ZN(n8802)
         );
  NOR4_X1 U10573 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8800) );
  NOR4_X1 U10574 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8799) );
  NOR4_X1 U10575 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n8798) );
  NOR4_X1 U10576 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n8797) );
  NAND4_X1 U10577 ( .A1(n8800), .A2(n8799), .A3(n8798), .A4(n8797), .ZN(n8801)
         );
  OAI21_X1 U10578 ( .B1(n8802), .B2(n8801), .A(n10309), .ZN(n11175) );
  NAND3_X1 U10579 ( .A1(n11184), .A2(n11174), .A3(n11175), .ZN(n11121) );
  INV_X1 U10580 ( .A(n12401), .ZN(n8804) );
  NOR2_X1 U10581 ( .A1(n12349), .A2(n12197), .ZN(n8803) );
  NAND2_X1 U10582 ( .A1(n7374), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U10583 ( .A1(n8807), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U10584 ( .A1(n13755), .A2(n13565), .ZN(n11269) );
  NOR2_X1 U10585 ( .A1(n13549), .A2(n11269), .ZN(n8815) );
  NAND2_X1 U10586 ( .A1(n11176), .A2(n8815), .ZN(n11122) );
  OR2_X1 U10587 ( .A1(n11121), .A2(n11122), .ZN(n8813) );
  AND3_X1 U10588 ( .A1(n7567), .A2(n11635), .A3(n11175), .ZN(n11124) );
  NAND2_X1 U10589 ( .A1(n13388), .A2(n11426), .ZN(n11181) );
  XNOR2_X1 U10590 ( .A(n11181), .B(n13565), .ZN(n8810) );
  NAND2_X1 U10591 ( .A1(n13388), .A2(n13743), .ZN(n8809) );
  NAND2_X1 U10592 ( .A1(n8810), .A2(n8809), .ZN(n11258) );
  INV_X1 U10593 ( .A(n13565), .ZN(n11259) );
  AND3_X1 U10594 ( .A1(n11176), .A2(n11258), .A3(n16054), .ZN(n8811) );
  NAND2_X1 U10595 ( .A1(n11124), .A2(n8811), .ZN(n8812) );
  INV_X1 U10596 ( .A(n13550), .ZN(n11683) );
  OR2_X1 U10597 ( .A1(n11124), .A2(n11683), .ZN(n8814) );
  NAND2_X1 U10598 ( .A1(n8814), .A2(n11639), .ZN(n13354) );
  INV_X1 U10599 ( .A(n11258), .ZN(n8818) );
  NAND2_X1 U10600 ( .A1(n11121), .A2(n8815), .ZN(n8817) );
  INV_X1 U10601 ( .A(n13388), .ZN(n11268) );
  NAND2_X1 U10602 ( .A1(n11426), .A2(n13743), .ZN(n11179) );
  INV_X1 U10603 ( .A(n11179), .ZN(n13563) );
  OR2_X1 U10604 ( .A1(n13474), .A2(n13563), .ZN(n11180) );
  AND3_X1 U10605 ( .A1(n9751), .A2(n10625), .A3(n11180), .ZN(n8816) );
  OAI211_X1 U10606 ( .C1(n11124), .C2(n8818), .A(n8817), .B(n8816), .ZN(n8819)
         );
  NAND2_X1 U10607 ( .A1(n8819), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8822) );
  NOR2_X1 U10608 ( .A1(n13474), .A2(n11179), .ZN(n11117) );
  NAND2_X1 U10609 ( .A1(n11176), .A2(n11117), .ZN(n13564) );
  INV_X1 U10610 ( .A(n13564), .ZN(n8820) );
  NAND2_X1 U10611 ( .A1(n11121), .A2(n8820), .ZN(n8821) );
  NAND2_X1 U10612 ( .A1(n8822), .A2(n8821), .ZN(n13351) );
  NAND2_X1 U10613 ( .A1(n8823), .A2(n13757), .ZN(n13369) );
  NAND2_X1 U10614 ( .A1(n13365), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8826) );
  NAND2_X1 U10615 ( .A1(n8472), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8825) );
  NAND2_X1 U10616 ( .A1(n13364), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8824) );
  NAND4_X1 U10617 ( .A1(n13369), .A2(n8826), .A3(n8825), .A4(n8824), .ZN(
        n13572) );
  INV_X1 U10618 ( .A(n13572), .ZN(n13767) );
  OR2_X1 U10619 ( .A1(n11121), .A2(n13564), .ZN(n8829) );
  INV_X1 U10620 ( .A(n8829), .ZN(n8828) );
  INV_X1 U10621 ( .A(n8827), .ZN(n12963) );
  NAND2_X1 U10622 ( .A1(n12963), .A2(n13603), .ZN(n10629) );
  NAND2_X1 U10623 ( .A1(n10628), .A2(n10629), .ZN(n11265) );
  NAND2_X1 U10624 ( .A1(n8828), .A2(n11265), .ZN(n13335) );
  NOR2_X1 U10625 ( .A1(n8829), .A2(n11265), .ZN(n13318) );
  AOI22_X1 U10626 ( .A1(n13318), .A2(n13574), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n8830) );
  OAI21_X1 U10627 ( .B1(n13767), .B2(n13335), .A(n8830), .ZN(n8831) );
  AOI21_X1 U10628 ( .B1(n13776), .B2(n13351), .A(n8831), .ZN(n8832) );
  NAND2_X1 U10629 ( .A1(n8835), .A2(n8834), .ZN(P3_U3160) );
  NAND4_X1 U10630 ( .A1(n8839), .A2(n8838), .A3(n8837), .A4(n9197), .ZN(n8840)
         );
  NOR2_X1 U10631 ( .A1(n8959), .A2(n8840), .ZN(n8844) );
  NOR2_X1 U10632 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n8843) );
  NOR2_X1 U10633 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8842) );
  NOR2_X1 U10634 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), 
        .ZN(n8841) );
  INV_X1 U10635 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8861) );
  NAND2_X2 U10636 ( .A1(n8851), .A2(n9696), .ZN(n8886) );
  NAND2_X1 U10637 ( .A1(n8862), .A2(n8854), .ZN(n8857) );
  NAND2_X1 U10638 ( .A1(n8858), .A2(n8853), .ZN(n8859) );
  NOR2_X1 U10639 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n8864) );
  NOR2_X1 U10640 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n8863) );
  AND2_X1 U10641 ( .A1(n8864), .A2(n8863), .ZN(n8866) );
  NOR2_X1 U10642 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8865) );
  NAND4_X1 U10643 ( .A1(n8866), .A2(n7250), .A3(n7343), .A4(n8865), .ZN(n8867)
         );
  INV_X1 U10644 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10438) );
  INV_X1 U10645 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10443) );
  INV_X1 U10646 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10439) );
  INV_X1 U10647 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10440) );
  NAND2_X1 U10648 ( .A1(n10252), .A2(SI_0_), .ZN(n8877) );
  XNOR2_X1 U10649 ( .A(n8877), .B(n8876), .ZN(n14872) );
  INV_X1 U10650 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8878) );
  INV_X1 U10651 ( .A(n8881), .ZN(n8882) );
  NAND2_X1 U10652 ( .A1(n9645), .A2(n9077), .ZN(n8892) );
  NAND3_X1 U10653 ( .A1(n8891), .A2(n8892), .A3(n8245), .ZN(n8890) );
  NAND2_X1 U10654 ( .A1(n8886), .A2(n12410), .ZN(n8888) );
  NAND2_X1 U10655 ( .A1(n8888), .A2(n11734), .ZN(n8889) );
  NAND2_X1 U10656 ( .A1(n8890), .A2(n8889), .ZN(n8896) );
  INV_X1 U10657 ( .A(n8891), .ZN(n8894) );
  INV_X1 U10658 ( .A(n8892), .ZN(n8893) );
  NAND2_X1 U10659 ( .A1(n8894), .A2(n8893), .ZN(n8895) );
  INV_X1 U10660 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11880) );
  INV_X1 U10661 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8897) );
  INV_X1 U10662 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11876) );
  OR2_X1 U10663 ( .A1(n9334), .A2(n11876), .ZN(n8899) );
  NAND2_X1 U10664 ( .A1(n8942), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8898) );
  NAND2_X1 U10665 ( .A1(n14377), .A2(n7206), .ZN(n8910) );
  XNOR2_X1 U10666 ( .A(n8923), .B(SI_1_), .ZN(n8954) );
  XNOR2_X1 U10667 ( .A(n7216), .B(n8954), .ZN(n10246) );
  NAND2_X1 U10668 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8902) );
  MUX2_X1 U10669 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8902), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8904) );
  INV_X1 U10670 ( .A(n8903), .ZN(n8927) );
  NAND2_X1 U10671 ( .A1(n8904), .A2(n8927), .ZN(n10520) );
  OR2_X1 U10672 ( .A1(n8917), .A2(n8906), .ZN(n8907) );
  NAND2_X1 U10673 ( .A1(n8885), .A2(n11879), .ZN(n8909) );
  NAND2_X1 U10674 ( .A1(n8910), .A2(n8909), .ZN(n8935) );
  NAND2_X1 U10675 ( .A1(n8942), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8916) );
  INV_X1 U10676 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8911) );
  INV_X1 U10677 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8912) );
  OR2_X1 U10678 ( .A1(n9334), .A2(n8912), .ZN(n8914) );
  INV_X1 U10679 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10523) );
  OR2_X1 U10680 ( .A1(n7208), .A2(n10523), .ZN(n8913) );
  NAND4_X2 U10681 ( .A1(n8916), .A2(n8915), .A3(n8914), .A4(n8913), .ZN(n14375) );
  NAND2_X1 U10682 ( .A1(n8923), .A2(SI_1_), .ZN(n8952) );
  OAI21_X1 U10683 ( .B1(SI_2_), .B2(n8918), .A(n8923), .ZN(n8921) );
  INV_X1 U10684 ( .A(SI_2_), .ZN(n10282) );
  OAI21_X1 U10685 ( .B1(SI_1_), .B2(n10282), .A(n8919), .ZN(n8920) );
  NAND2_X1 U10686 ( .A1(n8921), .A2(n8920), .ZN(n8925) );
  INV_X1 U10687 ( .A(n7216), .ZN(n8922) );
  OAI211_X1 U10688 ( .C1(n8923), .C2(SI_1_), .A(n8922), .B(n10282), .ZN(n8924)
         );
  MUX2_X1 U10689 ( .A(n10243), .B(n10259), .S(n8926), .Z(n8949) );
  OR2_X1 U10690 ( .A1(n9599), .A2(n7254), .ZN(n8931) );
  NAND2_X1 U10691 ( .A1(n8927), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8928) );
  MUX2_X1 U10692 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8928), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n8929) );
  NAND2_X1 U10693 ( .A1(n8929), .A2(n8959), .ZN(n15544) );
  OR2_X1 U10694 ( .A1(n10428), .A2(n15544), .ZN(n8930) );
  NAND2_X1 U10695 ( .A1(n14375), .A2(n9077), .ZN(n8933) );
  NAND2_X1 U10696 ( .A1(n8885), .A2(n10587), .ZN(n8932) );
  NAND2_X1 U10697 ( .A1(n8933), .A2(n8932), .ZN(n8937) );
  OAI22_X1 U10698 ( .A1(n8936), .A2(n8935), .B1(n8938), .B2(n8937), .ZN(n8941)
         );
  INV_X1 U10699 ( .A(n9077), .ZN(n9636) );
  AOI22_X1 U10700 ( .A1(n14377), .A2(n9636), .B1(n9077), .B2(n11879), .ZN(
        n8934) );
  AOI21_X1 U10701 ( .B1(n8936), .B2(n8935), .A(n8934), .ZN(n8940) );
  NAND2_X1 U10702 ( .A1(n8938), .A2(n8937), .ZN(n8939) );
  NAND2_X1 U10703 ( .A1(n9547), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8948) );
  INV_X1 U10704 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8944) );
  OR2_X1 U10705 ( .A1(n9608), .A2(n8944), .ZN(n8947) );
  OR2_X1 U10706 ( .A1(n9624), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8946) );
  INV_X1 U10708 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10525) );
  OR2_X1 U10709 ( .A1(n7209), .A2(n10525), .ZN(n8945) );
  NAND2_X1 U10710 ( .A1(n14374), .A2(n7206), .ZN(n8963) );
  INV_X1 U10711 ( .A(n8949), .ZN(n8950) );
  NAND2_X1 U10712 ( .A1(n8951), .A2(n8950), .ZN(n8957) );
  NAND2_X1 U10713 ( .A1(n8955), .A2(SI_2_), .ZN(n8956) );
  XNOR2_X1 U10714 ( .A(n8969), .B(n8967), .ZN(n9901) );
  NAND2_X1 U10715 ( .A1(n9901), .A2(n9620), .ZN(n8961) );
  NAND2_X1 U10716 ( .A1(n8959), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8958) );
  MUX2_X1 U10717 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8958), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8960) );
  AND2_X1 U10718 ( .A1(n8960), .A2(n8973), .ZN(n14387) );
  NAND2_X1 U10719 ( .A1(n12099), .A2(n9615), .ZN(n8962) );
  NAND2_X1 U10720 ( .A1(n8963), .A2(n8962), .ZN(n8965) );
  AOI22_X1 U10721 ( .A1(n9615), .A2(n14374), .B1(n12099), .B2(n9077), .ZN(
        n8964) );
  NAND2_X1 U10722 ( .A1(n8970), .A2(SI_3_), .ZN(n8971) );
  MUX2_X1 U10723 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7215), .Z(n8989) );
  XNOR2_X1 U10724 ( .A(n8989), .B(SI_4_), .ZN(n8986) );
  XNOR2_X1 U10725 ( .A(n8988), .B(n8986), .ZN(n10241) );
  NAND2_X1 U10726 ( .A1(n10241), .A2(n9620), .ZN(n8976) );
  NAND2_X1 U10727 ( .A1(n8973), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8972) );
  MUX2_X1 U10728 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8972), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8974) );
  INV_X1 U10729 ( .A(n9194), .ZN(n8992) );
  NAND2_X1 U10730 ( .A1(n8974), .A2(n8992), .ZN(n10529) );
  INV_X1 U10731 ( .A(n10529), .ZN(n15553) );
  AOI22_X1 U10732 ( .A1(n9354), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9353), .B2(
        n15553), .ZN(n8975) );
  NAND2_X1 U10733 ( .A1(n11738), .A2(n9077), .ZN(n8983) );
  NAND2_X1 U10734 ( .A1(n8942), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8981) );
  INV_X1 U10735 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8977) );
  OR2_X1 U10736 ( .A1(n9608), .A2(n8977), .ZN(n8980) );
  NAND2_X1 U10737 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8999) );
  OAI21_X1 U10738 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8999), .ZN(n11739) );
  OR2_X1 U10739 ( .A1(n9624), .A2(n11739), .ZN(n8979) );
  INV_X1 U10740 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10530) );
  OR2_X1 U10741 ( .A1(n7208), .A2(n10530), .ZN(n8978) );
  NAND2_X1 U10742 ( .A1(n14373), .A2(n9636), .ZN(n8982) );
  INV_X1 U10743 ( .A(n14373), .ZN(n10830) );
  NAND2_X1 U10744 ( .A1(n11738), .A2(n9615), .ZN(n8984) );
  INV_X1 U10745 ( .A(n8986), .ZN(n8987) );
  NAND2_X1 U10746 ( .A1(n8988), .A2(n8987), .ZN(n8991) );
  NAND2_X1 U10747 ( .A1(n8989), .A2(SI_4_), .ZN(n8990) );
  MUX2_X1 U10748 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10252), .Z(n9014) );
  XNOR2_X1 U10749 ( .A(n9014), .B(SI_5_), .ZN(n9011) );
  XNOR2_X1 U10750 ( .A(n9013), .B(n9011), .ZN(n10250) );
  NAND2_X1 U10751 ( .A1(n10250), .A2(n9620), .ZN(n8995) );
  NAND2_X1 U10752 ( .A1(n8992), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8993) );
  XNOR2_X1 U10753 ( .A(n8993), .B(P2_IR_REG_5__SCAN_IN), .ZN(n15565) );
  AOI22_X1 U10754 ( .A1(n9354), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9353), .B2(
        n15565), .ZN(n8994) );
  NAND2_X1 U10755 ( .A1(n8995), .A2(n8994), .ZN(n14269) );
  NAND2_X1 U10756 ( .A1(n14269), .A2(n9615), .ZN(n9006) );
  NAND2_X1 U10757 ( .A1(n9547), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9004) );
  INV_X1 U10758 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8996) );
  OR2_X1 U10759 ( .A1(n9608), .A2(n8996), .ZN(n9003) );
  INV_X1 U10760 ( .A(n8999), .ZN(n8997) );
  NAND2_X1 U10761 ( .A1(n8997), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9025) );
  INV_X1 U10762 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U10763 ( .A1(n8999), .A2(n8998), .ZN(n9000) );
  NAND2_X1 U10764 ( .A1(n9025), .A2(n9000), .ZN(n14270) );
  OR2_X1 U10765 ( .A1(n9624), .A2(n14270), .ZN(n9002) );
  INV_X1 U10766 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11767) );
  OR2_X1 U10767 ( .A1(n7209), .A2(n11767), .ZN(n9001) );
  NAND4_X1 U10768 ( .A1(n9004), .A2(n9003), .A3(n9002), .A4(n9001), .ZN(n14372) );
  NAND2_X1 U10769 ( .A1(n14372), .A2(n9634), .ZN(n9005) );
  NAND2_X1 U10770 ( .A1(n9006), .A2(n9005), .ZN(n9008) );
  AOI22_X1 U10771 ( .A1(n14269), .A2(n9634), .B1(n9615), .B2(n14372), .ZN(
        n9007) );
  INV_X1 U10772 ( .A(n9011), .ZN(n9012) );
  NAND2_X1 U10773 ( .A1(n9013), .A2(n9012), .ZN(n9016) );
  NAND2_X1 U10774 ( .A1(n9014), .A2(SI_5_), .ZN(n9015) );
  NAND2_X1 U10775 ( .A1(n10269), .A2(n9620), .ZN(n9021) );
  INV_X1 U10776 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9017) );
  INV_X1 U10777 ( .A(n9041), .ZN(n9018) );
  NAND2_X1 U10778 ( .A1(n9018), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9019) );
  XNOR2_X1 U10779 ( .A(n9019), .B(P2_IR_REG_6__SCAN_IN), .ZN(n15577) );
  AOI22_X1 U10780 ( .A1(n9354), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9353), .B2(
        n15577), .ZN(n9020) );
  NAND2_X1 U10781 ( .A1(n11400), .A2(n9634), .ZN(n9032) );
  NAND2_X1 U10782 ( .A1(n9547), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9030) );
  INV_X1 U10783 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9022) );
  OR2_X1 U10784 ( .A1(n9608), .A2(n9022), .ZN(n9029) );
  INV_X1 U10785 ( .A(n9025), .ZN(n9023) );
  NAND2_X1 U10786 ( .A1(n9023), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9048) );
  INV_X1 U10787 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U10788 ( .A1(n9025), .A2(n9024), .ZN(n9026) );
  NAND2_X1 U10789 ( .A1(n9048), .A2(n9026), .ZN(n11776) );
  OR2_X1 U10790 ( .A1(n9624), .A2(n11776), .ZN(n9028) );
  INV_X1 U10791 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11775) );
  OR2_X1 U10792 ( .A1(n7209), .A2(n11775), .ZN(n9027) );
  NAND4_X1 U10793 ( .A1(n9030), .A2(n9029), .A3(n9028), .A4(n9027), .ZN(n14371) );
  NAND2_X1 U10794 ( .A1(n14371), .A2(n9615), .ZN(n9031) );
  INV_X1 U10795 ( .A(n14371), .ZN(n11396) );
  NAND2_X1 U10796 ( .A1(n11400), .A2(n9615), .ZN(n9033) );
  OAI21_X1 U10797 ( .B1(n11396), .B2(n9615), .A(n9033), .ZN(n9034) );
  NAND2_X1 U10798 ( .A1(n9038), .A2(SI_6_), .ZN(n9039) );
  MUX2_X1 U10799 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10252), .Z(n9063) );
  XNOR2_X1 U10800 ( .A(n9063), .B(SI_7_), .ZN(n9060) );
  XNOR2_X1 U10801 ( .A(n9062), .B(n9060), .ZN(n10276) );
  NAND2_X1 U10802 ( .A1(n10276), .A2(n9620), .ZN(n9044) );
  INV_X1 U10803 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9040) );
  NAND2_X1 U10804 ( .A1(n9041), .A2(n9040), .ZN(n9064) );
  NAND2_X1 U10805 ( .A1(n9064), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9042) );
  XNOR2_X1 U10806 ( .A(n9042), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14400) );
  AOI22_X1 U10807 ( .A1(n9354), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9353), .B2(
        n14400), .ZN(n9043) );
  NAND2_X1 U10808 ( .A1(n11510), .A2(n9615), .ZN(n9055) );
  NAND2_X1 U10809 ( .A1(n9547), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9053) );
  INV_X1 U10810 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9045) );
  OR2_X1 U10811 ( .A1(n9608), .A2(n9045), .ZN(n9052) );
  INV_X1 U10812 ( .A(n9048), .ZN(n9046) );
  NAND2_X1 U10813 ( .A1(n9046), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9069) );
  INV_X1 U10814 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U10815 ( .A1(n9048), .A2(n9047), .ZN(n9049) );
  NAND2_X1 U10816 ( .A1(n9069), .A2(n9049), .ZN(n11806) );
  OR2_X1 U10817 ( .A1(n9624), .A2(n11806), .ZN(n9051) );
  INV_X1 U10818 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11805) );
  OR2_X1 U10819 ( .A1(n7208), .A2(n11805), .ZN(n9050) );
  NAND4_X1 U10820 ( .A1(n9053), .A2(n9052), .A3(n9051), .A4(n9050), .ZN(n14370) );
  NAND2_X1 U10821 ( .A1(n14370), .A2(n9634), .ZN(n9054) );
  NAND2_X1 U10822 ( .A1(n9055), .A2(n9054), .ZN(n9057) );
  AOI22_X1 U10823 ( .A1(n11510), .A2(n9634), .B1(n9615), .B2(n14370), .ZN(
        n9056) );
  INV_X1 U10824 ( .A(n9060), .ZN(n9061) );
  MUX2_X1 U10825 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10252), .Z(n9088) );
  XNOR2_X1 U10826 ( .A(n9088), .B(SI_8_), .ZN(n9085) );
  XNOR2_X1 U10827 ( .A(n9087), .B(n9085), .ZN(n10297) );
  NAND2_X1 U10828 ( .A1(n10297), .A2(n9620), .ZN(n9066) );
  NAND2_X1 U10829 ( .A1(n9177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9092) );
  XNOR2_X1 U10830 ( .A(n9092), .B(P2_IR_REG_8__SCAN_IN), .ZN(n14415) );
  AOI22_X1 U10831 ( .A1(n9354), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n14415), 
        .B2(n9353), .ZN(n9065) );
  NAND2_X1 U10832 ( .A1(n16003), .A2(n9634), .ZN(n9076) );
  NAND2_X1 U10833 ( .A1(n9547), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9074) );
  INV_X1 U10834 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9067) );
  OR2_X1 U10835 ( .A1(n9608), .A2(n9067), .ZN(n9073) );
  NAND2_X1 U10836 ( .A1(n9069), .A2(n9068), .ZN(n9070) );
  NAND2_X1 U10837 ( .A1(n9098), .A2(n9070), .ZN(n11761) );
  OR2_X1 U10838 ( .A1(n9624), .A2(n11761), .ZN(n9072) );
  INV_X1 U10839 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11756) );
  OR2_X1 U10840 ( .A1(n7208), .A2(n11756), .ZN(n9071) );
  NAND4_X1 U10841 ( .A1(n9074), .A2(n9073), .A3(n9072), .A4(n9071), .ZN(n14369) );
  NAND2_X1 U10842 ( .A1(n14369), .A2(n9615), .ZN(n9075) );
  NAND2_X1 U10843 ( .A1(n9076), .A2(n9075), .ZN(n9081) );
  NAND2_X1 U10844 ( .A1(n9082), .A2(n9081), .ZN(n9080) );
  INV_X1 U10845 ( .A(n14369), .ZN(n11514) );
  NAND2_X1 U10846 ( .A1(n16003), .A2(n9615), .ZN(n9078) );
  OAI21_X1 U10847 ( .B1(n11514), .B2(n9615), .A(n9078), .ZN(n9079) );
  NAND2_X1 U10848 ( .A1(n9080), .A2(n9079), .ZN(n9084) );
  INV_X1 U10849 ( .A(n9085), .ZN(n9086) );
  NAND2_X1 U10850 ( .A1(n9088), .A2(SI_8_), .ZN(n9089) );
  NAND2_X2 U10851 ( .A1(n9090), .A2(n9089), .ZN(n9135) );
  MUX2_X1 U10852 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10252), .Z(n9136) );
  INV_X1 U10853 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U10854 ( .A1(n9092), .A2(n9091), .ZN(n9093) );
  NAND2_X1 U10855 ( .A1(n9093), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9113) );
  XNOR2_X1 U10856 ( .A(n9113), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U10857 ( .A1(n10576), .A2(n9353), .B1(n9354), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U10858 ( .A1(n11795), .A2(n9615), .ZN(n9105) );
  NAND2_X1 U10859 ( .A1(n9626), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9103) );
  INV_X1 U10860 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9096) );
  OR2_X1 U10861 ( .A1(n7494), .A2(n9096), .ZN(n9102) );
  INV_X1 U10862 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11369) );
  NAND2_X1 U10863 ( .A1(n9098), .A2(n11369), .ZN(n9099) );
  NAND2_X1 U10864 ( .A1(n9121), .A2(n9099), .ZN(n11366) );
  OR2_X1 U10865 ( .A1(n9624), .A2(n11366), .ZN(n9101) );
  INV_X1 U10866 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10519) );
  OR2_X1 U10867 ( .A1(n7209), .A2(n10519), .ZN(n9100) );
  NAND4_X1 U10868 ( .A1(n9103), .A2(n9102), .A3(n9101), .A4(n9100), .ZN(n14368) );
  NAND2_X1 U10869 ( .A1(n14368), .A2(n9634), .ZN(n9104) );
  NAND2_X1 U10870 ( .A1(n9105), .A2(n9104), .ZN(n9107) );
  AOI22_X1 U10871 ( .A1(n11795), .A2(n9634), .B1(n9615), .B2(n14368), .ZN(
        n9106) );
  INV_X1 U10872 ( .A(n9110), .ZN(n9111) );
  MUX2_X1 U10873 ( .A(n10426), .B(n10424), .S(n10252), .Z(n9138) );
  NAND2_X1 U10874 ( .A1(n10423), .A2(n9620), .ZN(n9118) );
  INV_X1 U10875 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U10876 ( .A1(n9113), .A2(n9112), .ZN(n9114) );
  NAND2_X1 U10877 ( .A1(n9114), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9115) );
  INV_X1 U10878 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9173) );
  NAND2_X1 U10879 ( .A1(n9115), .A2(n9173), .ZN(n9146) );
  OR2_X1 U10880 ( .A1(n9115), .A2(n9173), .ZN(n9116) );
  AOI22_X1 U10881 ( .A1(n14428), .A2(n9353), .B1(P1_DATAO_REG_10__SCAN_IN), 
        .B2(n9354), .ZN(n9117) );
  NAND2_X1 U10882 ( .A1(n12157), .A2(n9634), .ZN(n9128) );
  NAND2_X1 U10883 ( .A1(n9547), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9126) );
  INV_X1 U10884 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9119) );
  OR2_X1 U10885 ( .A1(n9608), .A2(n9119), .ZN(n9125) );
  NAND2_X1 U10886 ( .A1(n9121), .A2(n9120), .ZN(n9122) );
  NAND2_X1 U10887 ( .A1(n9152), .A2(n9122), .ZN(n12154) );
  OR2_X1 U10888 ( .A1(n9624), .A2(n12154), .ZN(n9124) );
  INV_X1 U10889 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n14429) );
  OR2_X1 U10890 ( .A1(n7209), .A2(n14429), .ZN(n9123) );
  NAND4_X1 U10891 ( .A1(n9126), .A2(n9125), .A3(n9124), .A4(n9123), .ZN(n14367) );
  NAND2_X1 U10892 ( .A1(n14367), .A2(n9615), .ZN(n9127) );
  NAND2_X1 U10893 ( .A1(n9128), .A2(n9127), .ZN(n9131) );
  NAND2_X1 U10894 ( .A1(n12157), .A2(n9615), .ZN(n9129) );
  OAI21_X1 U10895 ( .B1(n11720), .B2(n9615), .A(n9129), .ZN(n9130) );
  INV_X1 U10896 ( .A(n9131), .ZN(n9132) );
  INV_X1 U10897 ( .A(n9136), .ZN(n9133) );
  AOI22_X1 U10898 ( .A1(n13136), .A2(n9133), .B1(n9138), .B2(n13133), .ZN(
        n9134) );
  NAND2_X1 U10899 ( .A1(n9136), .A2(SI_9_), .ZN(n9137) );
  INV_X1 U10900 ( .A(n9137), .ZN(n9141) );
  NAND2_X1 U10901 ( .A1(n9137), .A2(n13133), .ZN(n9140) );
  INV_X1 U10902 ( .A(n9138), .ZN(n9139) );
  AOI22_X1 U10903 ( .A1(n9141), .A2(SI_10_), .B1(n9140), .B2(n9139), .ZN(n9142) );
  MUX2_X1 U10904 ( .A(n10395), .B(n10397), .S(n10252), .Z(n9143) );
  NAND2_X1 U10905 ( .A1(n9143), .A2(n13130), .ZN(n9167) );
  INV_X1 U10906 ( .A(n9143), .ZN(n9144) );
  NAND2_X1 U10907 ( .A1(n9144), .A2(SI_11_), .ZN(n9145) );
  NAND2_X1 U10908 ( .A1(n9167), .A2(n9145), .ZN(n9165) );
  XNOR2_X1 U10909 ( .A(n9166), .B(n9165), .ZN(n10394) );
  INV_X4 U10910 ( .A(n9599), .ZN(n9620) );
  NAND2_X1 U10911 ( .A1(n10394), .A2(n9620), .ZN(n9149) );
  NAND2_X1 U10912 ( .A1(n9146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9147) );
  XNOR2_X1 U10913 ( .A(n9147), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U10914 ( .A1(n11080), .A2(n9353), .B1(P1_DATAO_REG_11__SCAN_IN), 
        .B2(n9354), .ZN(n9148) );
  NAND2_X1 U10915 ( .A1(n12091), .A2(n9615), .ZN(n9159) );
  NAND2_X1 U10916 ( .A1(n9547), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9157) );
  INV_X1 U10917 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9150) );
  OR2_X1 U10918 ( .A1(n9608), .A2(n9150), .ZN(n9156) );
  INV_X1 U10919 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11697) );
  NAND2_X1 U10920 ( .A1(n9152), .A2(n11697), .ZN(n9153) );
  NAND2_X1 U10921 ( .A1(n9204), .A2(n9153), .ZN(n11694) );
  OR2_X1 U10922 ( .A1(n9624), .A2(n11694), .ZN(n9155) );
  INV_X1 U10923 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11092) );
  OR2_X1 U10924 ( .A1(n7208), .A2(n11092), .ZN(n9154) );
  NAND4_X1 U10925 ( .A1(n9157), .A2(n9156), .A3(n9155), .A4(n9154), .ZN(n14366) );
  NAND2_X1 U10926 ( .A1(n14366), .A2(n9634), .ZN(n9158) );
  NAND2_X1 U10927 ( .A1(n9159), .A2(n9158), .ZN(n9161) );
  AOI22_X1 U10928 ( .A1(n12091), .A2(n9634), .B1(n9615), .B2(n14366), .ZN(
        n9160) );
  NOR2_X1 U10929 ( .A1(n9162), .A2(n9161), .ZN(n9163) );
  MUX2_X1 U10930 ( .A(n10422), .B(n10420), .S(n10252), .Z(n9168) );
  NAND2_X1 U10931 ( .A1(n9168), .A2(n13019), .ZN(n9191) );
  INV_X1 U10932 ( .A(n9168), .ZN(n9169) );
  NAND2_X1 U10933 ( .A1(n9169), .A2(SI_12_), .ZN(n9170) );
  OR2_X1 U10934 ( .A1(n9171), .A2(n8244), .ZN(n9172) );
  NAND2_X1 U10935 ( .A1(n9192), .A2(n9172), .ZN(n10419) );
  NAND2_X1 U10936 ( .A1(n10419), .A2(n9620), .ZN(n9180) );
  INV_X1 U10937 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9174) );
  NAND3_X1 U10938 ( .A1(n9175), .A2(n9174), .A3(n9173), .ZN(n9176) );
  OAI21_X1 U10939 ( .B1(n9177), .B2(n9176), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9178) );
  XNOR2_X1 U10940 ( .A(n9178), .B(P2_IR_REG_12__SCAN_IN), .ZN(n15626) );
  AOI22_X1 U10941 ( .A1(n9353), .A2(n15626), .B1(n9354), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U10942 ( .A1(n12179), .A2(n9634), .ZN(n9188) );
  NAND2_X1 U10943 ( .A1(n9626), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9186) );
  INV_X1 U10944 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9181) );
  OR2_X1 U10945 ( .A1(n7494), .A2(n9181), .ZN(n9185) );
  XNOR2_X1 U10946 ( .A(n9204), .B(n12288), .ZN(n12108) );
  OR2_X1 U10947 ( .A1(n9624), .A2(n12108), .ZN(n9184) );
  INV_X1 U10948 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9182) );
  OR2_X1 U10949 ( .A1(n7209), .A2(n9182), .ZN(n9183) );
  NAND4_X1 U10950 ( .A1(n9186), .A2(n9185), .A3(n9184), .A4(n9183), .ZN(n14365) );
  NAND2_X1 U10951 ( .A1(n14365), .A2(n9615), .ZN(n9187) );
  NAND2_X1 U10952 ( .A1(n9188), .A2(n9187), .ZN(n9190) );
  AOI22_X1 U10953 ( .A1(n12179), .A2(n9615), .B1(n14365), .B2(n9634), .ZN(
        n9189) );
  MUX2_X1 U10954 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10252), .Z(n9224) );
  XNOR2_X1 U10955 ( .A(n9224), .B(n13121), .ZN(n9221) );
  XNOR2_X1 U10956 ( .A(n9223), .B(n9221), .ZN(n10603) );
  NAND2_X1 U10957 ( .A1(n10603), .A2(n9620), .ZN(n9201) );
  AND2_X1 U10958 ( .A1(n9194), .A2(n9193), .ZN(n9198) );
  INV_X1 U10959 ( .A(n9198), .ZN(n9195) );
  NAND2_X1 U10960 ( .A1(n9195), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9196) );
  MUX2_X1 U10961 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9196), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n9199) );
  NAND2_X1 U10962 ( .A1(n9198), .A2(n9197), .ZN(n9249) );
  NAND2_X1 U10963 ( .A1(n9199), .A2(n9249), .ZN(n11098) );
  INV_X1 U10964 ( .A(n11098), .ZN(n15609) );
  AOI22_X1 U10965 ( .A1(n9354), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9353), 
        .B2(n15609), .ZN(n9200) );
  NAND2_X1 U10966 ( .A1(n12192), .A2(n9615), .ZN(n9211) );
  NAND2_X1 U10967 ( .A1(n9626), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9209) );
  INV_X1 U10968 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9202) );
  OR2_X1 U10969 ( .A1(n7494), .A2(n9202), .ZN(n9208) );
  INV_X1 U10970 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9203) );
  OAI21_X1 U10971 ( .B1(n9204), .B2(n12288), .A(n9203), .ZN(n9205) );
  NAND2_X1 U10972 ( .A1(n9205), .A2(n9230), .ZN(n12187) );
  OR2_X1 U10973 ( .A1(n9624), .A2(n12187), .ZN(n9207) );
  INV_X1 U10974 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12131) );
  OR2_X1 U10975 ( .A1(n7209), .A2(n12131), .ZN(n9206) );
  NAND4_X1 U10976 ( .A1(n9209), .A2(n9208), .A3(n9207), .A4(n9206), .ZN(n14364) );
  NAND2_X1 U10977 ( .A1(n14364), .A2(n9634), .ZN(n9210) );
  NAND2_X1 U10978 ( .A1(n9211), .A2(n9210), .ZN(n9216) );
  NAND2_X1 U10979 ( .A1(n12192), .A2(n9634), .ZN(n9212) );
  NAND2_X1 U10980 ( .A1(n9214), .A2(n9213), .ZN(n9220) );
  INV_X1 U10981 ( .A(n9215), .ZN(n9218) );
  INV_X1 U10982 ( .A(n9216), .ZN(n9217) );
  NAND2_X1 U10983 ( .A1(n9218), .A2(n9217), .ZN(n9219) );
  INV_X1 U10984 ( .A(n9221), .ZN(n9222) );
  NAND2_X1 U10985 ( .A1(n9224), .A2(SI_13_), .ZN(n9225) );
  XNOR2_X1 U10986 ( .A(n9274), .B(SI_14_), .ZN(n9241) );
  MUX2_X1 U10987 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10252), .Z(n9275) );
  XNOR2_X1 U10988 ( .A(n9241), .B(n9275), .ZN(n10926) );
  NAND2_X1 U10989 ( .A1(n10926), .A2(n9620), .ZN(n9228) );
  NAND2_X1 U10990 ( .A1(n9249), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9226) );
  XNOR2_X1 U10991 ( .A(n9226), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U10992 ( .A1(n9354), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9353), 
        .B2(n11558), .ZN(n9227) );
  NAND2_X1 U10993 ( .A1(n16111), .A2(n9634), .ZN(n9238) );
  INV_X1 U10994 ( .A(n9230), .ZN(n9229) );
  INV_X1 U10995 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U10996 ( .A1(n9230), .A2(n12270), .ZN(n9231) );
  NAND2_X1 U10997 ( .A1(n9257), .A2(n9231), .ZN(n12269) );
  OR2_X1 U10998 ( .A1(n12269), .A2(n9624), .ZN(n9236) );
  INV_X1 U10999 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9232) );
  OR2_X1 U11000 ( .A1(n9608), .A2(n9232), .ZN(n9235) );
  INV_X1 U11001 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11086) );
  OR2_X1 U11002 ( .A1(n7494), .A2(n11086), .ZN(n9234) );
  INV_X1 U11003 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n12122) );
  OR2_X1 U11004 ( .A1(n7208), .A2(n12122), .ZN(n9233) );
  NAND4_X1 U11005 ( .A1(n9236), .A2(n9235), .A3(n9234), .A4(n9233), .ZN(n14363) );
  NAND2_X1 U11006 ( .A1(n14363), .A2(n9615), .ZN(n9237) );
  NAND2_X1 U11007 ( .A1(n9238), .A2(n9237), .ZN(n9240) );
  AOI22_X1 U11008 ( .A1(n16111), .A2(n9615), .B1(n14363), .B2(n9634), .ZN(
        n9239) );
  INV_X1 U11009 ( .A(n9241), .ZN(n9242) );
  NAND2_X1 U11010 ( .A1(n9242), .A2(n9275), .ZN(n9244) );
  NAND2_X1 U11011 ( .A1(n9274), .A2(SI_14_), .ZN(n9243) );
  NAND2_X1 U11012 ( .A1(n9244), .A2(n9243), .ZN(n9248) );
  MUX2_X1 U11013 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n10252), .Z(n9245) );
  INV_X1 U11014 ( .A(n9245), .ZN(n9246) );
  NAND2_X1 U11015 ( .A1(n9246), .A2(n13122), .ZN(n9276) );
  NAND2_X1 U11016 ( .A1(n9278), .A2(n9276), .ZN(n9247) );
  NAND2_X1 U11017 ( .A1(n11012), .A2(n9620), .ZN(n9254) );
  NAND2_X1 U11018 ( .A1(n9251), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9250) );
  MUX2_X1 U11019 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9250), .S(
        P2_IR_REG_15__SCAN_IN), .Z(n9252) );
  AND2_X1 U11020 ( .A1(n9252), .A2(n9281), .ZN(n12322) );
  AOI22_X1 U11021 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n9354), .B1(n12322), 
        .B2(n9353), .ZN(n9253) );
  NAND2_X2 U11022 ( .A1(n9254), .A2(n9253), .ZN(n14359) );
  NAND2_X1 U11023 ( .A1(n14359), .A2(n9636), .ZN(n9266) );
  INV_X1 U11024 ( .A(n9257), .ZN(n9255) );
  INV_X1 U11025 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9256) );
  NAND2_X1 U11026 ( .A1(n9257), .A2(n9256), .ZN(n9258) );
  NAND2_X1 U11027 ( .A1(n9285), .A2(n9258), .ZN(n14350) );
  NOR2_X1 U11028 ( .A1(n14350), .A2(n9624), .ZN(n9264) );
  INV_X1 U11029 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9260) );
  NAND2_X1 U11030 ( .A1(n9626), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9259) );
  OAI21_X1 U11031 ( .B1(n9260), .B2(n7494), .A(n9259), .ZN(n9263) );
  INV_X1 U11032 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9261) );
  NOR2_X1 U11033 ( .A1(n7209), .A2(n9261), .ZN(n9262) );
  NAND2_X1 U11034 ( .A1(n14362), .A2(n9634), .ZN(n9265) );
  NAND2_X1 U11035 ( .A1(n9266), .A2(n9265), .ZN(n9269) );
  INV_X1 U11036 ( .A(n14362), .ZN(n12425) );
  NAND2_X1 U11037 ( .A1(n14359), .A2(n9634), .ZN(n9267) );
  OAI21_X1 U11038 ( .B1(n12425), .B2(n9634), .A(n9267), .ZN(n9268) );
  INV_X1 U11039 ( .A(n9268), .ZN(n9271) );
  INV_X1 U11040 ( .A(n9275), .ZN(n9273) );
  NOR2_X1 U11041 ( .A1(n9275), .A2(SI_14_), .ZN(n9279) );
  INV_X1 U11042 ( .A(n9276), .ZN(n9277) );
  MUX2_X1 U11043 ( .A(n10925), .B(n10923), .S(n10252), .Z(n9294) );
  XNOR2_X1 U11044 ( .A(n9294), .B(SI_16_), .ZN(n9293) );
  XNOR2_X1 U11045 ( .A(n9298), .B(n9293), .ZN(n10922) );
  NAND2_X1 U11046 ( .A1(n10922), .A2(n9620), .ZN(n9284) );
  NAND2_X1 U11047 ( .A1(n9281), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9282) );
  XNOR2_X1 U11048 ( .A(n9282), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15595) );
  AOI22_X1 U11049 ( .A1(n9353), .A2(n15595), .B1(n9354), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n9283) );
  NAND2_X1 U11050 ( .A1(n14808), .A2(n9634), .ZN(n9290) );
  NAND2_X1 U11051 ( .A1(n9285), .A2(n15589), .ZN(n9286) );
  NAND2_X1 U11052 ( .A1(n9310), .A2(n9286), .ZN(n12539) );
  AOI22_X1 U11053 ( .A1(n9547), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n9626), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n9288) );
  INV_X1 U11054 ( .A(n7208), .ZN(n9625) );
  NAND2_X1 U11055 ( .A1(n9625), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9287) );
  OAI211_X1 U11056 ( .C1(n12539), .C2(n9624), .A(n9288), .B(n9287), .ZN(n14463) );
  NAND2_X1 U11057 ( .A1(n14463), .A2(n9615), .ZN(n9289) );
  NAND2_X1 U11058 ( .A1(n9290), .A2(n9289), .ZN(n9292) );
  INV_X1 U11059 ( .A(n9294), .ZN(n9295) );
  NAND2_X1 U11060 ( .A1(n9295), .A2(SI_16_), .ZN(n9296) );
  MUX2_X1 U11061 ( .A(n11038), .B(n11040), .S(n10252), .Z(n9299) );
  INV_X1 U11062 ( .A(n9299), .ZN(n9300) );
  NAND2_X1 U11063 ( .A1(n9300), .A2(SI_17_), .ZN(n9301) );
  NAND2_X1 U11064 ( .A1(n9324), .A2(n9301), .ZN(n9302) );
  NAND2_X1 U11065 ( .A1(n9303), .A2(n9302), .ZN(n9304) );
  NAND2_X1 U11066 ( .A1(n9325), .A2(n9304), .ZN(n11037) );
  NAND2_X1 U11067 ( .A1(n11037), .A2(n9620), .ZN(n9307) );
  NAND2_X1 U11068 ( .A1(n9305), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9327) );
  XNOR2_X1 U11069 ( .A(n9327), .B(P2_IR_REG_17__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U11070 ( .A1(n9354), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9353), 
        .B2(n12337), .ZN(n9306) );
  INV_X1 U11071 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n12335) );
  INV_X1 U11072 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U11073 ( .A1(n9310), .A2(n9309), .ZN(n9311) );
  NAND2_X1 U11074 ( .A1(n9332), .A2(n9311), .ZN(n14719) );
  OR2_X1 U11075 ( .A1(n14719), .A2(n9624), .ZN(n9313) );
  AOI22_X1 U11076 ( .A1(n9625), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9626), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n9312) );
  OAI211_X1 U11077 ( .C1(n7494), .C2(n12335), .A(n9313), .B(n9312), .ZN(n14466) );
  AND2_X1 U11078 ( .A1(n14466), .A2(n9634), .ZN(n9314) );
  INV_X1 U11079 ( .A(n9320), .ZN(n9315) );
  INV_X1 U11080 ( .A(n14466), .ZN(n14495) );
  NAND2_X1 U11081 ( .A1(n14723), .A2(n9634), .ZN(n9316) );
  NAND2_X1 U11082 ( .A1(n9318), .A2(n9317), .ZN(n9323) );
  INV_X1 U11083 ( .A(n9319), .ZN(n9321) );
  NAND2_X1 U11084 ( .A1(n9321), .A2(n9320), .ZN(n9322) );
  INV_X1 U11085 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11321) );
  MUX2_X1 U11086 ( .A(n11323), .B(n11321), .S(n7215), .Z(n9373) );
  XNOR2_X1 U11087 ( .A(n9345), .B(n9373), .ZN(n11320) );
  NAND2_X1 U11088 ( .A1(n11320), .A2(n9620), .ZN(n9331) );
  NAND2_X1 U11089 ( .A1(n9327), .A2(n9326), .ZN(n9328) );
  NAND2_X1 U11090 ( .A1(n9328), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9329) );
  XNOR2_X1 U11091 ( .A(n9329), .B(P2_IR_REG_18__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U11092 ( .A1(n9354), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9353), 
        .B2(n11319), .ZN(n9330) );
  NAND2_X1 U11093 ( .A1(n14698), .A2(n9634), .ZN(n9342) );
  INV_X1 U11094 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U11095 ( .A1(n9332), .A2(n12340), .ZN(n9333) );
  AND2_X1 U11096 ( .A1(n9359), .A2(n9333), .ZN(n14696) );
  NAND2_X1 U11097 ( .A1(n14696), .A2(n9546), .ZN(n9340) );
  INV_X1 U11098 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9337) );
  NAND2_X1 U11099 ( .A1(n9626), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9336) );
  NAND2_X1 U11100 ( .A1(n9547), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9335) );
  OAI211_X1 U11101 ( .C1(n7209), .C2(n9337), .A(n9336), .B(n9335), .ZN(n9338)
         );
  INV_X1 U11102 ( .A(n9338), .ZN(n9339) );
  NAND2_X1 U11103 ( .A1(n9340), .A2(n9339), .ZN(n14497) );
  NAND2_X1 U11104 ( .A1(n14497), .A2(n9615), .ZN(n9341) );
  NAND2_X1 U11105 ( .A1(n9342), .A2(n9341), .ZN(n9344) );
  AOI22_X1 U11106 ( .A1(n14698), .A2(n9615), .B1(n14497), .B2(n9634), .ZN(
        n9343) );
  INV_X1 U11107 ( .A(n9373), .ZN(n9376) );
  NAND2_X1 U11108 ( .A1(n9345), .A2(n9376), .ZN(n9348) );
  INV_X1 U11109 ( .A(n9375), .ZN(n9346) );
  NAND2_X1 U11110 ( .A1(n9346), .A2(SI_18_), .ZN(n9347) );
  NAND2_X1 U11111 ( .A1(n9348), .A2(n9347), .ZN(n9352) );
  MUX2_X1 U11112 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n7215), .Z(n9349) );
  NAND2_X1 U11113 ( .A1(n9349), .A2(SI_19_), .ZN(n9379) );
  INV_X1 U11114 ( .A(n9349), .ZN(n9350) );
  NAND2_X1 U11115 ( .A1(n9350), .A2(n13092), .ZN(n9377) );
  NAND2_X1 U11116 ( .A1(n9379), .A2(n9377), .ZN(n9351) );
  NAND2_X1 U11117 ( .A1(n11421), .A2(n9620), .ZN(n9356) );
  AOI22_X1 U11118 ( .A1(n9354), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n12410), 
        .B2(n9353), .ZN(n9355) );
  NAND2_X2 U11119 ( .A1(n9356), .A2(n9355), .ZN(n14686) );
  NAND2_X1 U11120 ( .A1(n14686), .A2(n9615), .ZN(n9367) );
  INV_X1 U11121 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11122 ( .A1(n9359), .A2(n9358), .ZN(n9360) );
  NAND2_X1 U11123 ( .A1(n9386), .A2(n9360), .ZN(n14683) );
  OR2_X1 U11124 ( .A1(n14683), .A2(n9624), .ZN(n9365) );
  INV_X1 U11125 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14684) );
  NAND2_X1 U11126 ( .A1(n9547), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U11127 ( .A1(n9626), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9361) );
  OAI211_X1 U11128 ( .C1(n14684), .C2(n7209), .A(n9362), .B(n9361), .ZN(n9363)
         );
  INV_X1 U11129 ( .A(n9363), .ZN(n9364) );
  NAND2_X1 U11130 ( .A1(n9365), .A2(n9364), .ZN(n14470) );
  NAND2_X1 U11131 ( .A1(n14470), .A2(n9634), .ZN(n9366) );
  NAND2_X1 U11132 ( .A1(n9367), .A2(n9366), .ZN(n9369) );
  AOI22_X1 U11133 ( .A1(n14686), .A2(n9634), .B1(n9615), .B2(n14470), .ZN(
        n9368) );
  NOR2_X1 U11134 ( .A1(n9370), .A2(n9369), .ZN(n9371) );
  OAI21_X1 U11135 ( .B1(n13093), .B2(n9373), .A(n9379), .ZN(n9374) );
  NOR2_X1 U11136 ( .A1(n9376), .A2(SI_18_), .ZN(n9380) );
  INV_X1 U11137 ( .A(n9377), .ZN(n9378) );
  AOI21_X1 U11138 ( .B1(n9380), .B2(n9379), .A(n9378), .ZN(n9381) );
  MUX2_X1 U11139 ( .A(n11325), .B(n11428), .S(n10252), .Z(n9402) );
  XNOR2_X1 U11140 ( .A(n9402), .B(SI_20_), .ZN(n9383) );
  XNOR2_X1 U11141 ( .A(n7441), .B(n9383), .ZN(n11324) );
  NAND2_X1 U11142 ( .A1(n11324), .A2(n9620), .ZN(n9385) );
  OR2_X1 U11143 ( .A1(n9621), .A2(n11428), .ZN(n9384) );
  NAND2_X1 U11144 ( .A1(n14789), .A2(n9634), .ZN(n9394) );
  NAND2_X1 U11145 ( .A1(n9386), .A2(n14304), .ZN(n9387) );
  NAND2_X1 U11146 ( .A1(n9410), .A2(n9387), .ZN(n14663) );
  OR2_X1 U11147 ( .A1(n14663), .A2(n9624), .ZN(n9392) );
  INV_X1 U11148 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n14664) );
  NAND2_X1 U11149 ( .A1(n9547), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U11150 ( .A1(n9626), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9388) );
  OAI211_X1 U11151 ( .C1(n14664), .C2(n7208), .A(n9389), .B(n9388), .ZN(n9390)
         );
  INV_X1 U11152 ( .A(n9390), .ZN(n9391) );
  NAND2_X1 U11153 ( .A1(n14474), .A2(n9615), .ZN(n9393) );
  NAND2_X1 U11154 ( .A1(n9394), .A2(n9393), .ZN(n9398) );
  INV_X1 U11155 ( .A(n14474), .ZN(n14505) );
  NAND2_X1 U11156 ( .A1(n14789), .A2(n9615), .ZN(n9395) );
  INV_X1 U11157 ( .A(n9398), .ZN(n9399) );
  NAND2_X1 U11158 ( .A1(n9400), .A2(n9399), .ZN(n9401) );
  MUX2_X1 U11159 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10252), .Z(n9404) );
  OAI21_X1 U11160 ( .B1(SI_21_), .B2(n9404), .A(n9424), .ZN(n9405) );
  NAND2_X1 U11161 ( .A1(n9406), .A2(n9405), .ZN(n9407) );
  NAND2_X1 U11162 ( .A1(n9425), .A2(n9407), .ZN(n11418) );
  OR2_X1 U11163 ( .A1(n11418), .A2(n9599), .ZN(n9409) );
  OR2_X1 U11164 ( .A1(n9621), .A2(n11376), .ZN(n9408) );
  NAND2_X1 U11165 ( .A1(n14784), .A2(n9615), .ZN(n9419) );
  INV_X1 U11166 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n14244) );
  NAND2_X1 U11167 ( .A1(n9410), .A2(n14244), .ZN(n9411) );
  AND2_X1 U11168 ( .A1(n9434), .A2(n9411), .ZN(n14653) );
  NAND2_X1 U11169 ( .A1(n14653), .A2(n9546), .ZN(n9417) );
  INV_X1 U11170 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U11171 ( .A1(n9547), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n9413) );
  NAND2_X1 U11172 ( .A1(n9626), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9412) );
  OAI211_X1 U11173 ( .C1(n9414), .C2(n7209), .A(n9413), .B(n9412), .ZN(n9415)
         );
  INV_X1 U11174 ( .A(n9415), .ZN(n9416) );
  NAND2_X1 U11175 ( .A1(n14507), .A2(n9634), .ZN(n9418) );
  NAND2_X1 U11176 ( .A1(n9419), .A2(n9418), .ZN(n9422) );
  INV_X1 U11177 ( .A(n14507), .ZN(n14314) );
  NAND2_X1 U11178 ( .A1(n14784), .A2(n9634), .ZN(n9420) );
  OAI21_X1 U11179 ( .B1(n14314), .B2(n9634), .A(n9420), .ZN(n9421) );
  INV_X1 U11180 ( .A(n9422), .ZN(n9423) );
  MUX2_X1 U11181 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10252), .Z(n9426) );
  INV_X1 U11182 ( .A(n9752), .ZN(n9428) );
  INV_X1 U11183 ( .A(n9426), .ZN(n9427) );
  NAND2_X1 U11184 ( .A1(n9428), .A2(n9427), .ZN(n9429) );
  NAND2_X1 U11185 ( .A1(n9451), .A2(n9429), .ZN(n11872) );
  OR2_X1 U11186 ( .A1(n9621), .A2(n11873), .ZN(n9430) );
  NAND2_X1 U11187 ( .A1(n14778), .A2(n9634), .ZN(n9443) );
  INV_X1 U11188 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U11189 ( .A1(n9434), .A2(n9433), .ZN(n9435) );
  NAND2_X1 U11190 ( .A1(n9457), .A2(n9435), .ZN(n14636) );
  OR2_X1 U11191 ( .A1(n14636), .A2(n9624), .ZN(n9441) );
  INV_X1 U11192 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9438) );
  NAND2_X1 U11193 ( .A1(n9547), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9437) );
  NAND2_X1 U11194 ( .A1(n9626), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9436) );
  OAI211_X1 U11195 ( .C1(n9438), .C2(n7209), .A(n9437), .B(n9436), .ZN(n9439)
         );
  INV_X1 U11196 ( .A(n9439), .ZN(n9440) );
  NAND2_X1 U11197 ( .A1(n14476), .A2(n9615), .ZN(n9442) );
  NAND2_X1 U11198 ( .A1(n9443), .A2(n9442), .ZN(n9446) );
  AOI22_X1 U11199 ( .A1(n14778), .A2(n9615), .B1(n14476), .B2(n9634), .ZN(
        n9444) );
  AOI21_X1 U11200 ( .B1(n9447), .B2(n9446), .A(n9444), .ZN(n9445) );
  NOR2_X1 U11201 ( .A1(n9447), .A2(n9446), .ZN(n9448) );
  MUX2_X1 U11202 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10252), .Z(n9470) );
  XNOR2_X1 U11203 ( .A(n9470), .B(SI_23_), .ZN(n9452) );
  NAND2_X1 U11204 ( .A1(n12611), .A2(n9620), .ZN(n9454) );
  OR2_X1 U11205 ( .A1(n9621), .A2(n11954), .ZN(n9453) );
  NAND2_X1 U11206 ( .A1(n14769), .A2(n9615), .ZN(n9466) );
  INV_X1 U11207 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9456) );
  NAND2_X1 U11208 ( .A1(n9457), .A2(n9456), .ZN(n9458) );
  NAND2_X1 U11209 ( .A1(n9477), .A2(n9458), .ZN(n14621) );
  OR2_X1 U11210 ( .A1(n14621), .A2(n9624), .ZN(n9464) );
  INV_X1 U11211 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U11212 ( .A1(n9547), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U11213 ( .A1(n9626), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9459) );
  OAI211_X1 U11214 ( .C1(n9461), .C2(n7209), .A(n9460), .B(n9459), .ZN(n9462)
         );
  INV_X1 U11215 ( .A(n9462), .ZN(n9463) );
  NAND2_X1 U11216 ( .A1(n9464), .A2(n9463), .ZN(n14478) );
  NAND2_X1 U11217 ( .A1(n14478), .A2(n9634), .ZN(n9465) );
  INV_X1 U11218 ( .A(n14478), .ZN(n14512) );
  NAND2_X1 U11219 ( .A1(n14769), .A2(n9634), .ZN(n9467) );
  OAI21_X1 U11220 ( .B1(n14512), .B2(n9634), .A(n9467), .ZN(n9468) );
  NAND2_X1 U11221 ( .A1(n9471), .A2(SI_23_), .ZN(n9472) );
  MUX2_X1 U11222 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10252), .Z(n9488) );
  XNOR2_X1 U11223 ( .A(n9488), .B(SI_24_), .ZN(n9474) );
  NAND2_X1 U11224 ( .A1(n12598), .A2(n9620), .ZN(n9476) );
  OR2_X1 U11225 ( .A1(n9621), .A2(n12201), .ZN(n9475) );
  NAND2_X1 U11226 ( .A1(n14609), .A2(n9634), .ZN(n9486) );
  INV_X1 U11227 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n14291) );
  NAND2_X1 U11228 ( .A1(n9477), .A2(n14291), .ZN(n9478) );
  AND2_X1 U11229 ( .A1(n9498), .A2(n9478), .ZN(n14608) );
  NAND2_X1 U11230 ( .A1(n14608), .A2(n9546), .ZN(n9484) );
  INV_X1 U11231 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n9481) );
  NAND2_X1 U11232 ( .A1(n9547), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U11233 ( .A1(n9626), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9479) );
  OAI211_X1 U11234 ( .C1(n9481), .C2(n7208), .A(n9480), .B(n9479), .ZN(n9482)
         );
  INV_X1 U11235 ( .A(n9482), .ZN(n9483) );
  NAND2_X1 U11236 ( .A1(n14480), .A2(n9615), .ZN(n9485) );
  AOI22_X1 U11237 ( .A1(n14609), .A2(n9615), .B1(n14480), .B2(n9634), .ZN(
        n9487) );
  OAI21_X1 U11238 ( .B1(n9489), .B2(SI_24_), .A(n9488), .ZN(n9491) );
  NAND2_X1 U11239 ( .A1(n9489), .A2(SI_24_), .ZN(n9490) );
  NAND2_X1 U11240 ( .A1(n9491), .A2(n9490), .ZN(n9517) );
  MUX2_X1 U11241 ( .A(n12589), .B(n8113), .S(n10252), .Z(n9492) );
  NAND2_X1 U11242 ( .A1(n9492), .A2(n12348), .ZN(n9518) );
  INV_X1 U11243 ( .A(n9492), .ZN(n9493) );
  NAND2_X1 U11244 ( .A1(n9493), .A2(SI_25_), .ZN(n9494) );
  NAND2_X1 U11245 ( .A1(n9518), .A2(n9494), .ZN(n9516) );
  NAND2_X1 U11246 ( .A1(n12588), .A2(n9620), .ZN(n9496) );
  OR2_X1 U11247 ( .A1(n9621), .A2(n8113), .ZN(n9495) );
  NAND2_X1 U11248 ( .A1(n14759), .A2(n9615), .ZN(n9506) );
  INV_X1 U11249 ( .A(n9498), .ZN(n9497) );
  INV_X1 U11250 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n14258) );
  NAND2_X1 U11251 ( .A1(n9498), .A2(n14258), .ZN(n9499) );
  NAND2_X1 U11252 ( .A1(n9523), .A2(n9499), .ZN(n14589) );
  OR2_X1 U11253 ( .A1(n14589), .A2(n9624), .ZN(n9504) );
  INV_X1 U11254 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n14588) );
  NAND2_X1 U11255 ( .A1(n9547), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U11256 ( .A1(n9626), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9500) );
  OAI211_X1 U11257 ( .C1(n14588), .C2(n7208), .A(n9501), .B(n9500), .ZN(n9502)
         );
  INV_X1 U11258 ( .A(n9502), .ZN(n9503) );
  NAND2_X1 U11259 ( .A1(n14482), .A2(n9634), .ZN(n9505) );
  NAND2_X1 U11260 ( .A1(n9506), .A2(n9505), .ZN(n9511) );
  NAND2_X1 U11261 ( .A1(n9510), .A2(n9511), .ZN(n9509) );
  AOI22_X1 U11262 ( .A1(n14759), .A2(n9634), .B1(n9615), .B2(n14482), .ZN(
        n9507) );
  INV_X1 U11263 ( .A(n9507), .ZN(n9508) );
  INV_X1 U11264 ( .A(n9510), .ZN(n9513) );
  INV_X1 U11265 ( .A(n9511), .ZN(n9512) );
  INV_X1 U11266 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12617) );
  MUX2_X1 U11267 ( .A(n12617), .B(n12452), .S(n10252), .Z(n9538) );
  XNOR2_X1 U11268 ( .A(n9538), .B(SI_26_), .ZN(n9535) );
  XNOR2_X1 U11269 ( .A(n9537), .B(n9535), .ZN(n12616) );
  NAND2_X1 U11270 ( .A1(n12616), .A2(n9620), .ZN(n9521) );
  OR2_X1 U11271 ( .A1(n9621), .A2(n12452), .ZN(n9520) );
  INV_X1 U11272 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9522) );
  NAND2_X1 U11273 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  INV_X1 U11274 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U11275 ( .A1(n9626), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U11276 ( .A1(n9547), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9525) );
  OAI211_X1 U11277 ( .C1(n7209), .C2(n9527), .A(n9526), .B(n9525), .ZN(n9528)
         );
  OAI22_X1 U11278 ( .A1(n14573), .A2(n9615), .B1(n14484), .B2(n9634), .ZN(
        n9530) );
  NAND2_X1 U11279 ( .A1(n9529), .A2(n9530), .ZN(n9534) );
  INV_X1 U11280 ( .A(n9529), .ZN(n9532) );
  INV_X1 U11281 ( .A(n9530), .ZN(n9531) );
  INV_X1 U11282 ( .A(n9535), .ZN(n9536) );
  INV_X1 U11283 ( .A(n9538), .ZN(n9539) );
  NAND2_X1 U11284 ( .A1(n9539), .A2(SI_26_), .ZN(n9540) );
  MUX2_X1 U11285 ( .A(n15511), .B(n14870), .S(n7215), .Z(n9541) );
  NAND2_X1 U11286 ( .A1(n9541), .A2(n13101), .ZN(n9555) );
  INV_X1 U11287 ( .A(n9541), .ZN(n9542) );
  NAND2_X1 U11288 ( .A1(n9542), .A2(SI_27_), .ZN(n9543) );
  NAND2_X1 U11289 ( .A1(n9555), .A2(n9543), .ZN(n9553) );
  NAND2_X1 U11290 ( .A1(n14867), .A2(n9620), .ZN(n9545) );
  OR2_X1 U11291 ( .A1(n9621), .A2(n14870), .ZN(n9544) );
  XNOR2_X1 U11292 ( .A(n9583), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n14205) );
  NAND2_X1 U11293 ( .A1(n14205), .A2(n9546), .ZN(n9552) );
  INV_X1 U11294 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n14556) );
  NAND2_X1 U11295 ( .A1(n9547), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U11296 ( .A1(n9626), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9548) );
  OAI211_X1 U11297 ( .C1(n14556), .C2(n7209), .A(n9549), .B(n9548), .ZN(n9550)
         );
  INV_X1 U11298 ( .A(n9550), .ZN(n9551) );
  AOI22_X1 U11299 ( .A1(n14563), .A2(n9615), .B1(n14520), .B2(n9634), .ZN(
        n9642) );
  INV_X1 U11300 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12671) );
  MUX2_X1 U11301 ( .A(n12671), .B(n14865), .S(n10252), .Z(n9556) );
  NAND2_X1 U11302 ( .A1(n9556), .A2(n14156), .ZN(n9559) );
  INV_X1 U11303 ( .A(n9556), .ZN(n9557) );
  NAND2_X1 U11304 ( .A1(n9557), .A2(SI_28_), .ZN(n9558) );
  INV_X1 U11305 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12579) );
  MUX2_X1 U11306 ( .A(n15507), .B(n12579), .S(n10252), .Z(n9560) );
  XNOR2_X1 U11307 ( .A(n9560), .B(SI_29_), .ZN(n9618) );
  NAND2_X1 U11308 ( .A1(n9619), .A2(n9618), .ZN(n9562) );
  INV_X1 U11309 ( .A(SI_29_), .ZN(n14151) );
  NAND2_X1 U11310 ( .A1(n9560), .A2(n14151), .ZN(n9561) );
  MUX2_X1 U11311 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10252), .Z(n9563) );
  NAND2_X1 U11312 ( .A1(n9563), .A2(SI_30_), .ZN(n9564) );
  OAI21_X1 U11313 ( .B1(n9563), .B2(SI_30_), .A(n9564), .ZN(n9595) );
  NAND2_X1 U11314 ( .A1(n9598), .A2(n9564), .ZN(n9567) );
  MUX2_X1 U11315 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7215), .Z(n9565) );
  XNOR2_X1 U11316 ( .A(n9565), .B(SI_31_), .ZN(n9566) );
  NAND2_X1 U11317 ( .A1(n14851), .A2(n9620), .ZN(n9569) );
  INV_X1 U11318 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14854) );
  OR2_X1 U11319 ( .A1(n9621), .A2(n14854), .ZN(n9568) );
  INV_X1 U11320 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9570) );
  OR2_X1 U11321 ( .A1(n7494), .A2(n9570), .ZN(n9575) );
  INV_X1 U11322 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n14450) );
  OR2_X1 U11323 ( .A1(n7209), .A2(n14450), .ZN(n9574) );
  INV_X1 U11324 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9572) );
  OR2_X1 U11325 ( .A1(n9608), .A2(n9572), .ZN(n9573) );
  AND3_X1 U11326 ( .A1(n9575), .A2(n9574), .A3(n9573), .ZN(n9604) );
  XNOR2_X1 U11327 ( .A(n14730), .B(n9604), .ZN(n9677) );
  NAND2_X1 U11328 ( .A1(n14862), .A2(n9620), .ZN(n9581) );
  OR2_X1 U11329 ( .A1(n9621), .A2(n14865), .ZN(n9580) );
  INV_X1 U11330 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n14206) );
  INV_X1 U11331 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9582) );
  OAI21_X1 U11332 ( .B1(n9583), .B2(n14206), .A(n9582), .ZN(n9586) );
  INV_X1 U11333 ( .A(n9583), .ZN(n9585) );
  AND2_X1 U11334 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n9584) );
  NAND2_X1 U11335 ( .A1(n9585), .A2(n9584), .ZN(n14488) );
  NAND2_X1 U11336 ( .A1(n9586), .A2(n14488), .ZN(n14543) );
  INV_X1 U11337 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n14542) );
  NAND2_X1 U11338 ( .A1(n9547), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9588) );
  NAND2_X1 U11339 ( .A1(n9626), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9587) );
  OAI211_X1 U11340 ( .C1(n14542), .C2(n7209), .A(n9588), .B(n9587), .ZN(n9589)
         );
  INV_X1 U11341 ( .A(n9589), .ZN(n9590) );
  AND2_X1 U11342 ( .A1(n14526), .A2(n9615), .ZN(n9592) );
  AOI21_X1 U11343 ( .B1(n14545), .B2(n9634), .A(n9592), .ZN(n9680) );
  NAND2_X1 U11344 ( .A1(n14545), .A2(n9615), .ZN(n9594) );
  NAND2_X1 U11345 ( .A1(n14526), .A2(n9634), .ZN(n9593) );
  NAND2_X1 U11346 ( .A1(n9594), .A2(n9593), .ZN(n9678) );
  NAND2_X1 U11347 ( .A1(n9596), .A2(n9595), .ZN(n9597) );
  OR2_X1 U11348 ( .A1(n14859), .A2(n9599), .ZN(n9601) );
  INV_X1 U11349 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14858) );
  OR2_X1 U11350 ( .A1(n9621), .A2(n14858), .ZN(n9600) );
  NAND2_X1 U11351 ( .A1(n9710), .A2(n12410), .ZN(n10477) );
  INV_X1 U11352 ( .A(n10477), .ZN(n9603) );
  NAND2_X1 U11353 ( .A1(n10467), .A2(n12414), .ZN(n10649) );
  NAND2_X1 U11354 ( .A1(n10649), .A2(n10475), .ZN(n9602) );
  AOI21_X1 U11355 ( .B1(n9603), .B2(n10467), .A(n9602), .ZN(n9612) );
  INV_X1 U11356 ( .A(n9604), .ZN(n14454) );
  NAND2_X1 U11357 ( .A1(n14454), .A2(n9634), .ZN(n9684) );
  INV_X1 U11358 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9605) );
  OR2_X1 U11359 ( .A1(n7494), .A2(n9605), .ZN(n9611) );
  INV_X1 U11360 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n14458) );
  OR2_X1 U11361 ( .A1(n7208), .A2(n14458), .ZN(n9610) );
  INV_X1 U11362 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9607) );
  OR2_X1 U11363 ( .A1(n9608), .A2(n9607), .ZN(n9609) );
  AND3_X1 U11364 ( .A1(n9611), .A2(n9610), .A3(n9609), .ZN(n9614) );
  AOI21_X1 U11365 ( .B1(n9612), .B2(n9684), .A(n9614), .ZN(n9613) );
  AOI21_X1 U11366 ( .B1(n14461), .B2(n9615), .A(n9613), .ZN(n9674) );
  NAND2_X1 U11367 ( .A1(n14461), .A2(n9634), .ZN(n9617) );
  INV_X1 U11368 ( .A(n9614), .ZN(n14528) );
  NAND2_X1 U11369 ( .A1(n14528), .A2(n9636), .ZN(n9616) );
  NAND2_X1 U11370 ( .A1(n9617), .A2(n9616), .ZN(n9673) );
  NAND2_X1 U11371 ( .A1(n9674), .A2(n9673), .ZN(n9688) );
  NAND2_X1 U11372 ( .A1(n12825), .A2(n9620), .ZN(n9623) );
  OR2_X1 U11373 ( .A1(n9621), .A2(n12579), .ZN(n9622) );
  OR2_X1 U11374 ( .A1(n14488), .A2(n9624), .ZN(n9633) );
  INV_X1 U11375 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U11376 ( .A1(n9625), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9628) );
  NAND2_X1 U11377 ( .A1(n9626), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9627) );
  OAI211_X1 U11378 ( .C1(n9630), .C2(n7494), .A(n9628), .B(n9627), .ZN(n9631)
         );
  INV_X1 U11379 ( .A(n9631), .ZN(n9632) );
  NAND2_X1 U11380 ( .A1(n9633), .A2(n9632), .ZN(n14361) );
  AND2_X1 U11381 ( .A1(n14361), .A2(n9634), .ZN(n9635) );
  AOI21_X1 U11382 ( .B1(n14736), .B2(n9615), .A(n9635), .ZN(n9672) );
  NAND2_X1 U11383 ( .A1(n14736), .A2(n9634), .ZN(n9638) );
  NAND2_X1 U11384 ( .A1(n14361), .A2(n9615), .ZN(n9637) );
  NAND2_X1 U11385 ( .A1(n9638), .A2(n9637), .ZN(n9671) );
  NAND2_X1 U11386 ( .A1(n9672), .A2(n9671), .ZN(n9679) );
  OAI211_X1 U11387 ( .C1(n9680), .C2(n9678), .A(n9688), .B(n9679), .ZN(n9639)
         );
  AOI22_X1 U11388 ( .A1(n14563), .A2(n9634), .B1(n9615), .B2(n14520), .ZN(
        n9640) );
  INV_X1 U11389 ( .A(n9640), .ZN(n9641) );
  XNOR2_X1 U11390 ( .A(n14461), .B(n14528), .ZN(n9660) );
  INV_X1 U11391 ( .A(n14526), .ZN(n9643) );
  NAND2_X1 U11392 ( .A1(n14545), .A2(n9643), .ZN(n9644) );
  XNOR2_X1 U11393 ( .A(n14609), .B(n14515), .ZN(n14514) );
  XNOR2_X1 U11394 ( .A(n14769), .B(n14478), .ZN(n14617) );
  XNOR2_X1 U11395 ( .A(n14784), .B(n14507), .ZN(n14646) );
  XNOR2_X1 U11396 ( .A(n14723), .B(n14466), .ZN(n14493) );
  XNOR2_X1 U11397 ( .A(n12192), .B(n12184), .ZN(n12012) );
  XNOR2_X1 U11398 ( .A(n12157), .B(n11720), .ZN(n12144) );
  XNOR2_X1 U11399 ( .A(n12179), .B(n14365), .ZN(n11855) );
  INV_X1 U11400 ( .A(n14370), .ZN(n11511) );
  XNOR2_X1 U11401 ( .A(n11510), .B(n11511), .ZN(n11399) );
  XNOR2_X1 U11402 ( .A(n11400), .B(n14371), .ZN(n11394) );
  XNOR2_X1 U11403 ( .A(n14375), .B(n10587), .ZN(n10594) );
  INV_X1 U11404 ( .A(n10775), .ZN(n10496) );
  NAND2_X1 U11405 ( .A1(n10683), .A2(n9646), .ZN(n11156) );
  NAND4_X1 U11406 ( .A1(n7425), .A2(n10594), .A3(n10646), .A4(n11156), .ZN(
        n9647) );
  XNOR2_X1 U11407 ( .A(n14269), .B(n14372), .ZN(n11048) );
  XNOR2_X1 U11408 ( .A(n11738), .B(n14373), .ZN(n10828) );
  NAND4_X1 U11409 ( .A1(n11394), .A2(n9648), .A3(n11048), .A4(n10828), .ZN(
        n9649) );
  NOR2_X1 U11410 ( .A1(n11399), .A2(n9649), .ZN(n9650) );
  XNOR2_X1 U11411 ( .A(n12091), .B(n14366), .ZN(n11858) );
  XNOR2_X1 U11412 ( .A(n16003), .B(n14369), .ZN(n11513) );
  NAND4_X1 U11413 ( .A1(n11855), .A2(n9650), .A3(n11858), .A4(n11513), .ZN(
        n9651) );
  INV_X1 U11414 ( .A(n14368), .ZN(n11716) );
  OR3_X1 U11415 ( .A1(n12144), .A2(n9651), .A3(n11713), .ZN(n9652) );
  NOR2_X1 U11416 ( .A1(n12012), .A2(n9652), .ZN(n9653) );
  XNOR2_X1 U11417 ( .A(n14808), .B(n14463), .ZN(n12421) );
  XNOR2_X1 U11418 ( .A(n16111), .B(n14363), .ZN(n12127) );
  NAND4_X1 U11419 ( .A1(n14493), .A2(n9653), .A3(n12421), .A4(n12127), .ZN(
        n9654) );
  XNOR2_X1 U11420 ( .A(n14359), .B(n12425), .ZN(n12357) );
  NOR2_X1 U11421 ( .A1(n9654), .A2(n12357), .ZN(n9655) );
  XNOR2_X1 U11422 ( .A(n14698), .B(n14497), .ZN(n14468) );
  XNOR2_X1 U11423 ( .A(n14789), .B(n14474), .ZN(n14669) );
  AND4_X1 U11424 ( .A1(n14646), .A2(n9655), .A3(n14468), .A4(n14669), .ZN(
        n9656) );
  XNOR2_X1 U11425 ( .A(n14778), .B(n14476), .ZN(n14630) );
  XNOR2_X1 U11426 ( .A(n14686), .B(n14470), .ZN(n14676) );
  NAND4_X1 U11427 ( .A1(n14617), .A2(n9656), .A3(n14630), .A4(n14676), .ZN(
        n9657) );
  NOR2_X1 U11428 ( .A1(n14514), .A2(n9657), .ZN(n9658) );
  XNOR2_X1 U11429 ( .A(n14759), .B(n14482), .ZN(n14581) );
  INV_X1 U11430 ( .A(n14484), .ZN(n14517) );
  XNOR2_X1 U11431 ( .A(n14755), .B(n14517), .ZN(n14576) );
  AND4_X1 U11432 ( .A1(n14486), .A2(n9658), .A3(n14581), .A4(n14576), .ZN(
        n9659) );
  XNOR2_X1 U11433 ( .A(n14736), .B(n14361), .ZN(n14524) );
  XNOR2_X1 U11434 ( .A(n14563), .B(n14520), .ZN(n14552) );
  NAND4_X1 U11435 ( .A1(n9660), .A2(n9659), .A3(n14524), .A4(n14552), .ZN(
        n9661) );
  OR2_X1 U11436 ( .A1(n9677), .A2(n9661), .ZN(n9711) );
  NAND2_X1 U11437 ( .A1(n9696), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9663) );
  INV_X1 U11438 ( .A(n10761), .ZN(n10427) );
  NAND2_X1 U11439 ( .A1(n10427), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11952) );
  NAND2_X1 U11440 ( .A1(n11375), .A2(n12410), .ZN(n9664) );
  NOR2_X1 U11441 ( .A1(n11952), .A2(n9664), .ZN(n9665) );
  NAND2_X1 U11442 ( .A1(n9711), .A2(n9665), .ZN(n9717) );
  INV_X1 U11443 ( .A(n11952), .ZN(n9712) );
  NAND2_X1 U11444 ( .A1(n10646), .A2(n11375), .ZN(n9666) );
  AND2_X1 U11445 ( .A1(n9712), .A2(n9666), .ZN(n9690) );
  AOI21_X1 U11446 ( .B1(n8886), .B2(n10467), .A(n12414), .ZN(n9667) );
  NAND2_X1 U11447 ( .A1(n9690), .A2(n9667), .ZN(n9693) );
  NAND2_X1 U11448 ( .A1(n9668), .A2(n8247), .ZN(n9723) );
  MUX2_X1 U11449 ( .A(n14454), .B(n9615), .S(n14730), .Z(n9670) );
  NAND2_X1 U11450 ( .A1(n14454), .A2(n9615), .ZN(n9669) );
  NAND2_X1 U11451 ( .A1(n9670), .A2(n9669), .ZN(n9676) );
  OAI22_X1 U11452 ( .A1(n9674), .A2(n9673), .B1(n9672), .B2(n9671), .ZN(n9675)
         );
  NAND2_X1 U11453 ( .A1(n9676), .A2(n9675), .ZN(n9683) );
  INV_X1 U11454 ( .A(n9677), .ZN(n9681) );
  NAND4_X1 U11455 ( .A1(n9681), .A2(n9680), .A3(n9679), .A4(n9678), .ZN(n9682)
         );
  NAND2_X1 U11456 ( .A1(n9683), .A2(n9682), .ZN(n9689) );
  AND2_X1 U11457 ( .A1(n9615), .A2(n14454), .ZN(n9686) );
  AND2_X1 U11458 ( .A1(n9684), .A2(n9634), .ZN(n9685) );
  MUX2_X1 U11459 ( .A(n9686), .B(n9685), .S(n14730), .Z(n9687) );
  AOI21_X1 U11460 ( .B1(n9689), .B2(n9688), .A(n9687), .ZN(n9718) );
  INV_X1 U11461 ( .A(n11734), .ZN(n10658) );
  OAI21_X1 U11462 ( .B1(n9710), .B2(n10658), .A(n12410), .ZN(n9691) );
  INV_X1 U11463 ( .A(n9718), .ZN(n9695) );
  INV_X1 U11464 ( .A(n9693), .ZN(n9694) );
  NAND2_X1 U11465 ( .A1(n9695), .A2(n9694), .ZN(n9716) );
  NAND2_X1 U11466 ( .A1(n9705), .A2(n9704), .ZN(n9698) );
  OR2_X1 U11467 ( .A1(n9701), .A2(n9700), .ZN(n9702) );
  INV_X1 U11468 ( .A(n14868), .ZN(n10434) );
  INV_X1 U11469 ( .A(n9707), .ZN(n9708) );
  INV_X1 U11470 ( .A(n10649), .ZN(n10484) );
  NAND4_X1 U11471 ( .A1(n15525), .A2(n10434), .A3(n14525), .A4(n10484), .ZN(
        n9709) );
  OAI211_X1 U11472 ( .C1(n9710), .C2(n11952), .A(n9709), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9715) );
  INV_X1 U11473 ( .A(n9711), .ZN(n9713) );
  NAND4_X1 U11474 ( .A1(n9713), .A2(n9712), .A3(n12414), .A4(n11375), .ZN(
        n9714) );
  AOI21_X1 U11475 ( .B1(n9718), .B2(n11430), .A(n9717), .ZN(n9719) );
  INV_X1 U11476 ( .A(n9719), .ZN(n9720) );
  NAND3_X1 U11477 ( .A1(n9723), .A2(n9722), .A3(n9721), .ZN(P2_U3328) );
  NOR2_X1 U11478 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), 
        .ZN(n9724) );
  NAND4_X1 U11479 ( .A1(n9728), .A2(n9727), .A3(n9781), .A4(n9782), .ZN(n9729)
         );
  INV_X2 U11480 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n15634) );
  INV_X1 U11481 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9845) );
  OAI21_X1 U11482 ( .B1(n9784), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9733) );
  XNOR2_X1 U11483 ( .A(n9733), .B(n9734), .ZN(n10264) );
  NAND2_X1 U11484 ( .A1(n9754), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U11485 ( .A1(n9743), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9744) );
  INV_X1 U11486 ( .A(n12255), .ZN(n9748) );
  MUX2_X1 U11487 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9745), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9746) );
  NAND2_X1 U11488 ( .A1(n9746), .A2(n9743), .ZN(n12198) );
  INV_X1 U11489 ( .A(n12198), .ZN(n9747) );
  INV_X1 U11490 ( .A(n10226), .ZN(n9863) );
  INV_X1 U11491 ( .A(n9749), .ZN(n9750) );
  NOR2_X4 U11492 ( .A1(n9751), .A2(n10308), .ZN(P3_U3897) );
  NAND2_X1 U11493 ( .A1(n9752), .A2(n8315), .ZN(n9753) );
  XNOR2_X1 U11494 ( .A(n9753), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15514) );
  MUX2_X1 U11495 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9759), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n9760) );
  NAND2_X1 U11496 ( .A1(n9761), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9762) );
  MUX2_X1 U11497 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9762), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9764) );
  NAND2_X1 U11498 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9936) );
  NOR2_X1 U11499 ( .A1(n9936), .A2(n9935), .ZN(n9959) );
  NAND2_X1 U11500 ( .A1(n9959), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9977) );
  INV_X1 U11501 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9976) );
  AND2_X1 U11502 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n9765) );
  NAND2_X1 U11503 ( .A1(n10057), .A2(n9765), .ZN(n10079) );
  INV_X1 U11504 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10078) );
  INV_X1 U11505 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9816) );
  NAND2_X1 U11506 ( .A1(n10163), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10180) );
  INV_X1 U11507 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10179) );
  INV_X1 U11508 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n15018) );
  NAND2_X1 U11509 ( .A1(n9791), .A2(n10232), .ZN(n9766) );
  INV_X1 U11510 ( .A(n10220), .ZN(n10221) );
  NAND2_X1 U11511 ( .A1(n9766), .A2(n10221), .ZN(n15261) );
  XNOR2_X2 U11512 ( .A(n9769), .B(n9768), .ZN(n12936) );
  INV_X1 U11513 ( .A(n9773), .ZN(n9771) );
  NOR2_X2 U11514 ( .A1(n12936), .A2(n9771), .ZN(n9871) );
  OR2_X1 U11515 ( .A1(n15261), .A2(n10183), .ZN(n9779) );
  INV_X1 U11516 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9776) );
  NOR2_X2 U11517 ( .A1(n12936), .A2(n9773), .ZN(n9870) );
  NAND2_X1 U11518 ( .A1(n12829), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9775) );
  AND2_X2 U11519 ( .A1(n12936), .A2(n9773), .ZN(n9840) );
  NAND2_X1 U11520 ( .A1(n12833), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9774) );
  OAI211_X1 U11521 ( .C1(n9893), .C2(n9776), .A(n9775), .B(n9774), .ZN(n9777)
         );
  INV_X1 U11522 ( .A(n9777), .ZN(n9778) );
  INV_X1 U11523 ( .A(n7404), .ZN(n10154) );
  OAI22_X1 U11524 ( .A1(n15439), .A2(n9958), .B1(n14969), .B2(n10154), .ZN(
        n9787) );
  NAND2_X1 U11525 ( .A1(n9823), .A2(n9781), .ZN(n9827) );
  XNOR2_X1 U11526 ( .A(n9787), .B(n14954), .ZN(n14885) );
  NAND2_X2 U11527 ( .A1(n12849), .A2(n11419), .ZN(n15974) );
  AND2_X2 U11528 ( .A1(n7219), .A2(n15974), .ZN(n9887) );
  INV_X1 U11529 ( .A(n9887), .ZN(n10153) );
  OAI22_X1 U11530 ( .A1(n15439), .A2(n10154), .B1(n14969), .B2(n10153), .ZN(
        n14884) );
  XNOR2_X1 U11531 ( .A(n14885), .B(n14884), .ZN(n10218) );
  OR2_X1 U11532 ( .A1(n11418), .A2(n9846), .ZN(n9789) );
  INV_X1 U11533 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11420) );
  OR2_X1 U11534 ( .A1(n9902), .A2(n11420), .ZN(n9788) );
  OR2_X1 U11535 ( .A1(n9804), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9790) );
  NAND2_X1 U11536 ( .A1(n9791), .A2(n9790), .ZN(n15270) );
  OR2_X1 U11537 ( .A1(n15270), .A2(n10183), .ZN(n9797) );
  INV_X1 U11538 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9794) );
  NAND2_X1 U11539 ( .A1(n12829), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9793) );
  NAND2_X1 U11540 ( .A1(n9840), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9792) );
  OAI211_X1 U11541 ( .C1(n9893), .C2(n9794), .A(n9793), .B(n9792), .ZN(n9795)
         );
  INV_X1 U11542 ( .A(n9795), .ZN(n9796) );
  AOI22_X1 U11543 ( .A1(n15444), .A2(n9798), .B1(n14953), .B2(n15259), .ZN(
        n10196) );
  INV_X1 U11544 ( .A(n10196), .ZN(n10198) );
  NAND2_X1 U11545 ( .A1(n15444), .A2(n14905), .ZN(n9800) );
  NAND2_X1 U11546 ( .A1(n15259), .A2(n7404), .ZN(n9799) );
  NAND2_X1 U11547 ( .A1(n9800), .A2(n9799), .ZN(n9801) );
  XNOR2_X1 U11548 ( .A(n9801), .B(n14954), .ZN(n10197) );
  NAND2_X1 U11549 ( .A1(n11324), .A2(n7232), .ZN(n9803) );
  OR2_X1 U11550 ( .A1(n9902), .A2(n11325), .ZN(n9802) );
  AND2_X1 U11551 ( .A1(n10182), .A2(n15018), .ZN(n9805) );
  OR2_X1 U11552 ( .A1(n9805), .A2(n9804), .ZN(n15295) );
  AOI22_X1 U11553 ( .A1(n12833), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n12829), 
        .B2(P1_REG2_REG_20__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U11554 ( .A1(n12834), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9806) );
  OAI211_X1 U11555 ( .C1(n15295), .C2(n10183), .A(n9807), .B(n9806), .ZN(
        n15061) );
  AND2_X1 U11556 ( .A1(n15061), .A2(n14953), .ZN(n9808) );
  AOI21_X1 U11557 ( .B1(n15299), .B2(n7404), .A(n9808), .ZN(n10193) );
  INV_X1 U11558 ( .A(n10193), .ZN(n10195) );
  NAND2_X1 U11559 ( .A1(n15299), .A2(n14905), .ZN(n9810) );
  NAND2_X1 U11560 ( .A1(n15061), .A2(n7404), .ZN(n9809) );
  NAND2_X1 U11561 ( .A1(n9810), .A2(n9809), .ZN(n9811) );
  XNOR2_X1 U11562 ( .A(n9811), .B(n14954), .ZN(n10194) );
  NAND2_X1 U11563 ( .A1(n11037), .A2(n7232), .ZN(n9815) );
  NAND2_X1 U11564 ( .A1(n9827), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9812) );
  MUX2_X1 U11565 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9812), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n9813) );
  AND2_X1 U11566 ( .A1(n9813), .A2(n7253), .ZN(n15124) );
  AOI22_X1 U11567 ( .A1(n10176), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10175), 
        .B2(n15124), .ZN(n9814) );
  AND2_X1 U11568 ( .A1(n9834), .A2(n9816), .ZN(n9817) );
  OR2_X1 U11569 ( .A1(n9817), .A2(n10163), .ZN(n15342) );
  NAND2_X1 U11570 ( .A1(n12834), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U11571 ( .A1(n12833), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9818) );
  AND2_X1 U11572 ( .A1(n9819), .A2(n9818), .ZN(n9821) );
  NAND2_X1 U11573 ( .A1(n12829), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9820) );
  OAI211_X1 U11574 ( .C1(n15342), .C2(n10183), .A(n9821), .B(n9820), .ZN(
        n15064) );
  AOI22_X1 U11575 ( .A1(n15474), .A2(n14905), .B1(n7404), .B2(n15064), .ZN(
        n9822) );
  XOR2_X1 U11576 ( .A(n14954), .B(n9822), .Z(n14994) );
  INV_X1 U11577 ( .A(n14994), .ZN(n10159) );
  INV_X1 U11578 ( .A(n15064), .ZN(n15360) );
  OAI22_X1 U11579 ( .A1(n15345), .A2(n10154), .B1(n15360), .B2(n10153), .ZN(
        n10158) );
  INV_X1 U11580 ( .A(n10158), .ZN(n14993) );
  NAND2_X1 U11581 ( .A1(n10922), .A2(n7232), .ZN(n9831) );
  INV_X1 U11582 ( .A(n9823), .ZN(n9824) );
  NAND2_X1 U11583 ( .A1(n9824), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9825) );
  MUX2_X1 U11584 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9825), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9826) );
  INV_X1 U11585 ( .A(n9826), .ZN(n9829) );
  INV_X1 U11586 ( .A(n9827), .ZN(n9828) );
  NOR2_X1 U11587 ( .A1(n9829), .A2(n9828), .ZN(n15106) );
  AOI22_X1 U11588 ( .A1(n10176), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n10175), 
        .B2(n15106), .ZN(n9830) );
  NAND2_X1 U11589 ( .A1(n12834), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U11590 ( .A1(n9840), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U11591 ( .A1(n10144), .A2(n9832), .ZN(n9833) );
  AND2_X1 U11592 ( .A1(n9834), .A2(n9833), .ZN(n15361) );
  NAND2_X1 U11593 ( .A1(n7213), .A2(n15361), .ZN(n9836) );
  NAND2_X1 U11594 ( .A1(n12829), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9835) );
  NAND4_X1 U11595 ( .A1(n9838), .A2(n9837), .A3(n9836), .A4(n9835), .ZN(n15375) );
  AOI22_X1 U11596 ( .A1(n16133), .A2(n7404), .B1(n14953), .B2(n15375), .ZN(
        n10157) );
  AOI22_X1 U11597 ( .A1(n16133), .A2(n14905), .B1(n7404), .B2(n15375), .ZN(
        n9839) );
  XNOR2_X1 U11598 ( .A(n9839), .B(n14954), .ZN(n10156) );
  NAND2_X1 U11599 ( .A1(n9872), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9844) );
  NAND2_X1 U11600 ( .A1(n9840), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9843) );
  NAND2_X1 U11601 ( .A1(n9871), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U11602 ( .A1(n9870), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9841) );
  NAND2_X1 U11603 ( .A1(n10902), .A2(n9798), .ZN(n9848) );
  NAND2_X1 U11604 ( .A1(n15634), .A2(n9845), .ZN(n9878) );
  NAND2_X1 U11605 ( .A1(n12674), .A2(n7219), .ZN(n9847) );
  AND2_X1 U11606 ( .A1(n12674), .A2(n9798), .ZN(n9850) );
  NAND2_X1 U11607 ( .A1(n9852), .A2(n9851), .ZN(n9869) );
  NAND2_X1 U11608 ( .A1(n9853), .A2(n9869), .ZN(n10791) );
  INV_X1 U11609 ( .A(n10791), .ZN(n9868) );
  NAND2_X1 U11610 ( .A1(n9871), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9857) );
  NAND2_X1 U11611 ( .A1(n9840), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U11612 ( .A1(n9872), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U11613 ( .A1(n10907), .A2(n9798), .ZN(n9862) );
  NOR2_X1 U11614 ( .A1(n10252), .A2(n10253), .ZN(n9859) );
  XNOR2_X1 U11615 ( .A(n9859), .B(n9858), .ZN(n15515) );
  MUX2_X1 U11616 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15515), .S(n7230), .Z(n15878)
         );
  INV_X1 U11617 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15880) );
  NOR2_X1 U11618 ( .A1(n10226), .A2(n15880), .ZN(n9860) );
  AOI21_X1 U11619 ( .B1(n15878), .B2(n7219), .A(n9860), .ZN(n9861) );
  NAND2_X1 U11620 ( .A1(n10907), .A2(n9887), .ZN(n9865) );
  AOI22_X1 U11621 ( .A1(n15878), .A2(n9798), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n9863), .ZN(n9864) );
  INV_X1 U11622 ( .A(n10794), .ZN(n9867) );
  NAND2_X1 U11623 ( .A1(n9870), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U11624 ( .A1(n9872), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U11625 ( .A1(n15074), .A2(n9798), .ZN(n9885) );
  NAND2_X1 U11626 ( .A1(n9878), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9877) );
  MUX2_X1 U11627 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9877), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n9881) );
  INV_X1 U11628 ( .A(n9878), .ZN(n9880) );
  NAND2_X1 U11629 ( .A1(n9880), .A2(n9879), .ZN(n9993) );
  NAND2_X1 U11630 ( .A1(n9881), .A2(n9993), .ZN(n10351) );
  OR2_X1 U11631 ( .A1(n7236), .A2(n10243), .ZN(n9882) );
  OAI211_X2 U11632 ( .C1(n7421), .C2(n10351), .A(n9883), .B(n9882), .ZN(n12690) );
  NAND2_X1 U11633 ( .A1(n12690), .A2(n7219), .ZN(n9884) );
  NAND2_X1 U11634 ( .A1(n9885), .A2(n9884), .ZN(n9886) );
  AND2_X1 U11635 ( .A1(n12690), .A2(n9798), .ZN(n9888) );
  AOI21_X1 U11636 ( .B1(n15074), .B2(n9887), .A(n9888), .ZN(n9890) );
  INV_X1 U11637 ( .A(n9889), .ZN(n9891) );
  NAND2_X1 U11638 ( .A1(n9891), .A2(n9890), .ZN(n9892) );
  NAND2_X1 U11639 ( .A1(n9840), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9898) );
  NAND2_X1 U11640 ( .A1(n9872), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9897) );
  NAND2_X1 U11641 ( .A1(n9870), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9896) );
  INV_X1 U11642 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9912) );
  NAND2_X1 U11643 ( .A1(n7211), .A2(n9912), .ZN(n9895) );
  NAND4_X2 U11644 ( .A1(n9898), .A2(n9897), .A3(n9896), .A4(n9895), .ZN(n15073) );
  NAND2_X1 U11645 ( .A1(n15073), .A2(n9798), .ZN(n9905) );
  NAND2_X1 U11646 ( .A1(n9993), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9899) );
  MUX2_X1 U11647 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9899), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9900) );
  NAND2_X1 U11648 ( .A1(n9900), .A2(n9920), .ZN(n10390) );
  OR2_X1 U11649 ( .A1(n9902), .A2(n10244), .ZN(n9903) );
  NAND2_X1 U11650 ( .A1(n15906), .A2(n7219), .ZN(n9904) );
  NAND2_X1 U11651 ( .A1(n9905), .A2(n9904), .ZN(n9906) );
  XNOR2_X1 U11652 ( .A(n9906), .B(n14954), .ZN(n9910) );
  AND2_X1 U11653 ( .A1(n15906), .A2(n7404), .ZN(n9907) );
  AOI21_X1 U11654 ( .B1(n15073), .B2(n14953), .A(n9907), .ZN(n9908) );
  XNOR2_X1 U11655 ( .A(n9910), .B(n9908), .ZN(n14938) );
  INV_X1 U11656 ( .A(n9908), .ZN(n9909) );
  NAND2_X1 U11657 ( .A1(n9910), .A2(n9909), .ZN(n9930) );
  NAND2_X1 U11658 ( .A1(n12834), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9918) );
  NAND2_X1 U11659 ( .A1(n12833), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9917) );
  INV_X1 U11660 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9911) );
  NAND2_X1 U11661 ( .A1(n9912), .A2(n9911), .ZN(n9913) );
  AND2_X1 U11662 ( .A1(n9913), .A2(n9936), .ZN(n11354) );
  INV_X1 U11663 ( .A(n11354), .ZN(n9914) );
  NAND2_X1 U11664 ( .A1(n9870), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9915) );
  NAND2_X1 U11665 ( .A1(n9920), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9919) );
  MUX2_X1 U11666 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9919), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n9923) );
  INV_X1 U11667 ( .A(n9920), .ZN(n9922) );
  INV_X1 U11668 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9921) );
  NAND2_X1 U11669 ( .A1(n9922), .A2(n9921), .ZN(n9944) );
  NAND2_X1 U11670 ( .A1(n9923), .A2(n9944), .ZN(n10356) );
  NAND2_X1 U11671 ( .A1(n7232), .A2(n10241), .ZN(n9925) );
  OR2_X1 U11672 ( .A1(n9902), .A2(n10242), .ZN(n9924) );
  OAI211_X1 U11673 ( .C1(n7421), .C2(n10356), .A(n9925), .B(n9924), .ZN(n12703) );
  AOI22_X1 U11674 ( .A1(n15072), .A2(n14953), .B1(n7404), .B2(n12703), .ZN(
        n9931) );
  AND2_X1 U11675 ( .A1(n9930), .A2(n9931), .ZN(n9926) );
  NAND2_X1 U11676 ( .A1(n15072), .A2(n7404), .ZN(n9928) );
  NAND2_X1 U11677 ( .A1(n12703), .A2(n14905), .ZN(n9927) );
  NAND2_X1 U11678 ( .A1(n9928), .A2(n9927), .ZN(n9929) );
  NAND2_X1 U11679 ( .A1(n11283), .A2(n11285), .ZN(n9934) );
  NAND2_X1 U11680 ( .A1(n14936), .A2(n9930), .ZN(n9933) );
  INV_X1 U11681 ( .A(n9931), .ZN(n9932) );
  NAND2_X1 U11682 ( .A1(n9933), .A2(n9932), .ZN(n11282) );
  NAND2_X1 U11683 ( .A1(n9934), .A2(n11282), .ZN(n11295) );
  NAND2_X1 U11684 ( .A1(n12833), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9942) );
  NAND2_X1 U11685 ( .A1(n9870), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9941) );
  AND2_X1 U11686 ( .A1(n9936), .A2(n9935), .ZN(n9937) );
  NOR2_X1 U11687 ( .A1(n9959), .A2(n9937), .ZN(n11571) );
  INV_X1 U11688 ( .A(n11571), .ZN(n9938) );
  NAND2_X1 U11689 ( .A1(n12834), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9939) );
  NAND4_X1 U11690 ( .A1(n9942), .A2(n9941), .A3(n9940), .A4(n9939), .ZN(n15071) );
  NAND2_X1 U11691 ( .A1(n15071), .A2(n7404), .ZN(n9949) );
  NAND2_X1 U11692 ( .A1(n10250), .A2(n7232), .ZN(n9947) );
  NAND2_X1 U11693 ( .A1(n9944), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9943) );
  MUX2_X1 U11694 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9943), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9945) );
  AOI22_X1 U11695 ( .A1(n10176), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10175), 
        .B2(n10368), .ZN(n9946) );
  NAND2_X1 U11696 ( .A1(n9947), .A2(n9946), .ZN(n12709) );
  NAND2_X1 U11697 ( .A1(n12709), .A2(n14905), .ZN(n9948) );
  NAND2_X1 U11698 ( .A1(n9949), .A2(n9948), .ZN(n9950) );
  XNOR2_X1 U11699 ( .A(n9950), .B(n10188), .ZN(n9951) );
  AOI22_X1 U11700 ( .A1(n15071), .A2(n14953), .B1(n12709), .B2(n7404), .ZN(
        n9952) );
  INV_X1 U11701 ( .A(n9951), .ZN(n9954) );
  INV_X1 U11702 ( .A(n9952), .ZN(n9953) );
  NAND2_X1 U11703 ( .A1(n9954), .A2(n9953), .ZN(n11293) );
  NAND2_X1 U11704 ( .A1(n10269), .A2(n7232), .ZN(n9957) );
  NAND2_X1 U11705 ( .A1(n9972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9955) );
  XNOR2_X1 U11706 ( .A(n9955), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U11707 ( .A1(n10176), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10175), 
        .B2(n10402), .ZN(n9956) );
  NAND2_X1 U11708 ( .A1(n12716), .A2(n14905), .ZN(n9966) );
  NAND2_X1 U11709 ( .A1(n12834), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U11710 ( .A1(n12833), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9963) );
  OR2_X1 U11711 ( .A1(n9959), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9960) );
  AND2_X1 U11712 ( .A1(n9977), .A2(n9960), .ZN(n11607) );
  NAND2_X1 U11713 ( .A1(n7213), .A2(n11607), .ZN(n9962) );
  NAND2_X1 U11714 ( .A1(n12829), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9961) );
  NAND4_X1 U11715 ( .A1(n9964), .A2(n9963), .A3(n9962), .A4(n9961), .ZN(n15070) );
  NAND2_X1 U11716 ( .A1(n15070), .A2(n7404), .ZN(n9965) );
  NAND2_X1 U11717 ( .A1(n9966), .A2(n9965), .ZN(n9967) );
  XNOR2_X1 U11718 ( .A(n9967), .B(n14954), .ZN(n9968) );
  AOI22_X1 U11719 ( .A1(n12716), .A2(n7404), .B1(n15070), .B2(n14953), .ZN(
        n9969) );
  XNOR2_X1 U11720 ( .A(n9968), .B(n9969), .ZN(n11378) );
  INV_X1 U11721 ( .A(n9968), .ZN(n9970) );
  OR2_X1 U11722 ( .A1(n9970), .A2(n9969), .ZN(n9971) );
  NAND2_X1 U11723 ( .A1(n10276), .A2(n7232), .ZN(n9975) );
  OAI21_X1 U11724 ( .B1(n9972), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9973) );
  XNOR2_X1 U11725 ( .A(n9973), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U11726 ( .A1(n10176), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10175), 
        .B2(n10614), .ZN(n9974) );
  NAND2_X1 U11727 ( .A1(n12725), .A2(n14905), .ZN(n9984) );
  NAND2_X1 U11728 ( .A1(n12834), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U11729 ( .A1(n12833), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U11730 ( .A1(n9977), .A2(n9976), .ZN(n9978) );
  AND2_X1 U11731 ( .A1(n10000), .A2(n9978), .ZN(n11460) );
  NAND2_X1 U11732 ( .A1(n7213), .A2(n11460), .ZN(n9980) );
  NAND2_X1 U11733 ( .A1(n12829), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9979) );
  NAND4_X1 U11734 ( .A1(n9982), .A2(n9981), .A3(n9980), .A4(n9979), .ZN(n15069) );
  NAND2_X1 U11735 ( .A1(n15069), .A2(n7404), .ZN(n9983) );
  NAND2_X1 U11736 ( .A1(n9984), .A2(n9983), .ZN(n9985) );
  XNOR2_X1 U11737 ( .A(n9985), .B(n14954), .ZN(n9989) );
  AND2_X1 U11738 ( .A1(n15069), .A2(n14953), .ZN(n9986) );
  AOI21_X1 U11739 ( .B1(n12725), .B2(n7404), .A(n9986), .ZN(n9987) );
  XNOR2_X1 U11740 ( .A(n9989), .B(n9987), .ZN(n11455) );
  INV_X1 U11741 ( .A(n9987), .ZN(n9988) );
  NAND2_X1 U11742 ( .A1(n9989), .A2(n9988), .ZN(n9990) );
  NAND2_X1 U11743 ( .A1(n10297), .A2(n7232), .ZN(n9998) );
  INV_X1 U11744 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9991) );
  NAND2_X1 U11745 ( .A1(n9992), .A2(n9991), .ZN(n9994) );
  OAI21_X1 U11746 ( .B1(n9994), .B2(n9993), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9995) );
  MUX2_X1 U11747 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9995), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n9996) );
  AND2_X1 U11748 ( .A1(n9996), .A2(n10035), .ZN(n11159) );
  AOI22_X1 U11749 ( .A1(n10176), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10175), 
        .B2(n11159), .ZN(n9997) );
  NAND2_X1 U11750 ( .A1(n15992), .A2(n14905), .ZN(n10007) );
  NAND2_X1 U11751 ( .A1(n12833), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10005) );
  NAND2_X1 U11752 ( .A1(n12829), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10004) );
  NAND2_X1 U11753 ( .A1(n10000), .A2(n9999), .ZN(n10001) );
  NAND2_X1 U11754 ( .A1(n7212), .A2(n7252), .ZN(n10003) );
  NAND2_X1 U11755 ( .A1(n12834), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10002) );
  NAND4_X1 U11756 ( .A1(n10005), .A2(n10004), .A3(n10003), .A4(n10002), .ZN(
        n15068) );
  NAND2_X1 U11757 ( .A1(n15068), .A2(n7404), .ZN(n10006) );
  NAND2_X1 U11758 ( .A1(n10007), .A2(n10006), .ZN(n10008) );
  XNOR2_X1 U11759 ( .A(n10008), .B(n10188), .ZN(n10012) );
  AND2_X1 U11760 ( .A1(n15068), .A2(n14953), .ZN(n10009) );
  AOI21_X1 U11761 ( .B1(n15992), .B2(n7404), .A(n10009), .ZN(n10011) );
  XNOR2_X1 U11762 ( .A(n10012), .B(n10011), .ZN(n11667) );
  NAND2_X1 U11763 ( .A1(n10012), .A2(n10011), .ZN(n10013) );
  INV_X1 U11764 ( .A(n11847), .ZN(n10029) );
  NAND2_X1 U11765 ( .A1(n10380), .A2(n7232), .ZN(n10016) );
  NAND2_X1 U11766 ( .A1(n10035), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10014) );
  XNOR2_X1 U11767 ( .A(n10014), .B(P1_IR_REG_9__SCAN_IN), .ZN(n15088) );
  AOI22_X1 U11768 ( .A1(n10176), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10175), 
        .B2(n15088), .ZN(n10015) );
  NAND2_X1 U11769 ( .A1(n16019), .A2(n14905), .ZN(n10025) );
  NAND2_X1 U11770 ( .A1(n12834), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U11771 ( .A1(n12833), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10022) );
  AND2_X1 U11772 ( .A1(n10018), .A2(n10017), .ZN(n10019) );
  NOR2_X1 U11773 ( .A1(n10057), .A2(n10019), .ZN(n11922) );
  NAND2_X1 U11774 ( .A1(n7212), .A2(n11922), .ZN(n10021) );
  NAND2_X1 U11775 ( .A1(n12829), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10020) );
  NAND4_X1 U11776 ( .A1(n10023), .A2(n10022), .A3(n10021), .A4(n10020), .ZN(
        n16029) );
  NAND2_X1 U11777 ( .A1(n16029), .A2(n7404), .ZN(n10024) );
  NAND2_X1 U11778 ( .A1(n10025), .A2(n10024), .ZN(n10026) );
  XNOR2_X1 U11779 ( .A(n10026), .B(n10188), .ZN(n10030) );
  AND2_X1 U11780 ( .A1(n16029), .A2(n14953), .ZN(n10027) );
  AOI21_X1 U11781 ( .B1(n16019), .B2(n7404), .A(n10027), .ZN(n10031) );
  XNOR2_X1 U11782 ( .A(n10030), .B(n10031), .ZN(n11846) );
  INV_X1 U11783 ( .A(n10030), .ZN(n10033) );
  INV_X1 U11784 ( .A(n10031), .ZN(n10032) );
  NAND2_X1 U11785 ( .A1(n10033), .A2(n10032), .ZN(n10034) );
  OR2_X1 U11786 ( .A1(n10035), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n10038) );
  NAND2_X1 U11787 ( .A1(n10038), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10036) );
  MUX2_X1 U11788 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10036), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n10037) );
  INV_X1 U11789 ( .A(n10037), .ZN(n10039) );
  NOR2_X1 U11790 ( .A1(n10039), .A2(n10074), .ZN(n11236) );
  AOI22_X1 U11791 ( .A1(n10176), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10175), 
        .B2(n11236), .ZN(n10040) );
  NAND2_X1 U11792 ( .A1(n16031), .A2(n14905), .ZN(n10047) );
  NAND2_X1 U11793 ( .A1(n12834), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10045) );
  NAND2_X1 U11794 ( .A1(n12833), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10044) );
  INV_X1 U11795 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10041) );
  XNOR2_X1 U11796 ( .A(n10057), .B(n10041), .ZN(n12081) );
  NAND2_X1 U11797 ( .A1(n7213), .A2(n12081), .ZN(n10043) );
  NAND2_X1 U11798 ( .A1(n12829), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10042) );
  NAND4_X1 U11799 ( .A1(n10045), .A2(n10044), .A3(n10043), .A4(n10042), .ZN(
        n15067) );
  NAND2_X1 U11800 ( .A1(n15067), .A2(n7404), .ZN(n10046) );
  NAND2_X1 U11801 ( .A1(n10047), .A2(n10046), .ZN(n10048) );
  XNOR2_X1 U11802 ( .A(n10048), .B(n14954), .ZN(n10052) );
  AND2_X1 U11803 ( .A1(n15067), .A2(n14953), .ZN(n10049) );
  AOI21_X1 U11804 ( .B1(n16031), .B2(n7404), .A(n10049), .ZN(n10050) );
  XNOR2_X1 U11805 ( .A(n10052), .B(n10050), .ZN(n12079) );
  NAND2_X1 U11806 ( .A1(n12080), .A2(n12079), .ZN(n12078) );
  INV_X1 U11807 ( .A(n10050), .ZN(n10051) );
  NAND2_X1 U11808 ( .A1(n10052), .A2(n10051), .ZN(n10053) );
  INV_X1 U11809 ( .A(n12260), .ZN(n10070) );
  NAND2_X1 U11810 ( .A1(n10394), .A2(n7232), .ZN(n10056) );
  INV_X1 U11811 ( .A(n10074), .ZN(n10138) );
  NAND2_X1 U11812 ( .A1(n10138), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10054) );
  XNOR2_X1 U11813 ( .A(n10054), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U11814 ( .A1(n10176), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10175), 
        .B2(n11464), .ZN(n10055) );
  NAND2_X1 U11815 ( .A1(n12744), .A2(n14905), .ZN(n10066) );
  NAND2_X1 U11816 ( .A1(n12834), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10064) );
  NAND2_X1 U11817 ( .A1(n12833), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U11818 ( .A1(n10057), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10059) );
  INV_X1 U11819 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10058) );
  NAND2_X1 U11820 ( .A1(n10059), .A2(n10058), .ZN(n10060) );
  AND2_X1 U11821 ( .A1(n10060), .A2(n10079), .ZN(n12262) );
  NAND2_X1 U11822 ( .A1(n7213), .A2(n12262), .ZN(n10062) );
  NAND2_X1 U11823 ( .A1(n12829), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10061) );
  NAND4_X1 U11824 ( .A1(n10064), .A2(n10063), .A3(n10062), .A4(n10061), .ZN(
        n15066) );
  NAND2_X1 U11825 ( .A1(n15066), .A2(n7404), .ZN(n10065) );
  NAND2_X1 U11826 ( .A1(n10066), .A2(n10065), .ZN(n10067) );
  XNOR2_X1 U11827 ( .A(n10067), .B(n10188), .ZN(n10072) );
  AND2_X1 U11828 ( .A1(n15066), .A2(n14953), .ZN(n10068) );
  AOI21_X1 U11829 ( .B1(n12744), .B2(n7404), .A(n10068), .ZN(n10071) );
  XNOR2_X1 U11830 ( .A(n10072), .B(n10071), .ZN(n12261) );
  INV_X1 U11831 ( .A(n12261), .ZN(n10069) );
  NAND2_X1 U11832 ( .A1(n10072), .A2(n10071), .ZN(n10073) );
  NAND2_X1 U11833 ( .A1(n10419), .A2(n7232), .ZN(n10077) );
  NAND2_X1 U11834 ( .A1(n10074), .A2(n10136), .ZN(n10075) );
  NAND2_X1 U11835 ( .A1(n10075), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10095) );
  XNOR2_X1 U11836 ( .A(n10095), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U11837 ( .A1(n10176), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10175), 
        .B2(n11474), .ZN(n10076) );
  NAND2_X1 U11838 ( .A1(n12747), .A2(n14905), .ZN(n10086) );
  NAND2_X1 U11839 ( .A1(n12834), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10084) );
  NAND2_X1 U11840 ( .A1(n9840), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U11841 ( .A1(n10079), .A2(n10078), .ZN(n10080) );
  AND2_X1 U11842 ( .A1(n10102), .A2(n10080), .ZN(n12549) );
  NAND2_X1 U11843 ( .A1(n7213), .A2(n12549), .ZN(n10082) );
  NAND2_X1 U11844 ( .A1(n12829), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10081) );
  NAND4_X1 U11845 ( .A1(n10084), .A2(n10083), .A3(n10082), .A4(n10081), .ZN(
        n15065) );
  NAND2_X1 U11846 ( .A1(n15065), .A2(n7404), .ZN(n10085) );
  NAND2_X1 U11847 ( .A1(n10086), .A2(n10085), .ZN(n10087) );
  XNOR2_X1 U11848 ( .A(n10087), .B(n10188), .ZN(n10090) );
  AND2_X1 U11849 ( .A1(n15065), .A2(n14953), .ZN(n10088) );
  AOI21_X1 U11850 ( .B1(n12747), .B2(n7404), .A(n10088), .ZN(n10091) );
  XNOR2_X1 U11851 ( .A(n10090), .B(n10091), .ZN(n12556) );
  INV_X1 U11852 ( .A(n10090), .ZN(n10093) );
  INV_X1 U11853 ( .A(n10091), .ZN(n10092) );
  NAND2_X1 U11854 ( .A1(n10093), .A2(n10092), .ZN(n10094) );
  NAND2_X1 U11855 ( .A1(n10603), .A2(n7232), .ZN(n10100) );
  INV_X1 U11856 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10134) );
  NAND2_X1 U11857 ( .A1(n10095), .A2(n10134), .ZN(n10096) );
  NAND2_X1 U11858 ( .A1(n10096), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10097) );
  INV_X1 U11859 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10135) );
  NAND2_X1 U11860 ( .A1(n10097), .A2(n10135), .ZN(n10116) );
  OR2_X1 U11861 ( .A1(n10097), .A2(n10135), .ZN(n10098) );
  AOI22_X1 U11862 ( .A1(n10176), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n10175), 
        .B2(n11837), .ZN(n10099) );
  NAND2_X1 U11863 ( .A1(n12751), .A2(n14905), .ZN(n10109) );
  NAND2_X1 U11864 ( .A1(n12833), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10107) );
  NAND2_X1 U11865 ( .A1(n12834), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10106) );
  AND2_X1 U11866 ( .A1(n10102), .A2(n10101), .ZN(n10103) );
  NOR2_X1 U11867 ( .A1(n10120), .A2(n10103), .ZN(n12379) );
  NAND2_X1 U11868 ( .A1(n7213), .A2(n12379), .ZN(n10105) );
  NAND2_X1 U11869 ( .A1(n12829), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10104) );
  NAND4_X1 U11870 ( .A1(n10107), .A2(n10106), .A3(n10105), .A4(n10104), .ZN(
        n16086) );
  NAND2_X1 U11871 ( .A1(n16086), .A2(n7404), .ZN(n10108) );
  NAND2_X1 U11872 ( .A1(n10109), .A2(n10108), .ZN(n10110) );
  XNOR2_X1 U11873 ( .A(n10110), .B(n14954), .ZN(n10114) );
  AND2_X1 U11874 ( .A1(n16086), .A2(n14953), .ZN(n10111) );
  AOI21_X1 U11875 ( .B1(n12751), .B2(n7404), .A(n10111), .ZN(n10112) );
  XNOR2_X1 U11876 ( .A(n10114), .B(n10112), .ZN(n12509) );
  INV_X1 U11877 ( .A(n10112), .ZN(n10113) );
  NAND2_X1 U11878 ( .A1(n10114), .A2(n10113), .ZN(n10115) );
  NAND2_X1 U11879 ( .A1(n10926), .A2(n7232), .ZN(n10119) );
  NAND2_X1 U11880 ( .A1(n10116), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10117) );
  XNOR2_X1 U11881 ( .A(n10117), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U11882 ( .A1(n10176), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n10175), 
        .B2(n12488), .ZN(n10118) );
  NAND2_X1 U11883 ( .A1(n12755), .A2(n14905), .ZN(n10127) );
  NAND2_X1 U11884 ( .A1(n12833), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U11885 ( .A1(n12834), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n10124) );
  NAND2_X1 U11886 ( .A1(n12829), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10123) );
  NOR2_X1 U11887 ( .A1(n10120), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10121) );
  OR2_X1 U11888 ( .A1(n10142), .A2(n10121), .ZN(n16097) );
  INV_X1 U11889 ( .A(n16097), .ZN(n12439) );
  NAND2_X1 U11890 ( .A1(n7212), .A2(n12439), .ZN(n10122) );
  NAND4_X1 U11891 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n15374) );
  NAND2_X1 U11892 ( .A1(n15374), .A2(n7404), .ZN(n10126) );
  NAND2_X1 U11893 ( .A1(n10127), .A2(n10126), .ZN(n10128) );
  XNOR2_X1 U11894 ( .A(n10128), .B(n14954), .ZN(n10130) );
  AND2_X1 U11895 ( .A1(n15374), .A2(n14953), .ZN(n10129) );
  AOI21_X1 U11896 ( .B1(n12755), .B2(n7404), .A(n10129), .ZN(n10131) );
  XNOR2_X1 U11897 ( .A(n10130), .B(n10131), .ZN(n16085) );
  INV_X1 U11898 ( .A(n10130), .ZN(n10132) );
  NAND2_X1 U11899 ( .A1(n11012), .A2(n7232), .ZN(n10141) );
  INV_X1 U11900 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10133) );
  NAND4_X1 U11901 ( .A1(n10136), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(
        n10137) );
  OAI21_X1 U11902 ( .B1(n10138), .B2(n10137), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10139) );
  XNOR2_X1 U11903 ( .A(n10139), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U11904 ( .A1(n10176), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10175), 
        .B2(n12483), .ZN(n10140) );
  NAND2_X1 U11905 ( .A1(n12834), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n10148) );
  NAND2_X1 U11906 ( .A1(n12833), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n10147) );
  OR2_X1 U11907 ( .A1(n10142), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10143) );
  AND2_X1 U11908 ( .A1(n10144), .A2(n10143), .ZN(n15048) );
  NAND2_X1 U11909 ( .A1(n7212), .A2(n15048), .ZN(n10146) );
  NAND2_X1 U11910 ( .A1(n12829), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n10145) );
  NAND4_X1 U11911 ( .A1(n10148), .A2(n10147), .A3(n10146), .A4(n10145), .ZN(
        n16088) );
  AOI22_X1 U11912 ( .A1(n15386), .A2(n14905), .B1(n7404), .B2(n16088), .ZN(
        n10149) );
  XOR2_X1 U11913 ( .A(n14954), .B(n10149), .Z(n10151) );
  INV_X1 U11914 ( .A(n10151), .ZN(n10150) );
  INV_X1 U11915 ( .A(n15386), .ZN(n16124) );
  INV_X1 U11916 ( .A(n16088), .ZN(n15358) );
  OAI22_X1 U11917 ( .A1(n16124), .A2(n10154), .B1(n15358), .B2(n10153), .ZN(
        n15047) );
  XNOR2_X1 U11918 ( .A(n10156), .B(n10157), .ZN(n14986) );
  NAND2_X1 U11919 ( .A1(n11320), .A2(n7232), .ZN(n10162) );
  NAND2_X1 U11920 ( .A1(n7253), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10160) );
  XNOR2_X1 U11921 ( .A(n10160), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15138) );
  AOI22_X1 U11922 ( .A1(n10176), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10175), 
        .B2(n15138), .ZN(n10161) );
  NAND2_X1 U11923 ( .A1(n15466), .A2(n14905), .ZN(n10168) );
  OR2_X1 U11924 ( .A1(n10163), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10164) );
  NAND2_X1 U11925 ( .A1(n10180), .A2(n10164), .ZN(n15328) );
  AOI22_X1 U11926 ( .A1(n12834), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n12833), 
        .B2(P1_REG1_REG_18__SCAN_IN), .ZN(n10166) );
  NAND2_X1 U11927 ( .A1(n12829), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n10165) );
  OAI211_X1 U11928 ( .C1(n15328), .C2(n10183), .A(n10166), .B(n10165), .ZN(
        n15063) );
  NAND2_X1 U11929 ( .A1(n15063), .A2(n7404), .ZN(n10167) );
  NAND2_X1 U11930 ( .A1(n10168), .A2(n10167), .ZN(n10169) );
  XNOR2_X1 U11931 ( .A(n10169), .B(n10188), .ZN(n10172) );
  AND2_X1 U11932 ( .A1(n15063), .A2(n14953), .ZN(n10170) );
  AOI21_X1 U11933 ( .B1(n15466), .B2(n7404), .A(n10170), .ZN(n10171) );
  NAND2_X1 U11934 ( .A1(n10172), .A2(n10171), .ZN(n10173) );
  OAI21_X1 U11935 ( .B1(n10172), .B2(n10171), .A(n10173), .ZN(n15025) );
  INV_X1 U11936 ( .A(n10173), .ZN(n10174) );
  NAND2_X1 U11937 ( .A1(n11421), .A2(n7232), .ZN(n10178) );
  AOI22_X1 U11938 ( .A1(n10176), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10175), 
        .B2(n15150), .ZN(n10177) );
  NAND2_X1 U11939 ( .A1(n15460), .A2(n14905), .ZN(n10187) );
  INV_X1 U11940 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n15312) );
  NAND2_X1 U11941 ( .A1(n10180), .A2(n10179), .ZN(n10181) );
  NAND2_X1 U11942 ( .A1(n10182), .A2(n10181), .ZN(n15311) );
  OR2_X1 U11943 ( .A1(n15311), .A2(n10183), .ZN(n10185) );
  AOI22_X1 U11944 ( .A1(n12834), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n9840), 
        .B2(P1_REG1_REG_19__SCAN_IN), .ZN(n10184) );
  OAI211_X1 U11945 ( .C1(n9772), .C2(n15312), .A(n10185), .B(n10184), .ZN(
        n15062) );
  NAND2_X1 U11946 ( .A1(n15062), .A2(n7404), .ZN(n10186) );
  NAND2_X1 U11947 ( .A1(n10187), .A2(n10186), .ZN(n10189) );
  XNOR2_X1 U11948 ( .A(n10189), .B(n10188), .ZN(n10192) );
  AND2_X1 U11949 ( .A1(n15062), .A2(n14953), .ZN(n10190) );
  AOI21_X1 U11950 ( .B1(n15460), .B2(n7404), .A(n10190), .ZN(n10191) );
  NOR2_X1 U11951 ( .A1(n10192), .A2(n10191), .ZN(n14944) );
  NAND2_X1 U11952 ( .A1(n10192), .A2(n10191), .ZN(n14943) );
  XOR2_X1 U11953 ( .A(n10193), .B(n10194), .Z(n15014) );
  XNOR2_X1 U11954 ( .A(n10197), .B(n10196), .ZN(n14967) );
  NAND3_X1 U11955 ( .A1(n12255), .A2(P1_B_REG_SCAN_IN), .A3(n12198), .ZN(
        n10199) );
  OAI211_X1 U11956 ( .C1(P1_B_REG_SCAN_IN), .C2(n12198), .A(n10200), .B(n10199), .ZN(n15494) );
  INV_X1 U11957 ( .A(n10200), .ZN(n12455) );
  NAND2_X1 U11958 ( .A1(n12455), .A2(n12255), .ZN(n15496) );
  OAI21_X1 U11959 ( .B1(n15494), .B2(P1_D_REG_1__SCAN_IN), .A(n15496), .ZN(
        n10898) );
  NOR4_X1 U11960 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10209) );
  NOR4_X1 U11961 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10208) );
  NOR4_X1 U11962 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10204) );
  NOR4_X1 U11963 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10203) );
  NOR4_X1 U11964 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10202) );
  NOR4_X1 U11965 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10201) );
  NAND4_X1 U11966 ( .A1(n10204), .A2(n10203), .A3(n10202), .A4(n10201), .ZN(
        n10205) );
  NOR4_X1 U11967 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n10206), .A4(n10205), .ZN(n10207) );
  AND3_X1 U11968 ( .A1(n10209), .A2(n10208), .A3(n10207), .ZN(n10210) );
  NOR2_X1 U11969 ( .A1(n15494), .A2(n10210), .ZN(n10897) );
  NOR2_X1 U11970 ( .A1(n10898), .A2(n10897), .ZN(n11017) );
  INV_X1 U11971 ( .A(n15494), .ZN(n10212) );
  INV_X1 U11972 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U11973 ( .A1(n10212), .A2(n10211), .ZN(n10213) );
  NAND2_X1 U11974 ( .A1(n12455), .A2(n12198), .ZN(n15497) );
  NAND2_X1 U11975 ( .A1(n11017), .A2(n10917), .ZN(n10219) );
  INV_X1 U11976 ( .A(n10219), .ZN(n10230) );
  NAND2_X1 U11977 ( .A1(n10214), .A2(n10226), .ZN(n10263) );
  NAND2_X1 U11978 ( .A1(n7228), .A2(n12838), .ZN(n10227) );
  AND2_X1 U11979 ( .A1(n11027), .A2(n11419), .ZN(n15879) );
  INV_X1 U11980 ( .A(n10265), .ZN(n12851) );
  NAND2_X1 U11981 ( .A1(n16123), .A2(n12851), .ZN(n10215) );
  NOR2_X1 U11982 ( .A1(n10263), .A2(n10215), .ZN(n10216) );
  AOI211_X1 U11983 ( .C1(n10218), .C2(n10217), .A(n15042), .B(n14887), .ZN(
        n10238) );
  NAND2_X1 U11984 ( .A1(n10219), .A2(n11018), .ZN(n10449) );
  INV_X1 U11985 ( .A(n10263), .ZN(n15495) );
  AND2_X1 U11986 ( .A1(n11300), .A2(n16134), .ZN(n15040) );
  INV_X1 U11987 ( .A(n15040), .ZN(n16091) );
  NOR2_X1 U11988 ( .A1(n15439), .A2(n16091), .ZN(n10237) );
  NAND2_X1 U11989 ( .A1(n12833), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n10225) );
  NAND2_X1 U11990 ( .A1(n12834), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n10224) );
  INV_X1 U11991 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14931) );
  NAND2_X1 U11992 ( .A1(n10220), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n12593) );
  AOI21_X1 U11993 ( .B1(n14931), .B2(n10221), .A(n12580), .ZN(n14930) );
  NAND2_X1 U11994 ( .A1(n7212), .A2(n14930), .ZN(n10223) );
  NAND2_X1 U11995 ( .A1(n12829), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n10222) );
  NAND4_X1 U11996 ( .A1(n10225), .A2(n10224), .A3(n10223), .A4(n10222), .ZN(
        n15257) );
  INV_X1 U11997 ( .A(n15257), .ZN(n12615) );
  AND2_X1 U11998 ( .A1(n10226), .A2(n10264), .ZN(n10229) );
  NAND2_X1 U11999 ( .A1(n10265), .A2(n10227), .ZN(n10228) );
  AND2_X1 U12000 ( .A1(n10229), .A2(n10228), .ZN(n10233) );
  AND2_X1 U12001 ( .A1(n10233), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12911) );
  AND2_X1 U12002 ( .A1(n10230), .A2(n12911), .ZN(n15020) );
  NAND2_X1 U12003 ( .A1(n15020), .A2(n15376), .ZN(n15036) );
  OAI22_X1 U12004 ( .A1(n12615), .A2(n15036), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10232), .ZN(n10236) );
  INV_X1 U12005 ( .A(n15259), .ZN(n12780) );
  INV_X1 U12006 ( .A(n10231), .ZN(n10332) );
  AND2_X2 U12007 ( .A1(n10332), .A2(n10265), .ZN(n16030) );
  NAND2_X1 U12008 ( .A1(n15020), .A2(n16030), .ZN(n15049) );
  NAND2_X1 U12009 ( .A1(n10449), .A2(n10233), .ZN(n10234) );
  OAI22_X1 U12010 ( .A1(n12780), .A2(n15049), .B1(n16098), .B2(n15261), .ZN(
        n10235) );
  OR4_X1 U12011 ( .A1(n10238), .A2(n10237), .A3(n10236), .A4(n10235), .ZN(
        P1_U3235) );
  INV_X1 U12012 ( .A(n10729), .ZN(n10706) );
  NAND2_X1 U12013 ( .A1(n10706), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10239) );
  OAI21_X1 U12014 ( .B1(n10240), .B2(P3_STATE_REG_SCAN_IN), .A(n10239), .ZN(
        P3_U3294) );
  NAND2_X1 U12015 ( .A1(n10252), .A2(n7201), .ZN(n15512) );
  AND2_X1 U12016 ( .A1(n8315), .A2(P1_U3086), .ZN(n11949) );
  INV_X2 U12017 ( .A(n11949), .ZN(n15510) );
  OAI222_X1 U12018 ( .A1(n15512), .A2(n7646), .B1(n15510), .B2(n10246), .C1(
        n10331), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U12019 ( .A(n10241), .ZN(n10247) );
  OAI222_X1 U12020 ( .A1(n11951), .A2(n10242), .B1(n15510), .B2(n10247), .C1(
        P1_U3086), .C2(n10356), .ZN(P1_U3351) );
  OAI222_X1 U12021 ( .A1(n11951), .A2(n10243), .B1(n15510), .B2(n7254), .C1(
        n7201), .C2(n10351), .ZN(P1_U3353) );
  OAI222_X1 U12022 ( .A1(n11951), .A2(n10244), .B1(n15510), .B2(n10249), .C1(
        n7201), .C2(n10390), .ZN(P1_U3352) );
  AND2_X1 U12023 ( .A1(n10252), .A2(P2_U3088), .ZN(n14861) );
  INV_X2 U12024 ( .A(n14861), .ZN(n14869) );
  NAND2_X1 U12025 ( .A1(n8315), .A2(P2_U3088), .ZN(n14866) );
  INV_X1 U12026 ( .A(n14866), .ZN(n10258) );
  NOR2_X1 U12027 ( .A1(n10520), .A2(P2_U3088), .ZN(n15529) );
  AOI21_X1 U12028 ( .B1(n10258), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n15529), 
        .ZN(n10245) );
  OAI21_X1 U12029 ( .B1(n10246), .B2(n14869), .A(n10245), .ZN(P2_U3326) );
  INV_X1 U12030 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10248) );
  OAI222_X1 U12031 ( .A1(n14866), .A2(n10248), .B1(n14869), .B2(n10247), .C1(
        P2_U3088), .C2(n10529), .ZN(P2_U3323) );
  OAI222_X1 U12032 ( .A1(n14866), .A2(n8056), .B1(n14869), .B2(n10249), .C1(
        P2_U3088), .C2(n8055), .ZN(P2_U3324) );
  INV_X1 U12033 ( .A(n10250), .ZN(n10261) );
  INV_X1 U12034 ( .A(n10368), .ZN(n10344) );
  OAI222_X1 U12035 ( .A1(n11951), .A2(n10251), .B1(n15510), .B2(n10261), .C1(
        P1_U3086), .C2(n10344), .ZN(P1_U3350) );
  NOR2_X1 U12036 ( .A1(n10252), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14148) );
  INV_X2 U12037 ( .A(n14148), .ZN(n14158) );
  OAI222_X1 U12038 ( .A1(P3_U3151), .A2(n10717), .B1(n14158), .B2(n10254), 
        .C1(n10253), .C2(n14155), .ZN(P3_U3295) );
  OAI222_X1 U12039 ( .A1(n11499), .A2(P3_U3151), .B1(n14158), .B2(n10256), 
        .C1(n10255), .C2(n14155), .ZN(P3_U3287) );
  OAI222_X1 U12040 ( .A1(n12026), .A2(P3_U3151), .B1(n14158), .B2(n10257), 
        .C1(n13136), .C2(n14155), .ZN(P3_U3286) );
  OAI222_X1 U12041 ( .A1(n14871), .A2(n10259), .B1(n14869), .B2(n7254), .C1(
        P2_U3088), .C2(n15544), .ZN(P2_U3325) );
  INV_X1 U12042 ( .A(n15565), .ZN(n10260) );
  OAI222_X1 U12043 ( .A1(n14871), .A2(n10262), .B1(n14869), .B2(n10261), .C1(
        P2_U3088), .C2(n10260), .ZN(P2_U3322) );
  OR2_X1 U12044 ( .A1(n10264), .A2(P1_U3086), .ZN(n12913) );
  AND2_X1 U12045 ( .A1(n10263), .A2(n12913), .ZN(n10321) );
  INV_X1 U12046 ( .A(n10321), .ZN(n10268) );
  NAND2_X1 U12047 ( .A1(n10265), .A2(n10264), .ZN(n10266) );
  NAND2_X1 U12048 ( .A1(n7229), .A2(n10266), .ZN(n10322) );
  AND2_X1 U12049 ( .A1(n10268), .A2(n10322), .ZN(n15639) );
  NOR2_X1 U12050 ( .A1(n15639), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12051 ( .A(n10269), .ZN(n10272) );
  INV_X1 U12052 ( .A(n15577), .ZN(n10270) );
  OAI222_X1 U12053 ( .A1(n14866), .A2(n10271), .B1(n14869), .B2(n10272), .C1(
        P2_U3088), .C2(n10270), .ZN(P2_U3321) );
  INV_X1 U12054 ( .A(n10402), .ZN(n10406) );
  OAI222_X1 U12055 ( .A1(n11951), .A2(n10273), .B1(n15510), .B2(n10272), .C1(
        n7201), .C2(n10406), .ZN(P1_U3349) );
  INV_X1 U12056 ( .A(n10274), .ZN(n10275) );
  OAI222_X1 U12057 ( .A1(n15834), .A2(P3_U3151), .B1(n14158), .B2(n10275), 
        .C1(n13133), .C2(n14155), .ZN(P3_U3285) );
  INV_X1 U12058 ( .A(n10276), .ZN(n10284) );
  AOI22_X1 U12059 ( .A1(n10614), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n15503), .ZN(n10277) );
  OAI21_X1 U12060 ( .B1(n10284), .B2(n15510), .A(n10277), .ZN(P1_U3348) );
  OAI222_X1 U12061 ( .A1(n14158), .A2(n10279), .B1(n14155), .B2(n10278), .C1(
        P3_U3151), .C2(n11340), .ZN(P3_U3289) );
  INV_X1 U12062 ( .A(n10811), .ZN(n10853) );
  INV_X1 U12063 ( .A(n10280), .ZN(n10281) );
  OAI222_X1 U12064 ( .A1(P3_U3151), .A2(n10853), .B1(n14155), .B2(n10282), 
        .C1(n14158), .C2(n10281), .ZN(P3_U3293) );
  INV_X1 U12065 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10285) );
  INV_X1 U12066 ( .A(n14400), .ZN(n10283) );
  OAI222_X1 U12067 ( .A1(n14866), .A2(n10285), .B1(n14869), .B2(n10284), .C1(
        P2_U3088), .C2(n10283), .ZN(P2_U3320) );
  INV_X1 U12068 ( .A(n10286), .ZN(n10288) );
  INV_X1 U12069 ( .A(SI_5_), .ZN(n10287) );
  OAI222_X1 U12070 ( .A1(n10977), .A2(P3_U3151), .B1(n14158), .B2(n10288), 
        .C1(n10287), .C2(n14155), .ZN(P3_U3290) );
  INV_X1 U12071 ( .A(n10289), .ZN(n10291) );
  INV_X1 U12072 ( .A(SI_7_), .ZN(n10290) );
  OAI222_X1 U12073 ( .A1(n11498), .A2(P3_U3151), .B1(n14158), .B2(n10291), 
        .C1(n10290), .C2(n14155), .ZN(P3_U3288) );
  OAI222_X1 U12074 ( .A1(P3_U3151), .A2(n10974), .B1(n14158), .B2(n10293), 
        .C1(n10292), .C2(n14155), .ZN(P3_U3291) );
  INV_X1 U12075 ( .A(n10294), .ZN(n10296) );
  INV_X1 U12076 ( .A(SI_3_), .ZN(n10295) );
  OAI222_X1 U12077 ( .A1(P3_U3151), .A2(n7763), .B1(n14158), .B2(n10296), .C1(
        n10295), .C2(n14155), .ZN(P3_U3292) );
  INV_X1 U12078 ( .A(n10297), .ZN(n10300) );
  INV_X1 U12079 ( .A(n11159), .ZN(n11164) );
  OAI222_X1 U12080 ( .A1(n11951), .A2(n10298), .B1(n15510), .B2(n10300), .C1(
        P1_U3086), .C2(n11164), .ZN(P1_U3347) );
  INV_X1 U12081 ( .A(n14415), .ZN(n10299) );
  OAI222_X1 U12082 ( .A1(n14866), .A2(n10301), .B1(n14869), .B2(n10300), .C1(
        P2_U3088), .C2(n10299), .ZN(P2_U3319) );
  NAND2_X1 U12083 ( .A1(n11635), .A2(n14143), .ZN(n10302) );
  OAI21_X1 U12084 ( .B1(n10303), .B2(n14143), .A(n10302), .ZN(P3_U3377) );
  OAI21_X1 U12085 ( .B1(P2_U3947), .B2(n9858), .A(n10304), .ZN(P2_U3531) );
  INV_X1 U12086 ( .A(n10305), .ZN(n10306) );
  OAI222_X1 U12087 ( .A1(P3_U3151), .A2(n15855), .B1(n14155), .B2(n13130), 
        .C1(n14158), .C2(n10306), .ZN(P3_U3284) );
  OAI222_X1 U12088 ( .A1(n12051), .A2(P3_U3151), .B1(n14158), .B2(n10307), 
        .C1(n13019), .C2(n14155), .ZN(P3_U3283) );
  INV_X1 U12089 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10310) );
  NOR2_X1 U12090 ( .A1(n10547), .A2(n10310), .ZN(P3_U3260) );
  INV_X1 U12091 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10311) );
  NOR2_X1 U12092 ( .A1(n10547), .A2(n10311), .ZN(P3_U3251) );
  INV_X1 U12093 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10312) );
  NOR2_X1 U12094 ( .A1(n10547), .A2(n10312), .ZN(P3_U3259) );
  INV_X1 U12095 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10313) );
  NOR2_X1 U12096 ( .A1(n10547), .A2(n10313), .ZN(P3_U3247) );
  INV_X1 U12097 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10314) );
  NOR2_X1 U12098 ( .A1(n10547), .A2(n10314), .ZN(P3_U3248) );
  INV_X1 U12099 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10315) );
  NOR2_X1 U12100 ( .A1(n10547), .A2(n10315), .ZN(P3_U3261) );
  INV_X1 U12101 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10316) );
  NOR2_X1 U12102 ( .A1(n10547), .A2(n10316), .ZN(P3_U3246) );
  INV_X1 U12103 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10317) );
  NOR2_X1 U12104 ( .A1(n10547), .A2(n10317), .ZN(P3_U3249) );
  INV_X1 U12105 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10318) );
  NOR2_X1 U12106 ( .A1(n10547), .A2(n10318), .ZN(P3_U3250) );
  INV_X1 U12107 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10319) );
  NOR2_X1 U12108 ( .A1(n10547), .A2(n10319), .ZN(P3_U3258) );
  INV_X1 U12109 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10320) );
  NOR2_X1 U12110 ( .A1(n10547), .A2(n10320), .ZN(P3_U3253) );
  OR2_X1 U12111 ( .A1(n10322), .A2(n10321), .ZN(n15641) );
  INV_X1 U12112 ( .A(n10331), .ZN(n10347) );
  INV_X1 U12113 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11024) );
  OAI22_X1 U12114 ( .A1(n15656), .A2(n15664), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11024), .ZN(n10330) );
  NAND2_X1 U12115 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10328) );
  INV_X1 U12116 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10921) );
  INV_X1 U12117 ( .A(n10324), .ZN(n10327) );
  AND2_X1 U12118 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10323) );
  NAND2_X1 U12119 ( .A1(n10324), .A2(n10323), .ZN(n10338) );
  INV_X1 U12120 ( .A(n10338), .ZN(n10326) );
  INV_X1 U12121 ( .A(n15641), .ZN(n10325) );
  NAND2_X1 U12122 ( .A1(n10325), .A2(n15508), .ZN(n15145) );
  AOI211_X1 U12123 ( .C1(n10328), .C2(n10327), .A(n10326), .B(n15145), .ZN(
        n10329) );
  AOI211_X1 U12124 ( .C1(n15147), .C2(n10347), .A(n10330), .B(n10329), .ZN(
        n10336) );
  AND2_X1 U12125 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10334) );
  INV_X1 U12126 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11022) );
  MUX2_X1 U12127 ( .A(n11022), .B(P1_REG2_REG_1__SCAN_IN), .S(n10331), .Z(
        n10333) );
  NOR2_X1 U12128 ( .A1(n15641), .A2(n15508), .ZN(n15149) );
  AND2_X1 U12129 ( .A1(n15149), .A2(n10332), .ZN(n15143) );
  NAND2_X1 U12130 ( .A1(n10333), .A2(n10334), .ZN(n10349) );
  OAI211_X1 U12131 ( .C1(n10334), .C2(n10333), .A(n15143), .B(n10349), .ZN(
        n10335) );
  NAND2_X1 U12132 ( .A1(n10336), .A2(n10335), .ZN(P1_U3244) );
  INV_X1 U12133 ( .A(n10356), .ZN(n10742) );
  INV_X1 U12134 ( .A(n10390), .ZN(n10354) );
  INV_X1 U12135 ( .A(n10351), .ZN(n10783) );
  NAND2_X1 U12136 ( .A1(n10347), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10337) );
  NAND2_X1 U12137 ( .A1(n10338), .A2(n10337), .ZN(n10781) );
  INV_X1 U12138 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n11011) );
  MUX2_X1 U12139 ( .A(n11011), .B(P1_REG1_REG_2__SCAN_IN), .S(n10351), .Z(
        n10782) );
  NAND2_X1 U12140 ( .A1(n10781), .A2(n10782), .ZN(n10780) );
  INV_X1 U12141 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10339) );
  MUX2_X1 U12142 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10339), .S(n10390), .Z(
        n10386) );
  XOR2_X1 U12143 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10356), .Z(n10740) );
  NOR2_X1 U12144 ( .A1(n10741), .A2(n10740), .ZN(n10739) );
  AOI21_X1 U12145 ( .B1(n10742), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10739), .ZN(
        n10342) );
  INV_X1 U12146 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10340) );
  MUX2_X1 U12147 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10340), .S(n10368), .Z(
        n10341) );
  NAND2_X1 U12148 ( .A1(n10342), .A2(n10341), .ZN(n10365) );
  OAI21_X1 U12149 ( .B1(n10342), .B2(n10341), .A(n10365), .ZN(n10346) );
  INV_X1 U12150 ( .A(n15145), .ZN(n15652) );
  NAND2_X1 U12151 ( .A1(n7201), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11297) );
  NAND2_X1 U12152 ( .A1(n15639), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n10343) );
  OAI211_X1 U12153 ( .C1(n15647), .C2(n10344), .A(n11297), .B(n10343), .ZN(
        n10345) );
  AOI21_X1 U12154 ( .B1(n10346), .B2(n15652), .A(n10345), .ZN(n10364) );
  NAND2_X1 U12155 ( .A1(n10347), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10348) );
  NAND2_X1 U12156 ( .A1(n10349), .A2(n10348), .ZN(n10779) );
  XNOR2_X1 U12157 ( .A(n10351), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n10778) );
  INV_X1 U12158 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10350) );
  NOR2_X1 U12159 ( .A1(n10351), .A2(n10350), .ZN(n10352) );
  AOI21_X1 U12160 ( .B1(n10779), .B2(n10778), .A(n10352), .ZN(n10384) );
  INV_X1 U12161 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10353) );
  MUX2_X1 U12162 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10353), .S(n10390), .Z(
        n10383) );
  OR2_X1 U12163 ( .A1(n10384), .A2(n10383), .ZN(n10736) );
  NAND2_X1 U12164 ( .A1(n10354), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10735) );
  INV_X1 U12165 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10355) );
  MUX2_X1 U12166 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10355), .S(n10356), .Z(
        n10734) );
  AOI21_X1 U12167 ( .B1(n10736), .B2(n10735), .A(n10734), .ZN(n10738) );
  INV_X1 U12168 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10359) );
  MUX2_X1 U12169 ( .A(n10359), .B(P1_REG2_REG_5__SCAN_IN), .S(n10368), .Z(
        n10358) );
  NOR2_X1 U12170 ( .A1(n10356), .A2(n10355), .ZN(n10361) );
  INV_X1 U12171 ( .A(n10361), .ZN(n10357) );
  NAND2_X1 U12172 ( .A1(n10358), .A2(n10357), .ZN(n10362) );
  MUX2_X1 U12173 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10359), .S(n10368), .Z(
        n10360) );
  OAI21_X1 U12174 ( .B1(n10738), .B2(n10361), .A(n10360), .ZN(n10372) );
  OAI211_X1 U12175 ( .C1(n10738), .C2(n10362), .A(n15143), .B(n10372), .ZN(
        n10363) );
  NAND2_X1 U12176 ( .A1(n10364), .A2(n10363), .ZN(P1_U3248) );
  XNOR2_X1 U12177 ( .A(n10402), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10367) );
  OAI21_X1 U12178 ( .B1(n10368), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10365), .ZN(
        n10366) );
  NOR2_X1 U12179 ( .A1(n10366), .A2(n10367), .ZN(n10401) );
  AOI211_X1 U12180 ( .C1(n10367), .C2(n10366), .A(n15145), .B(n10401), .ZN(
        n10379) );
  NAND2_X1 U12181 ( .A1(n10368), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10371) );
  INV_X1 U12182 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10369) );
  MUX2_X1 U12183 ( .A(n10369), .B(P1_REG2_REG_6__SCAN_IN), .S(n10402), .Z(
        n10370) );
  AOI21_X1 U12184 ( .B1(n10372), .B2(n10371), .A(n10370), .ZN(n10413) );
  INV_X1 U12185 ( .A(n10413), .ZN(n10374) );
  NAND3_X1 U12186 ( .A1(n10372), .A2(n10371), .A3(n10370), .ZN(n10373) );
  NAND3_X1 U12187 ( .A1(n15143), .A2(n10374), .A3(n10373), .ZN(n10377) );
  INV_X1 U12188 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n11380) );
  NOR2_X1 U12189 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11380), .ZN(n10375) );
  AOI21_X1 U12190 ( .B1(n15639), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10375), .ZN(
        n10376) );
  OAI211_X1 U12191 ( .C1(n15647), .C2(n10406), .A(n10377), .B(n10376), .ZN(
        n10378) );
  OR2_X1 U12192 ( .A1(n10379), .A2(n10378), .ZN(P1_U3249) );
  INV_X1 U12193 ( .A(n10380), .ZN(n10398) );
  AOI22_X1 U12194 ( .A1(n15088), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n15503), .ZN(n10381) );
  OAI21_X1 U12195 ( .B1(n10398), .B2(n15510), .A(n10381), .ZN(P1_U3346) );
  INV_X1 U12196 ( .A(n10736), .ZN(n10382) );
  AOI211_X1 U12197 ( .C1(n10384), .C2(n10383), .A(n10382), .B(n15649), .ZN(
        n10393) );
  AOI211_X1 U12198 ( .C1(n10387), .C2(n10386), .A(n10385), .B(n15145), .ZN(
        n10392) );
  NOR2_X1 U12199 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9912), .ZN(n10388) );
  AOI21_X1 U12200 ( .B1(n15639), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n10388), .ZN(
        n10389) );
  OAI21_X1 U12201 ( .B1(n15647), .B2(n10390), .A(n10389), .ZN(n10391) );
  OR3_X1 U12202 ( .A1(n10393), .A2(n10392), .A3(n10391), .ZN(P1_U3246) );
  INV_X1 U12203 ( .A(n10394), .ZN(n10396) );
  INV_X1 U12204 ( .A(n11464), .ZN(n11468) );
  OAI222_X1 U12205 ( .A1(n11951), .A2(n10395), .B1(n15510), .B2(n10396), .C1(
        n7201), .C2(n11468), .ZN(P1_U3344) );
  INV_X1 U12206 ( .A(n11080), .ZN(n11093) );
  OAI222_X1 U12207 ( .A1(n14871), .A2(n10397), .B1(n14869), .B2(n10396), .C1(
        P2_U3088), .C2(n11093), .ZN(P2_U3316) );
  INV_X1 U12208 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10399) );
  INV_X1 U12209 ( .A(n10576), .ZN(n10542) );
  OAI222_X1 U12210 ( .A1(n14871), .A2(n10399), .B1(n14869), .B2(n10398), .C1(
        P2_U3088), .C2(n10542), .ZN(P2_U3318) );
  OAI222_X1 U12211 ( .A1(P3_U3151), .A2(n13608), .B1(n14155), .B2(n13121), 
        .C1(n14158), .C2(n10400), .ZN(P3_U3282) );
  INV_X1 U12212 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10403) );
  MUX2_X1 U12213 ( .A(n10403), .B(P1_REG1_REG_7__SCAN_IN), .S(n10614), .Z(
        n10404) );
  AOI211_X1 U12214 ( .C1(n10405), .C2(n10404), .A(n15145), .B(n10613), .ZN(
        n10418) );
  INV_X1 U12215 ( .A(n10614), .ZN(n10416) );
  NOR2_X1 U12216 ( .A1(n10406), .A2(n10369), .ZN(n10411) );
  INV_X1 U12217 ( .A(n10411), .ZN(n10409) );
  INV_X1 U12218 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10407) );
  MUX2_X1 U12219 ( .A(n10407), .B(P1_REG2_REG_7__SCAN_IN), .S(n10614), .Z(
        n10408) );
  NAND2_X1 U12220 ( .A1(n10409), .A2(n10408), .ZN(n10412) );
  MUX2_X1 U12221 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10407), .S(n10614), .Z(
        n10410) );
  OAI21_X1 U12222 ( .B1(n10413), .B2(n10411), .A(n10410), .ZN(n10611) );
  OAI211_X1 U12223 ( .C1(n10413), .C2(n10412), .A(n15143), .B(n10611), .ZN(
        n10415) );
  AND2_X1 U12224 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11459) );
  AOI21_X1 U12225 ( .B1(n15639), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n11459), .ZN(
        n10414) );
  OAI211_X1 U12226 ( .C1(n15647), .C2(n10416), .A(n10415), .B(n10414), .ZN(
        n10417) );
  OR2_X1 U12227 ( .A1(n10418), .A2(n10417), .ZN(P1_U3250) );
  INV_X1 U12228 ( .A(n10419), .ZN(n10421) );
  INV_X1 U12229 ( .A(n15626), .ZN(n11095) );
  OAI222_X1 U12230 ( .A1(n14871), .A2(n10420), .B1(n14869), .B2(n10421), .C1(
        P2_U3088), .C2(n11095), .ZN(P2_U3315) );
  INV_X1 U12231 ( .A(n11474), .ZN(n11835) );
  OAI222_X1 U12232 ( .A1(n11951), .A2(n10422), .B1(n15510), .B2(n10421), .C1(
        P1_U3086), .C2(n11835), .ZN(P1_U3343) );
  INV_X1 U12233 ( .A(n10423), .ZN(n10425) );
  INV_X1 U12234 ( .A(n14428), .ZN(n14420) );
  OAI222_X1 U12235 ( .A1(n14871), .A2(n10424), .B1(n14869), .B2(n10425), .C1(
        P2_U3088), .C2(n14420), .ZN(P2_U3317) );
  INV_X1 U12236 ( .A(n11236), .ZN(n11241) );
  OAI222_X1 U12237 ( .A1(n11951), .A2(n10426), .B1(n15510), .B2(n10425), .C1(
        P1_U3086), .C2(n11241), .ZN(P1_U3345) );
  OR2_X1 U12238 ( .A1(n10762), .A2(n10427), .ZN(n10431) );
  NAND2_X1 U12239 ( .A1(n10655), .A2(n10761), .ZN(n10429) );
  NAND2_X1 U12240 ( .A1(n10429), .A2(n10428), .ZN(n10430) );
  NAND2_X1 U12241 ( .A1(n10431), .A2(n10430), .ZN(n15530) );
  OR2_X1 U12242 ( .A1(n9707), .A2(P2_U3088), .ZN(n14863) );
  INV_X1 U12243 ( .A(n14863), .ZN(n10432) );
  INV_X1 U12244 ( .A(n10435), .ZN(n10433) );
  OR2_X1 U12245 ( .A1(n10433), .A2(n10434), .ZN(n15622) );
  NAND2_X1 U12246 ( .A1(n15611), .A2(n10439), .ZN(n10437) );
  AND2_X1 U12247 ( .A1(n9707), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10436) );
  NAND2_X1 U12248 ( .A1(n15530), .A2(n10436), .ZN(n15543) );
  OAI211_X1 U12249 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15622), .A(n10437), .B(
        n15543), .ZN(n10442) );
  INV_X1 U12250 ( .A(n15611), .ZN(n15630) );
  OAI22_X1 U12251 ( .A1(n15630), .A2(n10439), .B1(n10438), .B2(n15622), .ZN(
        n10441) );
  MUX2_X1 U12252 ( .A(n10442), .B(n10441), .S(n10440), .Z(n10446) );
  INV_X1 U12253 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10444) );
  OAI22_X1 U12254 ( .A1(n15616), .A2(n10444), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10443), .ZN(n10445) );
  OR2_X1 U12255 ( .A1(n10446), .A2(n10445), .ZN(P2_U3214) );
  INV_X1 U12256 ( .A(n15878), .ZN(n11060) );
  XOR2_X1 U12257 ( .A(n10448), .B(n10447), .Z(n10731) );
  NAND2_X1 U12258 ( .A1(n10731), .A2(n16093), .ZN(n10451) );
  INV_X1 U12259 ( .A(n15036), .ZN(n16089) );
  NAND2_X1 U12260 ( .A1(n10449), .A2(n12911), .ZN(n10990) );
  AOI22_X1 U12261 ( .A1(n16089), .A2(n15075), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10990), .ZN(n10450) );
  OAI211_X1 U12262 ( .C1(n16091), .C2(n11060), .A(n10451), .B(n10450), .ZN(
        P1_U3232) );
  NOR4_X1 U12263 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n10460) );
  NOR4_X1 U12264 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n10455) );
  NOR4_X1 U12265 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n10454) );
  NOR4_X1 U12266 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n10453) );
  NOR4_X1 U12267 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n10452) );
  NAND4_X1 U12268 ( .A1(n10455), .A2(n10454), .A3(n10453), .A4(n10452), .ZN(
        n10456) );
  NOR4_X1 U12269 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        n10457), .A4(n10456), .ZN(n10459) );
  NOR4_X1 U12270 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n10458) );
  NAND3_X1 U12271 ( .A1(n10460), .A2(n10459), .A3(n10458), .ZN(n10463) );
  XNOR2_X1 U12272 ( .A(n12199), .B(P2_B_REG_SCAN_IN), .ZN(n10461) );
  NAND2_X1 U12273 ( .A1(n12256), .A2(n10461), .ZN(n10462) );
  AND2_X1 U12274 ( .A1(n10463), .A2(n15519), .ZN(n10645) );
  AND2_X1 U12275 ( .A1(n10655), .A2(n10649), .ZN(n10651) );
  INV_X1 U12276 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15518) );
  NAND2_X1 U12277 ( .A1(n15519), .A2(n15518), .ZN(n10466) );
  INV_X1 U12278 ( .A(n12256), .ZN(n10464) );
  OR2_X1 U12279 ( .A1(n12451), .A2(n10464), .ZN(n10465) );
  NAND2_X1 U12280 ( .A1(n10466), .A2(n10465), .ZN(n11730) );
  AND2_X1 U12281 ( .A1(n11730), .A2(n15525), .ZN(n15517) );
  INV_X2 U12282 ( .A(n10697), .ZN(n14716) );
  AND2_X1 U12283 ( .A1(n15517), .A2(n10652), .ZN(n10469) );
  AND2_X1 U12284 ( .A1(n11733), .A2(n10469), .ZN(n10945) );
  INV_X1 U12285 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15523) );
  NAND2_X1 U12286 ( .A1(n15519), .A2(n15523), .ZN(n10472) );
  INV_X1 U12287 ( .A(n12199), .ZN(n10470) );
  INV_X1 U12288 ( .A(n15524), .ZN(n10473) );
  INV_X1 U12289 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10505) );
  NAND2_X1 U12290 ( .A1(n7425), .A2(n10493), .ZN(n10491) );
  OR2_X1 U12291 ( .A1(n14377), .A2(n10679), .ZN(n10474) );
  NAND2_X1 U12292 ( .A1(n10491), .A2(n10474), .ZN(n10595) );
  XNOR2_X1 U12293 ( .A(n10595), .B(n10594), .ZN(n10479) );
  NAND2_X1 U12294 ( .A1(n10646), .A2(n10475), .ZN(n10476) );
  INV_X1 U12295 ( .A(n14377), .ZN(n10478) );
  INV_X1 U12296 ( .A(n14374), .ZN(n10695) );
  NAND2_X1 U12297 ( .A1(n10655), .A2(n9707), .ZN(n14453) );
  OAI22_X1 U12298 ( .A1(n10478), .A2(n14313), .B1(n10695), .B2(n14453), .ZN(
        n10654) );
  AOI21_X1 U12299 ( .B1(n10479), .B2(n14710), .A(n10654), .ZN(n11828) );
  OR2_X1 U12300 ( .A1(n14377), .A2(n11879), .ZN(n10480) );
  NAND2_X1 U12301 ( .A1(n10488), .A2(n10480), .ZN(n10482) );
  INV_X1 U12302 ( .A(n10594), .ZN(n10481) );
  OAI21_X1 U12303 ( .B1(n10482), .B2(n10481), .A(n10589), .ZN(n11825) );
  XNOR2_X1 U12304 ( .A(n11734), .B(n8886), .ZN(n10483) );
  INV_X1 U12305 ( .A(n16006), .ZN(n16153) );
  INV_X1 U12306 ( .A(n10587), .ZN(n11822) );
  NOR2_X2 U12307 ( .A1(n10484), .A2(n10774), .ZN(n16112) );
  NAND2_X1 U12308 ( .A1(n10499), .A2(n11822), .ZN(n10591) );
  OAI211_X1 U12309 ( .C1(n10499), .C2(n11822), .A(n14716), .B(n10591), .ZN(
        n11821) );
  OAI21_X1 U12310 ( .B1(n11822), .B2(n16149), .A(n11821), .ZN(n10485) );
  AOI21_X1 U12311 ( .B1(n11825), .B2(n16153), .A(n10485), .ZN(n10486) );
  NAND2_X1 U12312 ( .A1(n11828), .A2(n10486), .ZN(n10948) );
  NAND2_X1 U12313 ( .A1(n16156), .A2(n10948), .ZN(n10487) );
  OAI21_X1 U12314 ( .B1(n16156), .B2(n10505), .A(n10487), .ZN(P2_U3501) );
  INV_X1 U12315 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10503) );
  INV_X1 U12316 ( .A(n10488), .ZN(n10489) );
  AOI21_X1 U12317 ( .B1(n10490), .B2(n7425), .A(n10489), .ZN(n11884) );
  OAI21_X1 U12318 ( .B1(n10493), .B2(n7425), .A(n10491), .ZN(n10495) );
  INV_X1 U12319 ( .A(n14375), .ZN(n10598) );
  OAI22_X1 U12320 ( .A1(n10494), .A2(n14313), .B1(n10598), .B2(n14453), .ZN(
        n10672) );
  AOI21_X1 U12321 ( .B1(n10495), .B2(n14710), .A(n10672), .ZN(n11881) );
  NAND2_X1 U12322 ( .A1(n10496), .A2(n11879), .ZN(n10497) );
  NAND2_X1 U12323 ( .A1(n10497), .A2(n14716), .ZN(n10498) );
  OR2_X1 U12324 ( .A1(n10499), .A2(n10498), .ZN(n11877) );
  INV_X1 U12325 ( .A(n11877), .ZN(n10500) );
  AOI21_X1 U12326 ( .B1(n16112), .B2(n11879), .A(n10500), .ZN(n10501) );
  OAI211_X1 U12327 ( .C1(n11884), .C2(n16006), .A(n11881), .B(n10501), .ZN(
        n10946) );
  NAND2_X1 U12328 ( .A1(n16156), .A2(n10946), .ZN(n10502) );
  OAI21_X1 U12329 ( .B1(n16156), .B2(n10503), .A(n10502), .ZN(P2_U3500) );
  MUX2_X1 U12330 ( .A(n9096), .B(P2_REG1_REG_9__SCAN_IN), .S(n10576), .Z(
        n10518) );
  MUX2_X1 U12331 ( .A(n10503), .B(P2_REG1_REG_1__SCAN_IN), .S(n10520), .Z(
        n15528) );
  AND2_X1 U12332 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15527) );
  NAND2_X1 U12333 ( .A1(n15528), .A2(n15527), .ZN(n15526) );
  INV_X1 U12334 ( .A(n10520), .ZN(n10521) );
  NAND2_X1 U12335 ( .A1(n10521), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10504) );
  NAND2_X1 U12336 ( .A1(n15526), .A2(n10504), .ZN(n15541) );
  MUX2_X1 U12337 ( .A(n10505), .B(P2_REG1_REG_2__SCAN_IN), .S(n15544), .Z(
        n15542) );
  NAND2_X1 U12338 ( .A1(n15541), .A2(n15542), .ZN(n15540) );
  INV_X1 U12339 ( .A(n15544), .ZN(n10524) );
  NAND2_X1 U12340 ( .A1(n10524), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10506) );
  NAND2_X1 U12341 ( .A1(n15540), .A2(n10506), .ZN(n14379) );
  INV_X1 U12342 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10602) );
  MUX2_X1 U12343 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10602), .S(n14387), .Z(
        n14380) );
  NAND2_X1 U12344 ( .A1(n14379), .A2(n14380), .ZN(n14378) );
  NAND2_X1 U12345 ( .A1(n14387), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10507) );
  NAND2_X1 U12346 ( .A1(n14378), .A2(n10507), .ZN(n15555) );
  INV_X1 U12347 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10703) );
  MUX2_X1 U12348 ( .A(n10703), .B(P2_REG1_REG_4__SCAN_IN), .S(n10529), .Z(
        n15556) );
  NAND2_X1 U12349 ( .A1(n15555), .A2(n15556), .ZN(n15554) );
  NAND2_X1 U12350 ( .A1(n15553), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10508) );
  NAND2_X1 U12351 ( .A1(n15554), .A2(n10508), .ZN(n15567) );
  INV_X1 U12352 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10509) );
  XNOR2_X1 U12353 ( .A(n15565), .B(n10509), .ZN(n15568) );
  NAND2_X1 U12354 ( .A1(n15567), .A2(n15568), .ZN(n15566) );
  NAND2_X1 U12355 ( .A1(n15565), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10510) );
  NAND2_X1 U12356 ( .A1(n15566), .A2(n10510), .ZN(n15579) );
  INV_X1 U12357 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10511) );
  XNOR2_X1 U12358 ( .A(n15577), .B(n10511), .ZN(n15580) );
  NAND2_X1 U12359 ( .A1(n15579), .A2(n15580), .ZN(n15578) );
  NAND2_X1 U12360 ( .A1(n15577), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10512) );
  NAND2_X1 U12361 ( .A1(n15578), .A2(n10512), .ZN(n14393) );
  INV_X1 U12362 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n11412) );
  MUX2_X1 U12363 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n11412), .S(n14400), .Z(
        n14394) );
  NAND2_X1 U12364 ( .A1(n14393), .A2(n14394), .ZN(n14392) );
  NAND2_X1 U12365 ( .A1(n14400), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10513) );
  NAND2_X1 U12366 ( .A1(n14392), .A2(n10513), .ZN(n14406) );
  INV_X1 U12367 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10514) );
  XNOR2_X1 U12368 ( .A(n14415), .B(n10514), .ZN(n14407) );
  NAND2_X1 U12369 ( .A1(n14406), .A2(n14407), .ZN(n14405) );
  NAND2_X1 U12370 ( .A1(n14415), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10515) );
  NAND2_X1 U12371 ( .A1(n14405), .A2(n10515), .ZN(n10517) );
  OR2_X1 U12372 ( .A1(n10517), .A2(n10518), .ZN(n10578) );
  INV_X1 U12373 ( .A(n10578), .ZN(n10516) );
  AOI21_X1 U12374 ( .B1(n10518), .B2(n10517), .A(n10516), .ZN(n10546) );
  INV_X1 U12375 ( .A(n15616), .ZN(n15619) );
  MUX2_X1 U12376 ( .A(n10519), .B(P2_REG2_REG_9__SCAN_IN), .S(n10576), .Z(
        n10540) );
  MUX2_X1 U12377 ( .A(n11880), .B(P2_REG2_REG_1__SCAN_IN), .S(n10520), .Z(
        n15535) );
  AND2_X1 U12378 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15536) );
  NAND2_X1 U12379 ( .A1(n15535), .A2(n15536), .ZN(n15534) );
  NAND2_X1 U12380 ( .A1(n10521), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10522) );
  NAND2_X1 U12381 ( .A1(n15534), .A2(n10522), .ZN(n15549) );
  MUX2_X1 U12382 ( .A(n10523), .B(P2_REG2_REG_2__SCAN_IN), .S(n15544), .Z(
        n15548) );
  NAND2_X1 U12383 ( .A1(n15549), .A2(n15548), .ZN(n15547) );
  NAND2_X1 U12384 ( .A1(n10524), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n14382) );
  NAND2_X1 U12385 ( .A1(n15547), .A2(n14382), .ZN(n10527) );
  MUX2_X1 U12386 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10525), .S(n14387), .Z(
        n10526) );
  NAND2_X1 U12387 ( .A1(n10527), .A2(n10526), .ZN(n14384) );
  NAND2_X1 U12388 ( .A1(n14387), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10528) );
  NAND2_X1 U12389 ( .A1(n14384), .A2(n10528), .ZN(n15561) );
  MUX2_X1 U12390 ( .A(n10530), .B(P2_REG2_REG_4__SCAN_IN), .S(n10529), .Z(
        n15560) );
  NAND2_X1 U12391 ( .A1(n15561), .A2(n15560), .ZN(n15559) );
  NAND2_X1 U12392 ( .A1(n15553), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10531) );
  NAND2_X1 U12393 ( .A1(n15559), .A2(n10531), .ZN(n15573) );
  MUX2_X1 U12394 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11767), .S(n15565), .Z(
        n15572) );
  NAND2_X1 U12395 ( .A1(n15573), .A2(n15572), .ZN(n15571) );
  NAND2_X1 U12396 ( .A1(n15565), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10532) );
  NAND2_X1 U12397 ( .A1(n15571), .A2(n10532), .ZN(n15585) );
  MUX2_X1 U12398 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11775), .S(n15577), .Z(
        n15584) );
  NAND2_X1 U12399 ( .A1(n15585), .A2(n15584), .ZN(n15583) );
  NAND2_X1 U12400 ( .A1(n15577), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n14396) );
  NAND2_X1 U12401 ( .A1(n15583), .A2(n14396), .ZN(n10534) );
  MUX2_X1 U12402 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11805), .S(n14400), .Z(
        n10533) );
  NAND2_X1 U12403 ( .A1(n10534), .A2(n10533), .ZN(n14410) );
  NAND2_X1 U12404 ( .A1(n14400), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n14409) );
  NAND2_X1 U12405 ( .A1(n14410), .A2(n14409), .ZN(n10536) );
  MUX2_X1 U12406 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11756), .S(n14415), .Z(
        n10535) );
  NAND2_X1 U12407 ( .A1(n10536), .A2(n10535), .ZN(n14412) );
  NAND2_X1 U12408 ( .A1(n14415), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10537) );
  NAND2_X1 U12409 ( .A1(n14412), .A2(n10537), .ZN(n10539) );
  OR2_X1 U12410 ( .A1(n10539), .A2(n10540), .ZN(n10569) );
  INV_X1 U12411 ( .A(n10569), .ZN(n10538) );
  AOI21_X1 U12412 ( .B1(n10540), .B2(n10539), .A(n10538), .ZN(n10541) );
  OAI22_X1 U12413 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11369), .B1(n10541), .B2(
        n15630), .ZN(n10544) );
  NOR2_X1 U12414 ( .A1(n15543), .A2(n10542), .ZN(n10543) );
  AOI211_X1 U12415 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n15619), .A(n10544), .B(
        n10543), .ZN(n10545) );
  OAI21_X1 U12416 ( .B1(n10546), .B2(n15622), .A(n10545), .ZN(P2_U3223) );
  CLKBUF_X1 U12417 ( .A(n10547), .Z(n10567) );
  INV_X1 U12418 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10548) );
  NOR2_X1 U12419 ( .A1(n10567), .A2(n10548), .ZN(P3_U3263) );
  INV_X1 U12420 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10549) );
  NOR2_X1 U12421 ( .A1(n10567), .A2(n10549), .ZN(P3_U3257) );
  INV_X1 U12422 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10550) );
  NOR2_X1 U12423 ( .A1(n10567), .A2(n10550), .ZN(P3_U3262) );
  INV_X1 U12424 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10551) );
  NOR2_X1 U12425 ( .A1(n10567), .A2(n10551), .ZN(P3_U3255) );
  INV_X1 U12426 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10552) );
  NOR2_X1 U12427 ( .A1(n10567), .A2(n10552), .ZN(P3_U3256) );
  INV_X1 U12428 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10553) );
  NOR2_X1 U12429 ( .A1(n10567), .A2(n10553), .ZN(P3_U3254) );
  INV_X1 U12430 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10554) );
  NOR2_X1 U12431 ( .A1(n10567), .A2(n10554), .ZN(P3_U3252) );
  INV_X1 U12432 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10555) );
  NOR2_X1 U12433 ( .A1(n10567), .A2(n10555), .ZN(P3_U3239) );
  INV_X1 U12434 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10556) );
  NOR2_X1 U12435 ( .A1(n10567), .A2(n10556), .ZN(P3_U3236) );
  INV_X1 U12436 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10557) );
  NOR2_X1 U12437 ( .A1(n10567), .A2(n10557), .ZN(P3_U3245) );
  INV_X1 U12438 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10558) );
  NOR2_X1 U12439 ( .A1(n10567), .A2(n10558), .ZN(P3_U3244) );
  INV_X1 U12440 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10559) );
  NOR2_X1 U12441 ( .A1(n10567), .A2(n10559), .ZN(P3_U3243) );
  INV_X1 U12442 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10560) );
  NOR2_X1 U12443 ( .A1(n10567), .A2(n10560), .ZN(P3_U3237) );
  INV_X1 U12444 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10561) );
  NOR2_X1 U12445 ( .A1(n10567), .A2(n10561), .ZN(P3_U3234) );
  INV_X1 U12446 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10562) );
  NOR2_X1 U12447 ( .A1(n10567), .A2(n10562), .ZN(P3_U3242) );
  INV_X1 U12448 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10563) );
  NOR2_X1 U12449 ( .A1(n10567), .A2(n10563), .ZN(P3_U3240) );
  INV_X1 U12450 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10564) );
  NOR2_X1 U12451 ( .A1(n10567), .A2(n10564), .ZN(P3_U3241) );
  INV_X1 U12452 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10565) );
  NOR2_X1 U12453 ( .A1(n10567), .A2(n10565), .ZN(P3_U3235) );
  INV_X1 U12454 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10566) );
  NOR2_X1 U12455 ( .A1(n10567), .A2(n10566), .ZN(P3_U3238) );
  OR2_X1 U12456 ( .A1(n10576), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10568) );
  NAND2_X1 U12457 ( .A1(n10569), .A2(n10568), .ZN(n14427) );
  MUX2_X1 U12458 ( .A(n14429), .B(P2_REG2_REG_10__SCAN_IN), .S(n14428), .Z(
        n10570) );
  OR2_X1 U12459 ( .A1(n14427), .A2(n10570), .ZN(n14430) );
  NAND2_X1 U12460 ( .A1(n14428), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10571) );
  NAND2_X1 U12461 ( .A1(n14430), .A2(n10571), .ZN(n10573) );
  MUX2_X1 U12462 ( .A(n11092), .B(P2_REG2_REG_11__SCAN_IN), .S(n11080), .Z(
        n10572) );
  NOR2_X1 U12463 ( .A1(n10573), .A2(n10572), .ZN(n11091) );
  AOI21_X1 U12464 ( .B1(n10573), .B2(n10572), .A(n11091), .ZN(n10586) );
  AND2_X1 U12465 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10575) );
  NOR2_X1 U12466 ( .A1(n15543), .A2(n11093), .ZN(n10574) );
  AOI211_X1 U12467 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n15619), .A(n10575), 
        .B(n10574), .ZN(n10585) );
  OR2_X1 U12468 ( .A1(n10576), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10577) );
  NAND2_X1 U12469 ( .A1(n10578), .A2(n10577), .ZN(n14424) );
  INV_X1 U12470 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10579) );
  MUX2_X1 U12471 ( .A(n10579), .B(P2_REG1_REG_10__SCAN_IN), .S(n14428), .Z(
        n14423) );
  OR2_X1 U12472 ( .A1(n14424), .A2(n14423), .ZN(n14425) );
  NAND2_X1 U12473 ( .A1(n14428), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10580) );
  NAND2_X1 U12474 ( .A1(n14425), .A2(n10580), .ZN(n10583) );
  INV_X1 U12475 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10581) );
  MUX2_X1 U12476 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10581), .S(n11080), .Z(
        n10582) );
  NAND2_X1 U12477 ( .A1(n10583), .A2(n10582), .ZN(n11082) );
  OAI211_X1 U12478 ( .C1(n10583), .C2(n10582), .A(n11082), .B(n15602), .ZN(
        n10584) );
  OAI211_X1 U12479 ( .C1(n10586), .C2(n15630), .A(n10585), .B(n10584), .ZN(
        P2_U3225) );
  OR2_X1 U12480 ( .A1(n14375), .A2(n10587), .ZN(n10588) );
  NAND2_X1 U12481 ( .A1(n10589), .A2(n10588), .ZN(n10590) );
  AOI21_X1 U12482 ( .B1(n10591), .B2(n12099), .A(n14633), .ZN(n10592) );
  OR2_X1 U12483 ( .A1(n10591), .A2(n12099), .ZN(n10698) );
  NAND2_X1 U12484 ( .A1(n10592), .A2(n10698), .ZN(n12103) );
  OAI21_X1 U12485 ( .B1(n10844), .B2(n16149), .A(n12103), .ZN(n10593) );
  AOI21_X1 U12486 ( .B1(n12105), .B2(n16153), .A(n10593), .ZN(n10600) );
  NAND2_X1 U12487 ( .A1(n10595), .A2(n10594), .ZN(n10597) );
  OR2_X1 U12488 ( .A1(n14375), .A2(n11822), .ZN(n10596) );
  XNOR2_X1 U12489 ( .A(n10692), .B(n10691), .ZN(n10599) );
  OAI22_X1 U12490 ( .A1(n10598), .A2(n14313), .B1(n10830), .B2(n14453), .ZN(
        n10842) );
  AOI21_X1 U12491 ( .B1(n10599), .B2(n14710), .A(n10842), .ZN(n12107) );
  NAND2_X1 U12492 ( .A1(n10600), .A2(n12107), .ZN(n10952) );
  NAND2_X1 U12493 ( .A1(n10952), .A2(n16156), .ZN(n10601) );
  OAI21_X1 U12494 ( .B1(n16156), .B2(n10602), .A(n10601), .ZN(P2_U3502) );
  INV_X1 U12495 ( .A(n10603), .ZN(n10604) );
  OAI222_X1 U12496 ( .A1(P2_U3088), .A2(n11098), .B1(n14869), .B2(n10604), 
        .C1(n8101), .C2(n14871), .ZN(P2_U3314) );
  INV_X1 U12497 ( .A(n11837), .ZN(n15096) );
  OAI222_X1 U12498 ( .A1(n11951), .A2(n10605), .B1(n15510), .B2(n10604), .C1(
        n15096), .C2(n7201), .ZN(P1_U3342) );
  INV_X1 U12499 ( .A(n13656), .ZN(n13634) );
  INV_X1 U12500 ( .A(n10606), .ZN(n10607) );
  OAI222_X1 U12501 ( .A1(P3_U3151), .A2(n13634), .B1(n14155), .B2(n13124), 
        .C1(n14158), .C2(n10607), .ZN(P3_U3281) );
  OAI222_X1 U12502 ( .A1(P3_U3151), .A2(n13657), .B1(n14155), .B2(n13122), 
        .C1(n14158), .C2(n10608), .ZN(P3_U3280) );
  NAND2_X1 U12503 ( .A1(n10614), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10610) );
  INV_X1 U12504 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11163) );
  MUX2_X1 U12505 ( .A(n11163), .B(P1_REG2_REG_8__SCAN_IN), .S(n11159), .Z(
        n10609) );
  AOI21_X1 U12506 ( .B1(n10611), .B2(n10610), .A(n10609), .ZN(n15087) );
  NAND3_X1 U12507 ( .A1(n10611), .A2(n10610), .A3(n10609), .ZN(n10612) );
  NAND2_X1 U12508 ( .A1(n15143), .A2(n10612), .ZN(n10623) );
  INV_X1 U12509 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10615) );
  MUX2_X1 U12510 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10615), .S(n11159), .Z(
        n10616) );
  OAI21_X1 U12511 ( .B1(n10617), .B2(n10616), .A(n11158), .ZN(n10618) );
  NAND2_X1 U12512 ( .A1(n10618), .A2(n15652), .ZN(n10622) );
  AND2_X1 U12513 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10620) );
  NOR2_X1 U12514 ( .A1(n15647), .A2(n11164), .ZN(n10619) );
  AOI211_X1 U12515 ( .C1(n15639), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10620), .B(
        n10619), .ZN(n10621) );
  OAI211_X1 U12516 ( .C1(n15087), .C2(n10623), .A(n10622), .B(n10621), .ZN(
        P1_U3251) );
  INV_X1 U12517 ( .A(n11176), .ZN(n10624) );
  OR2_X1 U12518 ( .A1(n10625), .A2(P3_U3151), .ZN(n13568) );
  NAND2_X1 U12519 ( .A1(n10624), .A2(n13568), .ZN(n10636) );
  INV_X1 U12520 ( .A(n10625), .ZN(n10626) );
  OR2_X1 U12521 ( .A1(n13474), .A2(n10626), .ZN(n10627) );
  AND2_X1 U12522 ( .A1(n7204), .A2(n10627), .ZN(n10635) );
  NAND2_X1 U12523 ( .A1(n10636), .A2(n10635), .ZN(n10638) );
  NAND2_X1 U12524 ( .A1(P3_U3897), .A2(n8827), .ZN(n15843) );
  NOR3_X1 U12525 ( .A1(n7465), .A2(n13722), .A3(n15863), .ZN(n10643) );
  INV_X1 U12526 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10632) );
  INV_X1 U12527 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10631) );
  MUX2_X1 U12528 ( .A(n10632), .B(n10631), .S(n10630), .Z(n10633) );
  INV_X1 U12529 ( .A(n10633), .ZN(n10634) );
  NAND2_X1 U12530 ( .A1(n10633), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10710) );
  INV_X1 U12531 ( .A(n10710), .ZN(n10712) );
  AOI21_X1 U12532 ( .B1(n10717), .B2(n10634), .A(n10712), .ZN(n10642) );
  INV_X1 U12533 ( .A(n10635), .ZN(n10637) );
  AOI22_X1 U12534 ( .A1(n15521), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10641) );
  INV_X1 U12535 ( .A(n10638), .ZN(n10639) );
  NAND2_X1 U12536 ( .A1(n13754), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10640) );
  OAI211_X1 U12537 ( .C1(n10643), .C2(n10642), .A(n10641), .B(n10640), .ZN(
        P3_U3182) );
  OR2_X1 U12538 ( .A1(n15524), .A2(n11730), .ZN(n10644) );
  NOR2_X1 U12539 ( .A1(n10645), .A2(n10644), .ZN(n10650) );
  NAND2_X1 U12540 ( .A1(n10650), .A2(n15525), .ZN(n10657) );
  NAND2_X1 U12541 ( .A1(n10468), .A2(n10646), .ZN(n11737) );
  OR2_X1 U12542 ( .A1(n10657), .A2(n11737), .ZN(n10648) );
  INV_X1 U12543 ( .A(n10652), .ZN(n10647) );
  INV_X1 U12544 ( .A(n10650), .ZN(n10653) );
  AOI21_X1 U12545 ( .B1(n10653), .B2(n10652), .A(n10651), .ZN(n10763) );
  NAND2_X1 U12546 ( .A1(n10763), .A2(n15525), .ZN(n10681) );
  AOI22_X1 U12547 ( .A1(n14348), .A2(n10654), .B1(n10681), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n10671) );
  OR2_X1 U12548 ( .A1(n16112), .A2(n10655), .ZN(n10656) );
  XNOR2_X1 U12549 ( .A(n14229), .B(n11822), .ZN(n10659) );
  NAND2_X1 U12550 ( .A1(n14375), .A2(n10697), .ZN(n10660) );
  NAND2_X1 U12551 ( .A1(n10659), .A2(n10660), .ZN(n10748) );
  XNOR2_X1 U12552 ( .A(n10679), .B(n10662), .ZN(n10663) );
  NAND2_X1 U12553 ( .A1(n14377), .A2(n10697), .ZN(n10664) );
  NAND2_X1 U12554 ( .A1(n10663), .A2(n10664), .ZN(n10667) );
  OR2_X1 U12555 ( .A1(n10683), .A2(n14716), .ZN(n10680) );
  NAND2_X1 U12556 ( .A1(n7214), .A2(n10775), .ZN(n10666) );
  NAND2_X1 U12557 ( .A1(n10673), .A2(n10667), .ZN(n10668) );
  NAND2_X1 U12558 ( .A1(n14311), .A2(n10669), .ZN(n10670) );
  OAI211_X1 U12559 ( .C1(n11822), .C2(n14309), .A(n10671), .B(n10670), .ZN(
        P2_U3209) );
  AOI22_X1 U12560 ( .A1(n14348), .A2(n10672), .B1(n10681), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10678) );
  OAI21_X1 U12561 ( .B1(n10675), .B2(n10674), .A(n10673), .ZN(n10676) );
  NAND2_X1 U12562 ( .A1(n14311), .A2(n10676), .ZN(n10677) );
  OAI211_X1 U12563 ( .C1(n10679), .C2(n14309), .A(n10678), .B(n10677), .ZN(
        P2_U3194) );
  AOI21_X1 U12564 ( .B1(n14311), .B2(n10680), .A(n14358), .ZN(n10686) );
  NAND2_X1 U12565 ( .A1(n14377), .A2(n14338), .ZN(n10772) );
  INV_X1 U12566 ( .A(n10772), .ZN(n10682) );
  AOI22_X1 U12567 ( .A1(n14348), .A2(n10682), .B1(n10681), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10685) );
  NOR2_X1 U12568 ( .A1(n14353), .A2(n14716), .ZN(n14330) );
  OAI211_X1 U12569 ( .C1(n10686), .C2(n10775), .A(n10685), .B(n10684), .ZN(
        P2_U3204) );
  OR2_X1 U12570 ( .A1(n14374), .A2(n12099), .ZN(n10687) );
  NAND2_X1 U12571 ( .A1(n10688), .A2(n10687), .ZN(n10690) );
  INV_X1 U12572 ( .A(n10828), .ZN(n10689) );
  NAND2_X1 U12573 ( .A1(n10690), .A2(n10689), .ZN(n10826) );
  OAI21_X1 U12574 ( .B1(n10690), .B2(n10689), .A(n10826), .ZN(n11747) );
  INV_X1 U12575 ( .A(n11747), .ZN(n10701) );
  NAND2_X1 U12576 ( .A1(n10692), .A2(n10691), .ZN(n10694) );
  OR2_X1 U12577 ( .A1(n14374), .A2(n10844), .ZN(n10693) );
  XNOR2_X1 U12578 ( .A(n10829), .B(n10828), .ZN(n10696) );
  INV_X1 U12579 ( .A(n14372), .ZN(n11050) );
  OAI22_X1 U12580 ( .A1(n10695), .A2(n14313), .B1(n11050), .B2(n14453), .ZN(
        n10765) );
  AOI21_X1 U12581 ( .B1(n10696), .B2(n14710), .A(n10765), .ZN(n11749) );
  AOI21_X1 U12582 ( .B1(n10698), .B2(n11738), .A(n14633), .ZN(n10699) );
  AND2_X1 U12583 ( .A1(n10699), .A2(n10827), .ZN(n11742) );
  AOI21_X1 U12584 ( .B1(n16112), .B2(n11738), .A(n11742), .ZN(n10700) );
  OAI211_X1 U12585 ( .C1(n10701), .C2(n16006), .A(n11749), .B(n10700), .ZN(
        n10950) );
  NAND2_X1 U12586 ( .A1(n10950), .A2(n16156), .ZN(n10702) );
  OAI21_X1 U12587 ( .B1(n16156), .B2(n10703), .A(n10702), .ZN(P2_U3503) );
  INV_X1 U12588 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10705) );
  INV_X1 U12589 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10704) );
  MUX2_X1 U12590 ( .A(n10705), .B(n10704), .S(n10630), .Z(n10707) );
  NAND2_X1 U12591 ( .A1(n10707), .A2(n10706), .ZN(n10817) );
  INV_X1 U12592 ( .A(n10707), .ZN(n10708) );
  NAND2_X1 U12593 ( .A1(n10708), .A2(n10729), .ZN(n10709) );
  NAND2_X1 U12594 ( .A1(n10817), .A2(n10709), .ZN(n10711) );
  INV_X1 U12595 ( .A(n10711), .ZN(n10713) );
  OAI21_X1 U12596 ( .B1(n10713), .B2(n10712), .A(n10818), .ZN(n10727) );
  AND2_X1 U12597 ( .A1(n10717), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10714) );
  NAND2_X1 U12598 ( .A1(n10718), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10803) );
  OAI21_X1 U12599 ( .B1(n10729), .B2(n10714), .A(n10803), .ZN(n10715) );
  OR2_X1 U12600 ( .A1(n10715), .A2(n10705), .ZN(n10804) );
  NAND2_X1 U12601 ( .A1(n10715), .A2(n10705), .ZN(n10716) );
  AND2_X1 U12602 ( .A1(n10804), .A2(n10716), .ZN(n10725) );
  AND2_X1 U12603 ( .A1(n10717), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10719) );
  NAND2_X1 U12604 ( .A1(n10718), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10798) );
  OAI21_X1 U12605 ( .B1(n10729), .B2(n10719), .A(n10798), .ZN(n10720) );
  OR2_X1 U12606 ( .A1(n10720), .A2(n10704), .ZN(n10799) );
  NAND2_X1 U12607 ( .A1(n10720), .A2(n10704), .ZN(n10721) );
  NAND2_X1 U12608 ( .A1(n10799), .A2(n10721), .ZN(n10722) );
  NAND2_X1 U12609 ( .A1(n13722), .A2(n10722), .ZN(n10724) );
  AOI22_X1 U12610 ( .A1(n15521), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10723) );
  OAI211_X1 U12611 ( .C1(n10725), .C2(n15872), .A(n10724), .B(n10723), .ZN(
        n10726) );
  AOI21_X1 U12612 ( .B1(n15863), .B2(n10727), .A(n10726), .ZN(n10728) );
  OAI21_X1 U12613 ( .B1(n10729), .B2(n15856), .A(n10728), .ZN(P3_U3183) );
  INV_X1 U12614 ( .A(n15508), .ZN(n15633) );
  NOR2_X1 U12615 ( .A1(n15508), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10730) );
  OR2_X1 U12616 ( .A1(n10231), .A2(n10730), .ZN(n15632) );
  NOR3_X1 U12617 ( .A1(n10731), .A2(n15633), .A3(n15632), .ZN(n10733) );
  INV_X2 U12618 ( .A(P1_U4016), .ZN(n15076) );
  NOR2_X1 U12619 ( .A1(n15632), .A2(n15508), .ZN(n10732) );
  MUX2_X1 U12620 ( .A(n10732), .B(n15632), .S(n15634), .Z(n15638) );
  NOR3_X1 U12621 ( .A1(n10733), .A2(n15076), .A3(n15638), .ZN(n10787) );
  AND3_X1 U12622 ( .A1(n10736), .A2(n10735), .A3(n10734), .ZN(n10737) );
  NOR3_X1 U12623 ( .A1(n15649), .A2(n10738), .A3(n10737), .ZN(n10747) );
  AOI211_X1 U12624 ( .C1(n10741), .C2(n10740), .A(n10739), .B(n15145), .ZN(
        n10746) );
  INV_X1 U12625 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10744) );
  NAND2_X1 U12626 ( .A1(n15147), .A2(n10742), .ZN(n10743) );
  NAND2_X1 U12627 ( .A1(n7201), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n11289) );
  OAI211_X1 U12628 ( .C1(n15656), .C2(n10744), .A(n10743), .B(n11289), .ZN(
        n10745) );
  OR4_X1 U12629 ( .A1(n10787), .A2(n10747), .A3(n10746), .A4(n10745), .ZN(
        P1_U3247) );
  NAND2_X1 U12630 ( .A1(n10749), .A2(n10748), .ZN(n10841) );
  INV_X1 U12631 ( .A(n10841), .ZN(n10753) );
  XNOR2_X1 U12632 ( .A(n14229), .B(n12099), .ZN(n10751) );
  AND2_X1 U12633 ( .A1(n14374), .A2(n14633), .ZN(n10750) );
  XNOR2_X1 U12634 ( .A(n10751), .B(n10750), .ZN(n10840) );
  XNOR2_X1 U12635 ( .A(n11738), .B(n14188), .ZN(n10754) );
  NAND2_X1 U12636 ( .A1(n14373), .A2(n14633), .ZN(n10755) );
  NAND2_X1 U12637 ( .A1(n10754), .A2(n10755), .ZN(n10930) );
  INV_X1 U12638 ( .A(n10754), .ZN(n10757) );
  INV_X1 U12639 ( .A(n10755), .ZN(n10756) );
  NAND2_X1 U12640 ( .A1(n10757), .A2(n10756), .ZN(n10758) );
  AND2_X1 U12641 ( .A1(n10930), .A2(n10758), .ZN(n10759) );
  OAI21_X1 U12642 ( .B1(n10760), .B2(n10759), .A(n10931), .ZN(n10769) );
  NAND3_X1 U12643 ( .A1(n10763), .A2(n10762), .A3(n10761), .ZN(n10764) );
  AOI22_X1 U12644 ( .A1(n14348), .A2(n10765), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10767) );
  NAND2_X1 U12645 ( .A1(n14358), .A2(n11738), .ZN(n10766) );
  OAI211_X1 U12646 ( .C1(n14351), .C2(n11739), .A(n10767), .B(n10766), .ZN(
        n10768) );
  AOI21_X1 U12647 ( .B1(n14311), .B2(n10769), .A(n10768), .ZN(n10770) );
  INV_X1 U12648 ( .A(n10770), .ZN(P2_U3202) );
  NAND2_X1 U12649 ( .A1(n16156), .A2(n16041), .ZN(n14816) );
  INV_X1 U12650 ( .A(n11156), .ZN(n15886) );
  OAI21_X1 U12651 ( .B1(n14803), .B2(n14710), .A(n15886), .ZN(n10773) );
  NAND2_X1 U12652 ( .A1(n10773), .A2(n10772), .ZN(n15883) );
  NOR2_X1 U12653 ( .A1(n10775), .A2(n10774), .ZN(n15885) );
  NOR2_X1 U12654 ( .A1(n15883), .A2(n15885), .ZN(n11153) );
  NOR2_X1 U12655 ( .A1(n16155), .A2(n11153), .ZN(n10776) );
  AOI21_X1 U12656 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n16155), .A(n10776), .ZN(
        n10777) );
  OAI21_X1 U12657 ( .B1(n11156), .B2(n14816), .A(n10777), .ZN(P2_U3499) );
  XOR2_X1 U12658 ( .A(n10779), .B(n10778), .Z(n10789) );
  OAI21_X1 U12659 ( .B1(n10782), .B2(n10781), .A(n10780), .ZN(n10786) );
  AOI22_X1 U12660 ( .A1(n15639), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n7201), .ZN(n10785) );
  NAND2_X1 U12661 ( .A1(n15147), .A2(n10783), .ZN(n10784) );
  OAI211_X1 U12662 ( .C1(n15145), .C2(n10786), .A(n10785), .B(n10784), .ZN(
        n10788) );
  AOI211_X1 U12663 ( .C1(n15143), .C2(n10789), .A(n10788), .B(n10787), .ZN(
        n10790) );
  INV_X1 U12664 ( .A(n10790), .ZN(P1_U3245) );
  INV_X1 U12665 ( .A(n10792), .ZN(n10793) );
  AOI21_X1 U12666 ( .B1(n10794), .B2(n10791), .A(n10793), .ZN(n10797) );
  AOI22_X1 U12667 ( .A1(n16089), .A2(n15074), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10990), .ZN(n10796) );
  INV_X1 U12668 ( .A(n15049), .ZN(n16087) );
  AOI22_X1 U12669 ( .A1(n15040), .A2(n12674), .B1(n16087), .B2(n10907), .ZN(
        n10795) );
  OAI211_X1 U12670 ( .C1(n10797), .C2(n15042), .A(n10796), .B(n10795), .ZN(
        P1_U3222) );
  INV_X1 U12671 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15896) );
  NAND2_X1 U12672 ( .A1(n10799), .A2(n10798), .ZN(n10800) );
  OAI21_X1 U12673 ( .B1(n10801), .B2(n10800), .A(n7435), .ZN(n10810) );
  INV_X1 U12674 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n13079) );
  NAND2_X1 U12675 ( .A1(n15521), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10802) );
  OAI21_X1 U12676 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n13079), .A(n10802), .ZN(
        n10809) );
  INV_X1 U12677 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11687) );
  MUX2_X1 U12678 ( .A(n11687), .B(P3_REG2_REG_2__SCAN_IN), .S(n10811), .Z(
        n10806) );
  NAND2_X1 U12679 ( .A1(n10804), .A2(n10803), .ZN(n10805) );
  NAND2_X1 U12680 ( .A1(n10806), .A2(n10805), .ZN(n10849) );
  OAI21_X1 U12681 ( .B1(n10806), .B2(n10805), .A(n10849), .ZN(n10807) );
  AND2_X1 U12682 ( .A1(n7465), .A2(n10807), .ZN(n10808) );
  AOI211_X1 U12683 ( .C1(n13722), .C2(n10810), .A(n10809), .B(n10808), .ZN(
        n10824) );
  INV_X1 U12684 ( .A(n10818), .ZN(n10816) );
  INV_X1 U12685 ( .A(n10817), .ZN(n10815) );
  MUX2_X1 U12686 ( .A(n11687), .B(n15896), .S(n10630), .Z(n10812) );
  NAND2_X1 U12687 ( .A1(n10812), .A2(n10811), .ZN(n10867) );
  INV_X1 U12688 ( .A(n10812), .ZN(n10813) );
  NAND2_X1 U12689 ( .A1(n10813), .A2(n10853), .ZN(n10814) );
  AND2_X1 U12690 ( .A1(n10867), .A2(n10814), .ZN(n10819) );
  NOR3_X1 U12691 ( .A1(n10816), .A2(n10815), .A3(n10819), .ZN(n10822) );
  NAND2_X1 U12692 ( .A1(n10818), .A2(n10817), .ZN(n10820) );
  NAND2_X1 U12693 ( .A1(n10820), .A2(n10819), .ZN(n10868) );
  INV_X1 U12694 ( .A(n10868), .ZN(n10821) );
  OAI21_X1 U12695 ( .B1(n10822), .B2(n10821), .A(n15863), .ZN(n10823) );
  OAI211_X1 U12696 ( .C1(n15856), .C2(n10853), .A(n10824), .B(n10823), .ZN(
        P3_U3184) );
  OR2_X1 U12697 ( .A1(n11738), .A2(n14373), .ZN(n10825) );
  XNOR2_X1 U12698 ( .A(n11042), .B(n11048), .ZN(n11773) );
  AOI211_X1 U12699 ( .C1(n14269), .C2(n10827), .A(n14633), .B(n11056), .ZN(
        n11770) );
  AOI21_X1 U12700 ( .B1(n16112), .B2(n14269), .A(n11770), .ZN(n10835) );
  NAND2_X1 U12701 ( .A1(n11738), .A2(n10830), .ZN(n10831) );
  XNOR2_X1 U12702 ( .A(n11049), .B(n11048), .ZN(n10834) );
  NAND2_X1 U12703 ( .A1(n14373), .A2(n14525), .ZN(n10833) );
  NAND2_X1 U12704 ( .A1(n14371), .A2(n14338), .ZN(n10832) );
  NAND2_X1 U12705 ( .A1(n10833), .A2(n10832), .ZN(n14268) );
  AOI21_X1 U12706 ( .B1(n10834), .B2(n14710), .A(n14268), .ZN(n11766) );
  OAI211_X1 U12707 ( .C1(n11773), .C2(n16006), .A(n10835), .B(n11766), .ZN(
        n10954) );
  NAND2_X1 U12708 ( .A1(n10954), .A2(n16156), .ZN(n10836) );
  OAI21_X1 U12709 ( .B1(n16156), .B2(n10509), .A(n10836), .ZN(P2_U3504) );
  INV_X1 U12710 ( .A(n13688), .ZN(n13695) );
  INV_X1 U12711 ( .A(SI_16_), .ZN(n10839) );
  INV_X1 U12712 ( .A(n10837), .ZN(n10838) );
  OAI222_X1 U12713 ( .A1(P3_U3151), .A2(n13695), .B1(n14155), .B2(n10839), 
        .C1(n14158), .C2(n10838), .ZN(P3_U3279) );
  XNOR2_X1 U12714 ( .A(n10841), .B(n10840), .ZN(n10847) );
  INV_X1 U12715 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n14385) );
  AOI22_X1 U12716 ( .A1(n14348), .A2(n10842), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10843) );
  OAI21_X1 U12717 ( .B1(n10844), .B2(n14309), .A(n10843), .ZN(n10845) );
  AOI21_X1 U12718 ( .B1(n14339), .B2(n14385), .A(n10845), .ZN(n10846) );
  OAI21_X1 U12719 ( .B1(n10847), .B2(n14353), .A(n10846), .ZN(P2_U3190) );
  INV_X1 U12720 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10852) );
  NAND2_X1 U12721 ( .A1(n10853), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10848) );
  INV_X1 U12722 ( .A(n10878), .ZN(n10850) );
  AOI21_X1 U12723 ( .B1(n10852), .B2(n10851), .A(n10850), .ZN(n10859) );
  OAI21_X1 U12724 ( .B1(n10854), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10884), .ZN(
        n10855) );
  NAND2_X1 U12725 ( .A1(n13722), .A2(n10855), .ZN(n10858) );
  NOR2_X1 U12726 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10856), .ZN(n11210) );
  AOI21_X1 U12727 ( .B1(n15521), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n11210), .ZN(
        n10857) );
  OAI211_X1 U12728 ( .C1(n10859), .C2(n15872), .A(n10858), .B(n10857), .ZN(
        n10871) );
  NAND2_X1 U12729 ( .A1(n10868), .A2(n10867), .ZN(n10864) );
  INV_X1 U12730 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10860) );
  MUX2_X1 U12731 ( .A(n10852), .B(n10860), .S(n10630), .Z(n10861) );
  NAND2_X1 U12732 ( .A1(n10861), .A2(n10872), .ZN(n10890) );
  INV_X1 U12733 ( .A(n10861), .ZN(n10862) );
  NAND2_X1 U12734 ( .A1(n10862), .A2(n7763), .ZN(n10863) );
  AND2_X1 U12735 ( .A1(n10890), .A2(n10863), .ZN(n10865) );
  NAND2_X1 U12736 ( .A1(n10864), .A2(n10865), .ZN(n10891) );
  INV_X1 U12737 ( .A(n10865), .ZN(n10866) );
  NAND3_X1 U12738 ( .A1(n10868), .A2(n10867), .A3(n10866), .ZN(n10869) );
  AOI21_X1 U12739 ( .B1(n10891), .B2(n10869), .A(n15843), .ZN(n10870) );
  AOI211_X1 U12740 ( .C1(n13754), .C2(n10872), .A(n10871), .B(n10870), .ZN(
        n10873) );
  INV_X1 U12741 ( .A(n10873), .ZN(P3_U3185) );
  INV_X1 U12742 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11644) );
  MUX2_X1 U12743 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n11644), .S(n10974), .Z(
        n10875) );
  NAND2_X1 U12744 ( .A1(n10874), .A2(n10875), .ZN(n10976) );
  INV_X1 U12745 ( .A(n10875), .ZN(n10877) );
  NAND3_X1 U12746 ( .A1(n10878), .A2(n10877), .A3(n10876), .ZN(n10879) );
  AOI21_X1 U12747 ( .B1(n10976), .B2(n10879), .A(n15872), .ZN(n10889) );
  INV_X1 U12748 ( .A(n10880), .ZN(n10882) );
  INV_X1 U12749 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10881) );
  MUX2_X1 U12750 ( .A(n10881), .B(P3_REG1_REG_4__SCAN_IN), .S(n10974), .Z(
        n10883) );
  NAND3_X1 U12751 ( .A1(n10884), .A2(n10883), .A3(n10882), .ZN(n10885) );
  AOI21_X1 U12752 ( .B1(n7378), .B2(n10885), .A(n15866), .ZN(n10888) );
  INV_X1 U12753 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n10886) );
  NOR2_X1 U12754 ( .A1(n15853), .A2(n10886), .ZN(n10887) );
  INV_X1 U12755 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n12993) );
  NOR2_X1 U12756 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12993), .ZN(n11390) );
  NOR4_X1 U12757 ( .A1(n10889), .A2(n10888), .A3(n10887), .A4(n11390), .ZN(
        n10896) );
  NAND2_X1 U12758 ( .A1(n10891), .A2(n10890), .ZN(n10893) );
  MUX2_X1 U12759 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n10630), .Z(n10962) );
  INV_X1 U12760 ( .A(n10974), .ZN(n10963) );
  XNOR2_X1 U12761 ( .A(n10962), .B(n10963), .ZN(n10892) );
  NAND2_X1 U12762 ( .A1(n10893), .A2(n10892), .ZN(n10966) );
  OAI21_X1 U12763 ( .B1(n10893), .B2(n10892), .A(n10966), .ZN(n10894) );
  NAND2_X1 U12764 ( .A1(n10894), .A2(n15863), .ZN(n10895) );
  OAI211_X1 U12765 ( .C1(n15856), .C2(n10974), .A(n10896), .B(n10895), .ZN(
        P3_U3186) );
  INV_X1 U12766 ( .A(n10897), .ZN(n10899) );
  AND3_X1 U12767 ( .A1(n10899), .A2(n10898), .A3(n11018), .ZN(n10900) );
  AND2_X1 U12768 ( .A1(n10900), .A2(n12911), .ZN(n10918) );
  INV_X1 U12769 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10916) );
  OR2_X1 U12770 ( .A1(n7228), .A2(n11027), .ZN(n10901) );
  NAND2_X1 U12771 ( .A1(n8048), .A2(n7620), .ZN(n12675) );
  NAND2_X1 U12772 ( .A1(n15075), .A2(n12674), .ZN(n10905) );
  INV_X1 U12773 ( .A(n10907), .ZN(n10906) );
  NAND2_X1 U12774 ( .A1(n10906), .A2(n15878), .ZN(n11062) );
  XNOR2_X1 U12775 ( .A(n12683), .B(n11062), .ZN(n11036) );
  NAND2_X1 U12776 ( .A1(n10907), .A2(n15878), .ZN(n10908) );
  OAI21_X1 U12777 ( .B1(n10909), .B2(n10908), .A(n10993), .ZN(n11034) );
  OR2_X1 U12778 ( .A1(n12676), .A2(n12672), .ZN(n10910) );
  NAND2_X1 U12779 ( .A1(n14954), .A2(n10910), .ZN(n11020) );
  NAND2_X1 U12780 ( .A1(n15150), .A2(n12849), .ZN(n16021) );
  NAND2_X1 U12781 ( .A1(n12674), .A2(n15878), .ZN(n10911) );
  AND3_X1 U12782 ( .A1(n11005), .A2(n15445), .A3(n10911), .ZN(n11026) );
  NAND2_X1 U12783 ( .A1(n15074), .A2(n15376), .ZN(n11023) );
  NAND2_X1 U12784 ( .A1(n10907), .A2(n16030), .ZN(n10912) );
  OAI211_X1 U12785 ( .C1(n10903), .C2(n16123), .A(n11023), .B(n10912), .ZN(
        n10913) );
  AOI211_X1 U12786 ( .C1(n11034), .C2(n16139), .A(n11026), .B(n10913), .ZN(
        n10914) );
  OAI21_X1 U12787 ( .B1(n16136), .B2(n11036), .A(n10914), .ZN(n10919) );
  NAND2_X1 U12788 ( .A1(n10919), .A2(n16147), .ZN(n10915) );
  OAI21_X1 U12789 ( .B1(n16147), .B2(n10916), .A(n10915), .ZN(P1_U3462) );
  AND2_X2 U12790 ( .A1(n10918), .A2(n10917), .ZN(n16143) );
  NAND2_X1 U12791 ( .A1(n10919), .A2(n16143), .ZN(n10920) );
  OAI21_X1 U12792 ( .B1(n16143), .B2(n10921), .A(n10920), .ZN(P1_U3529) );
  INV_X1 U12793 ( .A(n15595), .ZN(n12319) );
  INV_X1 U12794 ( .A(n10922), .ZN(n10924) );
  OAI222_X1 U12795 ( .A1(P2_U3088), .A2(n12319), .B1(n14869), .B2(n10924), 
        .C1(n10923), .C2(n14871), .ZN(P2_U3311) );
  INV_X1 U12796 ( .A(n15106), .ZN(n15110) );
  OAI222_X1 U12797 ( .A1(n15512), .A2(n10925), .B1(n15510), .B2(n10924), .C1(
        n15110), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12798 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10927) );
  INV_X1 U12799 ( .A(n10926), .ZN(n10928) );
  INV_X1 U12800 ( .A(n11558), .ZN(n11102) );
  OAI222_X1 U12801 ( .A1(n14871), .A2(n10927), .B1(n14869), .B2(n10928), .C1(
        P2_U3088), .C2(n11102), .ZN(P2_U3313) );
  INV_X1 U12802 ( .A(n12488), .ZN(n12482) );
  OAI222_X1 U12803 ( .A1(n11951), .A2(n10929), .B1(n15510), .B2(n10928), .C1(
        n7201), .C2(n12482), .ZN(P1_U3341) );
  XNOR2_X1 U12804 ( .A(n14269), .B(n14188), .ZN(n10932) );
  NAND2_X1 U12805 ( .A1(n14372), .A2(n14633), .ZN(n10933) );
  NAND2_X1 U12806 ( .A1(n10932), .A2(n10933), .ZN(n10937) );
  INV_X1 U12807 ( .A(n10932), .ZN(n10935) );
  INV_X1 U12808 ( .A(n10933), .ZN(n10934) );
  NAND2_X1 U12809 ( .A1(n10935), .A2(n10934), .ZN(n10936) );
  AND2_X1 U12810 ( .A1(n10937), .A2(n10936), .ZN(n14265) );
  XNOR2_X1 U12811 ( .A(n11400), .B(n14188), .ZN(n11216) );
  NAND2_X1 U12812 ( .A1(n14371), .A2(n14633), .ZN(n11217) );
  XNOR2_X1 U12813 ( .A(n11216), .B(n11217), .ZN(n11215) );
  XNOR2_X1 U12814 ( .A(n11214), .B(n11215), .ZN(n10944) );
  INV_X1 U12815 ( .A(n11776), .ZN(n10941) );
  NAND2_X1 U12816 ( .A1(n14372), .A2(n14525), .ZN(n10939) );
  NAND2_X1 U12817 ( .A1(n14370), .A2(n14338), .ZN(n10938) );
  AND2_X1 U12818 ( .A1(n10939), .A2(n10938), .ZN(n11053) );
  NAND2_X1 U12819 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n15587) );
  OAI21_X1 U12820 ( .B1(n14341), .B2(n11053), .A(n15587), .ZN(n10940) );
  AOI21_X1 U12821 ( .B1(n10941), .B2(n14339), .A(n10940), .ZN(n10943) );
  NAND2_X1 U12822 ( .A1(n14358), .A2(n11400), .ZN(n10942) );
  OAI211_X1 U12823 ( .C1(n10944), .C2(n14353), .A(n10943), .B(n10942), .ZN(
        P2_U3211) );
  NAND2_X1 U12824 ( .A1(n16160), .A2(n10946), .ZN(n10947) );
  OAI21_X1 U12825 ( .B1(n16160), .B2(n8897), .A(n10947), .ZN(P2_U3433) );
  NAND2_X1 U12826 ( .A1(n16160), .A2(n10948), .ZN(n10949) );
  OAI21_X1 U12827 ( .B1(n16160), .B2(n8911), .A(n10949), .ZN(P2_U3436) );
  NAND2_X1 U12828 ( .A1(n10950), .A2(n16160), .ZN(n10951) );
  OAI21_X1 U12829 ( .B1(n16160), .B2(n8977), .A(n10951), .ZN(P2_U3442) );
  NAND2_X1 U12830 ( .A1(n10952), .A2(n16160), .ZN(n10953) );
  OAI21_X1 U12831 ( .B1(n16160), .B2(n8944), .A(n10953), .ZN(P2_U3439) );
  NAND2_X1 U12832 ( .A1(n10954), .A2(n16160), .ZN(n10955) );
  OAI21_X1 U12833 ( .B1(n16160), .B2(n8996), .A(n10955), .ZN(P2_U3445) );
  NOR2_X1 U12834 ( .A1(n13351), .A2(P3_U3151), .ZN(n11190) );
  INV_X1 U12835 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n12574) );
  NAND2_X1 U12836 ( .A1(n13588), .A2(n12575), .ZN(n13382) );
  INV_X1 U12837 ( .A(n13382), .ZN(n10956) );
  NOR2_X1 U12838 ( .A1(n11264), .A2(n10956), .ZN(n13524) );
  INV_X1 U12839 ( .A(n13524), .ZN(n10958) );
  OAI22_X1 U12840 ( .A1(n11674), .A2(n13335), .B1(n12575), .B2(n13354), .ZN(
        n10957) );
  AOI21_X1 U12841 ( .B1(n10958), .B2(n13343), .A(n10957), .ZN(n10959) );
  OAI21_X1 U12842 ( .B1(n11190), .B2(n12574), .A(n10959), .ZN(P3_U3172) );
  INV_X1 U12843 ( .A(n10960), .ZN(n10961) );
  OAI222_X1 U12844 ( .A1(P3_U3151), .A2(n13710), .B1(n14155), .B2(n13119), 
        .C1(n14158), .C2(n10961), .ZN(P3_U3278) );
  INV_X1 U12845 ( .A(n10962), .ZN(n10964) );
  NAND2_X1 U12846 ( .A1(n10964), .A2(n10963), .ZN(n10965) );
  NAND2_X1 U12847 ( .A1(n10966), .A2(n10965), .ZN(n11131) );
  MUX2_X1 U12848 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n10630), .Z(n10967) );
  NAND2_X1 U12849 ( .A1(n10967), .A2(n10977), .ZN(n11130) );
  INV_X1 U12850 ( .A(n10967), .ZN(n10968) );
  NAND2_X1 U12851 ( .A1(n10968), .A2(n7780), .ZN(n11132) );
  NAND2_X1 U12852 ( .A1(n11130), .A2(n11132), .ZN(n10969) );
  XNOR2_X1 U12853 ( .A(n11131), .B(n10969), .ZN(n10983) );
  INV_X1 U12854 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10971) );
  AOI21_X1 U12855 ( .B1(n10971), .B2(n10970), .A(n11144), .ZN(n10973) );
  NOR2_X1 U12856 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8391), .ZN(n11480) );
  AOI21_X1 U12857 ( .B1(n15521), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11480), .ZN(
        n10972) );
  OAI21_X1 U12858 ( .B1(n10973), .B2(n15866), .A(n10972), .ZN(n10981) );
  NAND2_X1 U12859 ( .A1(n10974), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10975) );
  INV_X1 U12860 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11660) );
  NAND2_X1 U12861 ( .A1(n10978), .A2(n11660), .ZN(n10979) );
  AOI21_X1 U12862 ( .B1(n11140), .B2(n10979), .A(n15872), .ZN(n10980) );
  AOI211_X1 U12863 ( .C1(n13754), .C2(n7780), .A(n10981), .B(n10980), .ZN(
        n10982) );
  OAI21_X1 U12864 ( .B1(n10983), .B2(n15843), .A(n10982), .ZN(P3_U3187) );
  NAND2_X1 U12865 ( .A1(n15075), .A2(n16030), .ZN(n10985) );
  NAND2_X1 U12866 ( .A1(n15073), .A2(n15376), .ZN(n10984) );
  AND2_X1 U12867 ( .A1(n10985), .A2(n10984), .ZN(n11002) );
  OAI21_X1 U12868 ( .B1(n10988), .B2(n10987), .A(n10986), .ZN(n10989) );
  NAND2_X1 U12869 ( .A1(n10989), .A2(n16093), .ZN(n10992) );
  AOI22_X1 U12870 ( .A1(n15040), .A2(n12690), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10990), .ZN(n10991) );
  OAI211_X1 U12871 ( .C1(n11002), .C2(n15026), .A(n10992), .B(n10991), .ZN(
        P1_U3237) );
  INV_X1 U12872 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n11008) );
  INV_X1 U12873 ( .A(n12690), .ZN(n12691) );
  NAND2_X1 U12874 ( .A1(n15074), .A2(n12691), .ZN(n10995) );
  OAI21_X1 U12875 ( .B1(n10996), .B2(n11001), .A(n11197), .ZN(n10997) );
  INV_X1 U12876 ( .A(n10997), .ZN(n11111) );
  NAND2_X1 U12877 ( .A1(n12683), .A2(n10998), .ZN(n11000) );
  NAND2_X1 U12878 ( .A1(n10904), .A2(n12674), .ZN(n10999) );
  INV_X1 U12879 ( .A(n11001), .ZN(n12854) );
  INV_X1 U12880 ( .A(n11002), .ZN(n11003) );
  AOI21_X1 U12881 ( .B1(n11004), .B2(n16119), .A(n11003), .ZN(n11116) );
  AOI211_X1 U12882 ( .C1(n12690), .C2(n11005), .A(n15974), .B(n11199), .ZN(
        n11114) );
  AOI21_X1 U12883 ( .B1(n16134), .B2(n12690), .A(n11114), .ZN(n11006) );
  OAI211_X1 U12884 ( .C1(n11111), .C2(n15469), .A(n11116), .B(n11006), .ZN(
        n11009) );
  NAND2_X1 U12885 ( .A1(n11009), .A2(n16147), .ZN(n11007) );
  OAI21_X1 U12886 ( .B1(n16147), .B2(n11008), .A(n11007), .ZN(P1_U3465) );
  NAND2_X1 U12887 ( .A1(n11009), .A2(n16143), .ZN(n11010) );
  OAI21_X1 U12888 ( .B1(n16143), .B2(n11011), .A(n11010), .ZN(P1_U3530) );
  INV_X1 U12889 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11013) );
  INV_X1 U12890 ( .A(n11012), .ZN(n11014) );
  INV_X1 U12891 ( .A(n12322), .ZN(n12328) );
  OAI222_X1 U12892 ( .A1(n14871), .A2(n11013), .B1(n14869), .B2(n11014), .C1(
        P2_U3088), .C2(n12328), .ZN(P2_U3312) );
  INV_X1 U12893 ( .A(n12483), .ZN(n15648) );
  OAI222_X1 U12894 ( .A1(n15512), .A2(n11015), .B1(n15510), .B2(n11014), .C1(
        n7201), .C2(n15648), .ZN(P1_U3340) );
  NAND3_X1 U12895 ( .A1(n11017), .A2(n12911), .A3(n11016), .ZN(n15169) );
  INV_X1 U12896 ( .A(n11018), .ZN(n11019) );
  NOR2_X1 U12897 ( .A1(n16001), .A2(n16136), .ZN(n15389) );
  INV_X1 U12898 ( .A(n15389), .ZN(n15371) );
  INV_X1 U12899 ( .A(n11020), .ZN(n11021) );
  INV_X1 U12900 ( .A(n15392), .ZN(n15355) );
  MUX2_X1 U12901 ( .A(n11023), .B(n11022), .S(n16001), .Z(n11032) );
  NAND2_X1 U12902 ( .A1(n7218), .A2(n16030), .ZN(n15173) );
  OAI22_X1 U12903 ( .A1(n15173), .A2(n10906), .B1(n11024), .B2(n15377), .ZN(
        n11025) );
  INV_X1 U12904 ( .A(n11025), .ZN(n11031) );
  NOR2_X2 U12905 ( .A1(n15169), .A2(n15150), .ZN(n15368) );
  NAND2_X1 U12906 ( .A1(n11026), .A2(n15368), .ZN(n11030) );
  NAND2_X1 U12907 ( .A1(n11419), .A2(n7620), .ZN(n12897) );
  INV_X1 U12908 ( .A(n12897), .ZN(n12887) );
  AND2_X1 U12909 ( .A1(n12887), .A2(n11027), .ZN(n11028) );
  OR2_X1 U12910 ( .A1(n15365), .A2(n10903), .ZN(n11029) );
  NAND4_X1 U12911 ( .A1(n11032), .A2(n11031), .A3(n11030), .A4(n11029), .ZN(
        n11033) );
  AOI21_X1 U12912 ( .B1(n15355), .B2(n11034), .A(n11033), .ZN(n11035) );
  OAI21_X1 U12913 ( .B1(n15371), .B2(n11036), .A(n11035), .ZN(P1_U3292) );
  INV_X1 U12914 ( .A(n11037), .ZN(n11039) );
  INV_X1 U12915 ( .A(n15124), .ZN(n15122) );
  OAI222_X1 U12916 ( .A1(n15512), .A2(n11038), .B1(n15510), .B2(n11039), .C1(
        P1_U3086), .C2(n15122), .ZN(P1_U3338) );
  INV_X1 U12917 ( .A(n12337), .ZN(n14440) );
  OAI222_X1 U12918 ( .A1(n14871), .A2(n11040), .B1(n14869), .B2(n11039), .C1(
        P2_U3088), .C2(n14440), .ZN(P2_U3310) );
  INV_X1 U12919 ( .A(n11048), .ZN(n11041) );
  NAND2_X1 U12920 ( .A1(n11042), .A2(n11041), .ZN(n11044) );
  OR2_X1 U12921 ( .A1(n14269), .A2(n14372), .ZN(n11043) );
  INV_X1 U12922 ( .A(n11394), .ZN(n11045) );
  OAI21_X1 U12923 ( .B1(n11046), .B2(n11045), .A(n11402), .ZN(n11047) );
  INV_X1 U12924 ( .A(n11047), .ZN(n11782) );
  NAND2_X1 U12925 ( .A1(n14269), .A2(n11050), .ZN(n11051) );
  NAND2_X1 U12926 ( .A1(n11052), .A2(n11051), .ZN(n11395) );
  XNOR2_X1 U12927 ( .A(n11395), .B(n11394), .ZN(n11055) );
  INV_X1 U12928 ( .A(n11053), .ZN(n11054) );
  AOI21_X1 U12929 ( .B1(n11055), .B2(n14710), .A(n11054), .ZN(n11774) );
  INV_X1 U12930 ( .A(n11056), .ZN(n11057) );
  INV_X1 U12931 ( .A(n11400), .ZN(n11777) );
  AOI211_X1 U12932 ( .C1(n11400), .C2(n11057), .A(n14633), .B(n11409), .ZN(
        n11779) );
  AOI21_X1 U12933 ( .B1(n16112), .B2(n11400), .A(n11779), .ZN(n11058) );
  OAI211_X1 U12934 ( .C1(n11782), .C2(n16006), .A(n11774), .B(n11058), .ZN(
        n11078) );
  NAND2_X1 U12935 ( .A1(n11078), .A2(n16156), .ZN(n11059) );
  OAI21_X1 U12936 ( .B1(n16156), .B2(n10511), .A(n11059), .ZN(P2_U3505) );
  INV_X1 U12937 ( .A(n12928), .ZN(n16026) );
  NAND2_X1 U12938 ( .A1(n10907), .A2(n11060), .ZN(n11061) );
  NAND2_X1 U12939 ( .A1(n11062), .A2(n11061), .ZN(n11064) );
  OAI21_X1 U12940 ( .B1(n16026), .B2(n16119), .A(n11064), .ZN(n11063) );
  OAI21_X1 U12941 ( .B1(n10904), .B2(n15359), .A(n11063), .ZN(n15877) );
  INV_X1 U12942 ( .A(n11064), .ZN(n15875) );
  NAND2_X1 U12943 ( .A1(n15150), .A2(n11065), .ZN(n12852) );
  INV_X1 U12944 ( .A(n12852), .ZN(n11066) );
  NAND2_X1 U12945 ( .A1(n7218), .A2(n11066), .ZN(n12932) );
  INV_X1 U12946 ( .A(n15365), .ZN(n15991) );
  AND2_X1 U12947 ( .A1(n15368), .A2(n15445), .ZN(n15347) );
  OAI21_X1 U12948 ( .B1(n15991), .B2(n15347), .A(n15878), .ZN(n11068) );
  AOI22_X1 U12949 ( .A1(n16001), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n15990), .ZN(n11067) );
  OAI211_X1 U12950 ( .C1(n15875), .C2(n12932), .A(n11068), .B(n11067), .ZN(
        n11069) );
  AOI21_X1 U12951 ( .B1(n7218), .B2(n15877), .A(n11069), .ZN(n11070) );
  INV_X1 U12952 ( .A(n11070), .ZN(P1_U3293) );
  INV_X1 U12953 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11787) );
  OAI21_X1 U12954 ( .B1(n11073), .B2(n11072), .A(n11071), .ZN(n11074) );
  NAND2_X1 U12955 ( .A1(n11074), .A2(n13343), .ZN(n11077) );
  OAI22_X1 U12956 ( .A1(n11905), .A2(n13335), .B1(n13380), .B2(n13354), .ZN(
        n11075) );
  AOI21_X1 U12957 ( .B1(n13318), .B2(n13588), .A(n11075), .ZN(n11076) );
  OAI211_X1 U12958 ( .C1(n11190), .C2(n11787), .A(n11077), .B(n11076), .ZN(
        P3_U3162) );
  NAND2_X1 U12959 ( .A1(n11078), .A2(n16160), .ZN(n11079) );
  OAI21_X1 U12960 ( .B1(n16117), .B2(n9022), .A(n11079), .ZN(P2_U3448) );
  NAND2_X1 U12961 ( .A1(n11080), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U12962 ( .A1(n11082), .A2(n11081), .ZN(n15621) );
  MUX2_X1 U12963 ( .A(n9181), .B(P2_REG1_REG_12__SCAN_IN), .S(n15626), .Z(
        n15620) );
  OR2_X1 U12964 ( .A1(n15626), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11083) );
  NAND2_X1 U12965 ( .A1(n11098), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11084) );
  OAI21_X1 U12966 ( .B1(n11098), .B2(P2_REG1_REG_13__SCAN_IN), .A(n11084), 
        .ZN(n15604) );
  NAND2_X1 U12967 ( .A1(n15605), .A2(n15604), .ZN(n15603) );
  NAND2_X1 U12968 ( .A1(n15609), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11085) );
  NAND2_X1 U12969 ( .A1(n15603), .A2(n11085), .ZN(n11090) );
  OR2_X1 U12970 ( .A1(n11558), .A2(n11086), .ZN(n11088) );
  NAND2_X1 U12971 ( .A1(n11558), .A2(n11086), .ZN(n11087) );
  NAND2_X1 U12972 ( .A1(n11088), .A2(n11087), .ZN(n11089) );
  OAI21_X1 U12973 ( .B1(n11090), .B2(n11089), .A(n15602), .ZN(n11107) );
  NOR2_X1 U12974 ( .A1(n11098), .A2(n12131), .ZN(n11097) );
  INV_X1 U12975 ( .A(n11097), .ZN(n11099) );
  AOI21_X1 U12976 ( .B1(n11093), .B2(n11092), .A(n11091), .ZN(n11094) );
  NOR2_X1 U12977 ( .A1(n15626), .A2(n11094), .ZN(n11096) );
  XOR2_X1 U12978 ( .A(n11095), .B(n11094), .Z(n15618) );
  NOR2_X1 U12979 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n15618), .ZN(n15617) );
  NOR2_X1 U12980 ( .A1(n11096), .A2(n15617), .ZN(n15613) );
  AOI21_X1 U12981 ( .B1(n12131), .B2(n11098), .A(n11097), .ZN(n15612) );
  NAND2_X1 U12982 ( .A1(n15613), .A2(n15612), .ZN(n15610) );
  NAND2_X1 U12983 ( .A1(n11099), .A2(n15610), .ZN(n11101) );
  AOI22_X1 U12984 ( .A1(n11558), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12122), 
        .B2(n11102), .ZN(n11100) );
  NAND2_X1 U12985 ( .A1(n11100), .A2(n11101), .ZN(n11552) );
  OAI211_X1 U12986 ( .C1(n11101), .C2(n11100), .A(n15611), .B(n11552), .ZN(
        n11106) );
  NOR2_X1 U12987 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12270), .ZN(n11104) );
  NOR2_X1 U12988 ( .A1(n15543), .A2(n11102), .ZN(n11103) );
  AOI211_X1 U12989 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n15619), .A(n11104), 
        .B(n11103), .ZN(n11105) );
  OAI211_X1 U12990 ( .C1(n11557), .C2(n11107), .A(n11106), .B(n11105), .ZN(
        P2_U3228) );
  INV_X1 U12991 ( .A(n13749), .ZN(n13716) );
  INV_X1 U12992 ( .A(n11108), .ZN(n11109) );
  OAI222_X1 U12993 ( .A1(P3_U3151), .A2(n13716), .B1(n14155), .B2(n13093), 
        .C1(n14158), .C2(n11109), .ZN(P3_U3277) );
  AOI22_X1 U12994 ( .A1(n16001), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n15990), .ZN(n11110) );
  OAI21_X1 U12995 ( .B1(n15365), .B2(n12691), .A(n11110), .ZN(n11113) );
  NOR2_X1 U12996 ( .A1(n11111), .A2(n15392), .ZN(n11112) );
  AOI211_X1 U12997 ( .C1(n11114), .C2(n15368), .A(n11113), .B(n11112), .ZN(
        n11115) );
  OAI21_X1 U12998 ( .B1(n16001), .B2(n11116), .A(n11115), .ZN(P1_U3291) );
  OR3_X1 U12999 ( .A1(n13524), .A2(n15940), .A3(n11117), .ZN(n11119) );
  NAND2_X1 U13000 ( .A1(n13586), .A2(n13996), .ZN(n11118) );
  NAND2_X1 U13001 ( .A1(n11119), .A2(n11118), .ZN(n12573) );
  NAND2_X1 U13002 ( .A1(n11176), .A2(n11258), .ZN(n11120) );
  OR2_X1 U13003 ( .A1(n11121), .A2(n11120), .ZN(n11126) );
  NAND2_X1 U13004 ( .A1(n13564), .A2(n11122), .ZN(n11123) );
  NAND2_X1 U13005 ( .A1(n11124), .A2(n11123), .ZN(n11125) );
  INV_X1 U13006 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11127) );
  OAI22_X1 U13007 ( .A1(n14142), .A2(n12575), .B1(n11127), .B2(n16065), .ZN(
        n11128) );
  AOI21_X1 U13008 ( .B1(n12573), .B2(n16065), .A(n11128), .ZN(n11129) );
  INV_X1 U13009 ( .A(n11129), .ZN(P3_U3390) );
  NAND2_X1 U13010 ( .A1(n11131), .A2(n11130), .ZN(n11133) );
  NAND2_X1 U13011 ( .A1(n11133), .A2(n11132), .ZN(n11327) );
  INV_X1 U13012 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11894) );
  INV_X1 U13013 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15944) );
  MUX2_X1 U13014 ( .A(n11894), .B(n15944), .S(n10630), .Z(n11134) );
  INV_X1 U13015 ( .A(n11340), .ZN(n11336) );
  AND2_X1 U13016 ( .A1(n11134), .A2(n11336), .ZN(n11326) );
  INV_X1 U13017 ( .A(n11326), .ZN(n11136) );
  INV_X1 U13018 ( .A(n11134), .ZN(n11135) );
  NAND2_X1 U13019 ( .A1(n11135), .A2(n11340), .ZN(n11328) );
  NAND2_X1 U13020 ( .A1(n11136), .A2(n11328), .ZN(n11137) );
  XNOR2_X1 U13021 ( .A(n11327), .B(n11137), .ZN(n11152) );
  XNOR2_X1 U13022 ( .A(n11340), .B(P3_REG2_REG_6__SCAN_IN), .ZN(n11139) );
  AOI21_X1 U13023 ( .B1(n11140), .B2(n11138), .A(n11139), .ZN(n11339) );
  INV_X1 U13024 ( .A(n11339), .ZN(n11142) );
  NAND3_X1 U13025 ( .A1(n11140), .A2(n11139), .A3(n11138), .ZN(n11141) );
  AOI21_X1 U13026 ( .B1(n11142), .B2(n11141), .A(n15872), .ZN(n11150) );
  XNOR2_X1 U13027 ( .A(n11340), .B(n15944), .ZN(n11143) );
  INV_X1 U13028 ( .A(n11335), .ZN(n11147) );
  NOR3_X1 U13029 ( .A1(n11145), .A2(n11144), .A3(n11143), .ZN(n11146) );
  OAI21_X1 U13030 ( .B1(n11147), .B2(n11146), .A(n13722), .ZN(n11148) );
  NAND2_X1 U13031 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n11939) );
  OAI211_X1 U13032 ( .C1(n15707), .C2(n15853), .A(n11148), .B(n11939), .ZN(
        n11149) );
  AOI211_X1 U13033 ( .C1(n13754), .C2(n11336), .A(n11150), .B(n11149), .ZN(
        n11151) );
  OAI21_X1 U13034 ( .B1(n11152), .B2(n15843), .A(n11151), .ZN(P3_U3188) );
  NAND2_X1 U13035 ( .A1(n16160), .A2(n16041), .ZN(n14849) );
  INV_X1 U13036 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n11154) );
  MUX2_X1 U13037 ( .A(n11154), .B(n11153), .S(n16117), .Z(n11155) );
  OAI21_X1 U13038 ( .B1(n11156), .B2(n14849), .A(n11155), .ZN(P2_U3430) );
  INV_X1 U13039 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11157) );
  MUX2_X1 U13040 ( .A(n11157), .B(P1_REG1_REG_10__SCAN_IN), .S(n11236), .Z(
        n11162) );
  OAI21_X1 U13041 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n11159), .A(n11158), .ZN(
        n15078) );
  INV_X1 U13042 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11160) );
  MUX2_X1 U13043 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n11160), .S(n15088), .Z(
        n15079) );
  NAND2_X1 U13044 ( .A1(n15078), .A2(n15079), .ZN(n15077) );
  OAI21_X1 U13045 ( .B1(n15088), .B2(P1_REG1_REG_9__SCAN_IN), .A(n15077), .ZN(
        n11161) );
  NOR2_X1 U13046 ( .A1(n11161), .A2(n11162), .ZN(n11235) );
  AOI211_X1 U13047 ( .C1(n11162), .C2(n11161), .A(n15145), .B(n11235), .ZN(
        n11173) );
  NOR2_X1 U13048 ( .A1(n11164), .A2(n11163), .ZN(n15082) );
  INV_X1 U13049 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11936) );
  MUX2_X1 U13050 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11936), .S(n15088), .Z(
        n11165) );
  OAI21_X1 U13051 ( .B1(n15087), .B2(n15082), .A(n11165), .ZN(n15085) );
  NAND2_X1 U13052 ( .A1(n15088), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n11167) );
  INV_X1 U13053 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11240) );
  MUX2_X1 U13054 ( .A(n11240), .B(P1_REG2_REG_10__SCAN_IN), .S(n11236), .Z(
        n11166) );
  AOI21_X1 U13055 ( .B1(n15085), .B2(n11167), .A(n11166), .ZN(n11247) );
  INV_X1 U13056 ( .A(n11247), .ZN(n11169) );
  NAND3_X1 U13057 ( .A1(n15085), .A2(n11167), .A3(n11166), .ZN(n11168) );
  NAND3_X1 U13058 ( .A1(n11169), .A2(n15143), .A3(n11168), .ZN(n11171) );
  AND2_X1 U13059 ( .A1(n7201), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n12085) );
  AOI21_X1 U13060 ( .B1(n15639), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n12085), 
        .ZN(n11170) );
  OAI211_X1 U13061 ( .C1(n15647), .C2(n11241), .A(n11171), .B(n11170), .ZN(
        n11172) );
  OR2_X1 U13062 ( .A1(n11173), .A2(n11172), .ZN(P1_U3253) );
  XNOR2_X1 U13063 ( .A(n11174), .B(n11635), .ZN(n11178) );
  AND2_X1 U13064 ( .A1(n11176), .A2(n11175), .ZN(n11177) );
  AND2_X1 U13065 ( .A1(n11178), .A2(n11177), .ZN(n11638) );
  NAND2_X1 U13066 ( .A1(n11179), .A2(n11269), .ZN(n11260) );
  NAND2_X1 U13067 ( .A1(n11260), .A2(n13388), .ZN(n11183) );
  AND2_X1 U13068 ( .A1(n11183), .A2(n13565), .ZN(n11632) );
  AND2_X1 U13069 ( .A1(n11632), .A2(n11180), .ZN(n11634) );
  NAND2_X1 U13070 ( .A1(n11181), .A2(n11259), .ZN(n11182) );
  NAND2_X1 U13071 ( .A1(n11183), .A2(n11182), .ZN(n11185) );
  MUX2_X1 U13072 ( .A(n11634), .B(n11185), .S(n11184), .Z(n11186) );
  OAI22_X1 U13073 ( .A1(n14083), .A2(n12575), .B1(n16061), .B2(n10631), .ZN(
        n11187) );
  AOI21_X1 U13074 ( .B1(n12573), .B2(n16061), .A(n11187), .ZN(n11188) );
  INV_X1 U13075 ( .A(n11188), .ZN(P3_U3459) );
  OAI22_X1 U13076 ( .A1(n11673), .A2(n13335), .B1(n13354), .B2(n11619), .ZN(
        n11192) );
  NOR2_X1 U13077 ( .A1(n11190), .A2(n13079), .ZN(n11191) );
  AOI211_X1 U13078 ( .C1(n13318), .C2(n13586), .A(n11192), .B(n11191), .ZN(
        n11193) );
  OAI21_X1 U13079 ( .B1(n11194), .B2(n13314), .A(n11193), .ZN(P3_U3177) );
  INV_X1 U13080 ( .A(n11195), .ZN(n11196) );
  OAI222_X1 U13081 ( .A1(P3_U3151), .A2(n13743), .B1(n14158), .B2(n11196), 
        .C1(n13092), .C2(n14155), .ZN(P3_U3276) );
  OR2_X1 U13082 ( .A1(n15074), .A2(n12690), .ZN(n12685) );
  NAND2_X1 U13083 ( .A1(n11197), .A2(n12685), .ZN(n11198) );
  NAND2_X1 U13084 ( .A1(n11198), .A2(n11202), .ZN(n11350) );
  OAI21_X1 U13085 ( .B1(n11198), .B2(n11202), .A(n11350), .ZN(n15911) );
  INV_X1 U13086 ( .A(n15906), .ZN(n11355) );
  OAI211_X1 U13087 ( .C1(n11199), .C2(n11355), .A(n11352), .B(n15445), .ZN(
        n15909) );
  OAI21_X1 U13088 ( .B1(n11355), .B2(n16123), .A(n15909), .ZN(n11204) );
  INV_X1 U13089 ( .A(n15072), .ZN(n11431) );
  NAND2_X1 U13090 ( .A1(n11201), .A2(n11200), .ZN(n11358) );
  XNOR2_X1 U13091 ( .A(n11358), .B(n11202), .ZN(n11203) );
  OAI222_X1 U13092 ( .A1(n15357), .A2(n10994), .B1(n15359), .B2(n11431), .C1(
        n16136), .C2(n11203), .ZN(n15905) );
  AOI211_X1 U13093 ( .C1(n16139), .C2(n15911), .A(n11204), .B(n15905), .ZN(
        n11254) );
  NAND2_X1 U13094 ( .A1(n16141), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n11205) );
  OAI21_X1 U13095 ( .B1(n11254), .B2(n16141), .A(n11205), .ZN(P1_U3531) );
  INV_X1 U13096 ( .A(n13351), .ZN(n12397) );
  OAI211_X1 U13097 ( .C1(n11208), .C2(n11207), .A(n11206), .B(n13343), .ZN(
        n11212) );
  INV_X1 U13098 ( .A(n13318), .ZN(n13349) );
  OAI22_X1 U13099 ( .A1(n13349), .A2(n11905), .B1(n11904), .B2(n13335), .ZN(
        n11209) );
  AOI211_X1 U13100 ( .C1(n12565), .C2(n11624), .A(n11210), .B(n11209), .ZN(
        n11211) );
  OAI211_X1 U13101 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12397), .A(n11212), .B(
        n11211), .ZN(P3_U3158) );
  INV_X1 U13102 ( .A(P3_U3897), .ZN(n13587) );
  NAND2_X1 U13103 ( .A1(n13587), .A2(P3_DATAO_REG_25__SCAN_IN), .ZN(n11213) );
  OAI21_X1 U13104 ( .B1(n13827), .B2(n13587), .A(n11213), .ZN(P3_U3516) );
  INV_X1 U13105 ( .A(n11510), .ZN(n11807) );
  INV_X1 U13106 ( .A(n11216), .ZN(n11219) );
  INV_X1 U13107 ( .A(n11217), .ZN(n11218) );
  XNOR2_X1 U13108 ( .A(n11510), .B(n14188), .ZN(n11220) );
  NAND2_X1 U13109 ( .A1(n14370), .A2(n14633), .ZN(n11221) );
  NAND2_X1 U13110 ( .A1(n11220), .A2(n11221), .ZN(n11308) );
  INV_X1 U13111 ( .A(n11220), .ZN(n11223) );
  INV_X1 U13112 ( .A(n11221), .ZN(n11222) );
  NAND2_X1 U13113 ( .A1(n11223), .A2(n11222), .ZN(n11224) );
  AND2_X1 U13114 ( .A1(n11308), .A2(n11224), .ZN(n11225) );
  OAI21_X1 U13115 ( .B1(n11226), .B2(n11225), .A(n11309), .ZN(n11227) );
  NAND2_X1 U13116 ( .A1(n11227), .A2(n14311), .ZN(n11234) );
  INV_X1 U13117 ( .A(n11806), .ZN(n11232) );
  NAND2_X1 U13118 ( .A1(n14371), .A2(n14525), .ZN(n11229) );
  NAND2_X1 U13119 ( .A1(n14369), .A2(n14338), .ZN(n11228) );
  NAND2_X1 U13120 ( .A1(n11229), .A2(n11228), .ZN(n11407) );
  INV_X1 U13121 ( .A(n11407), .ZN(n11230) );
  NAND2_X1 U13122 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n14398) );
  OAI21_X1 U13123 ( .B1(n14341), .B2(n11230), .A(n14398), .ZN(n11231) );
  AOI21_X1 U13124 ( .B1(n11232), .B2(n14339), .A(n11231), .ZN(n11233) );
  OAI211_X1 U13125 ( .C1(n11807), .C2(n14309), .A(n11234), .B(n11233), .ZN(
        P2_U3185) );
  INV_X1 U13126 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11237) );
  MUX2_X1 U13127 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11237), .S(n11464), .Z(
        n11238) );
  OAI21_X1 U13128 ( .B1(n11239), .B2(n11238), .A(n11463), .ZN(n11252) );
  NOR2_X1 U13129 ( .A1(n11241), .A2(n11240), .ZN(n11245) );
  INV_X1 U13130 ( .A(n11245), .ZN(n11243) );
  INV_X1 U13131 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11989) );
  MUX2_X1 U13132 ( .A(n11989), .B(P1_REG2_REG_11__SCAN_IN), .S(n11464), .Z(
        n11242) );
  NAND2_X1 U13133 ( .A1(n11243), .A2(n11242), .ZN(n11246) );
  MUX2_X1 U13134 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11989), .S(n11464), .Z(
        n11244) );
  OAI21_X1 U13135 ( .B1(n11247), .B2(n11245), .A(n11244), .ZN(n11467) );
  OAI211_X1 U13136 ( .C1(n11247), .C2(n11246), .A(n11467), .B(n15143), .ZN(
        n11250) );
  NAND2_X1 U13137 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n12263)
         );
  INV_X1 U13138 ( .A(n12263), .ZN(n11248) );
  AOI21_X1 U13139 ( .B1(n15639), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n11248), 
        .ZN(n11249) );
  OAI211_X1 U13140 ( .C1(n15647), .C2(n11468), .A(n11250), .B(n11249), .ZN(
        n11251) );
  AOI21_X1 U13141 ( .B1(n11252), .B2(n15652), .A(n11251), .ZN(n11253) );
  INV_X1 U13142 ( .A(n11253), .ZN(P1_U3254) );
  INV_X1 U13143 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n11256) );
  OR2_X1 U13144 ( .A1(n11254), .A2(n16144), .ZN(n11255) );
  OAI21_X1 U13145 ( .B1(n16147), .B2(n11256), .A(n11255), .ZN(P1_U3468) );
  AND2_X1 U13146 ( .A1(n16054), .A2(n13563), .ZN(n11257) );
  NAND2_X1 U13147 ( .A1(n11258), .A2(n11257), .ZN(n11262) );
  OR2_X1 U13148 ( .A1(n11260), .A2(n11259), .ZN(n11261) );
  OR2_X1 U13149 ( .A1(n13550), .A2(n13565), .ZN(n16011) );
  INV_X1 U13150 ( .A(n14058), .ZN(n14080) );
  OAI21_X1 U13151 ( .B1(n11263), .B2(n11264), .A(n11627), .ZN(n11791) );
  INV_X1 U13152 ( .A(n11265), .ZN(n11266) );
  INV_X1 U13153 ( .A(n13588), .ZN(n11276) );
  NAND2_X1 U13154 ( .A1(n11268), .A2(n11267), .ZN(n13560) );
  NAND2_X1 U13155 ( .A1(n13588), .A2(n11270), .ZN(n11272) );
  INV_X1 U13156 ( .A(n11272), .ZN(n11274) );
  INV_X1 U13157 ( .A(n11677), .ZN(n11273) );
  AOI21_X1 U13158 ( .B1(n11274), .B2(n11263), .A(n11273), .ZN(n11275) );
  OAI222_X1 U13159 ( .A1(n13944), .A2(n11905), .B1(n13946), .B2(n11276), .C1(
        n14002), .C2(n11275), .ZN(n11789) );
  AOI21_X1 U13160 ( .B1(n14080), .B2(n11791), .A(n11789), .ZN(n11281) );
  INV_X1 U13161 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n11277) );
  OAI22_X1 U13162 ( .A1(n14142), .A2(n13380), .B1(n11277), .B2(n16065), .ZN(
        n11278) );
  INV_X1 U13163 ( .A(n11278), .ZN(n11279) );
  OAI21_X1 U13164 ( .B1(n11281), .B2(n16062), .A(n11279), .ZN(P3_U3393) );
  INV_X1 U13165 ( .A(n14083), .ZN(n14063) );
  INV_X1 U13166 ( .A(n13380), .ZN(n11626) );
  AOI22_X1 U13167 ( .A1(n14063), .A2(n11626), .B1(n12991), .B2(
        P3_REG1_REG_1__SCAN_IN), .ZN(n11280) );
  OAI21_X1 U13168 ( .B1(n11281), .B2(n12991), .A(n11280), .ZN(P3_U3460) );
  NAND2_X1 U13169 ( .A1(n11282), .A2(n11283), .ZN(n11284) );
  XOR2_X1 U13170 ( .A(n11285), .B(n11284), .Z(n11292) );
  AND2_X1 U13171 ( .A1(n12703), .A2(n16134), .ZN(n15920) );
  NAND2_X1 U13172 ( .A1(n15071), .A2(n15376), .ZN(n11287) );
  NAND2_X1 U13173 ( .A1(n15073), .A2(n16030), .ZN(n11286) );
  AND2_X1 U13174 ( .A1(n11287), .A2(n11286), .ZN(n15922) );
  NAND2_X1 U13175 ( .A1(n14987), .A2(n11354), .ZN(n11288) );
  OAI211_X1 U13176 ( .C1(n15922), .C2(n15026), .A(n11289), .B(n11288), .ZN(
        n11290) );
  AOI21_X1 U13177 ( .B1(n11300), .B2(n15920), .A(n11290), .ZN(n11291) );
  OAI21_X1 U13178 ( .B1(n11292), .B2(n15042), .A(n11291), .ZN(P1_U3230) );
  NAND2_X1 U13179 ( .A1(n11294), .A2(n11293), .ZN(n11296) );
  XOR2_X1 U13180 ( .A(n11296), .B(n11295), .Z(n11302) );
  AND2_X1 U13181 ( .A1(n12709), .A2(n16134), .ZN(n15931) );
  INV_X1 U13182 ( .A(n15070), .ZN(n11445) );
  AOI22_X1 U13183 ( .A1(n11571), .A2(n14987), .B1(n16087), .B2(n15072), .ZN(
        n11298) );
  OAI211_X1 U13184 ( .C1(n11445), .C2(n15036), .A(n11298), .B(n11297), .ZN(
        n11299) );
  AOI21_X1 U13185 ( .B1(n11300), .B2(n15931), .A(n11299), .ZN(n11301) );
  OAI21_X1 U13186 ( .B1(n11302), .B2(n15042), .A(n11301), .ZN(P1_U3227) );
  INV_X1 U13187 ( .A(n16003), .ZN(n11762) );
  XNOR2_X1 U13188 ( .A(n16003), .B(n14188), .ZN(n11303) );
  NAND2_X1 U13189 ( .A1(n14369), .A2(n14633), .ZN(n11304) );
  NAND2_X1 U13190 ( .A1(n11303), .A2(n11304), .ZN(n11364) );
  INV_X1 U13191 ( .A(n11303), .ZN(n11306) );
  INV_X1 U13192 ( .A(n11304), .ZN(n11305) );
  NAND2_X1 U13193 ( .A1(n11306), .A2(n11305), .ZN(n11307) );
  AND2_X1 U13194 ( .A1(n11364), .A2(n11307), .ZN(n11311) );
  OAI21_X1 U13195 ( .B1(n11311), .B2(n11310), .A(n11365), .ZN(n11312) );
  NAND2_X1 U13196 ( .A1(n11312), .A2(n14311), .ZN(n11318) );
  INV_X1 U13197 ( .A(n11761), .ZN(n11316) );
  NAND2_X1 U13198 ( .A1(n14368), .A2(n14338), .ZN(n11314) );
  NAND2_X1 U13199 ( .A1(n14370), .A2(n14525), .ZN(n11313) );
  AND2_X1 U13200 ( .A1(n11314), .A2(n11313), .ZN(n11753) );
  NAND2_X1 U13201 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14413) );
  OAI21_X1 U13202 ( .B1(n14341), .B2(n11753), .A(n14413), .ZN(n11315) );
  AOI21_X1 U13203 ( .B1(n11316), .B2(n14339), .A(n11315), .ZN(n11317) );
  OAI211_X1 U13204 ( .C1(n11762), .C2(n14309), .A(n11318), .B(n11317), .ZN(
        P2_U3193) );
  INV_X1 U13205 ( .A(n11319), .ZN(n12409) );
  INV_X1 U13206 ( .A(n11320), .ZN(n11322) );
  OAI222_X1 U13207 ( .A1(P2_U3088), .A2(n12409), .B1(n14869), .B2(n11322), 
        .C1(n11321), .C2(n14871), .ZN(P2_U3309) );
  INV_X1 U13208 ( .A(n15138), .ZN(n15125) );
  OAI222_X1 U13209 ( .A1(n15512), .A2(n11323), .B1(n15510), .B2(n11322), .C1(
        n15125), .C2(n7201), .ZN(P1_U3337) );
  INV_X1 U13210 ( .A(n11324), .ZN(n11429) );
  OAI222_X1 U13211 ( .A1(n15512), .A2(n11325), .B1(n7201), .B2(n12838), .C1(
        n15510), .C2(n11429), .ZN(P1_U3335) );
  INV_X1 U13212 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n12071) );
  INV_X1 U13213 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n12140) );
  MUX2_X1 U13214 ( .A(n12071), .B(n12140), .S(n10630), .Z(n11329) );
  NAND2_X1 U13215 ( .A1(n11329), .A2(n11342), .ZN(n11484) );
  INV_X1 U13216 ( .A(n11329), .ZN(n11330) );
  NAND2_X1 U13217 ( .A1(n11330), .A2(n11498), .ZN(n11331) );
  NAND2_X1 U13218 ( .A1(n11484), .A2(n11331), .ZN(n11332) );
  OR2_X1 U13219 ( .A1(n11333), .A2(n11332), .ZN(n11485) );
  NAND2_X1 U13220 ( .A1(n11333), .A2(n11332), .ZN(n11334) );
  AOI21_X1 U13221 ( .B1(n11485), .B2(n11334), .A(n15843), .ZN(n11348) );
  OAI21_X1 U13222 ( .B1(n11336), .B2(n15944), .A(n11335), .ZN(n11497) );
  XNOR2_X1 U13223 ( .A(n11497), .B(n11498), .ZN(n11337) );
  AOI21_X1 U13224 ( .B1(n12140), .B2(n11337), .A(n11496), .ZN(n11338) );
  NOR2_X1 U13225 ( .A1(n11338), .A2(n15866), .ZN(n11347) );
  XNOR2_X1 U13226 ( .A(n11488), .B(n11342), .ZN(n11341) );
  NOR2_X1 U13227 ( .A1(n11341), .A2(n12071), .ZN(n11489) );
  AOI21_X1 U13228 ( .B1(n12071), .B2(n11341), .A(n11489), .ZN(n11345) );
  AND2_X1 U13229 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11817) );
  AOI21_X1 U13230 ( .B1(n15521), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11817), .ZN(
        n11344) );
  NAND2_X1 U13231 ( .A1(n13754), .A2(n11342), .ZN(n11343) );
  OAI211_X1 U13232 ( .C1(n11345), .C2(n15872), .A(n11344), .B(n11343), .ZN(
        n11346) );
  OR3_X1 U13233 ( .A1(n11348), .A2(n11347), .A3(n11346), .ZN(P3_U3189) );
  INV_X1 U13234 ( .A(n15073), .ZN(n11356) );
  NAND2_X1 U13235 ( .A1(n11356), .A2(n11355), .ZN(n11349) );
  NAND2_X1 U13236 ( .A1(n11350), .A2(n11349), .ZN(n11351) );
  NAND2_X1 U13237 ( .A1(n11351), .A2(n12856), .ZN(n11433) );
  OAI21_X1 U13238 ( .B1(n11351), .B2(n12856), .A(n11433), .ZN(n15927) );
  AOI21_X1 U13239 ( .B1(n11352), .B2(n12703), .A(n15974), .ZN(n11353) );
  NAND2_X1 U13240 ( .A1(n11353), .A2(n11568), .ZN(n15923) );
  INV_X1 U13241 ( .A(n15368), .ZN(n15993) );
  OAI22_X1 U13242 ( .A1(n15923), .A2(n15993), .B1(n11440), .B2(n15365), .ZN(
        n11362) );
  NOR2_X1 U13243 ( .A1(n15073), .A2(n11355), .ZN(n11357) );
  XNOR2_X1 U13244 ( .A(n11439), .B(n12856), .ZN(n11359) );
  NAND2_X1 U13245 ( .A1(n11359), .A2(n16119), .ZN(n15924) );
  OAI211_X1 U13246 ( .C1(n15377), .C2(n9914), .A(n15924), .B(n15922), .ZN(
        n11360) );
  MUX2_X1 U13247 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11360), .S(n7218), .Z(
        n11361) );
  AOI211_X1 U13248 ( .C1(n15355), .C2(n15927), .A(n11362), .B(n11361), .ZN(
        n11363) );
  INV_X1 U13249 ( .A(n11363), .ZN(P1_U3289) );
  NAND2_X1 U13250 ( .A1(n14368), .A2(n14633), .ZN(n11589) );
  XNOR2_X1 U13251 ( .A(n11588), .B(n11589), .ZN(n11593) );
  XNOR2_X1 U13252 ( .A(n11594), .B(n11593), .ZN(n11374) );
  INV_X1 U13253 ( .A(n11366), .ZN(n11796) );
  NAND2_X1 U13254 ( .A1(n14367), .A2(n14338), .ZN(n11368) );
  NAND2_X1 U13255 ( .A1(n14369), .A2(n14525), .ZN(n11367) );
  NAND2_X1 U13256 ( .A1(n11368), .A2(n11367), .ZN(n11515) );
  INV_X1 U13257 ( .A(n11515), .ZN(n11370) );
  OAI22_X1 U13258 ( .A1(n14341), .A2(n11370), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11369), .ZN(n11371) );
  AOI21_X1 U13259 ( .B1(n11796), .B2(n14339), .A(n11371), .ZN(n11373) );
  NAND2_X1 U13260 ( .A1(n11795), .A2(n14358), .ZN(n11372) );
  OAI211_X1 U13261 ( .C1(n11374), .C2(n14353), .A(n11373), .B(n11372), .ZN(
        P2_U3203) );
  OAI222_X1 U13262 ( .A1(n14871), .A2(n11376), .B1(n14869), .B2(n11418), .C1(
        n11375), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI211_X1 U13263 ( .C1(n11379), .C2(n11378), .A(n11377), .B(n16093), .ZN(
        n11384) );
  INV_X1 U13264 ( .A(n15071), .ZN(n11610) );
  NOR2_X1 U13265 ( .A1(n11610), .A2(n15049), .ZN(n11382) );
  INV_X1 U13266 ( .A(n15069), .ZN(n11927) );
  OAI22_X1 U13267 ( .A1(n11927), .A2(n15036), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11380), .ZN(n11381) );
  AOI211_X1 U13268 ( .C1(n14987), .C2(n11607), .A(n11382), .B(n11381), .ZN(
        n11383) );
  OAI211_X1 U13269 ( .C1(n15948), .C2(n16091), .A(n11384), .B(n11383), .ZN(
        P1_U3239) );
  INV_X1 U13270 ( .A(n11385), .ZN(n11386) );
  AOI21_X1 U13271 ( .B1(n11388), .B2(n11387), .A(n11386), .ZN(n11393) );
  OAI22_X1 U13272 ( .A1(n13349), .A2(n11673), .B1(n11886), .B2(n13335), .ZN(
        n11389) );
  AOI211_X1 U13273 ( .C1(n12565), .C2(n11650), .A(n11390), .B(n11389), .ZN(
        n11392) );
  NAND2_X1 U13274 ( .A1(n13351), .A2(n11642), .ZN(n11391) );
  OAI211_X1 U13275 ( .C1(n11393), .C2(n13314), .A(n11392), .B(n11391), .ZN(
        P3_U3170) );
  NAND2_X1 U13276 ( .A1(n11395), .A2(n11394), .ZN(n11398) );
  NAND2_X1 U13277 ( .A1(n11400), .A2(n11396), .ZN(n11397) );
  INV_X1 U13278 ( .A(n11399), .ZN(n11403) );
  XNOR2_X1 U13279 ( .A(n11403), .B(n11512), .ZN(n11408) );
  OR2_X1 U13280 ( .A1(n11400), .A2(n14371), .ZN(n11401) );
  NAND2_X1 U13281 ( .A1(n11404), .A2(n11403), .ZN(n11405) );
  NAND2_X1 U13282 ( .A1(n11508), .A2(n11405), .ZN(n11812) );
  NOR2_X1 U13283 ( .A1(n11812), .A2(n14807), .ZN(n11406) );
  AOI211_X1 U13284 ( .C1(n14710), .C2(n11408), .A(n11407), .B(n11406), .ZN(
        n11804) );
  INV_X1 U13285 ( .A(n11409), .ZN(n11410) );
  AOI211_X1 U13286 ( .C1(n11510), .C2(n11410), .A(n14633), .B(n11757), .ZN(
        n11809) );
  INV_X1 U13287 ( .A(n11809), .ZN(n11411) );
  OAI211_X1 U13288 ( .C1(n11807), .C2(n16149), .A(n11804), .B(n11411), .ZN(
        n11416) );
  OAI22_X1 U13289 ( .A1(n11812), .A2(n14816), .B1(n16156), .B2(n11412), .ZN(
        n11413) );
  AOI21_X1 U13290 ( .B1(n11416), .B2(n16156), .A(n11413), .ZN(n11414) );
  INV_X1 U13291 ( .A(n11414), .ZN(P2_U3506) );
  OAI22_X1 U13292 ( .A1(n11812), .A2(n14849), .B1(n16160), .B2(n9045), .ZN(
        n11415) );
  AOI21_X1 U13293 ( .B1(n11416), .B2(n16117), .A(n11415), .ZN(n11417) );
  INV_X1 U13294 ( .A(n11417), .ZN(P2_U3451) );
  OAI222_X1 U13295 ( .A1(n11951), .A2(n11420), .B1(P1_U3086), .B2(n11419), 
        .C1(n15510), .C2(n11418), .ZN(P1_U3334) );
  INV_X1 U13296 ( .A(n11421), .ZN(n11423) );
  OAI222_X1 U13297 ( .A1(n14871), .A2(n11422), .B1(n14869), .B2(n11423), .C1(
        P2_U3088), .C2(n12414), .ZN(P2_U3308) );
  OAI222_X1 U13298 ( .A1(n15512), .A2(n11424), .B1(n15510), .B2(n11423), .C1(
        n7228), .C2(P1_U3086), .ZN(P1_U3336) );
  INV_X1 U13299 ( .A(n11425), .ZN(n11427) );
  OAI222_X1 U13300 ( .A1(n14158), .A2(n11427), .B1(n14155), .B2(n13114), .C1(
        P3_U3151), .C2(n11426), .ZN(P3_U3275) );
  OAI222_X1 U13301 ( .A1(P2_U3088), .A2(n11430), .B1(n14869), .B2(n11429), 
        .C1(n11428), .C2(n14871), .ZN(P2_U3307) );
  NAND2_X1 U13302 ( .A1(n11431), .A2(n11440), .ZN(n11432) );
  NAND2_X1 U13303 ( .A1(n11433), .A2(n11432), .ZN(n11565) );
  XNOR2_X1 U13304 ( .A(n15071), .B(n12709), .ZN(n12860) );
  INV_X1 U13305 ( .A(n12860), .ZN(n11564) );
  NAND2_X1 U13306 ( .A1(n11565), .A2(n11564), .ZN(n11567) );
  INV_X1 U13307 ( .A(n12709), .ZN(n12710) );
  NAND2_X1 U13308 ( .A1(n11610), .A2(n12710), .ZN(n11434) );
  NAND2_X1 U13309 ( .A1(n11567), .A2(n11434), .ZN(n11603) );
  NAND2_X1 U13310 ( .A1(n12716), .A2(n15070), .ZN(n11435) );
  NAND2_X1 U13311 ( .A1(n11603), .A2(n11435), .ZN(n11437) );
  OR2_X1 U13312 ( .A1(n12716), .A2(n15070), .ZN(n11436) );
  NAND2_X1 U13313 ( .A1(n11437), .A2(n11436), .ZN(n11915) );
  XNOR2_X1 U13314 ( .A(n12725), .B(n15069), .ZN(n12859) );
  XNOR2_X1 U13315 ( .A(n11915), .B(n12859), .ZN(n15958) );
  INV_X1 U13316 ( .A(n12856), .ZN(n11438) );
  NAND2_X1 U13317 ( .A1(n11439), .A2(n11438), .ZN(n11442) );
  NAND2_X1 U13318 ( .A1(n15072), .A2(n11440), .ZN(n11441) );
  NAND2_X1 U13319 ( .A1(n11442), .A2(n11441), .ZN(n11573) );
  NAND2_X1 U13320 ( .A1(n11573), .A2(n12860), .ZN(n11444) );
  NAND2_X1 U13321 ( .A1(n12710), .A2(n15071), .ZN(n11443) );
  NAND2_X1 U13322 ( .A1(n11444), .A2(n11443), .ZN(n11609) );
  XNOR2_X1 U13323 ( .A(n12716), .B(n15070), .ZN(n12858) );
  OR2_X1 U13324 ( .A1(n11445), .A2(n12716), .ZN(n11446) );
  INV_X1 U13325 ( .A(n12859), .ZN(n11914) );
  XNOR2_X1 U13326 ( .A(n11926), .B(n11914), .ZN(n11448) );
  AOI22_X1 U13327 ( .A1(n15376), .A2(n15068), .B1(n15070), .B2(n16030), .ZN(
        n11457) );
  INV_X1 U13328 ( .A(n11457), .ZN(n11447) );
  AOI21_X1 U13329 ( .B1(n11448), .B2(n16119), .A(n11447), .ZN(n15956) );
  MUX2_X1 U13330 ( .A(n10407), .B(n15956), .S(n7218), .Z(n11453) );
  AND2_X1 U13331 ( .A1(n11604), .A2(n15948), .ZN(n11605) );
  NAND2_X1 U13332 ( .A1(n11605), .A2(n15957), .ZN(n15975) );
  OAI211_X1 U13333 ( .C1(n11605), .C2(n15957), .A(n15445), .B(n15975), .ZN(
        n15955) );
  INV_X1 U13334 ( .A(n15955), .ZN(n11451) );
  INV_X1 U13335 ( .A(n11460), .ZN(n11449) );
  OAI22_X1 U13336 ( .A1(n15957), .A2(n15365), .B1(n15377), .B2(n11449), .ZN(
        n11450) );
  AOI21_X1 U13337 ( .B1(n11451), .B2(n15368), .A(n11450), .ZN(n11452) );
  OAI211_X1 U13338 ( .C1(n15392), .C2(n15958), .A(n11453), .B(n11452), .ZN(
        P1_U3286) );
  OAI211_X1 U13339 ( .C1(n11456), .C2(n11455), .A(n11454), .B(n16093), .ZN(
        n11462) );
  NOR2_X1 U13340 ( .A1(n11457), .A2(n15026), .ZN(n11458) );
  AOI211_X1 U13341 ( .C1(n14987), .C2(n11460), .A(n11459), .B(n11458), .ZN(
        n11461) );
  OAI211_X1 U13342 ( .C1(n15957), .C2(n16091), .A(n11462), .B(n11461), .ZN(
        P1_U3213) );
  INV_X1 U13343 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n16073) );
  XOR2_X1 U13344 ( .A(n16073), .B(n11836), .Z(n11476) );
  INV_X1 U13345 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n11465) );
  NAND2_X1 U13346 ( .A1(n7201), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n12550) );
  OAI21_X1 U13347 ( .B1(n15656), .B2(n11465), .A(n12550), .ZN(n11473) );
  INV_X1 U13348 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11466) );
  MUX2_X1 U13349 ( .A(n11466), .B(P1_REG2_REG_12__SCAN_IN), .S(n11474), .Z(
        n11470) );
  OAI21_X1 U13350 ( .B1(n11989), .B2(n11468), .A(n11467), .ZN(n11469) );
  NOR2_X1 U13351 ( .A1(n11469), .A2(n11470), .ZN(n11829) );
  AOI21_X1 U13352 ( .B1(n11470), .B2(n11469), .A(n11829), .ZN(n11471) );
  NOR2_X1 U13353 ( .A1(n11471), .A2(n15649), .ZN(n11472) );
  AOI211_X1 U13354 ( .C1(n15147), .C2(n11474), .A(n11473), .B(n11472), .ZN(
        n11475) );
  OAI21_X1 U13355 ( .B1(n11476), .B2(n15145), .A(n11475), .ZN(P1_U3255) );
  XOR2_X1 U13356 ( .A(n11478), .B(n11477), .Z(n11483) );
  OAI22_X1 U13357 ( .A1(n13349), .A2(n11904), .B1(n13412), .B2(n13335), .ZN(
        n11479) );
  AOI211_X1 U13358 ( .C1(n12565), .C2(n11955), .A(n11480), .B(n11479), .ZN(
        n11482) );
  NAND2_X1 U13359 ( .A1(n13351), .A2(n11658), .ZN(n11481) );
  OAI211_X1 U13360 ( .C1(n11483), .C2(n13314), .A(n11482), .B(n11481), .ZN(
        P3_U3167) );
  NAND2_X1 U13361 ( .A1(n11485), .A2(n11484), .ZN(n11487) );
  MUX2_X1 U13362 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n10630), .Z(n11524) );
  INV_X1 U13363 ( .A(n11499), .ZN(n11525) );
  XNOR2_X1 U13364 ( .A(n11524), .B(n11525), .ZN(n11486) );
  NAND2_X1 U13365 ( .A1(n11487), .A2(n11486), .ZN(n11530) );
  OAI21_X1 U13366 ( .B1(n11487), .B2(n11486), .A(n11530), .ZN(n11505) );
  INV_X1 U13367 ( .A(n11488), .ZN(n11490) );
  NAND2_X1 U13368 ( .A1(n11499), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11533) );
  OAI21_X1 U13369 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11499), .A(n11533), .ZN(
        n11491) );
  NOR2_X1 U13370 ( .A1(n11492), .A2(n11491), .ZN(n11531) );
  AOI21_X1 U13371 ( .B1(n11492), .B2(n11491), .A(n11531), .ZN(n11495) );
  AND2_X1 U13372 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n12004) );
  AOI21_X1 U13373 ( .B1(n15521), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12004), .ZN(
        n11494) );
  NAND2_X1 U13374 ( .A1(n13754), .A2(n11525), .ZN(n11493) );
  OAI211_X1 U13375 ( .C1(n11495), .C2(n15872), .A(n11494), .B(n11493), .ZN(
        n11504) );
  NAND2_X1 U13376 ( .A1(n11499), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11538) );
  OAI21_X1 U13377 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n11499), .A(n11538), .ZN(
        n11500) );
  AOI21_X1 U13378 ( .B1(n11501), .B2(n11500), .A(n11536), .ZN(n11502) );
  NOR2_X1 U13379 ( .A1(n11502), .A2(n15866), .ZN(n11503) );
  AOI211_X1 U13380 ( .C1(n15863), .C2(n11505), .A(n11504), .B(n11503), .ZN(
        n11506) );
  INV_X1 U13381 ( .A(n11506), .ZN(P3_U3190) );
  AOI211_X1 U13382 ( .C1(n11795), .C2(n11758), .A(n14633), .B(n7709), .ZN(
        n11800) );
  NAND2_X1 U13383 ( .A1(n11510), .A2(n14370), .ZN(n11507) );
  NAND2_X1 U13384 ( .A1(n16003), .A2(n14369), .ZN(n11509) );
  XNOR2_X1 U13385 ( .A(n11702), .B(n11713), .ZN(n11803) );
  XNOR2_X1 U13386 ( .A(n11715), .B(n11713), .ZN(n11516) );
  AOI21_X1 U13387 ( .B1(n11516), .B2(n14710), .A(n11515), .ZN(n11517) );
  OAI21_X1 U13388 ( .B1(n11803), .B2(n14807), .A(n11517), .ZN(n11794) );
  AOI211_X1 U13389 ( .C1(n16112), .C2(n11795), .A(n11800), .B(n11794), .ZN(
        n11523) );
  INV_X1 U13390 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11518) );
  OAI22_X1 U13391 ( .A1(n11803), .A2(n14849), .B1(n16160), .B2(n11518), .ZN(
        n11519) );
  INV_X1 U13392 ( .A(n11519), .ZN(n11520) );
  OAI21_X1 U13393 ( .B1(n11523), .B2(n16157), .A(n11520), .ZN(P2_U3457) );
  INV_X1 U13394 ( .A(n11803), .ZN(n11521) );
  AOI22_X1 U13395 ( .A1(n11521), .A2(n12464), .B1(n16155), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11522) );
  OAI21_X1 U13396 ( .B1(n11523), .B2(n16155), .A(n11522), .ZN(P2_U3508) );
  MUX2_X1 U13397 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n10630), .Z(n12027) );
  XNOR2_X1 U13398 ( .A(n12027), .B(n7794), .ZN(n11528) );
  INV_X1 U13399 ( .A(n11524), .ZN(n11526) );
  NAND2_X1 U13400 ( .A1(n11526), .A2(n11525), .ZN(n11529) );
  AND2_X1 U13401 ( .A1(n11528), .A2(n11529), .ZN(n11527) );
  NAND2_X1 U13402 ( .A1(n11530), .A2(n11527), .ZN(n12029) );
  NAND2_X1 U13403 ( .A1(n12029), .A2(n15863), .ZN(n11549) );
  AOI21_X1 U13404 ( .B1(n11530), .B2(n11529), .A(n11528), .ZN(n11548) );
  INV_X1 U13405 ( .A(n11531), .ZN(n11532) );
  NAND2_X1 U13406 ( .A1(n11533), .A2(n11532), .ZN(n11534) );
  INV_X1 U13407 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12174) );
  AOI21_X1 U13408 ( .B1(n11535), .B2(n12174), .A(n12045), .ZN(n11545) );
  NOR2_X1 U13409 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8469), .ZN(n12236) );
  NAND2_X1 U13410 ( .A1(n11538), .A2(n11537), .ZN(n11540) );
  INV_X1 U13411 ( .A(n12057), .ZN(n11539) );
  OAI21_X1 U13412 ( .B1(n11540), .B2(n12026), .A(n11539), .ZN(n11541) );
  INV_X1 U13413 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n16015) );
  AOI21_X1 U13414 ( .B1(n11541), .B2(n16015), .A(n12056), .ZN(n11542) );
  NOR2_X1 U13415 ( .A1(n15866), .A2(n11542), .ZN(n11543) );
  AOI211_X1 U13416 ( .C1(n15521), .C2(P3_ADDR_REG_9__SCAN_IN), .A(n12236), .B(
        n11543), .ZN(n11544) );
  OAI21_X1 U13417 ( .B1(n11545), .B2(n15872), .A(n11544), .ZN(n11546) );
  AOI21_X1 U13418 ( .B1(n7794), .B2(n13754), .A(n11546), .ZN(n11547) );
  OAI21_X1 U13419 ( .B1(n11549), .B2(n11548), .A(n11547), .ZN(P3_U3191) );
  INV_X1 U13420 ( .A(n11550), .ZN(n11551) );
  OAI222_X1 U13421 ( .A1(n14158), .A2(n11551), .B1(n14155), .B2(n13112), .C1(
        P3_U3151), .C2(n13388), .ZN(P3_U3274) );
  NAND2_X1 U13422 ( .A1(n11558), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11553) );
  NAND2_X1 U13423 ( .A1(n11553), .A2(n11552), .ZN(n12321) );
  XOR2_X1 U13424 ( .A(n12321), .B(n12322), .Z(n11554) );
  NAND2_X1 U13425 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n11554), .ZN(n12323) );
  OAI211_X1 U13426 ( .C1(n11554), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15611), 
        .B(n12323), .ZN(n11563) );
  AND2_X1 U13427 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n11555) );
  AOI21_X1 U13428 ( .B1(n15627), .B2(n12322), .A(n11555), .ZN(n11556) );
  INV_X1 U13429 ( .A(n11556), .ZN(n11561) );
  AOI21_X1 U13430 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n11558), .A(n11557), 
        .ZN(n12329) );
  XNOR2_X1 U13431 ( .A(n12328), .B(n12329), .ZN(n11559) );
  NOR2_X1 U13432 ( .A1(n9260), .A2(n11559), .ZN(n12330) );
  AOI211_X1 U13433 ( .C1(n9260), .C2(n11559), .A(n12330), .B(n15622), .ZN(
        n11560) );
  AOI211_X1 U13434 ( .C1(n15619), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n11561), 
        .B(n11560), .ZN(n11562) );
  NAND2_X1 U13435 ( .A1(n11563), .A2(n11562), .ZN(P2_U3229) );
  INV_X1 U13436 ( .A(n12932), .ZN(n15996) );
  OR2_X1 U13437 ( .A1(n11565), .A2(n11564), .ZN(n11566) );
  NAND2_X1 U13438 ( .A1(n11567), .A2(n11566), .ZN(n15936) );
  INV_X1 U13439 ( .A(n11568), .ZN(n11570) );
  INV_X1 U13440 ( .A(n11604), .ZN(n11569) );
  OAI211_X1 U13441 ( .C1(n12710), .C2(n11570), .A(n11569), .B(n15445), .ZN(
        n15933) );
  AOI22_X1 U13442 ( .A1(n15991), .A2(n12709), .B1(n15990), .B2(n11571), .ZN(
        n11572) );
  OAI21_X1 U13443 ( .B1(n15933), .B2(n15993), .A(n11572), .ZN(n11578) );
  XNOR2_X1 U13444 ( .A(n11573), .B(n12860), .ZN(n11576) );
  NAND2_X1 U13445 ( .A1(n15936), .A2(n16026), .ZN(n11575) );
  AOI22_X1 U13446 ( .A1(n15376), .A2(n15070), .B1(n15072), .B2(n16030), .ZN(
        n11574) );
  OAI211_X1 U13447 ( .C1(n16136), .C2(n11576), .A(n11575), .B(n11574), .ZN(
        n15934) );
  MUX2_X1 U13448 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n15934), .S(n7218), .Z(
        n11577) );
  AOI211_X1 U13449 ( .C1(n15996), .C2(n15936), .A(n11578), .B(n11577), .ZN(
        n11579) );
  INV_X1 U13450 ( .A(n11579), .ZN(P1_U3288) );
  INV_X1 U13451 ( .A(n11580), .ZN(n11582) );
  OAI22_X1 U13452 ( .A1(n13565), .A2(P3_U3151), .B1(SI_22_), .B2(n14155), .ZN(
        n11581) );
  AOI21_X1 U13453 ( .B1(n11582), .B2(n14148), .A(n11581), .ZN(P3_U3273) );
  XNOR2_X1 U13454 ( .A(n12157), .B(n14188), .ZN(n11583) );
  NAND2_X1 U13455 ( .A1(n14367), .A2(n14633), .ZN(n11584) );
  NAND2_X1 U13456 ( .A1(n11583), .A2(n11584), .ZN(n11691) );
  INV_X1 U13457 ( .A(n11583), .ZN(n11586) );
  INV_X1 U13458 ( .A(n11584), .ZN(n11585) );
  NAND2_X1 U13459 ( .A1(n11586), .A2(n11585), .ZN(n11587) );
  AND2_X1 U13460 ( .A1(n11691), .A2(n11587), .ZN(n11596) );
  INV_X1 U13461 ( .A(n11588), .ZN(n11591) );
  INV_X1 U13462 ( .A(n11589), .ZN(n11590) );
  NAND2_X1 U13463 ( .A1(n11591), .A2(n11590), .ZN(n11592) );
  OAI21_X1 U13464 ( .B1(n11596), .B2(n11595), .A(n11692), .ZN(n11597) );
  NAND2_X1 U13465 ( .A1(n11597), .A2(n14311), .ZN(n11602) );
  NAND2_X1 U13466 ( .A1(n14366), .A2(n14338), .ZN(n11599) );
  NAND2_X1 U13467 ( .A1(n14368), .A2(n14525), .ZN(n11598) );
  NAND2_X1 U13468 ( .A1(n11599), .A2(n11598), .ZN(n12146) );
  AND2_X1 U13469 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n14422) );
  NOR2_X1 U13470 ( .A1(n14351), .A2(n12154), .ZN(n11600) );
  AOI211_X1 U13471 ( .C1(n14348), .C2(n12146), .A(n14422), .B(n11600), .ZN(
        n11601) );
  OAI211_X1 U13472 ( .C1(n7708), .C2(n14309), .A(n11602), .B(n11601), .ZN(
        P2_U3189) );
  XNOR2_X1 U13473 ( .A(n11603), .B(n12858), .ZN(n11614) );
  INV_X1 U13474 ( .A(n11614), .ZN(n15951) );
  OAI21_X1 U13475 ( .B1(n11604), .B2(n15948), .A(n15445), .ZN(n11606) );
  OR2_X1 U13476 ( .A1(n11606), .A2(n11605), .ZN(n15947) );
  AOI22_X1 U13477 ( .A1(n15991), .A2(n12716), .B1(n11607), .B2(n15990), .ZN(
        n11608) );
  OAI21_X1 U13478 ( .B1(n15947), .B2(n15993), .A(n11608), .ZN(n11616) );
  XOR2_X1 U13479 ( .A(n11609), .B(n12858), .Z(n11612) );
  OAI22_X1 U13480 ( .A1(n11927), .A2(n15359), .B1(n11610), .B2(n15357), .ZN(
        n11611) );
  AOI21_X1 U13481 ( .B1(n11612), .B2(n16119), .A(n11611), .ZN(n11613) );
  OAI21_X1 U13482 ( .B1(n11614), .B2(n12928), .A(n11613), .ZN(n15949) );
  MUX2_X1 U13483 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n15949), .S(n7218), .Z(
        n11615) );
  AOI211_X1 U13484 ( .C1(n15951), .C2(n15996), .A(n11616), .B(n11615), .ZN(
        n11617) );
  INV_X1 U13485 ( .A(n11617), .ZN(P1_U3287) );
  NAND2_X1 U13486 ( .A1(n11904), .A2(n11650), .ZN(n13400) );
  INV_X1 U13487 ( .A(n11650), .ZN(n15914) );
  NAND2_X1 U13488 ( .A1(n13583), .A2(n15914), .ZN(n13401) );
  NAND2_X1 U13489 ( .A1(n11674), .A2(n13380), .ZN(n11676) );
  NAND2_X1 U13490 ( .A1(n11677), .A2(n11676), .ZN(n11618) );
  NAND2_X1 U13491 ( .A1(n11620), .A2(n11682), .ZN(n13392) );
  INV_X1 U13492 ( .A(n11620), .ZN(n13585) );
  NAND2_X1 U13493 ( .A1(n13585), .A2(n11619), .ZN(n13384) );
  NAND2_X1 U13494 ( .A1(n11618), .A2(n13386), .ZN(n11675) );
  INV_X1 U13495 ( .A(n11624), .ZN(n15899) );
  AND2_X1 U13496 ( .A1(n15899), .A2(n11902), .ZN(n11621) );
  NAND2_X1 U13497 ( .A1(n13584), .A2(n11621), .ZN(n11622) );
  NAND2_X1 U13498 ( .A1(n11675), .A2(n11623), .ZN(n11901) );
  NAND2_X1 U13499 ( .A1(n13584), .A2(n11624), .ZN(n11625) );
  XNOR2_X1 U13500 ( .A(n11649), .B(n11648), .ZN(n11631) );
  NAND2_X1 U13501 ( .A1(n11674), .A2(n11626), .ZN(n13383) );
  NAND2_X1 U13502 ( .A1(n13391), .A2(n13523), .ZN(n11672) );
  NAND2_X1 U13503 ( .A1(n11672), .A2(n13392), .ZN(n11898) );
  NAND2_X1 U13504 ( .A1(n13584), .A2(n15899), .ZN(n13395) );
  NAND2_X1 U13505 ( .A1(n11898), .A2(n8243), .ZN(n11900) );
  OAI21_X1 U13506 ( .B1(n11628), .B2(n13528), .A(n11653), .ZN(n15917) );
  NAND2_X1 U13507 ( .A1(n15917), .A2(n13994), .ZN(n11630) );
  AOI22_X1 U13508 ( .A1(n13584), .A2(n13997), .B1(n13996), .B2(n13582), .ZN(
        n11629) );
  OAI211_X1 U13509 ( .C1(n14002), .C2(n11631), .A(n11630), .B(n11629), .ZN(
        n15915) );
  INV_X1 U13510 ( .A(n15915), .ZN(n11647) );
  NAND2_X1 U13511 ( .A1(n11635), .A2(n11632), .ZN(n11633) );
  OAI21_X1 U13512 ( .B1(n11635), .B2(n11634), .A(n11633), .ZN(n11636) );
  INV_X1 U13513 ( .A(n11636), .ZN(n11637) );
  NOR2_X1 U13514 ( .A1(n13388), .A2(n13550), .ZN(n11640) );
  OR2_X1 U13515 ( .A1(n16054), .A2(n11683), .ZN(n11786) );
  INV_X1 U13516 ( .A(n14006), .ZN(n13986) );
  AOI22_X1 U13517 ( .A1(n13986), .A2(n11650), .B1(n14004), .B2(n11642), .ZN(
        n11643) );
  OAI21_X1 U13518 ( .B1(n11644), .B2(n13966), .A(n11643), .ZN(n11645) );
  AOI21_X1 U13519 ( .B1(n15917), .B2(n14008), .A(n11645), .ZN(n11646) );
  OAI21_X1 U13520 ( .B1(n11647), .B2(n13963), .A(n11646), .ZN(P3_U3229) );
  NAND2_X1 U13521 ( .A1(n13583), .A2(n11650), .ZN(n11651) );
  INV_X1 U13522 ( .A(n11890), .ZN(n11887) );
  AOI21_X1 U13523 ( .B1(n13533), .B2(n11652), .A(n11887), .ZN(n11657) );
  AOI22_X1 U13524 ( .A1(n13996), .A2(n13581), .B1(n13583), .B2(n13997), .ZN(
        n11656) );
  NAND2_X1 U13525 ( .A1(n11653), .A2(n13400), .ZN(n11654) );
  NAND2_X1 U13526 ( .A1(n11654), .A2(n13533), .ZN(n11885) );
  OAI21_X1 U13527 ( .B1(n11654), .B2(n13533), .A(n11885), .ZN(n11689) );
  NAND2_X1 U13528 ( .A1(n11689), .A2(n13994), .ZN(n11655) );
  OAI211_X1 U13529 ( .C1(n11657), .C2(n14002), .A(n11656), .B(n11655), .ZN(
        n11688) );
  INV_X1 U13530 ( .A(n11688), .ZN(n11663) );
  AOI22_X1 U13531 ( .A1(n13986), .A2(n11955), .B1(n14004), .B2(n11658), .ZN(
        n11659) );
  OAI21_X1 U13532 ( .B1(n11660), .B2(n13966), .A(n11659), .ZN(n11661) );
  AOI21_X1 U13533 ( .B1(n11689), .B2(n14008), .A(n11661), .ZN(n11662) );
  OAI21_X1 U13534 ( .B1(n11663), .B2(n13963), .A(n11662), .ZN(P3_U3228) );
  INV_X1 U13535 ( .A(n11664), .ZN(n11665) );
  AOI21_X1 U13536 ( .B1(n11667), .B2(n11666), .A(n11665), .ZN(n11671) );
  AOI22_X1 U13537 ( .A1(n15376), .A2(n16029), .B1(n15069), .B2(n16030), .ZN(
        n15979) );
  AOI22_X1 U13538 ( .A1(n14987), .A2(n7252), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        n7201), .ZN(n11668) );
  OAI21_X1 U13539 ( .B1(n15979), .B2(n15026), .A(n11668), .ZN(n11669) );
  AOI21_X1 U13540 ( .B1(n15040), .B2(n15992), .A(n11669), .ZN(n11670) );
  OAI21_X1 U13541 ( .B1(n11671), .B2(n15042), .A(n11670), .ZN(P1_U3221) );
  OAI21_X1 U13542 ( .B1(n13391), .B2(n13523), .A(n11672), .ZN(n15895) );
  OAI22_X1 U13543 ( .A1(n11674), .A2(n13946), .B1(n11673), .B2(n13944), .ZN(
        n11680) );
  NAND3_X1 U13544 ( .A1(n13523), .A2(n11677), .A3(n11676), .ZN(n11678) );
  AOI21_X1 U13545 ( .B1(n11675), .B2(n11678), .A(n14002), .ZN(n11679) );
  AOI211_X1 U13546 ( .C1(n13994), .C2(n15895), .A(n11680), .B(n11679), .ZN(
        n11681) );
  INV_X1 U13547 ( .A(n11681), .ZN(n15893) );
  NAND2_X1 U13548 ( .A1(n11682), .A2(n15940), .ZN(n15892) );
  OAI22_X1 U13549 ( .A1(n15892), .A2(n11683), .B1(n13983), .B2(n13079), .ZN(
        n11684) );
  OAI21_X1 U13550 ( .B1(n15893), .B2(n11684), .A(n13966), .ZN(n11686) );
  NAND2_X1 U13551 ( .A1(n15895), .A2(n14008), .ZN(n11685) );
  OAI211_X1 U13552 ( .C1(n11687), .C2(n13966), .A(n11686), .B(n11685), .ZN(
        P3_U3231) );
  AOI21_X1 U13553 ( .B1(n16059), .B2(n11689), .A(n11688), .ZN(n11956) );
  AOI22_X1 U13554 ( .A1(n14124), .A2(n11955), .B1(P3_REG0_REG_5__SCAN_IN), 
        .B2(n16062), .ZN(n11690) );
  OAI21_X1 U13555 ( .B1(n11956), .B2(n16062), .A(n11690), .ZN(P3_U3405) );
  INV_X1 U13556 ( .A(n14366), .ZN(n12282) );
  NOR2_X1 U13557 ( .A1(n12282), .A2(n14716), .ZN(n12181) );
  XNOR2_X1 U13558 ( .A(n12091), .B(n14188), .ZN(n12283) );
  XOR2_X1 U13559 ( .A(n12181), .B(n12283), .Z(n11693) );
  XNOR2_X1 U13560 ( .A(n12284), .B(n11693), .ZN(n11701) );
  INV_X1 U13561 ( .A(n11694), .ZN(n12090) );
  NAND2_X1 U13562 ( .A1(n14365), .A2(n14338), .ZN(n11696) );
  NAND2_X1 U13563 ( .A1(n14367), .A2(n14525), .ZN(n11695) );
  AND2_X1 U13564 ( .A1(n11696), .A2(n11695), .ZN(n11723) );
  OAI22_X1 U13565 ( .A1(n14341), .A2(n11723), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11697), .ZN(n11698) );
  AOI21_X1 U13566 ( .B1(n12090), .B2(n14339), .A(n11698), .ZN(n11700) );
  NAND2_X1 U13567 ( .A1(n12091), .A2(n14358), .ZN(n11699) );
  OAI211_X1 U13568 ( .C1(n11701), .C2(n14353), .A(n11700), .B(n11699), .ZN(
        P2_U3208) );
  NAND2_X1 U13569 ( .A1(n11702), .A2(n11713), .ZN(n11704) );
  NAND2_X1 U13570 ( .A1(n11795), .A2(n14368), .ZN(n11703) );
  NAND2_X1 U13571 ( .A1(n12143), .A2(n12157), .ZN(n11705) );
  NAND2_X1 U13572 ( .A1(n11708), .A2(n11858), .ZN(n11709) );
  INV_X1 U13573 ( .A(n12091), .ZN(n11712) );
  NAND2_X1 U13574 ( .A1(n12152), .A2(n12091), .ZN(n11710) );
  NAND2_X1 U13575 ( .A1(n11710), .A2(n14716), .ZN(n11711) );
  OR2_X1 U13576 ( .A1(n11711), .A2(n11867), .ZN(n12094) );
  OAI21_X1 U13577 ( .B1(n11712), .B2(n16149), .A(n12094), .ZN(n11725) );
  OR2_X1 U13578 ( .A1(n11795), .A2(n11716), .ZN(n11717) );
  NAND2_X1 U13579 ( .A1(n11718), .A2(n11717), .ZN(n12145) );
  NOR2_X1 U13580 ( .A1(n12157), .A2(n11720), .ZN(n11719) );
  NAND2_X1 U13581 ( .A1(n12157), .A2(n11720), .ZN(n11721) );
  XOR2_X1 U13582 ( .A(n11858), .B(n11859), .Z(n11724) );
  OAI21_X1 U13583 ( .B1(n11724), .B2(n14679), .A(n11723), .ZN(n12089) );
  AOI211_X1 U13584 ( .C1(n14803), .C2(n12096), .A(n11725), .B(n12089), .ZN(
        n11729) );
  AOI22_X1 U13585 ( .A1(n12096), .A2(n12464), .B1(n16155), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11726) );
  OAI21_X1 U13586 ( .B1(n11729), .B2(n16155), .A(n11726), .ZN(P2_U3510) );
  INV_X1 U13587 ( .A(n14849), .ZN(n12462) );
  NOR2_X1 U13588 ( .A1(n16117), .A2(n9150), .ZN(n11727) );
  AOI21_X1 U13589 ( .B1(n12096), .B2(n12462), .A(n11727), .ZN(n11728) );
  OAI21_X1 U13590 ( .B1(n11729), .B2(n16157), .A(n11728), .ZN(P2_U3463) );
  INV_X1 U13591 ( .A(n11730), .ZN(n11731) );
  AND3_X1 U13592 ( .A1(n11731), .A2(n15525), .A3(n15524), .ZN(n11732) );
  NAND2_X1 U13593 ( .A1(n11733), .A2(n11732), .ZN(n11741) );
  INV_X2 U13594 ( .A(n14697), .ZN(n12155) );
  NAND2_X1 U13595 ( .A1(n11734), .A2(n12410), .ZN(n11735) );
  OR2_X1 U13596 ( .A1(n15891), .A2(n14807), .ZN(n11736) );
  INV_X1 U13597 ( .A(n11738), .ZN(n11745) );
  NOR2_X1 U13598 ( .A1(n14718), .A2(n11739), .ZN(n11740) );
  AOI21_X1 U13599 ( .B1(n14697), .B2(P2_REG2_REG_4__SCAN_IN), .A(n11740), .ZN(
        n11744) );
  NAND2_X1 U13600 ( .A1(n14667), .A2(n11742), .ZN(n11743) );
  OAI211_X1 U13601 ( .C1(n14661), .C2(n11745), .A(n11744), .B(n11743), .ZN(
        n11746) );
  AOI21_X1 U13602 ( .B1(n14642), .B2(n11747), .A(n11746), .ZN(n11748) );
  OAI21_X1 U13603 ( .B1(n14697), .B2(n11749), .A(n11748), .ZN(P2_U3261) );
  XNOR2_X1 U13604 ( .A(n11750), .B(n11751), .ZN(n16007) );
  XNOR2_X1 U13605 ( .A(n11752), .B(n11751), .ZN(n11755) );
  INV_X1 U13606 ( .A(n11753), .ZN(n11754) );
  AOI21_X1 U13607 ( .B1(n11755), .B2(n14710), .A(n11754), .ZN(n16005) );
  MUX2_X1 U13608 ( .A(n11756), .B(n16005), .S(n12155), .Z(n11765) );
  INV_X1 U13609 ( .A(n11757), .ZN(n11760) );
  INV_X1 U13610 ( .A(n11758), .ZN(n11759) );
  AOI211_X1 U13611 ( .C1(n16003), .C2(n11760), .A(n14633), .B(n11759), .ZN(
        n16002) );
  OAI22_X1 U13612 ( .A1(n14661), .A2(n11762), .B1(n11761), .B2(n14718), .ZN(
        n11763) );
  AOI21_X1 U13613 ( .B1(n16002), .B2(n14667), .A(n11763), .ZN(n11764) );
  OAI211_X1 U13614 ( .C1(n14728), .C2(n16007), .A(n11765), .B(n11764), .ZN(
        P2_U3257) );
  MUX2_X1 U13615 ( .A(n11767), .B(n11766), .S(n12155), .Z(n11772) );
  INV_X1 U13616 ( .A(n14269), .ZN(n11768) );
  OAI22_X1 U13617 ( .A1(n14661), .A2(n11768), .B1(n14270), .B2(n14718), .ZN(
        n11769) );
  AOI21_X1 U13618 ( .B1(n14667), .B2(n11770), .A(n11769), .ZN(n11771) );
  OAI211_X1 U13619 ( .C1(n14728), .C2(n11773), .A(n11772), .B(n11771), .ZN(
        P2_U3260) );
  MUX2_X1 U13620 ( .A(n11775), .B(n11774), .S(n12155), .Z(n11781) );
  OAI22_X1 U13621 ( .A1(n14661), .A2(n11777), .B1(n11776), .B2(n14718), .ZN(
        n11778) );
  AOI21_X1 U13622 ( .B1(n14667), .B2(n11779), .A(n11778), .ZN(n11780) );
  OAI211_X1 U13623 ( .C1(n14728), .C2(n11782), .A(n11781), .B(n11780), .ZN(
        P2_U3259) );
  NAND2_X1 U13624 ( .A1(n11783), .A2(n14148), .ZN(n11784) );
  OAI211_X1 U13625 ( .C1(n11785), .C2(n14155), .A(n11784), .B(n13568), .ZN(
        P3_U3272) );
  OAI22_X1 U13626 ( .A1(n13983), .A2(n11787), .B1(n13380), .B2(n11786), .ZN(
        n11788) );
  OAI21_X1 U13627 ( .B1(n11789), .B2(n11788), .A(n13966), .ZN(n11793) );
  NAND2_X1 U13628 ( .A1(n13966), .A2(n13994), .ZN(n11790) );
  INV_X1 U13629 ( .A(n13968), .ZN(n13981) );
  NAND2_X1 U13630 ( .A1(n11791), .A2(n13981), .ZN(n11792) );
  OAI211_X1 U13631 ( .C1(n10705), .C2(n13966), .A(n11793), .B(n11792), .ZN(
        P3_U3232) );
  NAND2_X1 U13632 ( .A1(n11794), .A2(n12155), .ZN(n11802) );
  INV_X1 U13633 ( .A(n11795), .ZN(n11798) );
  INV_X1 U13634 ( .A(n14718), .ZN(n15884) );
  AOI22_X1 U13635 ( .A1(n14697), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11796), 
        .B2(n15884), .ZN(n11797) );
  OAI21_X1 U13636 ( .B1(n11798), .B2(n14661), .A(n11797), .ZN(n11799) );
  AOI21_X1 U13637 ( .B1(n11800), .B2(n14667), .A(n11799), .ZN(n11801) );
  OAI211_X1 U13638 ( .C1(n11803), .C2(n12150), .A(n11802), .B(n11801), .ZN(
        P2_U3256) );
  MUX2_X1 U13639 ( .A(n11805), .B(n11804), .S(n12155), .Z(n11811) );
  OAI22_X1 U13640 ( .A1(n14661), .A2(n11807), .B1(n11806), .B2(n14718), .ZN(
        n11808) );
  AOI21_X1 U13641 ( .B1(n11809), .B2(n14667), .A(n11808), .ZN(n11810) );
  OAI211_X1 U13642 ( .C1(n11812), .C2(n12150), .A(n11811), .B(n11810), .ZN(
        P2_U3258) );
  INV_X1 U13643 ( .A(n12072), .ZN(n11820) );
  OAI211_X1 U13644 ( .C1(n11815), .C2(n11814), .A(n11813), .B(n13343), .ZN(
        n11819) );
  INV_X1 U13645 ( .A(n13420), .ZN(n12167) );
  OAI22_X1 U13646 ( .A1(n13349), .A2(n13412), .B1(n12234), .B2(n13335), .ZN(
        n11816) );
  AOI211_X1 U13647 ( .C1(n12565), .C2(n12167), .A(n11817), .B(n11816), .ZN(
        n11818) );
  OAI211_X1 U13648 ( .C1(n11820), .C2(n12397), .A(n11819), .B(n11818), .ZN(
        P3_U3153) );
  OAI22_X1 U13649 ( .A1(n14725), .A2(n11821), .B1(n8912), .B2(n14718), .ZN(
        n11824) );
  NOR2_X1 U13650 ( .A1(n14661), .A2(n11822), .ZN(n11823) );
  AOI211_X1 U13651 ( .C1(n15891), .C2(P2_REG2_REG_2__SCAN_IN), .A(n11824), .B(
        n11823), .ZN(n11827) );
  NAND2_X1 U13652 ( .A1(n14642), .A2(n11825), .ZN(n11826) );
  OAI211_X1 U13653 ( .C1(n15891), .C2(n11828), .A(n11827), .B(n11826), .ZN(
        P2_U3263) );
  AOI21_X1 U13654 ( .B1(n11466), .B2(n11835), .A(n11829), .ZN(n15101) );
  INV_X1 U13655 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n12380) );
  MUX2_X1 U13656 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n12380), .S(n11837), .Z(
        n15100) );
  NAND2_X1 U13657 ( .A1(n15101), .A2(n15100), .ZN(n15099) );
  NAND2_X1 U13658 ( .A1(n11837), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11832) );
  INV_X1 U13659 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11830) );
  MUX2_X1 U13660 ( .A(n11830), .B(P1_REG2_REG_14__SCAN_IN), .S(n12488), .Z(
        n11831) );
  AOI21_X1 U13661 ( .B1(n15099), .B2(n11832), .A(n11831), .ZN(n12487) );
  NAND3_X1 U13662 ( .A1(n15099), .A2(n11832), .A3(n11831), .ZN(n11833) );
  NAND2_X1 U13663 ( .A1(n11833), .A2(n15143), .ZN(n11845) );
  INV_X1 U13664 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U13665 ( .A1(n11836), .A2(n16073), .B1(n11835), .B2(n11834), .ZN(
        n15095) );
  MUX2_X1 U13666 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n11838), .S(n11837), .Z(
        n15094) );
  NAND2_X1 U13667 ( .A1(n15095), .A2(n15094), .ZN(n15093) );
  OAI21_X1 U13668 ( .B1(n11838), .B2(n15096), .A(n15093), .ZN(n11840) );
  INV_X1 U13669 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n16105) );
  MUX2_X1 U13670 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n16105), .S(n12488), .Z(
        n11839) );
  NAND2_X1 U13671 ( .A1(n11840), .A2(n11839), .ZN(n12481) );
  OAI211_X1 U13672 ( .C1(n11840), .C2(n11839), .A(n12481), .B(n15652), .ZN(
        n11844) );
  NAND2_X1 U13673 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n16095)
         );
  INV_X1 U13674 ( .A(n16095), .ZN(n11842) );
  NOR2_X1 U13675 ( .A1(n15647), .A2(n12482), .ZN(n11841) );
  AOI211_X1 U13676 ( .C1(n15639), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n11842), 
        .B(n11841), .ZN(n11843) );
  OAI211_X1 U13677 ( .C1(n12487), .C2(n11845), .A(n11844), .B(n11843), .ZN(
        P1_U3257) );
  INV_X1 U13678 ( .A(n16019), .ZN(n11924) );
  AOI21_X1 U13679 ( .B1(n11847), .B2(n11846), .A(n15042), .ZN(n11849) );
  NAND2_X1 U13680 ( .A1(n11849), .A2(n11848), .ZN(n11852) );
  AND2_X1 U13681 ( .A1(n7201), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n15081) );
  AOI22_X1 U13682 ( .A1(n16030), .A2(n15068), .B1(n15067), .B2(n15376), .ZN(
        n11933) );
  NOR2_X1 U13683 ( .A1(n11933), .A2(n15026), .ZN(n11850) );
  AOI211_X1 U13684 ( .C1(n14987), .C2(n11922), .A(n15081), .B(n11850), .ZN(
        n11851) );
  OAI211_X1 U13685 ( .C1(n11924), .C2(n16091), .A(n11852), .B(n11851), .ZN(
        P1_U3231) );
  NAND2_X1 U13686 ( .A1(n12091), .A2(n14366), .ZN(n11853) );
  OR2_X1 U13687 ( .A1(n11856), .A2(n11861), .ZN(n11857) );
  INV_X1 U13688 ( .A(n12179), .ZN(n12294) );
  NAND2_X1 U13689 ( .A1(n12091), .A2(n12282), .ZN(n11860) );
  AOI21_X1 U13690 ( .B1(n11862), .B2(n11861), .A(n14679), .ZN(n11866) );
  NAND2_X1 U13691 ( .A1(n14364), .A2(n14338), .ZN(n11864) );
  NAND2_X1 U13692 ( .A1(n14366), .A2(n14525), .ZN(n11863) );
  AND2_X1 U13693 ( .A1(n11864), .A2(n11863), .ZN(n12289) );
  INV_X1 U13694 ( .A(n12289), .ZN(n11865) );
  AOI21_X1 U13695 ( .B1(n11866), .B2(n12011), .A(n11865), .ZN(n12115) );
  OAI211_X1 U13696 ( .C1(n11867), .C2(n12294), .A(n14716), .B(n12019), .ZN(
        n12111) );
  OAI211_X1 U13697 ( .C1(n12294), .C2(n16149), .A(n12115), .B(n12111), .ZN(
        n11868) );
  AOI21_X1 U13698 ( .B1(n14803), .B2(n12113), .A(n11868), .ZN(n11875) );
  INV_X1 U13699 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11869) );
  NOR2_X1 U13700 ( .A1(n16117), .A2(n11869), .ZN(n11870) );
  AOI21_X1 U13701 ( .B1(n12113), .B2(n12462), .A(n11870), .ZN(n11871) );
  OAI21_X1 U13702 ( .B1(n11875), .B2(n16157), .A(n11871), .ZN(P2_U3466) );
  OAI222_X1 U13703 ( .A1(n14871), .A2(n11873), .B1(P2_U3088), .B2(n8886), .C1(
        n14869), .C2(n11872), .ZN(P2_U3305) );
  AOI22_X1 U13704 ( .A1(n12113), .A2(n12464), .B1(n16155), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n11874) );
  OAI21_X1 U13705 ( .B1(n11875), .B2(n16155), .A(n11874), .ZN(P2_U3511) );
  OAI22_X1 U13706 ( .A1(n14725), .A2(n11877), .B1(n11876), .B2(n14718), .ZN(
        n11878) );
  AOI21_X1 U13707 ( .B1(n14722), .B2(n11879), .A(n11878), .ZN(n11883) );
  MUX2_X1 U13708 ( .A(n11881), .B(n11880), .S(n15891), .Z(n11882) );
  OAI211_X1 U13709 ( .C1(n14728), .C2(n11884), .A(n11883), .B(n11882), .ZN(
        P2_U3264) );
  NAND2_X1 U13710 ( .A1(n11886), .A2(n11955), .ZN(n13403) );
  NAND2_X1 U13711 ( .A1(n13412), .A2(n13411), .ZN(n13414) );
  NAND2_X1 U13712 ( .A1(n13581), .A2(n15939), .ZN(n13415) );
  NAND2_X1 U13713 ( .A1(n13414), .A2(n13415), .ZN(n13526) );
  XNOR2_X1 U13714 ( .A(n11959), .B(n13526), .ZN(n15941) );
  INV_X1 U13715 ( .A(n15941), .ZN(n11897) );
  INV_X1 U13716 ( .A(n13580), .ZN(n12163) );
  OAI22_X1 U13717 ( .A1(n11886), .A2(n13946), .B1(n12163), .B2(n13944), .ZN(
        n11893) );
  NOR2_X1 U13718 ( .A1(n13582), .A2(n11955), .ZN(n11888) );
  OAI21_X1 U13719 ( .B1(n11887), .B2(n11888), .A(n13526), .ZN(n11891) );
  NOR2_X1 U13720 ( .A1(n13526), .A2(n11888), .ZN(n11889) );
  AND3_X1 U13721 ( .A1(n11962), .A2(n13970), .A3(n11891), .ZN(n11892) );
  AOI211_X1 U13722 ( .C1(n13994), .C2(n15941), .A(n11893), .B(n11892), .ZN(
        n15943) );
  MUX2_X1 U13723 ( .A(n11894), .B(n15943), .S(n13966), .Z(n11896) );
  AOI22_X1 U13724 ( .A1(n13986), .A2(n15939), .B1(n14004), .B2(n11947), .ZN(
        n11895) );
  OAI211_X1 U13725 ( .C1(n11897), .C2(n12254), .A(n11896), .B(n11895), .ZN(
        P3_U3227) );
  OR2_X1 U13726 ( .A1(n11898), .A2(n8243), .ZN(n11899) );
  NAND2_X1 U13727 ( .A1(n11900), .A2(n11899), .ZN(n15902) );
  OAI22_X1 U13728 ( .A1(n14006), .A2(n15899), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n13983), .ZN(n11912) );
  NAND2_X1 U13729 ( .A1(n15902), .A2(n13994), .ZN(n11910) );
  AND2_X1 U13730 ( .A1(n11901), .A2(n13970), .ZN(n11908) );
  NAND2_X1 U13731 ( .A1(n11675), .A2(n11902), .ZN(n11903) );
  NAND2_X1 U13732 ( .A1(n11903), .A2(n8243), .ZN(n11907) );
  OAI22_X1 U13733 ( .A1(n11905), .A2(n13946), .B1(n11904), .B2(n13944), .ZN(
        n11906) );
  AOI21_X1 U13734 ( .B1(n11908), .B2(n11907), .A(n11906), .ZN(n11909) );
  NAND2_X1 U13735 ( .A1(n11910), .A2(n11909), .ZN(n15900) );
  INV_X2 U13736 ( .A(n13966), .ZN(n13963) );
  MUX2_X1 U13737 ( .A(n15900), .B(P3_REG2_REG_3__SCAN_IN), .S(n13963), .Z(
        n11911) );
  AOI211_X1 U13738 ( .C1(n14008), .C2(n15902), .A(n11912), .B(n11911), .ZN(
        n11913) );
  INV_X1 U13739 ( .A(n11913), .ZN(P3_U3230) );
  XNOR2_X1 U13740 ( .A(n16019), .B(n16029), .ZN(n12864) );
  OR2_X1 U13741 ( .A1(n12725), .A2(n15069), .ZN(n11916) );
  INV_X1 U13742 ( .A(n15068), .ZN(n11931) );
  XNOR2_X1 U13743 ( .A(n15992), .B(n11931), .ZN(n15983) );
  NAND2_X1 U13744 ( .A1(n15992), .A2(n15068), .ZN(n11917) );
  NAND2_X1 U13745 ( .A1(n15973), .A2(n11917), .ZN(n11921) );
  INV_X1 U13746 ( .A(n11921), .ZN(n11919) );
  NAND2_X1 U13747 ( .A1(n11919), .A2(n11918), .ZN(n11978) );
  INV_X1 U13748 ( .A(n11978), .ZN(n11920) );
  AOI21_X1 U13749 ( .B1(n12864), .B2(n11921), .A(n11920), .ZN(n16022) );
  AOI211_X1 U13750 ( .C1(n16019), .C2(n15976), .A(n15974), .B(n11972), .ZN(
        n16018) );
  INV_X1 U13751 ( .A(n11922), .ZN(n11923) );
  OAI22_X1 U13752 ( .A1(n11924), .A2(n15365), .B1(n15377), .B2(n11923), .ZN(
        n11925) );
  AOI21_X1 U13753 ( .B1(n16018), .B2(n15368), .A(n11925), .ZN(n11938) );
  NAND2_X1 U13754 ( .A1(n12725), .A2(n11927), .ZN(n11928) );
  NAND2_X1 U13755 ( .A1(n11929), .A2(n11928), .ZN(n15982) );
  OR2_X1 U13756 ( .A1(n15992), .A2(n11931), .ZN(n11932) );
  XNOR2_X1 U13757 ( .A(n11968), .B(n12864), .ZN(n11934) );
  OAI21_X1 U13758 ( .B1(n11934), .B2(n16136), .A(n11933), .ZN(n16024) );
  INV_X1 U13759 ( .A(n16024), .ZN(n11935) );
  MUX2_X1 U13760 ( .A(n11936), .B(n11935), .S(n7218), .Z(n11937) );
  OAI211_X1 U13761 ( .C1(n16022), .C2(n15392), .A(n11938), .B(n11937), .ZN(
        P1_U3284) );
  INV_X1 U13762 ( .A(n13335), .ZN(n13346) );
  AOI22_X1 U13763 ( .A1(n13346), .A2(n13580), .B1(n13318), .B2(n13582), .ZN(
        n11940) );
  OAI211_X1 U13764 ( .C1(n13411), .C2(n13354), .A(n11940), .B(n11939), .ZN(
        n11946) );
  INV_X1 U13765 ( .A(n11941), .ZN(n11942) );
  AOI211_X1 U13766 ( .C1(n11944), .C2(n11943), .A(n13314), .B(n11942), .ZN(
        n11945) );
  AOI211_X1 U13767 ( .C1(n11947), .C2(n13351), .A(n11946), .B(n11945), .ZN(
        n11948) );
  INV_X1 U13768 ( .A(n11948), .ZN(P3_U3179) );
  INV_X1 U13769 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12612) );
  NAND2_X1 U13770 ( .A1(n12611), .A2(n11949), .ZN(n11950) );
  OAI211_X1 U13771 ( .C1(n12612), .C2(n11951), .A(n11950), .B(n12913), .ZN(
        P1_U3332) );
  NAND2_X1 U13772 ( .A1(n12611), .A2(n14861), .ZN(n11953) );
  OAI211_X1 U13773 ( .C1(n11954), .C2(n14866), .A(n11953), .B(n11952), .ZN(
        P2_U3304) );
  INV_X1 U13774 ( .A(n11955), .ZN(n13402) );
  MUX2_X1 U13775 ( .A(n10971), .B(n11956), .S(n16061), .Z(n11957) );
  OAI21_X1 U13776 ( .B1(n14083), .B2(n13402), .A(n11957), .ZN(P3_U3464) );
  NAND2_X1 U13777 ( .A1(n13581), .A2(n13411), .ZN(n11958) );
  NAND2_X1 U13778 ( .A1(n11959), .A2(n11958), .ZN(n11961) );
  NAND2_X1 U13779 ( .A1(n13412), .A2(n15939), .ZN(n11960) );
  XNOR2_X1 U13780 ( .A(n13580), .B(n13420), .ZN(n13529) );
  XNOR2_X1 U13781 ( .A(n12162), .B(n13529), .ZN(n12075) );
  INV_X1 U13782 ( .A(n12075), .ZN(n11966) );
  INV_X1 U13783 ( .A(n13529), .ZN(n12161) );
  XNOR2_X1 U13784 ( .A(n12166), .B(n12161), .ZN(n11964) );
  OAI22_X1 U13785 ( .A1(n13412), .A2(n13946), .B1(n12234), .B2(n13944), .ZN(
        n11963) );
  AOI21_X1 U13786 ( .B1(n11964), .B2(n13970), .A(n11963), .ZN(n11965) );
  OAI21_X1 U13787 ( .B1(n12075), .B2(n13885), .A(n11965), .ZN(n12069) );
  AOI21_X1 U13788 ( .B1(n16059), .B2(n11966), .A(n12069), .ZN(n12139) );
  AOI22_X1 U13789 ( .A1(n14124), .A2(n12167), .B1(P3_REG0_REG_7__SCAN_IN), 
        .B2(n16062), .ZN(n11967) );
  OAI21_X1 U13790 ( .B1(n12139), .B2(n16062), .A(n11967), .ZN(P3_U3411) );
  INV_X1 U13791 ( .A(n16029), .ZN(n12083) );
  OR2_X1 U13792 ( .A1(n16019), .A2(n12083), .ZN(n11969) );
  NAND2_X1 U13793 ( .A1(n11970), .A2(n11969), .ZN(n11981) );
  XNOR2_X1 U13794 ( .A(n11981), .B(n12737), .ZN(n16034) );
  AOI22_X1 U13795 ( .A1(n16001), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n12081), 
        .B2(n15990), .ZN(n11971) );
  OAI21_X1 U13796 ( .B1(n15173), .B2(n12083), .A(n11971), .ZN(n11976) );
  INV_X1 U13797 ( .A(n11972), .ZN(n11973) );
  INV_X1 U13798 ( .A(n16031), .ZN(n12088) );
  AND2_X2 U13799 ( .A1(n11972), .A2(n12088), .ZN(n12310) );
  AOI211_X1 U13800 ( .C1(n16031), .C2(n11973), .A(n15974), .B(n12310), .ZN(
        n11974) );
  AOI21_X1 U13801 ( .B1(n15376), .B2(n15066), .A(n11974), .ZN(n16033) );
  NOR2_X1 U13802 ( .A1(n16033), .A2(n15993), .ZN(n11975) );
  AOI211_X1 U13803 ( .C1(n15991), .C2(n16031), .A(n11976), .B(n11975), .ZN(
        n11980) );
  OR2_X1 U13804 ( .A1(n16019), .A2(n16029), .ZN(n11977) );
  NAND2_X1 U13805 ( .A1(n11978), .A2(n11977), .ZN(n11993) );
  XNOR2_X1 U13806 ( .A(n11993), .B(n12868), .ZN(n16036) );
  NAND2_X1 U13807 ( .A1(n16036), .A2(n15355), .ZN(n11979) );
  OAI211_X1 U13808 ( .C1(n16034), .C2(n15371), .A(n11980), .B(n11979), .ZN(
        P1_U3283) );
  INV_X1 U13809 ( .A(n15067), .ZN(n11982) );
  XNOR2_X1 U13810 ( .A(n12744), .B(n15066), .ZN(n12863) );
  INV_X1 U13811 ( .A(n12863), .ZN(n11984) );
  XNOR2_X1 U13812 ( .A(n12298), .B(n11984), .ZN(n11985) );
  NAND2_X1 U13813 ( .A1(n11985), .A2(n16119), .ZN(n11987) );
  AOI22_X1 U13814 ( .A1(n15376), .A2(n15065), .B1(n15067), .B2(n16030), .ZN(
        n11986) );
  NAND2_X1 U13815 ( .A1(n11987), .A2(n11986), .ZN(n16050) );
  INV_X1 U13816 ( .A(n16050), .ZN(n11998) );
  INV_X1 U13817 ( .A(n12262), .ZN(n11988) );
  OAI22_X1 U13818 ( .A1(n7218), .A2(n11989), .B1(n11988), .B2(n15377), .ZN(
        n11992) );
  XNOR2_X1 U13819 ( .A(n12310), .B(n12744), .ZN(n11990) );
  NAND2_X1 U13820 ( .A1(n11990), .A2(n15445), .ZN(n16047) );
  NOR2_X1 U13821 ( .A1(n16047), .A2(n15993), .ZN(n11991) );
  AOI211_X1 U13822 ( .C1(n15991), .C2(n12744), .A(n11992), .B(n11991), .ZN(
        n11997) );
  OR2_X1 U13823 ( .A1(n16031), .A2(n15067), .ZN(n11994) );
  NAND2_X1 U13824 ( .A1(n11995), .A2(n12863), .ZN(n16046) );
  NAND3_X1 U13825 ( .A1(n12302), .A2(n16046), .A3(n15355), .ZN(n11996) );
  OAI211_X1 U13826 ( .C1(n11998), .C2(n16001), .A(n11997), .B(n11996), .ZN(
        P1_U3282) );
  INV_X1 U13827 ( .A(n11999), .ZN(n12250) );
  OAI211_X1 U13828 ( .C1(n12002), .C2(n12001), .A(n12000), .B(n13343), .ZN(
        n12006) );
  OAI22_X1 U13829 ( .A1(n13349), .A2(n12163), .B1(n12392), .B2(n13335), .ZN(
        n12003) );
  AOI211_X1 U13830 ( .C1(n12565), .C2(n12165), .A(n12004), .B(n12003), .ZN(
        n12005) );
  OAI211_X1 U13831 ( .C1(n12250), .C2(n12397), .A(n12006), .B(n12005), .ZN(
        P3_U3161) );
  NAND2_X1 U13832 ( .A1(n12179), .A2(n14365), .ZN(n12007) );
  INV_X1 U13833 ( .A(n12012), .ZN(n12014) );
  OAI21_X1 U13834 ( .B1(n7361), .B2(n12012), .A(n12126), .ZN(n12136) );
  INV_X1 U13835 ( .A(n12192), .ZN(n12021) );
  INV_X1 U13836 ( .A(n14365), .ZN(n12009) );
  OR2_X1 U13837 ( .A1(n12179), .A2(n12009), .ZN(n12010) );
  NAND2_X1 U13838 ( .A1(n12011), .A2(n12010), .ZN(n12015) );
  INV_X1 U13839 ( .A(n12015), .ZN(n12013) );
  AOI21_X1 U13840 ( .B1(n12013), .B2(n12012), .A(n14679), .ZN(n12018) );
  NAND2_X1 U13841 ( .A1(n14365), .A2(n14525), .ZN(n12017) );
  NAND2_X1 U13842 ( .A1(n14363), .A2(n14338), .ZN(n12016) );
  NAND2_X1 U13843 ( .A1(n12017), .A2(n12016), .ZN(n12185) );
  AOI21_X1 U13844 ( .B1(n12018), .B2(n12117), .A(n12185), .ZN(n12138) );
  INV_X1 U13845 ( .A(n12019), .ZN(n12020) );
  OAI211_X1 U13846 ( .C1(n12020), .C2(n12021), .A(n14716), .B(n12120), .ZN(
        n12134) );
  OAI211_X1 U13847 ( .C1(n12021), .C2(n16149), .A(n12138), .B(n12134), .ZN(
        n12022) );
  AOI21_X1 U13848 ( .B1(n14803), .B2(n12136), .A(n12022), .ZN(n12077) );
  INV_X1 U13849 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n12023) );
  NOR2_X1 U13850 ( .A1(n16117), .A2(n12023), .ZN(n12024) );
  AOI21_X1 U13851 ( .B1(n12136), .B2(n12462), .A(n12024), .ZN(n12025) );
  OAI21_X1 U13852 ( .B1(n12077), .B2(n16157), .A(n12025), .ZN(P2_U3469) );
  NAND2_X1 U13853 ( .A1(n12027), .A2(n12026), .ZN(n12028) );
  NAND2_X1 U13854 ( .A1(n12029), .A2(n12028), .ZN(n15838) );
  INV_X1 U13855 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12216) );
  INV_X1 U13856 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12030) );
  MUX2_X1 U13857 ( .A(n12216), .B(n12030), .S(n10630), .Z(n12031) );
  NAND2_X1 U13858 ( .A1(n12031), .A2(n12058), .ZN(n12034) );
  INV_X1 U13859 ( .A(n12031), .ZN(n12032) );
  NAND2_X1 U13860 ( .A1(n12032), .A2(n15834), .ZN(n12033) );
  NAND2_X1 U13861 ( .A1(n12034), .A2(n12033), .ZN(n15837) );
  NAND2_X1 U13862 ( .A1(n15835), .A2(n12034), .ZN(n15862) );
  MUX2_X1 U13863 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n10630), .Z(n12035) );
  XNOR2_X1 U13864 ( .A(n12035), .B(n12036), .ZN(n15861) );
  NAND2_X1 U13865 ( .A1(n15862), .A2(n15861), .ZN(n15860) );
  INV_X1 U13866 ( .A(n12035), .ZN(n12037) );
  NAND2_X1 U13867 ( .A1(n12037), .A2(n12036), .ZN(n12043) );
  NAND2_X1 U13868 ( .A1(n12051), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n13605) );
  OR2_X1 U13869 ( .A1(n12051), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12038) );
  AND2_X1 U13870 ( .A1(n13605), .A2(n12038), .ZN(n12041) );
  NAND2_X1 U13871 ( .A1(n12051), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n13604) );
  OR2_X1 U13872 ( .A1(n12051), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12039) );
  NAND2_X1 U13873 ( .A1(n13604), .A2(n12039), .ZN(n12063) );
  INV_X1 U13874 ( .A(n12063), .ZN(n12040) );
  MUX2_X1 U13875 ( .A(n12041), .B(n12040), .S(n10630), .Z(n12042) );
  AOI21_X1 U13876 ( .B1(n15860), .B2(n12043), .A(n12042), .ZN(n12068) );
  AND2_X1 U13877 ( .A1(n12043), .A2(n12042), .ZN(n12044) );
  NAND2_X1 U13878 ( .A1(n15860), .A2(n12044), .ZN(n13607) );
  NAND2_X1 U13879 ( .A1(n13607), .A2(n15863), .ZN(n12067) );
  INV_X1 U13880 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n13174) );
  NOR2_X1 U13881 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13174), .ZN(n12563) );
  AOI22_X1 U13882 ( .A1(n12058), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n12216), 
        .B2(n15834), .ZN(n15832) );
  NAND2_X1 U13883 ( .A1(n12048), .A2(n15855), .ZN(n12047) );
  INV_X1 U13884 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n15852) );
  OAI21_X1 U13885 ( .B1(n12048), .B2(n15855), .A(n12047), .ZN(n15851) );
  OAI21_X1 U13886 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n12051), .A(n13605), 
        .ZN(n12049) );
  AOI21_X1 U13887 ( .B1(n12050), .B2(n12049), .A(n13589), .ZN(n12054) );
  INV_X1 U13888 ( .A(n12051), .ZN(n12052) );
  AOI22_X1 U13889 ( .A1(n13754), .A2(n12052), .B1(n15521), .B2(
        P3_ADDR_REG_12__SCAN_IN), .ZN(n12053) );
  OAI21_X1 U13890 ( .B1(n15872), .B2(n12054), .A(n12053), .ZN(n12055) );
  NOR2_X1 U13891 ( .A1(n12563), .A2(n12055), .ZN(n12066) );
  AOI22_X1 U13892 ( .A1(n12058), .A2(P3_REG1_REG_10__SCAN_IN), .B1(n12030), 
        .B2(n15834), .ZN(n15840) );
  INV_X1 U13893 ( .A(n12059), .ZN(n12061) );
  INV_X1 U13894 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n15858) );
  NOR2_X1 U13895 ( .A1(n12062), .A2(n12063), .ZN(n13595) );
  AND2_X1 U13896 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  OAI21_X1 U13897 ( .B1(n13595), .B2(n12064), .A(n13722), .ZN(n12065) );
  OAI211_X1 U13898 ( .C1(n12068), .C2(n12067), .A(n12066), .B(n12065), .ZN(
        P3_U3194) );
  INV_X1 U13899 ( .A(n12069), .ZN(n12070) );
  MUX2_X1 U13900 ( .A(n12071), .B(n12070), .S(n13966), .Z(n12074) );
  AOI22_X1 U13901 ( .A1(n13986), .A2(n12167), .B1(n14004), .B2(n12072), .ZN(
        n12073) );
  OAI211_X1 U13902 ( .C1(n12075), .C2(n12254), .A(n12074), .B(n12073), .ZN(
        P3_U3226) );
  AOI22_X1 U13903 ( .A1(n12136), .A2(n12464), .B1(n16155), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n12076) );
  OAI21_X1 U13904 ( .B1(n12077), .B2(n16155), .A(n12076), .ZN(P2_U3512) );
  OAI211_X1 U13905 ( .C1(n12080), .C2(n12079), .A(n12078), .B(n16093), .ZN(
        n12087) );
  INV_X1 U13906 ( .A(n12081), .ZN(n12082) );
  OAI22_X1 U13907 ( .A1(n12083), .A2(n15049), .B1(n12082), .B2(n16098), .ZN(
        n12084) );
  AOI211_X1 U13908 ( .C1(n16089), .C2(n15066), .A(n12085), .B(n12084), .ZN(
        n12086) );
  OAI211_X1 U13909 ( .C1(n12088), .C2(n16091), .A(n12087), .B(n12086), .ZN(
        P1_U3217) );
  INV_X1 U13910 ( .A(n12089), .ZN(n12098) );
  AOI22_X1 U13911 ( .A1(n14697), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n12090), 
        .B2(n15884), .ZN(n12093) );
  NAND2_X1 U13912 ( .A1(n14722), .A2(n12091), .ZN(n12092) );
  OAI211_X1 U13913 ( .C1(n12094), .C2(n14725), .A(n12093), .B(n12092), .ZN(
        n12095) );
  AOI21_X1 U13914 ( .B1(n12096), .B2(n14642), .A(n12095), .ZN(n12097) );
  OAI21_X1 U13915 ( .B1(n12098), .B2(n15891), .A(n12097), .ZN(P2_U3254) );
  NAND2_X1 U13916 ( .A1(n14722), .A2(n12099), .ZN(n12102) );
  NOR2_X1 U13917 ( .A1(n14718), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n12100) );
  AOI21_X1 U13918 ( .B1(n14697), .B2(P2_REG2_REG_3__SCAN_IN), .A(n12100), .ZN(
        n12101) );
  OAI211_X1 U13919 ( .C1(n12103), .C2(n14725), .A(n12102), .B(n12101), .ZN(
        n12104) );
  AOI21_X1 U13920 ( .B1(n14642), .B2(n12105), .A(n12104), .ZN(n12106) );
  OAI21_X1 U13921 ( .B1(n14697), .B2(n12107), .A(n12106), .ZN(P2_U3262) );
  INV_X1 U13922 ( .A(n12108), .ZN(n12291) );
  AOI22_X1 U13923 ( .A1(n14697), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n12291), 
        .B2(n15884), .ZN(n12110) );
  NAND2_X1 U13924 ( .A1(n12179), .A2(n14722), .ZN(n12109) );
  OAI211_X1 U13925 ( .C1(n12111), .C2(n14725), .A(n12110), .B(n12109), .ZN(
        n12112) );
  AOI21_X1 U13926 ( .B1(n12113), .B2(n14642), .A(n12112), .ZN(n12114) );
  OAI21_X1 U13927 ( .B1(n15891), .B2(n12115), .A(n12114), .ZN(P2_U3253) );
  OR2_X1 U13928 ( .A1(n12192), .A2(n12184), .ZN(n12116) );
  NAND2_X1 U13929 ( .A1(n12117), .A2(n12116), .ZN(n12351) );
  XNOR2_X1 U13930 ( .A(n12351), .B(n8076), .ZN(n12119) );
  AOI22_X1 U13931 ( .A1(n14362), .A2(n14338), .B1(n14364), .B2(n14525), .ZN(
        n12271) );
  INV_X1 U13932 ( .A(n12271), .ZN(n12118) );
  AOI21_X1 U13933 ( .B1(n12119), .B2(n14710), .A(n12118), .ZN(n16114) );
  AOI211_X1 U13934 ( .C1(n16111), .C2(n12120), .A(n14633), .B(n12359), .ZN(
        n16110) );
  INV_X1 U13935 ( .A(n16111), .ZN(n12121) );
  NOR2_X1 U13936 ( .A1(n12121), .A2(n14661), .ZN(n12124) );
  OAI22_X1 U13937 ( .A1(n12155), .A2(n12122), .B1(n12269), .B2(n14718), .ZN(
        n12123) );
  AOI211_X1 U13938 ( .C1(n16110), .C2(n14667), .A(n12124), .B(n12123), .ZN(
        n12130) );
  OR2_X1 U13939 ( .A1(n12192), .A2(n14364), .ZN(n12125) );
  NAND2_X1 U13940 ( .A1(n12128), .A2(n12127), .ZN(n16108) );
  NAND3_X1 U13941 ( .A1(n16109), .A2(n14642), .A3(n16108), .ZN(n12129) );
  OAI211_X1 U13942 ( .C1(n16114), .C2(n15891), .A(n12130), .B(n12129), .ZN(
        P2_U3251) );
  OAI22_X1 U13943 ( .A1(n12155), .A2(n12131), .B1(n12187), .B2(n14718), .ZN(
        n12132) );
  AOI21_X1 U13944 ( .B1(n12192), .B2(n14722), .A(n12132), .ZN(n12133) );
  OAI21_X1 U13945 ( .B1(n12134), .B2(n14725), .A(n12133), .ZN(n12135) );
  AOI21_X1 U13946 ( .B1(n12136), .B2(n14642), .A(n12135), .ZN(n12137) );
  OAI21_X1 U13947 ( .B1(n14697), .B2(n12138), .A(n12137), .ZN(P2_U3252) );
  MUX2_X1 U13948 ( .A(n12140), .B(n12139), .S(n16061), .Z(n12141) );
  OAI21_X1 U13949 ( .B1(n14083), .B2(n13420), .A(n12141), .ZN(P3_U3466) );
  INV_X1 U13950 ( .A(n12144), .ZN(n12142) );
  XNOR2_X1 U13951 ( .A(n12143), .B(n12142), .ZN(n16042) );
  NAND2_X1 U13952 ( .A1(n16042), .A2(n14803), .ZN(n12149) );
  XNOR2_X1 U13953 ( .A(n12145), .B(n12144), .ZN(n12147) );
  AOI21_X1 U13954 ( .B1(n12147), .B2(n14710), .A(n12146), .ZN(n12148) );
  INV_X1 U13955 ( .A(n12150), .ZN(n15887) );
  AOI21_X1 U13956 ( .B1(n12157), .B2(n12151), .A(n14633), .ZN(n12153) );
  NAND2_X1 U13957 ( .A1(n12153), .A2(n12152), .ZN(n16039) );
  OAI22_X1 U13958 ( .A1(n12155), .A2(n14429), .B1(n12154), .B2(n14718), .ZN(
        n12156) );
  AOI21_X1 U13959 ( .B1(n12157), .B2(n14722), .A(n12156), .ZN(n12158) );
  OAI21_X1 U13960 ( .B1(n16039), .B2(n14725), .A(n12158), .ZN(n12159) );
  AOI21_X1 U13961 ( .B1(n16042), .B2(n15887), .A(n12159), .ZN(n12160) );
  OAI21_X1 U13962 ( .B1(n16044), .B2(n15891), .A(n12160), .ZN(P2_U3255) );
  NAND2_X1 U13963 ( .A1(n12162), .A2(n12161), .ZN(n12164) );
  NAND2_X1 U13964 ( .A1(n12163), .A2(n12167), .ZN(n13421) );
  NAND2_X1 U13965 ( .A1(n12234), .A2(n12165), .ZN(n13426) );
  INV_X1 U13966 ( .A(n12234), .ZN(n13579) );
  INV_X1 U13967 ( .A(n12165), .ZN(n15964) );
  NAND2_X1 U13968 ( .A1(n13579), .A2(n15964), .ZN(n13430) );
  INV_X1 U13969 ( .A(n12237), .ZN(n16010) );
  NOR2_X1 U13970 ( .A1(n13578), .A2(n16010), .ZN(n13432) );
  OR2_X1 U13971 ( .A1(n7244), .A2(n13432), .ZN(n13522) );
  XNOR2_X1 U13972 ( .A(n12202), .B(n13522), .ZN(n16012) );
  NAND2_X1 U13973 ( .A1(n13580), .A2(n12167), .ZN(n12168) );
  NAND2_X1 U13974 ( .A1(n12234), .A2(n15964), .ZN(n12208) );
  NAND2_X1 U13975 ( .A1(n12243), .A2(n12208), .ZN(n12203) );
  XNOR2_X1 U13976 ( .A(n12203), .B(n13522), .ZN(n12171) );
  OAI22_X1 U13977 ( .A1(n12234), .A2(n13946), .B1(n12474), .B2(n13944), .ZN(
        n12170) );
  AOI21_X1 U13978 ( .B1(n12171), .B2(n13970), .A(n12170), .ZN(n12172) );
  OAI21_X1 U13979 ( .B1(n16012), .B2(n13885), .A(n12172), .ZN(n16014) );
  INV_X1 U13980 ( .A(n16014), .ZN(n12178) );
  INV_X1 U13981 ( .A(n16012), .ZN(n12176) );
  AOI22_X1 U13982 ( .A1(n13986), .A2(n12237), .B1(n14004), .B2(n12238), .ZN(
        n12173) );
  OAI21_X1 U13983 ( .B1(n12174), .B2(n13966), .A(n12173), .ZN(n12175) );
  AOI21_X1 U13984 ( .B1(n12176), .B2(n14008), .A(n12175), .ZN(n12177) );
  OAI21_X1 U13985 ( .B1(n12178), .B2(n13963), .A(n12177), .ZN(P3_U3224) );
  XNOR2_X1 U13986 ( .A(n12179), .B(n14229), .ZN(n12188) );
  INV_X1 U13987 ( .A(n12188), .ZN(n12183) );
  NAND2_X1 U13988 ( .A1(n14365), .A2(n14633), .ZN(n12182) );
  NAND2_X1 U13989 ( .A1(n12284), .A2(n12283), .ZN(n12280) );
  XNOR2_X1 U13990 ( .A(n12188), .B(n12182), .ZN(n12285) );
  OAI21_X1 U13991 ( .B1(n12284), .B2(n12283), .A(n12285), .ZN(n12180) );
  XNOR2_X1 U13992 ( .A(n12192), .B(n14229), .ZN(n12274) );
  NOR2_X1 U13993 ( .A1(n12184), .A2(n14716), .ZN(n12268) );
  INV_X1 U13994 ( .A(n12277), .ZN(n12194) );
  AOI22_X1 U13995 ( .A1(n14348), .A2(n12185), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12186) );
  OAI21_X1 U13996 ( .B1(n14351), .B2(n12187), .A(n12186), .ZN(n12191) );
  AOI22_X1 U13997 ( .A1(n12188), .A2(n14311), .B1(n14330), .B2(n14365), .ZN(
        n12189) );
  NOR3_X1 U13998 ( .A1(n12296), .A2(n12189), .A3(n7371), .ZN(n12190) );
  AOI211_X1 U13999 ( .C1(n12192), .C2(n14358), .A(n12191), .B(n12190), .ZN(
        n12193) );
  OAI21_X1 U14000 ( .B1(n14353), .B2(n12194), .A(n12193), .ZN(P2_U3206) );
  INV_X1 U14001 ( .A(n12195), .ZN(n12196) );
  OAI222_X1 U14002 ( .A1(n12197), .A2(P3_U3151), .B1(n14158), .B2(n12196), 
        .C1(n13005), .C2(n14155), .ZN(P3_U3271) );
  INV_X1 U14003 ( .A(n12598), .ZN(n12200) );
  OAI222_X1 U14004 ( .A1(n15512), .A2(n12599), .B1(n15510), .B2(n12200), .C1(
        n12198), .C2(n7201), .ZN(P1_U3331) );
  OAI222_X1 U14005 ( .A1(n14871), .A2(n12201), .B1(n14869), .B2(n12200), .C1(
        P2_U3088), .C2(n12199), .ZN(P2_U3303) );
  NAND2_X1 U14006 ( .A1(n12474), .A2(n12394), .ZN(n13435) );
  INV_X1 U14007 ( .A(n12474), .ZN(n13577) );
  INV_X1 U14008 ( .A(n12394), .ZN(n12226) );
  NAND2_X1 U14009 ( .A1(n13577), .A2(n12226), .ZN(n13428) );
  OAI21_X1 U14010 ( .B1(n7372), .B2(n12205), .A(n12369), .ZN(n12223) );
  INV_X1 U14011 ( .A(n12223), .ZN(n12221) );
  NAND2_X1 U14012 ( .A1(n13578), .A2(n12237), .ZN(n12210) );
  NAND2_X1 U14013 ( .A1(n12203), .A2(n12210), .ZN(n12204) );
  NAND2_X1 U14014 ( .A1(n12392), .A2(n16010), .ZN(n12206) );
  AND2_X1 U14015 ( .A1(n12204), .A2(n12206), .ZN(n12213) );
  INV_X1 U14016 ( .A(n12205), .ZN(n12207) );
  AND2_X1 U14017 ( .A1(n12207), .A2(n12206), .ZN(n12209) );
  AND2_X1 U14018 ( .A1(n12208), .A2(n12209), .ZN(n12212) );
  INV_X1 U14019 ( .A(n12209), .ZN(n12211) );
  OAI211_X1 U14020 ( .C1(n12213), .C2(n12207), .A(n13970), .B(n12367), .ZN(
        n12215) );
  AOI22_X1 U14021 ( .A1(n13998), .A2(n13996), .B1(n13997), .B2(n13578), .ZN(
        n12214) );
  NAND2_X1 U14022 ( .A1(n12215), .A2(n12214), .ZN(n12222) );
  NOR2_X1 U14023 ( .A1(n13966), .A2(n12216), .ZN(n12219) );
  INV_X1 U14024 ( .A(n12217), .ZN(n12398) );
  OAI22_X1 U14025 ( .A1(n14006), .A2(n12226), .B1(n12398), .B2(n13983), .ZN(
        n12218) );
  AOI211_X1 U14026 ( .C1(n12222), .C2(n13966), .A(n12219), .B(n12218), .ZN(
        n12220) );
  OAI21_X1 U14027 ( .B1(n12221), .B2(n13968), .A(n12220), .ZN(P3_U3223) );
  AOI21_X1 U14028 ( .B1(n12223), .B2(n14080), .A(n12222), .ZN(n12229) );
  AOI22_X1 U14029 ( .A1(n14063), .A2(n12394), .B1(n12991), .B2(
        P3_REG1_REG_10__SCAN_IN), .ZN(n12224) );
  OAI21_X1 U14030 ( .B1(n12229), .B2(n12991), .A(n12224), .ZN(P3_U3469) );
  INV_X1 U14031 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n12225) );
  OAI22_X1 U14032 ( .A1(n14142), .A2(n12226), .B1(n12225), .B2(n16065), .ZN(
        n12227) );
  INV_X1 U14033 ( .A(n12227), .ZN(n12228) );
  OAI21_X1 U14034 ( .B1(n12229), .B2(n16062), .A(n12228), .ZN(P3_U3420) );
  INV_X1 U14035 ( .A(n12230), .ZN(n12231) );
  AOI21_X1 U14036 ( .B1(n12233), .B2(n12232), .A(n12231), .ZN(n12241) );
  OAI22_X1 U14037 ( .A1(n13349), .A2(n12234), .B1(n12474), .B2(n13335), .ZN(
        n12235) );
  AOI211_X1 U14038 ( .C1(n12565), .C2(n12237), .A(n12236), .B(n12235), .ZN(
        n12240) );
  NAND2_X1 U14039 ( .A1(n13351), .A2(n12238), .ZN(n12239) );
  OAI211_X1 U14040 ( .C1(n12241), .C2(n13314), .A(n12240), .B(n12239), .ZN(
        P3_U3171) );
  XOR2_X1 U14041 ( .A(n13527), .B(n12242), .Z(n15965) );
  INV_X1 U14042 ( .A(n12243), .ZN(n12244) );
  AOI21_X1 U14043 ( .B1(n13527), .B2(n12245), .A(n12244), .ZN(n12249) );
  AOI22_X1 U14044 ( .A1(n13997), .A2(n13580), .B1(n13578), .B2(n13996), .ZN(
        n12248) );
  INV_X1 U14045 ( .A(n15965), .ZN(n12246) );
  NAND2_X1 U14046 ( .A1(n12246), .A2(n13994), .ZN(n12247) );
  OAI211_X1 U14047 ( .C1(n12249), .C2(n14002), .A(n12248), .B(n12247), .ZN(
        n15966) );
  NAND2_X1 U14048 ( .A1(n15966), .A2(n13966), .ZN(n12253) );
  OAI22_X1 U14049 ( .A1(n14006), .A2(n15964), .B1(n12250), .B2(n13983), .ZN(
        n12251) );
  AOI21_X1 U14050 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n13963), .A(n12251), .ZN(
        n12252) );
  OAI211_X1 U14051 ( .C1(n15965), .C2(n12254), .A(n12253), .B(n12252), .ZN(
        P3_U3225) );
  INV_X1 U14052 ( .A(n12588), .ZN(n12257) );
  OAI222_X1 U14053 ( .A1(n15512), .A2(n12589), .B1(n15510), .B2(n12257), .C1(
        n12255), .C2(P1_U3086), .ZN(P1_U3330) );
  OAI222_X1 U14054 ( .A1(n14871), .A2(n8113), .B1(n14869), .B2(n12257), .C1(
        P2_U3088), .C2(n12256), .ZN(P2_U3302) );
  INV_X1 U14055 ( .A(n12258), .ZN(n12259) );
  AOI21_X1 U14056 ( .B1(n12261), .B2(n12260), .A(n12259), .ZN(n12267) );
  INV_X1 U14057 ( .A(n15065), .ZN(n12512) );
  AOI22_X1 U14058 ( .A1(n14987), .A2(n12262), .B1(n16087), .B2(n15067), .ZN(
        n12264) );
  OAI211_X1 U14059 ( .C1(n12512), .C2(n15036), .A(n12264), .B(n12263), .ZN(
        n12265) );
  AOI21_X1 U14060 ( .B1(n12744), .B2(n15040), .A(n12265), .ZN(n12266) );
  OAI21_X1 U14061 ( .B1(n12267), .B2(n15042), .A(n12266), .ZN(P1_U3236) );
  XNOR2_X1 U14062 ( .A(n16111), .B(n14229), .ZN(n12534) );
  NAND2_X1 U14063 ( .A1(n14363), .A2(n14633), .ZN(n12532) );
  XNOR2_X1 U14064 ( .A(n12534), .B(n12532), .ZN(n12275) );
  NOR2_X1 U14065 ( .A1(n14351), .A2(n12269), .ZN(n12273) );
  OAI22_X1 U14066 ( .A1(n14341), .A2(n12271), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12270), .ZN(n12272) );
  AOI211_X1 U14067 ( .C1(n16111), .C2(n14358), .A(n12273), .B(n12272), .ZN(
        n12279) );
  AOI22_X1 U14068 ( .A1(n12274), .A2(n14311), .B1(n14330), .B2(n14364), .ZN(
        n12276) );
  OR3_X1 U14069 ( .A1(n12277), .A2(n12276), .A3(n12275), .ZN(n12278) );
  OAI211_X1 U14070 ( .C1(n12533), .C2(n14353), .A(n12279), .B(n12278), .ZN(
        P2_U3187) );
  INV_X1 U14071 ( .A(n14330), .ZN(n14296) );
  INV_X1 U14072 ( .A(n12280), .ZN(n12281) );
  OAI33_X1 U14073 ( .A1(n12284), .A2(n12283), .A3(n14353), .B1(n14296), .B2(
        n12282), .B3(n12281), .ZN(n12287) );
  INV_X1 U14074 ( .A(n12285), .ZN(n12286) );
  NAND2_X1 U14075 ( .A1(n12287), .A2(n12286), .ZN(n12293) );
  OAI22_X1 U14076 ( .A1(n14341), .A2(n12289), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12288), .ZN(n12290) );
  AOI21_X1 U14077 ( .B1(n12291), .B2(n14339), .A(n12290), .ZN(n12292) );
  OAI211_X1 U14078 ( .C1(n12294), .C2(n14309), .A(n12293), .B(n12292), .ZN(
        n12295) );
  AOI21_X1 U14079 ( .B1(n14311), .B2(n12296), .A(n12295), .ZN(n12297) );
  INV_X1 U14080 ( .A(n12297), .ZN(P2_U3196) );
  INV_X1 U14081 ( .A(n15066), .ZN(n12299) );
  NAND2_X1 U14082 ( .A1(n12747), .A2(n15065), .ZN(n12300) );
  NAND2_X1 U14083 ( .A1(n12385), .A2(n12300), .ZN(n12866) );
  XNOR2_X1 U14084 ( .A(n12375), .B(n12866), .ZN(n12308) );
  NAND2_X1 U14085 ( .A1(n12744), .A2(n15066), .ZN(n12301) );
  INV_X1 U14086 ( .A(n12866), .ZN(n12303) );
  NAND2_X1 U14087 ( .A1(n12304), .A2(n12866), .ZN(n12305) );
  NAND2_X1 U14088 ( .A1(n12386), .A2(n12305), .ZN(n16067) );
  NAND2_X1 U14089 ( .A1(n16067), .A2(n16026), .ZN(n12307) );
  AOI22_X1 U14090 ( .A1(n15376), .A2(n16086), .B1(n15066), .B2(n16030), .ZN(
        n12306) );
  OAI211_X1 U14091 ( .C1(n16136), .C2(n12308), .A(n12307), .B(n12306), .ZN(
        n16072) );
  INV_X1 U14092 ( .A(n16072), .ZN(n12316) );
  NOR2_X1 U14093 ( .A1(n12747), .A2(n12744), .ZN(n12309) );
  NAND2_X1 U14094 ( .A1(n12310), .A2(n12309), .ZN(n12381) );
  INV_X1 U14095 ( .A(n12381), .ZN(n12382) );
  INV_X1 U14096 ( .A(n12744), .ZN(n16049) );
  INV_X1 U14097 ( .A(n12747), .ZN(n16070) );
  AOI21_X1 U14098 ( .B1(n12310), .B2(n16049), .A(n16070), .ZN(n12311) );
  OR3_X1 U14099 ( .A1(n12382), .A2(n12311), .A3(n15974), .ZN(n16068) );
  AOI22_X1 U14100 ( .A1(n16001), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n12549), 
        .B2(n15990), .ZN(n12313) );
  NAND2_X1 U14101 ( .A1(n12747), .A2(n15991), .ZN(n12312) );
  OAI211_X1 U14102 ( .C1(n16068), .C2(n15993), .A(n12313), .B(n12312), .ZN(
        n12314) );
  AOI21_X1 U14103 ( .B1(n16067), .B2(n15996), .A(n12314), .ZN(n12315) );
  OAI21_X1 U14104 ( .B1(n12316), .B2(n16001), .A(n12315), .ZN(P1_U3281) );
  INV_X1 U14105 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14720) );
  NOR2_X1 U14106 ( .A1(n14440), .A2(n14720), .ZN(n12317) );
  AOI21_X1 U14107 ( .B1(n14720), .B2(n14440), .A(n12317), .ZN(n14444) );
  NAND2_X1 U14108 ( .A1(n15595), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n12325) );
  INV_X1 U14109 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12320) );
  INV_X1 U14110 ( .A(n12325), .ZN(n12318) );
  AOI21_X1 U14111 ( .B1(n12320), .B2(n12319), .A(n12318), .ZN(n15598) );
  NAND2_X1 U14112 ( .A1(n12322), .A2(n12321), .ZN(n12324) );
  NAND2_X1 U14113 ( .A1(n12324), .A2(n12323), .ZN(n15597) );
  NAND2_X1 U14114 ( .A1(n15598), .A2(n15597), .ZN(n15596) );
  NAND2_X1 U14115 ( .A1(n12325), .A2(n15596), .ZN(n14445) );
  NAND2_X1 U14116 ( .A1(n14444), .A2(n14445), .ZN(n14443) );
  INV_X1 U14117 ( .A(n14443), .ZN(n12326) );
  AOI21_X1 U14118 ( .B1(n12337), .B2(P2_REG2_REG_17__SCAN_IN), .A(n12326), 
        .ZN(n12408) );
  XNOR2_X1 U14119 ( .A(n12408), .B(n12409), .ZN(n12327) );
  NOR2_X1 U14120 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n12327), .ZN(n12407) );
  AOI21_X1 U14121 ( .B1(n12327), .B2(P2_REG2_REG_18__SCAN_IN), .A(n12407), 
        .ZN(n12345) );
  NOR2_X1 U14122 ( .A1(n12329), .A2(n12328), .ZN(n12331) );
  NOR2_X1 U14123 ( .A1(n12331), .A2(n12330), .ZN(n15592) );
  INV_X1 U14124 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n12333) );
  NAND2_X1 U14125 ( .A1(n15595), .A2(n12333), .ZN(n12332) );
  OAI21_X1 U14126 ( .B1(n15595), .B2(n12333), .A(n12332), .ZN(n12334) );
  INV_X1 U14127 ( .A(n12334), .ZN(n15591) );
  NOR2_X1 U14128 ( .A1(n15592), .A2(n15591), .ZN(n15590) );
  AOI21_X1 U14129 ( .B1(n15595), .B2(P2_REG1_REG_16__SCAN_IN), .A(n15590), 
        .ZN(n14437) );
  NOR2_X1 U14130 ( .A1(n12337), .A2(n12335), .ZN(n12336) );
  AOI21_X1 U14131 ( .B1(n12337), .B2(n12335), .A(n12336), .ZN(n14438) );
  NOR2_X1 U14132 ( .A1(n14437), .A2(n14438), .ZN(n14436) );
  AOI21_X1 U14133 ( .B1(n12337), .B2(P2_REG1_REG_17__SCAN_IN), .A(n14436), 
        .ZN(n12338) );
  NOR2_X1 U14134 ( .A1(n12338), .A2(n12409), .ZN(n12402) );
  AOI21_X1 U14135 ( .B1(n12338), .B2(n12409), .A(n12402), .ZN(n12339) );
  NAND2_X1 U14136 ( .A1(n12339), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n12404) );
  OAI211_X1 U14137 ( .C1(n12339), .C2(P2_REG1_REG_18__SCAN_IN), .A(n12404), 
        .B(n15602), .ZN(n12344) );
  NOR2_X1 U14138 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12340), .ZN(n12342) );
  NOR2_X1 U14139 ( .A1(n15543), .A2(n12409), .ZN(n12341) );
  AOI211_X1 U14140 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n15619), .A(n12342), 
        .B(n12341), .ZN(n12343) );
  OAI211_X1 U14141 ( .C1(n12345), .C2(n15630), .A(n12344), .B(n12343), .ZN(
        P2_U3232) );
  INV_X1 U14142 ( .A(n12346), .ZN(n12347) );
  OAI222_X1 U14143 ( .A1(P3_U3151), .A2(n12349), .B1(n14155), .B2(n12348), 
        .C1(n14158), .C2(n12347), .ZN(P3_U3270) );
  INV_X1 U14144 ( .A(n14363), .ZN(n12352) );
  NAND2_X1 U14145 ( .A1(n16111), .A2(n12352), .ZN(n12350) );
  NAND2_X1 U14146 ( .A1(n12351), .A2(n12350), .ZN(n12354) );
  OR2_X1 U14147 ( .A1(n16111), .A2(n12352), .ZN(n12353) );
  XOR2_X1 U14148 ( .A(n12424), .B(n12357), .Z(n12355) );
  AOI22_X1 U14149 ( .A1(n14463), .A2(n14338), .B1(n14525), .B2(n14363), .ZN(
        n14346) );
  OAI21_X1 U14150 ( .B1(n12355), .B2(n14679), .A(n14346), .ZN(n12458) );
  INV_X1 U14151 ( .A(n12458), .ZN(n12365) );
  NAND2_X1 U14152 ( .A1(n16111), .A2(n14363), .ZN(n12356) );
  OAI21_X1 U14153 ( .B1(n12358), .B2(n12357), .A(n12420), .ZN(n12465) );
  INV_X1 U14154 ( .A(n14359), .ZN(n12457) );
  OAI211_X1 U14155 ( .C1(n12457), .C2(n12359), .A(n14716), .B(n7360), .ZN(
        n12456) );
  NAND2_X1 U14156 ( .A1(n14697), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n12360) );
  OAI21_X1 U14157 ( .B1(n14718), .B2(n14350), .A(n12360), .ZN(n12361) );
  AOI21_X1 U14158 ( .B1(n14359), .B2(n14722), .A(n12361), .ZN(n12362) );
  OAI21_X1 U14159 ( .B1(n12456), .B2(n14725), .A(n12362), .ZN(n12363) );
  AOI21_X1 U14160 ( .B1(n12465), .B2(n14642), .A(n12363), .ZN(n12364) );
  OAI21_X1 U14161 ( .B1(n12365), .B2(n14697), .A(n12364), .ZN(P2_U3250) );
  NAND2_X1 U14162 ( .A1(n13577), .A2(n12394), .ZN(n12366) );
  NAND2_X1 U14163 ( .A1(n12367), .A2(n12366), .ZN(n12520) );
  INV_X1 U14164 ( .A(n13532), .ZN(n13441) );
  XNOR2_X1 U14165 ( .A(n12520), .B(n13441), .ZN(n12368) );
  OAI222_X1 U14166 ( .A1(n13944), .A2(n13309), .B1(n13946), .B2(n12474), .C1(
        n12368), .C2(n14002), .ZN(n12501) );
  INV_X1 U14167 ( .A(n12501), .ZN(n12374) );
  OAI21_X1 U14168 ( .B1(n12370), .B2(n13532), .A(n12516), .ZN(n12502) );
  AOI22_X1 U14169 ( .A1(n13963), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n14004), 
        .B2(n12477), .ZN(n12371) );
  OAI21_X1 U14170 ( .B1(n12507), .B2(n14006), .A(n12371), .ZN(n12372) );
  AOI21_X1 U14171 ( .B1(n12502), .B2(n13981), .A(n12372), .ZN(n12373) );
  OAI21_X1 U14172 ( .B1(n12374), .B2(n13963), .A(n12373), .ZN(P3_U3222) );
  OR2_X1 U14173 ( .A1(n12747), .A2(n12512), .ZN(n12376) );
  XNOR2_X1 U14174 ( .A(n12751), .B(n16086), .ZN(n12869) );
  XNOR2_X1 U14175 ( .A(n12437), .B(n12444), .ZN(n12378) );
  AOI222_X1 U14176 ( .A1(n16119), .A2(n12378), .B1(n15065), .B2(n16030), .C1(
        n15374), .C2(n15376), .ZN(n16077) );
  INV_X1 U14177 ( .A(n12379), .ZN(n12511) );
  OAI22_X1 U14178 ( .A1(n7218), .A2(n12380), .B1(n12511), .B2(n15377), .ZN(
        n12384) );
  INV_X1 U14179 ( .A(n12751), .ZN(n16078) );
  OAI211_X1 U14180 ( .C1(n12382), .C2(n16078), .A(n15445), .B(n12441), .ZN(
        n16076) );
  NOR2_X1 U14181 ( .A1(n16076), .A2(n15993), .ZN(n12383) );
  AOI211_X1 U14182 ( .C1(n15991), .C2(n12751), .A(n12384), .B(n12383), .ZN(
        n12388) );
  XNOR2_X1 U14183 ( .A(n12445), .B(n12444), .ZN(n16080) );
  NAND2_X1 U14184 ( .A1(n16080), .A2(n15355), .ZN(n12387) );
  OAI211_X1 U14185 ( .C1(n16077), .C2(n16001), .A(n12388), .B(n12387), .ZN(
        P1_U3280) );
  OAI211_X1 U14186 ( .C1(n7369), .C2(n12390), .A(n12389), .B(n13343), .ZN(
        n12396) );
  INV_X1 U14187 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n13166) );
  NOR2_X1 U14188 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13166), .ZN(n15847) );
  AOI21_X1 U14189 ( .B1(n13998), .B2(n13346), .A(n15847), .ZN(n12391) );
  OAI21_X1 U14190 ( .B1(n12392), .B2(n13349), .A(n12391), .ZN(n12393) );
  AOI21_X1 U14191 ( .B1(n12394), .B2(n12565), .A(n12393), .ZN(n12395) );
  OAI211_X1 U14192 ( .C1(n12398), .C2(n12397), .A(n12396), .B(n12395), .ZN(
        P3_U3157) );
  INV_X1 U14193 ( .A(n12399), .ZN(n12400) );
  OAI222_X1 U14194 ( .A1(n12401), .A2(P3_U3151), .B1(n14158), .B2(n12400), 
        .C1(n13103), .C2(n14155), .ZN(P3_U3269) );
  INV_X1 U14195 ( .A(n12402), .ZN(n12403) );
  NAND2_X1 U14196 ( .A1(n12404), .A2(n12403), .ZN(n12406) );
  INV_X1 U14197 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14797) );
  XNOR2_X1 U14198 ( .A(n12410), .B(n14797), .ZN(n12405) );
  XNOR2_X1 U14199 ( .A(n12406), .B(n12405), .ZN(n12418) );
  AOI21_X1 U14200 ( .B1(n12409), .B2(n12408), .A(n12407), .ZN(n12412) );
  MUX2_X1 U14201 ( .A(n14684), .B(P2_REG2_REG_19__SCAN_IN), .S(n12410), .Z(
        n12411) );
  XNOR2_X1 U14202 ( .A(n12412), .B(n12411), .ZN(n12416) );
  NAND2_X1 U14203 ( .A1(n15619), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n12413) );
  NAND2_X1 U14204 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14222)
         );
  OAI211_X1 U14205 ( .C1(n12414), .C2(n15543), .A(n12413), .B(n14222), .ZN(
        n12415) );
  AOI21_X1 U14206 ( .B1(n15611), .B2(n12416), .A(n12415), .ZN(n12417) );
  OAI21_X1 U14207 ( .B1(n12418), .B2(n15622), .A(n12417), .ZN(P2_U3233) );
  OR2_X1 U14208 ( .A1(n14359), .A2(n14362), .ZN(n12419) );
  OAI21_X1 U14209 ( .B1(n12422), .B2(n12427), .A(n14465), .ZN(n14850) );
  NOR2_X1 U14210 ( .A1(n14359), .A2(n12425), .ZN(n12423) );
  NAND2_X1 U14211 ( .A1(n14359), .A2(n12425), .ZN(n12426) );
  NAND2_X1 U14212 ( .A1(n12428), .A2(n12427), .ZN(n12429) );
  NAND3_X1 U14213 ( .A1(n14708), .A2(n14710), .A3(n12429), .ZN(n12431) );
  AND2_X1 U14214 ( .A1(n14362), .A2(n14525), .ZN(n12430) );
  AOI21_X1 U14215 ( .B1(n14466), .B2(n14338), .A(n12430), .ZN(n12540) );
  NAND2_X1 U14216 ( .A1(n12431), .A2(n12540), .ZN(n14812) );
  AOI21_X1 U14217 ( .B1(n7360), .B2(n14808), .A(n14633), .ZN(n12432) );
  NAND2_X1 U14218 ( .A1(n12432), .A2(n14714), .ZN(n14809) );
  OAI22_X1 U14219 ( .A1(n12155), .A2(n12320), .B1(n12539), .B2(n14718), .ZN(
        n12433) );
  AOI21_X1 U14220 ( .B1(n14808), .B2(n14722), .A(n12433), .ZN(n12434) );
  OAI21_X1 U14221 ( .B1(n14809), .B2(n14725), .A(n12434), .ZN(n12435) );
  AOI21_X1 U14222 ( .B1(n14812), .B2(n12155), .A(n12435), .ZN(n12436) );
  OAI21_X1 U14223 ( .B1(n14850), .B2(n14728), .A(n12436), .ZN(P2_U3249) );
  INV_X1 U14224 ( .A(n16086), .ZN(n12552) );
  OR2_X1 U14225 ( .A1(n12751), .A2(n12552), .ZN(n12438) );
  XOR2_X1 U14226 ( .A(n12602), .B(n12871), .Z(n16104) );
  INV_X1 U14227 ( .A(n16104), .ZN(n12450) );
  AOI22_X1 U14228 ( .A1(n15376), .A2(n16088), .B1(n16086), .B2(n16030), .ZN(
        n16099) );
  AOI22_X1 U14229 ( .A1(n16001), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n12439), 
        .B2(n15990), .ZN(n12440) );
  OAI21_X1 U14230 ( .B1(n16099), .B2(n16001), .A(n12440), .ZN(n12443) );
  OAI211_X1 U14231 ( .C1(n7737), .C2(n7738), .A(n15380), .B(n15445), .ZN(
        n16100) );
  NOR2_X1 U14232 ( .A1(n16100), .A2(n15993), .ZN(n12442) );
  AOI211_X1 U14233 ( .C1(n15991), .C2(n12755), .A(n12443), .B(n12442), .ZN(
        n12449) );
  OR2_X1 U14234 ( .A1(n12751), .A2(n16086), .ZN(n12446) );
  NAND2_X1 U14235 ( .A1(n12447), .A2(n12871), .ZN(n16101) );
  NAND3_X1 U14236 ( .A1(n7359), .A2(n16101), .A3(n15355), .ZN(n12448) );
  OAI211_X1 U14237 ( .C1(n12450), .C2(n15371), .A(n12449), .B(n12448), .ZN(
        P1_U3279) );
  INV_X1 U14238 ( .A(n12451), .ZN(n12453) );
  INV_X1 U14239 ( .A(n12616), .ZN(n12454) );
  OAI222_X1 U14240 ( .A1(P2_U3088), .A2(n12453), .B1(n14869), .B2(n12454), 
        .C1(n12452), .C2(n14871), .ZN(P2_U3301) );
  OAI222_X1 U14241 ( .A1(n12455), .A2(n7201), .B1(n15510), .B2(n12454), .C1(
        n12617), .C2(n15512), .ZN(P1_U3329) );
  OAI21_X1 U14242 ( .B1(n12457), .B2(n16149), .A(n12456), .ZN(n12459) );
  AOI211_X1 U14243 ( .C1(n14803), .C2(n12465), .A(n12459), .B(n12458), .ZN(
        n12467) );
  INV_X1 U14244 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n12460) );
  NOR2_X1 U14245 ( .A1(n16117), .A2(n12460), .ZN(n12461) );
  AOI21_X1 U14246 ( .B1(n12465), .B2(n12462), .A(n12461), .ZN(n12463) );
  OAI21_X1 U14247 ( .B1(n12467), .B2(n16157), .A(n12463), .ZN(P2_U3475) );
  AOI22_X1 U14248 ( .A1(n12465), .A2(n12464), .B1(n16155), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n12466) );
  OAI21_X1 U14249 ( .B1(n12467), .B2(n16155), .A(n12466), .ZN(P2_U3514) );
  OAI222_X1 U14250 ( .A1(n14158), .A2(n12468), .B1(n14155), .B2(n13101), .C1(
        P3_U3151), .C2(n10630), .ZN(P3_U3268) );
  OAI211_X1 U14251 ( .C1(n12471), .C2(n12470), .A(n12469), .B(n13343), .ZN(
        n12479) );
  NOR2_X1 U14252 ( .A1(n13354), .A2(n12507), .ZN(n12476) );
  NAND2_X1 U14253 ( .A1(n13346), .A2(n13576), .ZN(n12473) );
  AND2_X1 U14254 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n15870) );
  INV_X1 U14255 ( .A(n15870), .ZN(n12472) );
  OAI211_X1 U14256 ( .C1(n13349), .C2(n12474), .A(n12473), .B(n12472), .ZN(
        n12475) );
  AOI211_X1 U14257 ( .C1(n12477), .C2(n13351), .A(n12476), .B(n12475), .ZN(
        n12478) );
  NAND2_X1 U14258 ( .A1(n12479), .A2(n12478), .ZN(P3_U3176) );
  INV_X1 U14259 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n16142) );
  NOR2_X1 U14260 ( .A1(n15106), .A2(n16142), .ZN(n12480) );
  AOI21_X1 U14261 ( .B1(n15106), .B2(n16142), .A(n12480), .ZN(n12486) );
  OAI21_X1 U14262 ( .B1(n12482), .B2(n16105), .A(n12481), .ZN(n12484) );
  XNOR2_X1 U14263 ( .A(n12484), .B(n15648), .ZN(n15644) );
  INV_X1 U14264 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n16128) );
  NAND2_X1 U14265 ( .A1(n15644), .A2(n16128), .ZN(n15643) );
  OAI21_X1 U14266 ( .B1(n12484), .B2(n12483), .A(n15643), .ZN(n12485) );
  NOR2_X1 U14267 ( .A1(n12485), .A2(n12486), .ZN(n15105) );
  AOI211_X1 U14268 ( .C1(n12486), .C2(n12485), .A(n15145), .B(n15105), .ZN(
        n12500) );
  INV_X1 U14269 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12491) );
  MUX2_X1 U14270 ( .A(n12491), .B(P1_REG2_REG_16__SCAN_IN), .S(n15106), .Z(
        n12496) );
  AOI21_X1 U14271 ( .B1(n12488), .B2(P1_REG2_REG_14__SCAN_IN), .A(n12487), 
        .ZN(n12489) );
  NAND2_X1 U14272 ( .A1(n12489), .A2(n15648), .ZN(n12493) );
  XNOR2_X1 U14273 ( .A(n12489), .B(n15648), .ZN(n15646) );
  NOR2_X1 U14274 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15646), .ZN(n15645) );
  INV_X1 U14275 ( .A(n15645), .ZN(n12490) );
  NAND2_X1 U14276 ( .A1(n12493), .A2(n12490), .ZN(n12495) );
  AOI21_X1 U14277 ( .B1(n15110), .B2(n12491), .A(n15645), .ZN(n12492) );
  OAI211_X1 U14278 ( .C1(n15110), .C2(n12491), .A(n12493), .B(n12492), .ZN(
        n15109) );
  INV_X1 U14279 ( .A(n15109), .ZN(n12494) );
  AOI211_X1 U14280 ( .C1(n12496), .C2(n12495), .A(n15649), .B(n12494), .ZN(
        n12499) );
  NAND2_X1 U14281 ( .A1(n7201), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14988) );
  NAND2_X1 U14282 ( .A1(n15639), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n12497) );
  OAI211_X1 U14283 ( .C1(n15647), .C2(n15110), .A(n14988), .B(n12497), .ZN(
        n12498) );
  OR3_X1 U14284 ( .A1(n12500), .A2(n12499), .A3(n12498), .ZN(P1_U3259) );
  AOI21_X1 U14285 ( .B1(n14080), .B2(n12502), .A(n12501), .ZN(n12504) );
  MUX2_X1 U14286 ( .A(n15858), .B(n12504), .S(n16061), .Z(n12503) );
  OAI21_X1 U14287 ( .B1(n14083), .B2(n12507), .A(n12503), .ZN(P3_U3470) );
  INV_X1 U14288 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n12505) );
  MUX2_X1 U14289 ( .A(n12505), .B(n12504), .S(n16065), .Z(n12506) );
  OAI21_X1 U14290 ( .B1(n14142), .B2(n12507), .A(n12506), .ZN(P3_U3423) );
  OAI211_X1 U14291 ( .C1(n12510), .C2(n12509), .A(n12508), .B(n16093), .ZN(
        n12515) );
  AND2_X1 U14292 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(n7201), .ZN(n15098) );
  OAI22_X1 U14293 ( .A1(n12512), .A2(n15049), .B1(n16098), .B2(n12511), .ZN(
        n12513) );
  AOI211_X1 U14294 ( .C1(n16089), .C2(n15374), .A(n15098), .B(n12513), .ZN(
        n12514) );
  OAI211_X1 U14295 ( .C1(n16078), .C2(n16091), .A(n12515), .B(n12514), .ZN(
        P1_U3234) );
  NAND2_X1 U14296 ( .A1(n13309), .A2(n12564), .ZN(n13448) );
  NAND2_X1 U14297 ( .A1(n13576), .A2(n16055), .ZN(n13445) );
  NAND2_X1 U14298 ( .A1(n13993), .A2(n13992), .ZN(n13991) );
  NAND2_X1 U14299 ( .A1(n14141), .A2(n13995), .ZN(n13449) );
  OAI21_X1 U14300 ( .B1(n12517), .B2(n13447), .A(n12970), .ZN(n14079) );
  INV_X1 U14301 ( .A(n14079), .ZN(n12531) );
  NAND2_X1 U14302 ( .A1(n13576), .A2(n12564), .ZN(n12521) );
  NAND2_X1 U14303 ( .A1(n13990), .A2(n12521), .ZN(n12523) );
  NAND2_X1 U14304 ( .A1(n13309), .A2(n16055), .ZN(n12522) );
  NAND2_X1 U14305 ( .A1(n12523), .A2(n12522), .ZN(n12524) );
  INV_X1 U14306 ( .A(n12524), .ZN(n12525) );
  INV_X1 U14307 ( .A(n13447), .ZN(n13535) );
  OAI211_X1 U14308 ( .C1(n12525), .C2(n13535), .A(n13970), .B(n12938), .ZN(
        n12527) );
  AOI22_X1 U14309 ( .A1(n13959), .A2(n13996), .B1(n13997), .B2(n13576), .ZN(
        n12526) );
  NAND2_X1 U14310 ( .A1(n12527), .A2(n12526), .ZN(n14078) );
  AOI22_X1 U14311 ( .A1(n13963), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n14004), 
        .B2(n13312), .ZN(n12528) );
  OAI21_X1 U14312 ( .B1(n14141), .B2(n14006), .A(n12528), .ZN(n12529) );
  AOI21_X1 U14313 ( .B1(n14078), .B2(n13966), .A(n12529), .ZN(n12530) );
  OAI21_X1 U14314 ( .B1(n12531), .B2(n13968), .A(n12530), .ZN(P3_U3220) );
  INV_X1 U14315 ( .A(n12532), .ZN(n12535) );
  XNOR2_X1 U14316 ( .A(n14359), .B(n14229), .ZN(n12543) );
  AND2_X1 U14317 ( .A1(n14362), .A2(n14633), .ZN(n12536) );
  NAND2_X1 U14318 ( .A1(n12543), .A2(n12536), .ZN(n12537) );
  OAI21_X1 U14319 ( .B1(n12543), .B2(n12536), .A(n12537), .ZN(n14354) );
  INV_X1 U14320 ( .A(n12537), .ZN(n12538) );
  XNOR2_X1 U14321 ( .A(n14808), .B(n14188), .ZN(n14281) );
  NAND2_X1 U14322 ( .A1(n14463), .A2(n14633), .ZN(n14159) );
  XNOR2_X1 U14323 ( .A(n14281), .B(n14159), .ZN(n12545) );
  INV_X1 U14324 ( .A(n14164), .ZN(n14284) );
  NOR2_X1 U14325 ( .A1(n14351), .A2(n12539), .ZN(n12542) );
  OAI22_X1 U14326 ( .A1(n14341), .A2(n12540), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15589), .ZN(n12541) );
  AOI211_X1 U14327 ( .C1(n14808), .C2(n14358), .A(n12542), .B(n12541), .ZN(
        n12548) );
  NAND3_X1 U14328 ( .A1(n12543), .A2(n14330), .A3(n14362), .ZN(n12544) );
  OAI21_X1 U14329 ( .B1(n7895), .B2(n14353), .A(n12544), .ZN(n12546) );
  NAND2_X1 U14330 ( .A1(n12546), .A2(n12545), .ZN(n12547) );
  OAI211_X1 U14331 ( .C1(n14284), .C2(n14353), .A(n12548), .B(n12547), .ZN(
        P2_U3198) );
  AOI22_X1 U14332 ( .A1(n14987), .A2(n12549), .B1(n16087), .B2(n15066), .ZN(
        n12551) );
  OAI211_X1 U14333 ( .C1(n12552), .C2(n15036), .A(n12551), .B(n12550), .ZN(
        n12558) );
  INV_X1 U14334 ( .A(n12553), .ZN(n12554) );
  AOI211_X1 U14335 ( .C1(n12556), .C2(n12555), .A(n15042), .B(n12554), .ZN(
        n12557) );
  AOI211_X1 U14336 ( .C1(n15040), .C2(n12747), .A(n12558), .B(n12557), .ZN(
        n12559) );
  INV_X1 U14337 ( .A(n12559), .ZN(P1_U3224) );
  XNOR2_X1 U14338 ( .A(n12560), .B(n13576), .ZN(n12561) );
  XNOR2_X1 U14339 ( .A(n12562), .B(n12561), .ZN(n12571) );
  AOI21_X1 U14340 ( .B1(n13346), .B2(n13995), .A(n12563), .ZN(n12569) );
  NAND2_X1 U14341 ( .A1(n12565), .A2(n12564), .ZN(n12568) );
  NAND2_X1 U14342 ( .A1(n13998), .A2(n13318), .ZN(n12567) );
  NAND2_X1 U14343 ( .A1(n13351), .A2(n14003), .ZN(n12566) );
  NAND4_X1 U14344 ( .A1(n12569), .A2(n12568), .A3(n12567), .A4(n12566), .ZN(
        n12570) );
  AOI21_X1 U14345 ( .B1(n12571), .B2(n13343), .A(n12570), .ZN(n12572) );
  INV_X1 U14346 ( .A(n12572), .ZN(P3_U3164) );
  MUX2_X1 U14347 ( .A(n12573), .B(P3_REG2_REG_0__SCAN_IN), .S(n13963), .Z(
        n12577) );
  OAI22_X1 U14348 ( .A1(n14006), .A2(n12575), .B1(n13983), .B2(n12574), .ZN(
        n12576) );
  OR2_X1 U14349 ( .A1(n12577), .A2(n12576), .ZN(P3_U3233) );
  INV_X1 U14350 ( .A(n12825), .ZN(n15506) );
  OAI222_X1 U14351 ( .A1(n14871), .A2(n12579), .B1(n14869), .B2(n15506), .C1(
        n12578), .C2(P2_U3088), .ZN(P2_U3298) );
  NAND2_X1 U14352 ( .A1(n12833), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n12587) );
  NAND2_X1 U14353 ( .A1(n12829), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n12586) );
  INV_X1 U14354 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n12581) );
  NAND2_X1 U14355 ( .A1(n12580), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n12582) );
  NAND2_X1 U14356 ( .A1(n12581), .A2(n12582), .ZN(n12583) );
  NAND2_X1 U14357 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n12592), .ZN(n12621) );
  AND2_X1 U14358 ( .A1(n12583), .A2(n12621), .ZN(n15212) );
  NAND2_X1 U14359 ( .A1(n7212), .A2(n15212), .ZN(n12585) );
  NAND2_X1 U14360 ( .A1(n12834), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n12584) );
  NAND4_X1 U14361 ( .A1(n12587), .A2(n12586), .A3(n12585), .A4(n12584), .ZN(
        n15058) );
  NAND2_X1 U14362 ( .A1(n12588), .A2(n7232), .ZN(n12591) );
  OR2_X1 U14363 ( .A1(n9902), .A2(n12589), .ZN(n12590) );
  NAND2_X1 U14364 ( .A1(n12834), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n12597) );
  NAND2_X1 U14365 ( .A1(n12833), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n12596) );
  INV_X1 U14366 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n15007) );
  AOI21_X1 U14367 ( .B1(n15007), .B2(n12593), .A(n12592), .ZN(n15229) );
  NAND2_X1 U14368 ( .A1(n7213), .A2(n15229), .ZN(n12595) );
  NAND2_X1 U14369 ( .A1(n12829), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n12594) );
  NAND4_X1 U14370 ( .A1(n12597), .A2(n12596), .A3(n12595), .A4(n12594), .ZN(
        n15059) );
  INV_X1 U14371 ( .A(n15059), .ZN(n14929) );
  NAND2_X1 U14372 ( .A1(n12598), .A2(n7232), .ZN(n12601) );
  OR2_X1 U14373 ( .A1(n9902), .A2(n12599), .ZN(n12600) );
  INV_X1 U14374 ( .A(n15374), .ZN(n15050) );
  NAND2_X1 U14375 ( .A1(n12755), .A2(n15050), .ZN(n12603) );
  XNOR2_X1 U14376 ( .A(n15386), .B(n16088), .ZN(n12872) );
  OR2_X1 U14377 ( .A1(n15386), .A2(n15358), .ZN(n12605) );
  XNOR2_X1 U14378 ( .A(n16133), .B(n15375), .ZN(n15351) );
  INV_X1 U14379 ( .A(n15375), .ZN(n15340) );
  NAND2_X1 U14380 ( .A1(n16133), .A2(n15340), .ZN(n12606) );
  NAND2_X1 U14381 ( .A1(n12607), .A2(n12606), .ZN(n15335) );
  XNOR2_X1 U14382 ( .A(n15474), .B(n15064), .ZN(n15338) );
  XNOR2_X1 U14383 ( .A(n15466), .B(n15063), .ZN(n15322) );
  INV_X1 U14384 ( .A(n15322), .ZN(n15319) );
  NAND2_X1 U14385 ( .A1(n15323), .A2(n15322), .ZN(n15321) );
  INV_X1 U14386 ( .A(n15063), .ZN(n15341) );
  OR2_X1 U14387 ( .A1(n15466), .A2(n15341), .ZN(n12608) );
  AND2_X2 U14388 ( .A1(n15321), .A2(n12608), .ZN(n15304) );
  XNOR2_X1 U14389 ( .A(n15460), .B(n15062), .ZN(n15303) );
  INV_X1 U14390 ( .A(n15062), .ZN(n12609) );
  NAND2_X1 U14391 ( .A1(n15460), .A2(n12609), .ZN(n12610) );
  XNOR2_X1 U14392 ( .A(n15299), .B(n15061), .ZN(n15290) );
  INV_X1 U14393 ( .A(n15290), .ZN(n15282) );
  XNOR2_X1 U14394 ( .A(n15444), .B(n12780), .ZN(n15276) );
  XNOR2_X1 U14395 ( .A(n15439), .B(n14969), .ZN(n15254) );
  NAND2_X1 U14396 ( .A1(n12611), .A2(n7232), .ZN(n12614) );
  OR2_X1 U14397 ( .A1(n9902), .A2(n12612), .ZN(n12613) );
  XNOR2_X1 U14398 ( .A(n15433), .B(n12615), .ZN(n12877) );
  XNOR2_X1 U14399 ( .A(n15429), .B(n14929), .ZN(n15220) );
  INV_X1 U14400 ( .A(n15220), .ZN(n15223) );
  XNOR2_X1 U14401 ( .A(n15425), .B(n15191), .ZN(n15203) );
  NAND2_X1 U14402 ( .A1(n12616), .A2(n7232), .ZN(n12619) );
  OR2_X1 U14403 ( .A1(n9902), .A2(n12617), .ZN(n12618) );
  NAND2_X1 U14404 ( .A1(n12834), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n12626) );
  NAND2_X1 U14405 ( .A1(n12833), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n12625) );
  INV_X1 U14406 ( .A(n12621), .ZN(n12620) );
  INV_X1 U14407 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n15035) );
  NAND2_X1 U14408 ( .A1(n12621), .A2(n15035), .ZN(n12622) );
  NAND2_X1 U14409 ( .A1(n7213), .A2(n15195), .ZN(n12624) );
  NAND2_X1 U14410 ( .A1(n12829), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n12623) );
  NAND2_X1 U14411 ( .A1(n14867), .A2(n7232), .ZN(n12628) );
  OR2_X1 U14412 ( .A1(n9902), .A2(n15511), .ZN(n12627) );
  NAND2_X1 U14413 ( .A1(n12834), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n12632) );
  NAND2_X1 U14414 ( .A1(n12833), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n12631) );
  XNOR2_X1 U14415 ( .A(n12637), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n14922) );
  NAND2_X1 U14416 ( .A1(n7212), .A2(n14922), .ZN(n12630) );
  NAND2_X1 U14417 ( .A1(n12829), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n12629) );
  NAND2_X1 U14418 ( .A1(n14862), .A2(n7232), .ZN(n12634) );
  OR2_X1 U14419 ( .A1(n9902), .A2(n12671), .ZN(n12633) );
  NAND2_X1 U14420 ( .A1(n12834), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n12642) );
  NAND2_X1 U14421 ( .A1(n12833), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n12641) );
  INV_X1 U14422 ( .A(n12637), .ZN(n12636) );
  AND2_X1 U14423 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n12635) );
  NAND2_X1 U14424 ( .A1(n12636), .A2(n12635), .ZN(n12643) );
  INV_X1 U14425 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14919) );
  INV_X1 U14426 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n14959) );
  OAI21_X1 U14427 ( .B1(n12637), .B2(n14919), .A(n14959), .ZN(n12638) );
  NAND2_X1 U14428 ( .A1(n7213), .A2(n14960), .ZN(n12640) );
  NAND2_X1 U14429 ( .A1(n12829), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n12639) );
  NAND4_X1 U14430 ( .A1(n12642), .A2(n12641), .A3(n12640), .A4(n12639), .ZN(
        n15401) );
  XNOR2_X1 U14431 ( .A(n15408), .B(n15401), .ZN(n12880) );
  INV_X1 U14432 ( .A(n12880), .ZN(n12665) );
  XNOR2_X1 U14433 ( .A(n15179), .B(n12665), .ZN(n12651) );
  NAND2_X1 U14434 ( .A1(n12834), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n12647) );
  NAND2_X1 U14435 ( .A1(n12833), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n12646) );
  INV_X1 U14436 ( .A(n12643), .ZN(n15168) );
  NAND2_X1 U14437 ( .A1(n7212), .A2(n15168), .ZN(n12645) );
  NAND2_X1 U14438 ( .A1(n12829), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12644) );
  INV_X1 U14439 ( .A(n14962), .ZN(n15055) );
  NAND2_X1 U14440 ( .A1(n15055), .A2(n15376), .ZN(n12649) );
  NAND2_X1 U14441 ( .A1(n15056), .A2(n16030), .ZN(n12648) );
  AOI21_X2 U14442 ( .B1(n12651), .B2(n16119), .A(n12650), .ZN(n15411) );
  INV_X1 U14443 ( .A(n16133), .ZN(n15366) );
  NAND2_X1 U14444 ( .A1(n7271), .A2(n15345), .ZN(n15339) );
  OR2_X2 U14445 ( .A1(n15466), .A2(n15339), .ZN(n15326) );
  INV_X1 U14446 ( .A(n12930), .ZN(n12653) );
  NAND2_X1 U14447 ( .A1(n15176), .A2(n12930), .ZN(n15166) );
  INV_X1 U14448 ( .A(n15166), .ZN(n12652) );
  AOI21_X1 U14449 ( .B1(n15408), .B2(n12653), .A(n12652), .ZN(n15409) );
  AOI22_X1 U14450 ( .A1(n16001), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n14960), 
        .B2(n15990), .ZN(n12654) );
  OAI21_X1 U14451 ( .B1(n15176), .B2(n15365), .A(n12654), .ZN(n12668) );
  INV_X1 U14452 ( .A(n15413), .ZN(n14924) );
  INV_X1 U14453 ( .A(n15439), .ZN(n12664) );
  OR2_X1 U14454 ( .A1(n15386), .A2(n16088), .ZN(n12655) );
  OR2_X1 U14455 ( .A1(n16133), .A2(n15375), .ZN(n12656) );
  NAND2_X1 U14456 ( .A1(n15474), .A2(n15064), .ZN(n12658) );
  OR2_X1 U14457 ( .A1(n15466), .A2(n15063), .ZN(n12660) );
  AND2_X1 U14458 ( .A1(n15466), .A2(n15063), .ZN(n12659) );
  INV_X1 U14459 ( .A(n15303), .ZN(n15307) );
  OR2_X1 U14460 ( .A1(n15460), .A2(n15062), .ZN(n12661) );
  INV_X1 U14461 ( .A(n15061), .ZN(n15310) );
  INV_X1 U14462 ( .A(n15276), .ZN(n12663) );
  INV_X1 U14463 ( .A(n15254), .ZN(n15250) );
  NAND2_X1 U14464 ( .A1(n15251), .A2(n15250), .ZN(n15249) );
  INV_X1 U14465 ( .A(n15203), .ZN(n15208) );
  OAI21_X1 U14466 ( .B1(n12666), .B2(n12665), .A(n15164), .ZN(n15412) );
  NOR2_X1 U14467 ( .A1(n15412), .A2(n15392), .ZN(n12667) );
  OAI21_X1 U14468 ( .B1(n15411), .B2(n16001), .A(n12669), .ZN(P1_U3265) );
  INV_X1 U14469 ( .A(n14862), .ZN(n12670) );
  OAI222_X1 U14470 ( .A1(n15512), .A2(n12671), .B1(n15510), .B2(n12670), .C1(
        n10231), .C2(n7201), .ZN(P1_U3327) );
  MUX2_X1 U14471 ( .A(n15401), .B(n15408), .S(n12702), .Z(n12819) );
  INV_X1 U14472 ( .A(n12819), .ZN(n12823) );
  INV_X1 U14473 ( .A(n12673), .ZN(n12689) );
  MUX2_X1 U14474 ( .A(n15075), .B(n12674), .S(n12826), .Z(n12688) );
  NAND2_X1 U14475 ( .A1(n15878), .A2(n12702), .ZN(n12681) );
  MUX2_X1 U14476 ( .A(n8048), .B(n12675), .S(n12843), .Z(n12678) );
  OAI21_X1 U14477 ( .B1(n15878), .B2(n12676), .A(n12678), .ZN(n12677) );
  NAND2_X1 U14478 ( .A1(n10907), .A2(n12677), .ZN(n12680) );
  OR2_X1 U14479 ( .A1(n15878), .A2(n12678), .ZN(n12679) );
  OAI211_X1 U14480 ( .C1(n10907), .C2(n12681), .A(n12680), .B(n12679), .ZN(
        n12682) );
  NAND2_X1 U14481 ( .A1(n12683), .A2(n12682), .ZN(n12687) );
  NAND2_X1 U14482 ( .A1(n15074), .A2(n12690), .ZN(n12684) );
  NAND2_X1 U14483 ( .A1(n12685), .A2(n12684), .ZN(n12686) );
  OAI211_X1 U14484 ( .C1(n12689), .C2(n12688), .A(n12687), .B(n12686), .ZN(
        n12696) );
  OAI21_X1 U14485 ( .B1(n15074), .B2(n12743), .A(n12690), .ZN(n12694) );
  NAND2_X1 U14486 ( .A1(n15074), .A2(n12743), .ZN(n12692) );
  NAND2_X1 U14487 ( .A1(n12692), .A2(n12691), .ZN(n12693) );
  NAND2_X1 U14488 ( .A1(n12694), .A2(n12693), .ZN(n12695) );
  NAND3_X1 U14489 ( .A1(n12696), .A2(n12855), .A3(n12695), .ZN(n12701) );
  INV_X1 U14490 ( .A(n12697), .ZN(n12699) );
  AOI21_X1 U14491 ( .B1(n15073), .B2(n12826), .A(n15906), .ZN(n12698) );
  OR2_X1 U14492 ( .A1(n12699), .A2(n12698), .ZN(n12700) );
  NAND2_X1 U14493 ( .A1(n12701), .A2(n12700), .ZN(n12708) );
  MUX2_X1 U14494 ( .A(n15072), .B(n12703), .S(n12743), .Z(n12707) );
  NAND2_X1 U14495 ( .A1(n12708), .A2(n12707), .ZN(n12705) );
  MUX2_X1 U14496 ( .A(n15072), .B(n12703), .S(n12826), .Z(n12704) );
  NAND2_X1 U14497 ( .A1(n12705), .A2(n12704), .ZN(n12706) );
  OAI211_X1 U14498 ( .C1(n12708), .C2(n12707), .A(n12706), .B(n12860), .ZN(
        n12715) );
  OAI21_X1 U14499 ( .B1(n15071), .B2(n12826), .A(n12709), .ZN(n12713) );
  NAND2_X1 U14500 ( .A1(n15071), .A2(n12826), .ZN(n12711) );
  NAND2_X1 U14501 ( .A1(n12711), .A2(n12710), .ZN(n12712) );
  NAND2_X1 U14502 ( .A1(n12713), .A2(n12712), .ZN(n12714) );
  NAND2_X1 U14503 ( .A1(n12715), .A2(n12714), .ZN(n12719) );
  MUX2_X1 U14504 ( .A(n15070), .B(n12716), .S(n12743), .Z(n12720) );
  NAND2_X1 U14505 ( .A1(n12719), .A2(n12720), .ZN(n12718) );
  MUX2_X1 U14506 ( .A(n15070), .B(n12716), .S(n12826), .Z(n12717) );
  NAND2_X1 U14507 ( .A1(n12718), .A2(n12717), .ZN(n12724) );
  INV_X1 U14508 ( .A(n12719), .ZN(n12722) );
  INV_X1 U14509 ( .A(n12720), .ZN(n12721) );
  NAND2_X1 U14510 ( .A1(n12722), .A2(n12721), .ZN(n12723) );
  MUX2_X1 U14511 ( .A(n15069), .B(n12725), .S(n12743), .Z(n12726) );
  MUX2_X1 U14512 ( .A(n15068), .B(n15992), .S(n12743), .Z(n12731) );
  NAND2_X1 U14513 ( .A1(n12730), .A2(n12731), .ZN(n12729) );
  MUX2_X1 U14514 ( .A(n15068), .B(n15992), .S(n12826), .Z(n12728) );
  NAND2_X1 U14515 ( .A1(n12729), .A2(n12728), .ZN(n12735) );
  INV_X1 U14516 ( .A(n12730), .ZN(n12733) );
  INV_X1 U14517 ( .A(n12731), .ZN(n12732) );
  NAND2_X1 U14518 ( .A1(n12733), .A2(n12732), .ZN(n12734) );
  MUX2_X1 U14519 ( .A(n16029), .B(n16019), .S(n12826), .Z(n12738) );
  MUX2_X1 U14520 ( .A(n16029), .B(n16019), .S(n12743), .Z(n12736) );
  AND2_X1 U14521 ( .A1(n15067), .A2(n12743), .ZN(n12740) );
  OAI21_X1 U14522 ( .B1(n12743), .B2(n15067), .A(n16031), .ZN(n12739) );
  OAI21_X1 U14523 ( .B1(n12740), .B2(n16031), .A(n12739), .ZN(n12741) );
  MUX2_X1 U14524 ( .A(n15066), .B(n12744), .S(n12826), .Z(n12746) );
  MUX2_X1 U14525 ( .A(n15066), .B(n12744), .S(n12743), .Z(n12745) );
  MUX2_X1 U14526 ( .A(n15065), .B(n12747), .S(n12743), .Z(n12749) );
  MUX2_X1 U14527 ( .A(n15065), .B(n12747), .S(n12826), .Z(n12748) );
  INV_X1 U14528 ( .A(n12749), .ZN(n12750) );
  MUX2_X1 U14529 ( .A(n16086), .B(n12751), .S(n12826), .Z(n12754) );
  MUX2_X1 U14530 ( .A(n16086), .B(n12751), .S(n12743), .Z(n12752) );
  MUX2_X1 U14531 ( .A(n15374), .B(n12755), .S(n12743), .Z(n12757) );
  MUX2_X1 U14532 ( .A(n15374), .B(n12755), .S(n12826), .Z(n12756) );
  MUX2_X1 U14533 ( .A(n16088), .B(n15386), .S(n12826), .Z(n12761) );
  NAND2_X1 U14534 ( .A1(n12760), .A2(n12761), .ZN(n12759) );
  MUX2_X1 U14535 ( .A(n16088), .B(n15386), .S(n12702), .Z(n12758) );
  NAND2_X1 U14536 ( .A1(n12759), .A2(n12758), .ZN(n12765) );
  INV_X1 U14537 ( .A(n12760), .ZN(n12763) );
  INV_X1 U14538 ( .A(n12761), .ZN(n12762) );
  NAND2_X1 U14539 ( .A1(n12763), .A2(n12762), .ZN(n12764) );
  NAND2_X1 U14540 ( .A1(n12765), .A2(n12764), .ZN(n12768) );
  MUX2_X1 U14541 ( .A(n15375), .B(n16133), .S(n12702), .Z(n12767) );
  MUX2_X1 U14542 ( .A(n15375), .B(n16133), .S(n12826), .Z(n12766) );
  MUX2_X1 U14543 ( .A(n15064), .B(n15474), .S(n12826), .Z(n12770) );
  MUX2_X1 U14544 ( .A(n15474), .B(n15064), .S(n12826), .Z(n12769) );
  INV_X1 U14545 ( .A(n12770), .ZN(n12771) );
  MUX2_X1 U14546 ( .A(n15063), .B(n15466), .S(n12743), .Z(n12773) );
  MUX2_X1 U14547 ( .A(n15063), .B(n15466), .S(n12826), .Z(n12772) );
  INV_X1 U14548 ( .A(n12773), .ZN(n12774) );
  MUX2_X1 U14549 ( .A(n15062), .B(n15460), .S(n12826), .Z(n12777) );
  MUX2_X1 U14550 ( .A(n15062), .B(n15460), .S(n12743), .Z(n12775) );
  MUX2_X1 U14551 ( .A(n15061), .B(n15299), .S(n12743), .Z(n12779) );
  MUX2_X1 U14552 ( .A(n15061), .B(n15299), .S(n12826), .Z(n12778) );
  MUX2_X1 U14553 ( .A(n15444), .B(n15259), .S(n12702), .Z(n12782) );
  OAI21_X1 U14554 ( .B1(n12783), .B2(n12782), .A(n15254), .ZN(n12785) );
  MUX2_X1 U14555 ( .A(n15273), .B(n12780), .S(n12826), .Z(n12781) );
  AOI21_X1 U14556 ( .B1(n12783), .B2(n12782), .A(n12781), .ZN(n12784) );
  AND2_X1 U14557 ( .A1(n14969), .A2(n12826), .ZN(n12787) );
  OAI21_X1 U14558 ( .B1(n14969), .B2(n12826), .A(n15439), .ZN(n12786) );
  OAI21_X1 U14559 ( .B1(n12787), .B2(n15439), .A(n12786), .ZN(n12788) );
  MUX2_X1 U14560 ( .A(n15257), .B(n15433), .S(n12826), .Z(n12791) );
  MUX2_X1 U14561 ( .A(n15257), .B(n15433), .S(n12702), .Z(n12789) );
  INV_X1 U14562 ( .A(n12790), .ZN(n12793) );
  INV_X1 U14563 ( .A(n12791), .ZN(n12792) );
  NAND2_X1 U14564 ( .A1(n12793), .A2(n12792), .ZN(n12794) );
  NAND2_X1 U14565 ( .A1(n12795), .A2(n12794), .ZN(n12798) );
  MUX2_X1 U14566 ( .A(n15059), .B(n15429), .S(n12743), .Z(n12797) );
  MUX2_X1 U14567 ( .A(n15059), .B(n15429), .S(n12826), .Z(n12796) );
  MUX2_X1 U14568 ( .A(n15058), .B(n15425), .S(n12826), .Z(n12802) );
  MUX2_X1 U14569 ( .A(n15058), .B(n15425), .S(n12743), .Z(n12799) );
  NAND2_X1 U14570 ( .A1(n12800), .A2(n12799), .ZN(n12806) );
  INV_X1 U14571 ( .A(n12801), .ZN(n12804) );
  INV_X1 U14572 ( .A(n12802), .ZN(n12803) );
  NAND2_X1 U14573 ( .A1(n12804), .A2(n12803), .ZN(n12805) );
  NAND2_X1 U14574 ( .A1(n12806), .A2(n12805), .ZN(n12809) );
  MUX2_X1 U14575 ( .A(n15057), .B(n15420), .S(n12743), .Z(n12810) );
  NAND2_X1 U14576 ( .A1(n12809), .A2(n12810), .ZN(n12808) );
  MUX2_X1 U14577 ( .A(n15057), .B(n15420), .S(n12826), .Z(n12807) );
  NAND2_X1 U14578 ( .A1(n12808), .A2(n12807), .ZN(n12814) );
  INV_X1 U14579 ( .A(n12809), .ZN(n12812) );
  INV_X1 U14580 ( .A(n12810), .ZN(n12811) );
  MUX2_X1 U14581 ( .A(n15056), .B(n15413), .S(n12826), .Z(n12816) );
  MUX2_X1 U14582 ( .A(n15056), .B(n15413), .S(n12702), .Z(n12815) );
  INV_X1 U14583 ( .A(n12816), .ZN(n12817) );
  INV_X1 U14584 ( .A(n12820), .ZN(n12822) );
  MUX2_X1 U14585 ( .A(n15176), .B(n15177), .S(n12702), .Z(n12818) );
  AOI21_X1 U14586 ( .B1(n12820), .B2(n12819), .A(n12818), .ZN(n12821) );
  NOR2_X1 U14587 ( .A1(n9902), .A2(n15507), .ZN(n12824) );
  MUX2_X1 U14588 ( .A(n14962), .B(n15403), .S(n12826), .Z(n12827) );
  MUX2_X1 U14589 ( .A(n14962), .B(n15403), .S(n12702), .Z(n12828) );
  NAND2_X1 U14590 ( .A1(n12833), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12832) );
  NAND2_X1 U14591 ( .A1(n12829), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n12831) );
  NAND2_X1 U14592 ( .A1(n12834), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12830) );
  AND3_X1 U14593 ( .A1(n12832), .A2(n12831), .A3(n12830), .ZN(n12889) );
  NAND2_X1 U14594 ( .A1(n12833), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U14595 ( .A1(n12829), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12836) );
  NAND2_X1 U14596 ( .A1(n12834), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12835) );
  NAND3_X1 U14597 ( .A1(n12837), .A2(n12836), .A3(n12835), .ZN(n15400) );
  OAI21_X1 U14598 ( .B1(n15155), .B2(n12838), .A(n15400), .ZN(n12839) );
  INV_X1 U14599 ( .A(n12839), .ZN(n12842) );
  INV_X1 U14600 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13357) );
  OR2_X1 U14601 ( .A1(n9902), .A2(n13357), .ZN(n12840) );
  MUX2_X1 U14602 ( .A(n12842), .B(n15153), .S(n12702), .Z(n12901) );
  INV_X1 U14603 ( .A(n12901), .ZN(n12908) );
  OAI21_X1 U14604 ( .B1(n15155), .B2(n12843), .A(n15400), .ZN(n12844) );
  INV_X1 U14605 ( .A(n12844), .ZN(n12845) );
  MUX2_X1 U14606 ( .A(n15153), .B(n12845), .S(n12702), .Z(n12907) );
  NAND2_X1 U14607 ( .A1(n14851), .A2(n7232), .ZN(n12848) );
  INV_X1 U14608 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12846) );
  OR2_X1 U14609 ( .A1(n9902), .A2(n12846), .ZN(n12847) );
  XNOR2_X1 U14610 ( .A(n15156), .B(n12889), .ZN(n12883) );
  INV_X1 U14611 ( .A(n12883), .ZN(n12910) );
  INV_X1 U14612 ( .A(n12849), .ZN(n12850) );
  NAND2_X1 U14613 ( .A1(n12851), .A2(n12850), .ZN(n12853) );
  AND2_X1 U14614 ( .A1(n12853), .A2(n12852), .ZN(n12892) );
  INV_X1 U14615 ( .A(n12892), .ZN(n12898) );
  NOR2_X1 U14616 ( .A1(n12898), .A2(n12913), .ZN(n12909) );
  OAI211_X1 U14617 ( .C1(n12908), .C2(n12907), .A(n12910), .B(n12909), .ZN(
        n12919) );
  XNOR2_X1 U14618 ( .A(n15153), .B(n15400), .ZN(n12882) );
  NAND4_X1 U14619 ( .A1(n12855), .A2(n15875), .A3(n12854), .A4(n12683), .ZN(
        n12857) );
  NOR2_X1 U14620 ( .A1(n12857), .A2(n12856), .ZN(n12861) );
  NAND4_X1 U14621 ( .A1(n12861), .A2(n12860), .A3(n12859), .A4(n12858), .ZN(
        n12862) );
  NOR2_X1 U14622 ( .A1(n15983), .A2(n12862), .ZN(n12865) );
  NAND4_X1 U14623 ( .A1(n12866), .A2(n12865), .A3(n12864), .A4(n12863), .ZN(
        n12867) );
  NOR2_X1 U14624 ( .A1(n12868), .A2(n12867), .ZN(n12870) );
  AND4_X1 U14625 ( .A1(n15338), .A2(n12870), .A3(n15351), .A4(n12869), .ZN(
        n12873) );
  NAND4_X1 U14626 ( .A1(n15290), .A2(n12873), .A3(n12872), .A4(n12871), .ZN(
        n12874) );
  NOR2_X1 U14627 ( .A1(n15276), .A2(n12874), .ZN(n12875) );
  NAND4_X1 U14628 ( .A1(n15254), .A2(n12875), .A3(n15322), .A4(n15303), .ZN(
        n12876) );
  OR4_X1 U14629 ( .A1(n15203), .A2(n15220), .A3(n12877), .A4(n12876), .ZN(
        n12878) );
  NOR2_X1 U14630 ( .A1(n12879), .A2(n12878), .ZN(n12881) );
  NAND4_X1 U14631 ( .A1(n12882), .A2(n12881), .A3(n12923), .A4(n12880), .ZN(
        n12884) );
  XNOR2_X1 U14632 ( .A(n15167), .B(n14962), .ZN(n15182) );
  OR3_X1 U14633 ( .A1(n12884), .A2(n12883), .A3(n15182), .ZN(n12886) );
  XNOR2_X1 U14634 ( .A(n12886), .B(n7228), .ZN(n12888) );
  NAND2_X1 U14635 ( .A1(n15156), .A2(n12889), .ZN(n12891) );
  OR2_X1 U14636 ( .A1(n15156), .A2(n12889), .ZN(n12890) );
  MUX2_X1 U14637 ( .A(n12891), .B(n12890), .S(n12826), .Z(n12896) );
  XNOR2_X1 U14638 ( .A(n12896), .B(n12892), .ZN(n12893) );
  NAND2_X1 U14639 ( .A1(n12893), .A2(n12897), .ZN(n12894) );
  INV_X1 U14640 ( .A(n12907), .ZN(n12895) );
  NAND2_X1 U14641 ( .A1(n12895), .A2(n8001), .ZN(n12902) );
  INV_X1 U14642 ( .A(n12896), .ZN(n12906) );
  AND2_X1 U14643 ( .A1(n12898), .A2(n12897), .ZN(n12904) );
  INV_X1 U14644 ( .A(n12904), .ZN(n12899) );
  NOR2_X1 U14645 ( .A1(n12899), .A2(n12913), .ZN(n12900) );
  NAND2_X1 U14646 ( .A1(n12901), .A2(n12900), .ZN(n12905) );
  OAI22_X1 U14647 ( .A1(n12903), .A2(n12902), .B1(n12906), .B2(n12905), .ZN(
        n12917) );
  OR3_X1 U14648 ( .A1(n12906), .A2(n12907), .A3(n12905), .ZN(n12916) );
  NAND4_X1 U14649 ( .A1(n12910), .A2(n12909), .A3(n12908), .A4(n12907), .ZN(
        n12915) );
  NAND3_X1 U14650 ( .A1(n12911), .A2(n15633), .A3(n16030), .ZN(n12912) );
  OAI211_X1 U14651 ( .C1(n15513), .C2(n12913), .A(n12912), .B(P1_B_REG_SCAN_IN), .ZN(n12914) );
  OAI21_X1 U14652 ( .B1(n12920), .B2(n12919), .A(n12918), .ZN(P1_U3242) );
  AOI21_X1 U14653 ( .B1(n12923), .B2(n12922), .A(n12921), .ZN(n15417) );
  XNOR2_X1 U14654 ( .A(n12924), .B(n12923), .ZN(n12926) );
  OAI22_X1 U14655 ( .A1(n15177), .A2(n15359), .B1(n14918), .B2(n15357), .ZN(
        n12925) );
  AOI21_X1 U14656 ( .B1(n15413), .B2(n15192), .A(n12930), .ZN(n15414) );
  AOI22_X1 U14657 ( .A1(n16001), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14922), 
        .B2(n15990), .ZN(n12931) );
  OAI21_X1 U14658 ( .B1(n14924), .B2(n15365), .A(n12931), .ZN(n12934) );
  NOR2_X1 U14659 ( .A1(n15417), .A2(n12932), .ZN(n12933) );
  AOI211_X1 U14660 ( .C1(n15347), .C2(n15414), .A(n12934), .B(n12933), .ZN(
        n12935) );
  OAI21_X1 U14661 ( .B1(n15416), .B2(n16001), .A(n12935), .ZN(P1_U3266) );
  OAI222_X1 U14662 ( .A1(n15510), .A2(n14859), .B1(P1_U3086), .B2(n12936), 
        .C1(n13357), .C2(n15512), .ZN(P1_U3325) );
  INV_X1 U14663 ( .A(n14039), .ZN(n13862) );
  OR2_X1 U14664 ( .A1(n13987), .A2(n13348), .ZN(n13455) );
  NAND2_X1 U14665 ( .A1(n13987), .A2(n13348), .ZN(n13454) );
  NAND2_X1 U14666 ( .A1(n13455), .A2(n13454), .ZN(n13972) );
  NAND2_X1 U14667 ( .A1(n13987), .A2(n13959), .ZN(n12939) );
  NAND2_X1 U14668 ( .A1(n14133), .A2(n13974), .ZN(n13458) );
  NAND2_X1 U14669 ( .A1(n13459), .A2(n13458), .ZN(n13956) );
  OR2_X1 U14670 ( .A1(n14133), .A2(n13945), .ZN(n12940) );
  XNOR2_X1 U14671 ( .A(n13468), .B(n13958), .ZN(n13941) );
  OR2_X1 U14672 ( .A1(n13468), .A2(n13958), .ZN(n12941) );
  OR2_X1 U14673 ( .A1(n14123), .A2(n13943), .ZN(n13379) );
  NAND2_X1 U14674 ( .A1(n14123), .A2(n13943), .ZN(n13906) );
  NAND2_X1 U14675 ( .A1(n14054), .A2(n13899), .ZN(n12972) );
  NAND2_X1 U14676 ( .A1(n13378), .A2(n12972), .ZN(n13912) );
  NOR2_X1 U14677 ( .A1(n14051), .A2(n13915), .ZN(n12943) );
  INV_X1 U14678 ( .A(n14051), .ZN(n13903) );
  NAND2_X1 U14679 ( .A1(n14118), .A2(n13866), .ZN(n13476) );
  INV_X1 U14680 ( .A(n14118), .ZN(n12944) );
  NAND2_X1 U14681 ( .A1(n12944), .A2(n13900), .ZN(n13475) );
  NAND2_X1 U14682 ( .A1(n13476), .A2(n13475), .ZN(n13540) );
  AOI22_X2 U14683 ( .A1(n13879), .A2(n13540), .B1(n13866), .B2(n12944), .ZN(
        n13865) );
  NAND2_X1 U14684 ( .A1(n12977), .A2(n13857), .ZN(n12945) );
  OR2_X1 U14685 ( .A1(n14039), .A2(n13846), .ZN(n13375) );
  NAND2_X1 U14686 ( .A1(n14039), .A2(n13846), .ZN(n13376) );
  NAND2_X1 U14687 ( .A1(n13375), .A2(n13376), .ZN(n13855) );
  XNOR2_X1 U14688 ( .A(n14035), .B(n13826), .ZN(n13841) );
  INV_X1 U14689 ( .A(n14035), .ZN(n13246) );
  NAND2_X1 U14690 ( .A1(n14108), .A2(n13812), .ZN(n12948) );
  NAND2_X1 U14691 ( .A1(n12949), .A2(n13827), .ZN(n13491) );
  XNOR2_X1 U14692 ( .A(n13494), .B(n13813), .ZN(n12983) );
  NAND2_X1 U14693 ( .A1(n14096), .A2(n13574), .ZN(n13497) );
  NAND2_X1 U14694 ( .A1(n12950), .A2(n12951), .ZN(n13496) );
  NAND2_X1 U14695 ( .A1(n14865), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12953) );
  AND2_X2 U14696 ( .A1(n12954), .A2(n12953), .ZN(n12955) );
  XNOR2_X1 U14697 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12956) );
  INV_X1 U14698 ( .A(n12955), .ZN(n12958) );
  INV_X1 U14699 ( .A(n12956), .ZN(n12957) );
  NAND2_X1 U14700 ( .A1(n12958), .A2(n12957), .ZN(n12959) );
  NAND2_X1 U14701 ( .A1(n13210), .A2(n12959), .ZN(n14152) );
  OR2_X1 U14702 ( .A1(n12960), .A2(n14151), .ZN(n12961) );
  NAND2_X1 U14703 ( .A1(n12988), .A2(n13572), .ZN(n13551) );
  NAND2_X1 U14704 ( .A1(n13218), .A2(n13767), .ZN(n13515) );
  NAND2_X1 U14705 ( .A1(n13551), .A2(n13515), .ZN(n12987) );
  AND2_X1 U14706 ( .A1(n12963), .A2(P3_B_REG_SCAN_IN), .ZN(n12964) );
  NOR2_X1 U14707 ( .A1(n13944), .A2(n12964), .ZN(n13758) );
  NAND2_X1 U14708 ( .A1(n13365), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12967) );
  NAND2_X1 U14709 ( .A1(n13364), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n12966) );
  NAND2_X1 U14710 ( .A1(n8472), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12965) );
  NAND4_X1 U14711 ( .A1(n13369), .A2(n12967), .A3(n12966), .A4(n12965), .ZN(
        n13571) );
  INV_X1 U14712 ( .A(n13787), .ZN(n13573) );
  AOI22_X1 U14713 ( .A1(n13758), .A2(n13571), .B1(n13573), .B2(n13997), .ZN(
        n12968) );
  NAND2_X1 U14714 ( .A1(n12970), .A2(n13450), .ZN(n13978) );
  INV_X1 U14715 ( .A(n13972), .ZN(n13977) );
  NAND2_X1 U14716 ( .A1(n13978), .A2(n13977), .ZN(n13980) );
  INV_X1 U14717 ( .A(n13378), .ZN(n13892) );
  INV_X1 U14718 ( .A(n13521), .ZN(n12975) );
  INV_X1 U14719 ( .A(n13906), .ZN(n12971) );
  NAND2_X1 U14720 ( .A1(n13378), .A2(n12971), .ZN(n12973) );
  AND2_X1 U14721 ( .A1(n8229), .A2(n13893), .ZN(n12974) );
  NOR2_X1 U14722 ( .A1(n12977), .A2(n13880), .ZN(n13479) );
  INV_X1 U14723 ( .A(n13855), .ZN(n12978) );
  NAND2_X1 U14724 ( .A1(n13853), .A2(n12978), .ZN(n12979) );
  OR2_X1 U14725 ( .A1(n14035), .A2(n13826), .ZN(n13487) );
  NAND2_X1 U14726 ( .A1(n12980), .A2(n13812), .ZN(n13499) );
  NAND2_X1 U14727 ( .A1(n13809), .A2(n13811), .ZN(n12982) );
  OR2_X1 U14728 ( .A1(n13494), .A2(n13813), .ZN(n12984) );
  INV_X1 U14729 ( .A(n13496), .ZN(n13772) );
  NOR2_X1 U14730 ( .A1(n13771), .A2(n13772), .ZN(n12986) );
  INV_X1 U14731 ( .A(n12987), .ZN(n13546) );
  OAI22_X1 U14732 ( .A1(n12993), .A2(keyinput_52), .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .ZN(n12992) );
  AOI221_X1 U14733 ( .B1(n12993), .B2(keyinput_52), .C1(keyinput_51), .C2(
        P3_REG3_REG_24__SCAN_IN), .A(n12992), .ZN(n13076) );
  OAI22_X1 U14734 ( .A1(n8391), .A2(keyinput_49), .B1(n12995), .B2(keyinput_48), .ZN(n12994) );
  AOI221_X1 U14735 ( .B1(n8391), .B2(keyinput_49), .C1(keyinput_48), .C2(
        n12995), .A(n12994), .ZN(n13073) );
  INV_X1 U14736 ( .A(keyinput_47), .ZN(n13071) );
  INV_X1 U14737 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n13177) );
  INV_X1 U14738 ( .A(keyinput_46), .ZN(n13069) );
  XNOR2_X1 U14739 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n13057)
         );
  INV_X1 U14740 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15874) );
  INV_X1 U14741 ( .A(keyinput_23), .ZN(n13029) );
  INV_X1 U14742 ( .A(keyinput_22), .ZN(n13027) );
  INV_X1 U14743 ( .A(keyinput_21), .ZN(n13025) );
  INV_X1 U14744 ( .A(SI_17_), .ZN(n13119) );
  AOI22_X1 U14745 ( .A1(SI_19_), .A2(keyinput_13), .B1(n13093), .B2(
        keyinput_14), .ZN(n12996) );
  OAI221_X1 U14746 ( .B1(SI_19_), .B2(keyinput_13), .C1(n13093), .C2(
        keyinput_14), .A(n12996), .ZN(n13015) );
  INV_X1 U14747 ( .A(keyinput_12), .ZN(n13013) );
  INV_X1 U14748 ( .A(keyinput_11), .ZN(n13011) );
  OAI22_X1 U14749 ( .A1(SI_25_), .A2(keyinput_7), .B1(SI_26_), .B2(keyinput_6), 
        .ZN(n12997) );
  AOI221_X1 U14750 ( .B1(SI_25_), .B2(keyinput_7), .C1(keyinput_6), .C2(SI_26_), .A(n12997), .ZN(n13009) );
  XOR2_X1 U14751 ( .A(SI_30_), .B(keyinput_2), .Z(n13003) );
  AOI22_X1 U14752 ( .A1(SI_31_), .A2(keyinput_1), .B1(P3_WR_REG_SCAN_IN), .B2(
        keyinput_0), .ZN(n12998) );
  OAI221_X1 U14753 ( .B1(SI_31_), .B2(keyinput_1), .C1(P3_WR_REG_SCAN_IN), 
        .C2(keyinput_0), .A(n12998), .ZN(n13002) );
  OAI22_X1 U14754 ( .A1(n14151), .A2(keyinput_3), .B1(SI_27_), .B2(keyinput_5), 
        .ZN(n12999) );
  AOI221_X1 U14755 ( .B1(n14151), .B2(keyinput_3), .C1(keyinput_5), .C2(SI_27_), .A(n12999), .ZN(n13001) );
  XNOR2_X1 U14756 ( .A(SI_28_), .B(keyinput_4), .ZN(n13000) );
  OAI211_X1 U14757 ( .C1(n13003), .C2(n13002), .A(n13001), .B(n13000), .ZN(
        n13008) );
  XOR2_X1 U14758 ( .A(SI_23_), .B(keyinput_9), .Z(n13007) );
  AOI22_X1 U14759 ( .A1(keyinput_10), .A2(SI_22_), .B1(n13005), .B2(keyinput_8), .ZN(n13004) );
  OAI221_X1 U14760 ( .B1(keyinput_10), .B2(SI_22_), .C1(n13005), .C2(
        keyinput_8), .A(n13004), .ZN(n13006) );
  AOI211_X1 U14761 ( .C1(n13009), .C2(n13008), .A(n13007), .B(n13006), .ZN(
        n13010) );
  AOI221_X1 U14762 ( .B1(SI_21_), .B2(keyinput_11), .C1(n13112), .C2(n13011), 
        .A(n13010), .ZN(n13012) );
  AOI221_X1 U14763 ( .B1(SI_20_), .B2(keyinput_12), .C1(n13114), .C2(n13013), 
        .A(n13012), .ZN(n13014) );
  OAI22_X1 U14764 ( .A1(keyinput_15), .A2(n13119), .B1(n13015), .B2(n13014), 
        .ZN(n13016) );
  AOI21_X1 U14765 ( .B1(keyinput_15), .B2(n13119), .A(n13016), .ZN(n13023) );
  XNOR2_X1 U14766 ( .A(SI_16_), .B(keyinput_16), .ZN(n13022) );
  OAI22_X1 U14767 ( .A1(n13124), .A2(keyinput_18), .B1(n13122), .B2(
        keyinput_17), .ZN(n13017) );
  AOI221_X1 U14768 ( .B1(n13124), .B2(keyinput_18), .C1(keyinput_17), .C2(
        n13122), .A(n13017), .ZN(n13021) );
  OAI22_X1 U14769 ( .A1(n13019), .A2(keyinput_20), .B1(n13121), .B2(
        keyinput_19), .ZN(n13018) );
  AOI221_X1 U14770 ( .B1(n13019), .B2(keyinput_20), .C1(keyinput_19), .C2(
        n13121), .A(n13018), .ZN(n13020) );
  OAI211_X1 U14771 ( .C1(n13023), .C2(n13022), .A(n13021), .B(n13020), .ZN(
        n13024) );
  OAI221_X1 U14772 ( .B1(SI_11_), .B2(keyinput_21), .C1(n13130), .C2(n13025), 
        .A(n13024), .ZN(n13026) );
  OAI221_X1 U14773 ( .B1(SI_10_), .B2(keyinput_22), .C1(n13133), .C2(n13027), 
        .A(n13026), .ZN(n13028) );
  OAI221_X1 U14774 ( .B1(SI_9_), .B2(keyinput_23), .C1(n13136), .C2(n13029), 
        .A(n13028), .ZN(n13032) );
  INV_X1 U14775 ( .A(keyinput_24), .ZN(n13030) );
  MUX2_X1 U14776 ( .A(n13030), .B(keyinput_24), .S(SI_8_), .Z(n13031) );
  NAND2_X1 U14777 ( .A1(n13032), .A2(n13031), .ZN(n13035) );
  INV_X1 U14778 ( .A(keyinput_25), .ZN(n13033) );
  MUX2_X1 U14779 ( .A(n13033), .B(keyinput_25), .S(SI_7_), .Z(n13034) );
  NAND2_X1 U14780 ( .A1(n13035), .A2(n13034), .ZN(n13042) );
  INV_X1 U14781 ( .A(keyinput_26), .ZN(n13036) );
  MUX2_X1 U14782 ( .A(keyinput_26), .B(n13036), .S(SI_6_), .Z(n13041) );
  XOR2_X1 U14783 ( .A(SI_5_), .B(keyinput_27), .Z(n13039) );
  XOR2_X1 U14784 ( .A(SI_3_), .B(keyinput_29), .Z(n13038) );
  XNOR2_X1 U14785 ( .A(SI_4_), .B(keyinput_28), .ZN(n13037) );
  NAND3_X1 U14786 ( .A1(n13039), .A2(n13038), .A3(n13037), .ZN(n13040) );
  AOI21_X1 U14787 ( .B1(n13042), .B2(n13041), .A(n13040), .ZN(n13047) );
  INV_X1 U14788 ( .A(keyinput_30), .ZN(n13043) );
  MUX2_X1 U14789 ( .A(keyinput_30), .B(n13043), .S(SI_2_), .Z(n13046) );
  XOR2_X1 U14790 ( .A(SI_0_), .B(keyinput_32), .Z(n13045) );
  XNOR2_X1 U14791 ( .A(SI_1_), .B(keyinput_31), .ZN(n13044) );
  OAI211_X1 U14792 ( .C1(n13047), .C2(n13046), .A(n13045), .B(n13044), .ZN(
        n13048) );
  OAI21_X1 U14793 ( .B1(keyinput_33), .B2(n15874), .A(n13048), .ZN(n13049) );
  AOI21_X1 U14794 ( .B1(keyinput_33), .B2(n15874), .A(n13049), .ZN(n13055) );
  AOI22_X1 U14795 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput_35), .B1(
        P3_U3151), .B2(keyinput_34), .ZN(n13050) );
  OAI221_X1 U14796 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput_35), .C1(
        P3_U3151), .C2(keyinput_34), .A(n13050), .ZN(n13054) );
  INV_X1 U14797 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n13235) );
  OAI22_X1 U14798 ( .A1(n13052), .A2(keyinput_36), .B1(n13235), .B2(
        keyinput_37), .ZN(n13051) );
  AOI221_X1 U14799 ( .B1(n13052), .B2(keyinput_36), .C1(keyinput_37), .C2(
        n13235), .A(n13051), .ZN(n13053) );
  OAI21_X1 U14800 ( .B1(n13055), .B2(n13054), .A(n13053), .ZN(n13056) );
  AOI22_X1 U14801 ( .A1(n13057), .A2(n13056), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(keyinput_40), .ZN(n13058) );
  OAI21_X1 U14802 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .A(n13058), 
        .ZN(n13067) );
  INV_X1 U14803 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n13250) );
  AOI22_X1 U14804 ( .A1(keyinput_39), .A2(P3_REG3_REG_10__SCAN_IN), .B1(n13250), .B2(keyinput_41), .ZN(n13059) );
  OAI221_X1 U14805 ( .B1(keyinput_39), .B2(P3_REG3_REG_10__SCAN_IN), .C1(
        n13250), .C2(keyinput_41), .A(n13059), .ZN(n13066) );
  INV_X1 U14806 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n13061) );
  OAI22_X1 U14807 ( .A1(n13062), .A2(keyinput_43), .B1(n13061), .B2(
        keyinput_45), .ZN(n13060) );
  AOI221_X1 U14808 ( .B1(n13062), .B2(keyinput_43), .C1(keyinput_45), .C2(
        n13061), .A(n13060), .ZN(n13065) );
  OAI22_X1 U14809 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(keyinput_42), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(keyinput_44), .ZN(n13063) );
  AOI221_X1 U14810 ( .B1(P3_REG3_REG_28__SCAN_IN), .B2(keyinput_42), .C1(
        keyinput_44), .C2(P3_REG3_REG_1__SCAN_IN), .A(n13063), .ZN(n13064) );
  OAI211_X1 U14811 ( .C1(n13067), .C2(n13066), .A(n13065), .B(n13064), .ZN(
        n13068) );
  OAI221_X1 U14812 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(n13069), .C1(n13174), 
        .C2(keyinput_46), .A(n13068), .ZN(n13070) );
  OAI221_X1 U14813 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(n13071), .C1(n13177), 
        .C2(keyinput_47), .A(n13070), .ZN(n13072) );
  AOI22_X1 U14814 ( .A1(n13073), .A2(n13072), .B1(keyinput_50), .B2(
        P3_REG3_REG_17__SCAN_IN), .ZN(n13074) );
  OAI21_X1 U14815 ( .B1(keyinput_50), .B2(P3_REG3_REG_17__SCAN_IN), .A(n13074), 
        .ZN(n13075) );
  OAI211_X1 U14816 ( .C1(P3_REG3_REG_9__SCAN_IN), .C2(keyinput_53), .A(n13076), 
        .B(n13075), .ZN(n13077) );
  AOI21_X1 U14817 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .A(n13077), 
        .ZN(n13086) );
  AOI22_X1 U14818 ( .A1(keyinput_57), .A2(P3_REG3_REG_22__SCAN_IN), .B1(n13079), .B2(keyinput_59), .ZN(n13078) );
  OAI221_X1 U14819 ( .B1(keyinput_57), .B2(P3_REG3_REG_22__SCAN_IN), .C1(
        n13079), .C2(keyinput_59), .A(n13078), .ZN(n13085) );
  AOI22_X1 U14820 ( .A1(keyinput_58), .A2(P3_REG3_REG_11__SCAN_IN), .B1(n8546), 
        .B2(keyinput_56), .ZN(n13080) );
  OAI221_X1 U14821 ( .B1(keyinput_58), .B2(P3_REG3_REG_11__SCAN_IN), .C1(n8546), .C2(keyinput_56), .A(n13080), .ZN(n13084) );
  XNOR2_X1 U14822 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n13082)
         );
  XNOR2_X1 U14823 ( .A(keyinput_55), .B(P3_REG3_REG_20__SCAN_IN), .ZN(n13081)
         );
  NAND2_X1 U14824 ( .A1(n13082), .A2(n13081), .ZN(n13083) );
  NOR4_X1 U14825 ( .A1(n13086), .A2(n13085), .A3(n13084), .A4(n13083), .ZN(
        n13207) );
  INV_X1 U14826 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n13196) );
  OR2_X1 U14827 ( .A1(n13196), .A2(keyinput_61), .ZN(n13088) );
  AOI22_X1 U14828 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_60), .B1(n13196), .B2(keyinput_61), .ZN(n13087) );
  OAI211_X1 U14829 ( .C1(keyinput_60), .C2(P3_REG3_REG_18__SCAN_IN), .A(n13088), .B(n13087), .ZN(n13206) );
  XOR2_X1 U14830 ( .A(keyinput_116), .B(P3_REG3_REG_4__SCAN_IN), .Z(n13186) );
  AOI22_X1 U14831 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_112), .B1(
        P3_REG3_REG_5__SCAN_IN), .B2(keyinput_113), .ZN(n13089) );
  OAI221_X1 U14832 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_112), .C1(
        P3_REG3_REG_5__SCAN_IN), .C2(keyinput_113), .A(n13089), .ZN(n13180) );
  INV_X1 U14833 ( .A(keyinput_111), .ZN(n13178) );
  INV_X1 U14834 ( .A(keyinput_110), .ZN(n13175) );
  XOR2_X1 U14835 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_102), .Z(n13163)
         );
  OAI22_X1 U14836 ( .A1(P3_STATE_REG_SCAN_IN), .A2(keyinput_98), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput_99), .ZN(n13090) );
  AOI221_X1 U14837 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput_98), .C1(
        keyinput_99), .C2(P3_REG3_REG_7__SCAN_IN), .A(n13090), .ZN(n13161) );
  INV_X1 U14838 ( .A(keyinput_87), .ZN(n13137) );
  INV_X1 U14839 ( .A(keyinput_86), .ZN(n13134) );
  INV_X1 U14840 ( .A(keyinput_85), .ZN(n13131) );
  XNOR2_X1 U14841 ( .A(SI_16_), .B(keyinput_80), .ZN(n13128) );
  OAI22_X1 U14842 ( .A1(n13093), .A2(keyinput_78), .B1(n13092), .B2(
        keyinput_77), .ZN(n13091) );
  AOI221_X1 U14843 ( .B1(n13093), .B2(keyinput_78), .C1(keyinput_77), .C2(
        n13092), .A(n13091), .ZN(n13117) );
  INV_X1 U14844 ( .A(keyinput_76), .ZN(n13115) );
  INV_X1 U14845 ( .A(keyinput_75), .ZN(n13111) );
  OAI22_X1 U14846 ( .A1(n14151), .A2(keyinput_67), .B1(SI_28_), .B2(
        keyinput_68), .ZN(n13094) );
  AOI221_X1 U14847 ( .B1(n14151), .B2(keyinput_67), .C1(keyinput_68), .C2(
        SI_28_), .A(n13094), .ZN(n13099) );
  INV_X1 U14848 ( .A(SI_31_), .ZN(n14145) );
  INV_X1 U14849 ( .A(keyinput_65), .ZN(n13097) );
  OAI22_X1 U14850 ( .A1(SI_30_), .A2(keyinput_66), .B1(P3_WR_REG_SCAN_IN), 
        .B2(keyinput_64), .ZN(n13095) );
  AOI221_X1 U14851 ( .B1(SI_30_), .B2(keyinput_66), .C1(keyinput_64), .C2(
        P3_WR_REG_SCAN_IN), .A(n13095), .ZN(n13096) );
  OAI221_X1 U14852 ( .B1(SI_31_), .B2(keyinput_65), .C1(n14145), .C2(n13097), 
        .A(n13096), .ZN(n13098) );
  OAI211_X1 U14853 ( .C1(n13101), .C2(keyinput_69), .A(n13099), .B(n13098), 
        .ZN(n13100) );
  AOI21_X1 U14854 ( .B1(n13101), .B2(keyinput_69), .A(n13100), .ZN(n13109) );
  AOI22_X1 U14855 ( .A1(SI_25_), .A2(keyinput_71), .B1(n13103), .B2(
        keyinput_70), .ZN(n13102) );
  OAI221_X1 U14856 ( .B1(SI_25_), .B2(keyinput_71), .C1(n13103), .C2(
        keyinput_70), .A(n13102), .ZN(n13108) );
  OAI22_X1 U14857 ( .A1(n13105), .A2(keyinput_74), .B1(SI_24_), .B2(
        keyinput_72), .ZN(n13104) );
  AOI221_X1 U14858 ( .B1(n13105), .B2(keyinput_74), .C1(keyinput_72), .C2(
        SI_24_), .A(n13104), .ZN(n13107) );
  XNOR2_X1 U14859 ( .A(SI_23_), .B(keyinput_73), .ZN(n13106) );
  OAI211_X1 U14860 ( .C1(n13109), .C2(n13108), .A(n13107), .B(n13106), .ZN(
        n13110) );
  OAI221_X1 U14861 ( .B1(SI_21_), .B2(keyinput_75), .C1(n13112), .C2(n13111), 
        .A(n13110), .ZN(n13113) );
  OAI221_X1 U14862 ( .B1(SI_20_), .B2(n13115), .C1(n13114), .C2(keyinput_76), 
        .A(n13113), .ZN(n13116) );
  AOI22_X1 U14863 ( .A1(keyinput_79), .A2(n13119), .B1(n13117), .B2(n13116), 
        .ZN(n13118) );
  OAI21_X1 U14864 ( .B1(n13119), .B2(keyinput_79), .A(n13118), .ZN(n13127) );
  AOI22_X1 U14865 ( .A1(n13122), .A2(keyinput_81), .B1(n13121), .B2(
        keyinput_83), .ZN(n13120) );
  OAI221_X1 U14866 ( .B1(n13122), .B2(keyinput_81), .C1(n13121), .C2(
        keyinput_83), .A(n13120), .ZN(n13126) );
  AOI22_X1 U14867 ( .A1(SI_12_), .A2(keyinput_84), .B1(n13124), .B2(
        keyinput_82), .ZN(n13123) );
  OAI221_X1 U14868 ( .B1(SI_12_), .B2(keyinput_84), .C1(n13124), .C2(
        keyinput_82), .A(n13123), .ZN(n13125) );
  AOI211_X1 U14869 ( .C1(n13128), .C2(n13127), .A(n13126), .B(n13125), .ZN(
        n13129) );
  AOI221_X1 U14870 ( .B1(SI_11_), .B2(n13131), .C1(n13130), .C2(keyinput_85), 
        .A(n13129), .ZN(n13132) );
  AOI221_X1 U14871 ( .B1(SI_10_), .B2(n13134), .C1(n13133), .C2(keyinput_86), 
        .A(n13132), .ZN(n13135) );
  AOI221_X1 U14872 ( .B1(SI_9_), .B2(n13137), .C1(n13136), .C2(keyinput_87), 
        .A(n13135), .ZN(n13140) );
  INV_X1 U14873 ( .A(keyinput_88), .ZN(n13138) );
  MUX2_X1 U14874 ( .A(keyinput_88), .B(n13138), .S(SI_8_), .Z(n13139) );
  NOR2_X1 U14875 ( .A1(n13140), .A2(n13139), .ZN(n13143) );
  INV_X1 U14876 ( .A(keyinput_89), .ZN(n13141) );
  MUX2_X1 U14877 ( .A(keyinput_89), .B(n13141), .S(SI_7_), .Z(n13142) );
  NOR2_X1 U14878 ( .A1(n13143), .A2(n13142), .ZN(n13150) );
  INV_X1 U14879 ( .A(keyinput_90), .ZN(n13144) );
  MUX2_X1 U14880 ( .A(keyinput_90), .B(n13144), .S(SI_6_), .Z(n13149) );
  XOR2_X1 U14881 ( .A(SI_4_), .B(keyinput_92), .Z(n13147) );
  XOR2_X1 U14882 ( .A(SI_5_), .B(keyinput_91), .Z(n13146) );
  XNOR2_X1 U14883 ( .A(SI_3_), .B(keyinput_93), .ZN(n13145) );
  NOR3_X1 U14884 ( .A1(n13147), .A2(n13146), .A3(n13145), .ZN(n13148) );
  OAI21_X1 U14885 ( .B1(n13150), .B2(n13149), .A(n13148), .ZN(n13153) );
  INV_X1 U14886 ( .A(keyinput_94), .ZN(n13151) );
  MUX2_X1 U14887 ( .A(keyinput_94), .B(n13151), .S(SI_2_), .Z(n13152) );
  NAND2_X1 U14888 ( .A1(n13153), .A2(n13152), .ZN(n13156) );
  OAI22_X1 U14889 ( .A1(SI_1_), .A2(keyinput_95), .B1(SI_0_), .B2(keyinput_96), 
        .ZN(n13154) );
  AOI221_X1 U14890 ( .B1(SI_1_), .B2(keyinput_95), .C1(keyinput_96), .C2(SI_0_), .A(n13154), .ZN(n13155) );
  AOI22_X1 U14891 ( .A1(n13156), .A2(n13155), .B1(P3_RD_REG_SCAN_IN), .B2(
        keyinput_97), .ZN(n13157) );
  OAI21_X1 U14892 ( .B1(keyinput_97), .B2(P3_RD_REG_SCAN_IN), .A(n13157), .ZN(
        n13160) );
  AOI22_X1 U14893 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_100), .B1(
        n13235), .B2(keyinput_101), .ZN(n13158) );
  OAI221_X1 U14894 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_100), .C1(
        n13235), .C2(keyinput_101), .A(n13158), .ZN(n13159) );
  AOI21_X1 U14895 ( .B1(n13161), .B2(n13160), .A(n13159), .ZN(n13162) );
  OAI22_X1 U14896 ( .A1(n13163), .A2(n13162), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(keyinput_104), .ZN(n13164) );
  AOI21_X1 U14897 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .A(n13164), 
        .ZN(n13172) );
  OAI22_X1 U14898 ( .A1(n13166), .A2(keyinput_103), .B1(n13250), .B2(
        keyinput_105), .ZN(n13165) );
  AOI221_X1 U14899 ( .B1(n13166), .B2(keyinput_103), .C1(keyinput_105), .C2(
        n13250), .A(n13165), .ZN(n13171) );
  AOI22_X1 U14900 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_106), .ZN(n13167) );
  OAI221_X1 U14901 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_106), .A(n13167), .ZN(n13170)
         );
  AOI22_X1 U14902 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_109), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(keyinput_108), .ZN(n13168) );
  OAI221_X1 U14903 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .C1(
        P3_REG3_REG_1__SCAN_IN), .C2(keyinput_108), .A(n13168), .ZN(n13169) );
  AOI211_X1 U14904 ( .C1(n13172), .C2(n13171), .A(n13170), .B(n13169), .ZN(
        n13173) );
  AOI221_X1 U14905 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(n13175), .C1(n13174), 
        .C2(keyinput_110), .A(n13173), .ZN(n13176) );
  AOI221_X1 U14906 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(n13178), .C1(n13177), 
        .C2(keyinput_111), .A(n13176), .ZN(n13179) );
  OAI22_X1 U14907 ( .A1(keyinput_114), .A2(n13182), .B1(n13180), .B2(n13179), 
        .ZN(n13181) );
  AOI21_X1 U14908 ( .B1(keyinput_114), .B2(n13182), .A(n13181), .ZN(n13185) );
  AOI22_X1 U14909 ( .A1(n13293), .A2(keyinput_115), .B1(n8469), .B2(
        keyinput_117), .ZN(n13183) );
  OAI221_X1 U14910 ( .B1(n13293), .B2(keyinput_115), .C1(n8469), .C2(
        keyinput_117), .A(n13183), .ZN(n13184) );
  NOR3_X1 U14911 ( .A1(n13186), .A2(n13185), .A3(n13184), .ZN(n13194) );
  AOI22_X1 U14912 ( .A1(P3_REG3_REG_20__SCAN_IN), .A2(keyinput_119), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(keyinput_123), .ZN(n13187) );
  OAI221_X1 U14913 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(
        P3_REG3_REG_2__SCAN_IN), .C2(keyinput_123), .A(n13187), .ZN(n13193) );
  AOI22_X1 U14914 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_122), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_121), .ZN(n13188) );
  OAI221_X1 U14915 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_121), .A(n13188), .ZN(n13192)
         );
  XOR2_X1 U14916 ( .A(keyinput_120), .B(n8546), .Z(n13190) );
  XNOR2_X1 U14917 ( .A(keyinput_118), .B(P3_REG3_REG_0__SCAN_IN), .ZN(n13189)
         );
  NAND2_X1 U14918 ( .A1(n13190), .A2(n13189), .ZN(n13191) );
  NOR4_X1 U14919 ( .A1(n13194), .A2(n13193), .A3(n13192), .A4(n13191), .ZN(
        n13200) );
  AOI22_X1 U14920 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_124), .B1(
        n13196), .B2(keyinput_125), .ZN(n13195) );
  OAI221_X1 U14921 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .C1(
        n13196), .C2(keyinput_125), .A(n13195), .ZN(n13199) );
  OAI22_X1 U14922 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(keyinput_127), .B1(
        keyinput_126), .B2(P3_REG3_REG_26__SCAN_IN), .ZN(n13197) );
  AOI221_X1 U14923 ( .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_127), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_126), .A(n13197), .ZN(n13198)
         );
  OAI21_X1 U14924 ( .B1(n13200), .B2(n13199), .A(n13198), .ZN(n13205) );
  OAI22_X1 U14925 ( .A1(n13334), .A2(keyinput_62), .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_63), .ZN(n13203) );
  INV_X1 U14926 ( .A(keyinput_62), .ZN(n13201) );
  NOR2_X1 U14927 ( .A1(n13201), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n13202) );
  AOI211_X1 U14928 ( .C1(keyinput_63), .C2(P3_REG3_REG_15__SCAN_IN), .A(n13203), .B(n13202), .ZN(n13204) );
  OAI211_X1 U14929 ( .C1(n13207), .C2(n13206), .A(n13205), .B(n13204), .ZN(
        n13208) );
  INV_X1 U14930 ( .A(SI_30_), .ZN(n13372) );
  NAND2_X1 U14931 ( .A1(n15507), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13209) );
  NAND2_X1 U14932 ( .A1(n13210), .A2(n13209), .ZN(n13356) );
  XNOR2_X1 U14933 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n13355) );
  INV_X1 U14934 ( .A(n13355), .ZN(n13211) );
  XNOR2_X1 U14935 ( .A(n13356), .B(n13211), .ZN(n13371) );
  INV_X1 U14936 ( .A(n13371), .ZN(n13212) );
  NAND2_X1 U14937 ( .A1(n13214), .A2(n13966), .ZN(n13220) );
  INV_X1 U14938 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n13216) );
  INV_X1 U14939 ( .A(n13757), .ZN(n13215) );
  OAI22_X1 U14940 ( .A1(n13966), .A2(n13216), .B1(n13215), .B2(n13983), .ZN(
        n13217) );
  AOI21_X1 U14941 ( .B1(n13218), .B2(n13986), .A(n13217), .ZN(n13219) );
  OAI211_X1 U14942 ( .C1(n13221), .C2(n13968), .A(n13220), .B(n13219), .ZN(
        P3_U3204) );
  XNOR2_X1 U14943 ( .A(n13223), .B(n13222), .ZN(n13224) );
  NAND2_X1 U14944 ( .A1(n13224), .A2(n13343), .ZN(n13228) );
  AOI22_X1 U14945 ( .A1(n13575), .A2(n13318), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13225) );
  OAI21_X1 U14946 ( .B1(n13787), .B2(n13335), .A(n13225), .ZN(n13226) );
  AOI21_X1 U14947 ( .B1(n13792), .B2(n13351), .A(n13226), .ZN(n13227) );
  OAI211_X1 U14948 ( .C1(n14096), .C2(n13354), .A(n13228), .B(n13227), .ZN(
        P3_U3154) );
  INV_X1 U14949 ( .A(n13987), .ZN(n14137) );
  INV_X1 U14950 ( .A(n13229), .ZN(n13305) );
  INV_X1 U14951 ( .A(n13230), .ZN(n13232) );
  NOR3_X1 U14952 ( .A1(n13305), .A2(n13232), .A3(n13231), .ZN(n13234) );
  INV_X1 U14953 ( .A(n13341), .ZN(n13233) );
  OAI21_X1 U14954 ( .B1(n13234), .B2(n13233), .A(n13343), .ZN(n13240) );
  NOR2_X1 U14955 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13235), .ZN(n13631) );
  AOI21_X1 U14956 ( .B1(n13346), .B2(n13974), .A(n13631), .ZN(n13236) );
  OAI21_X1 U14957 ( .B1(n13237), .B2(n13349), .A(n13236), .ZN(n13238) );
  AOI21_X1 U14958 ( .B1(n13982), .B2(n13351), .A(n13238), .ZN(n13239) );
  OAI211_X1 U14959 ( .C1(n14137), .C2(n13354), .A(n13240), .B(n13239), .ZN(
        P3_U3155) );
  XNOR2_X1 U14960 ( .A(n13287), .B(n13286), .ZN(n13288) );
  XNOR2_X1 U14961 ( .A(n13288), .B(n12946), .ZN(n13241) );
  NAND2_X1 U14962 ( .A1(n13241), .A2(n13343), .ZN(n13245) );
  AOI22_X1 U14963 ( .A1(n13843), .A2(n13346), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13242) );
  OAI21_X1 U14964 ( .B1(n13846), .B2(n13349), .A(n13242), .ZN(n13243) );
  AOI21_X1 U14965 ( .B1(n13847), .B2(n13351), .A(n13243), .ZN(n13244) );
  OAI211_X1 U14966 ( .C1(n13246), .C2(n13354), .A(n13245), .B(n13244), .ZN(
        P3_U3156) );
  OAI211_X1 U14967 ( .C1(n13249), .C2(n13248), .A(n13247), .B(n13343), .ZN(
        n13254) );
  NOR2_X1 U14968 ( .A1(n13250), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13744) );
  AOI21_X1 U14969 ( .B1(n13346), .B2(n13866), .A(n13744), .ZN(n13251) );
  OAI21_X1 U14970 ( .B1(n13899), .B2(n13349), .A(n13251), .ZN(n13252) );
  AOI21_X1 U14971 ( .B1(n13901), .B2(n13351), .A(n13252), .ZN(n13253) );
  OAI211_X1 U14972 ( .C1(n13903), .C2(n13354), .A(n13254), .B(n13253), .ZN(
        P3_U3159) );
  OAI211_X1 U14973 ( .C1(n13257), .C2(n13256), .A(n13255), .B(n13343), .ZN(
        n13261) );
  AOI22_X1 U14974 ( .A1(n13318), .A2(n13866), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13258) );
  OAI21_X1 U14975 ( .B1(n13846), .B2(n13335), .A(n13258), .ZN(n13259) );
  AOI21_X1 U14976 ( .B1(n13872), .B2(n13351), .A(n13259), .ZN(n13260) );
  OAI211_X1 U14977 ( .C1(n14114), .C2(n13354), .A(n13261), .B(n13260), .ZN(
        P3_U3163) );
  XNOR2_X1 U14978 ( .A(n13263), .B(n13262), .ZN(n13264) );
  NAND2_X1 U14979 ( .A1(n13264), .A2(n13343), .ZN(n13268) );
  AOI22_X1 U14980 ( .A1(n13575), .A2(n13346), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13265) );
  OAI21_X1 U14981 ( .B1(n13812), .B2(n13349), .A(n13265), .ZN(n13266) );
  AOI21_X1 U14982 ( .B1(n13818), .B2(n13351), .A(n13266), .ZN(n13267) );
  OAI211_X1 U14983 ( .C1(n14104), .C2(n13354), .A(n13268), .B(n13267), .ZN(
        P3_U3165) );
  NAND2_X1 U14984 ( .A1(n13270), .A2(n13269), .ZN(n13271) );
  XNOR2_X1 U14985 ( .A(n13272), .B(n13271), .ZN(n13273) );
  NAND2_X1 U14986 ( .A1(n13273), .A2(n13343), .ZN(n13277) );
  NAND2_X1 U14987 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n13677)
         );
  NAND2_X1 U14988 ( .A1(n13318), .A2(n13974), .ZN(n13274) );
  OAI211_X1 U14989 ( .C1(n13943), .C2(n13335), .A(n13677), .B(n13274), .ZN(
        n13275) );
  AOI21_X1 U14990 ( .B1(n13947), .B2(n13351), .A(n13275), .ZN(n13276) );
  OAI211_X1 U14991 ( .C1(n14129), .C2(n13354), .A(n13277), .B(n13276), .ZN(
        P3_U3166) );
  INV_X1 U14992 ( .A(n14123), .ZN(n13285) );
  OAI211_X1 U14993 ( .C1(n13280), .C2(n13279), .A(n13278), .B(n13343), .ZN(
        n13284) );
  NAND2_X1 U14994 ( .A1(n13318), .A2(n13958), .ZN(n13281) );
  NAND2_X1 U14995 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13699)
         );
  OAI211_X1 U14996 ( .C1(n13899), .C2(n13335), .A(n13281), .B(n13699), .ZN(
        n13282) );
  AOI21_X1 U14997 ( .B1(n13927), .B2(n13351), .A(n13282), .ZN(n13283) );
  OAI211_X1 U14998 ( .C1(n13285), .C2(n13354), .A(n13284), .B(n13283), .ZN(
        P3_U3168) );
  OAI22_X1 U14999 ( .A1(n13288), .A2(n12946), .B1(n13287), .B2(n13286), .ZN(
        n13291) );
  XNOR2_X1 U15000 ( .A(n13289), .B(n13843), .ZN(n13290) );
  XNOR2_X1 U15001 ( .A(n13291), .B(n13290), .ZN(n13292) );
  NAND2_X1 U15002 ( .A1(n13292), .A2(n13343), .ZN(n13297) );
  OAI22_X1 U15003 ( .A1(n13827), .A2(n13335), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13293), .ZN(n13295) );
  NOR2_X1 U15004 ( .A1(n13349), .A2(n13826), .ZN(n13294) );
  AOI211_X1 U15005 ( .C1(n13832), .C2(n13351), .A(n13295), .B(n13294), .ZN(
        n13296) );
  OAI211_X1 U15006 ( .C1(n14108), .C2(n13354), .A(n13297), .B(n13296), .ZN(
        P3_U3169) );
  OAI211_X1 U15007 ( .C1(n13300), .C2(n13299), .A(n13298), .B(n13343), .ZN(
        n13304) );
  AOI22_X1 U15008 ( .A1(n13346), .A2(n13857), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13301) );
  OAI21_X1 U15009 ( .B1(n13881), .B2(n13349), .A(n13301), .ZN(n13302) );
  AOI21_X1 U15010 ( .B1(n13887), .B2(n13351), .A(n13302), .ZN(n13303) );
  OAI211_X1 U15011 ( .C1(n14118), .C2(n13354), .A(n13304), .B(n13303), .ZN(
        P3_U3173) );
  AOI21_X1 U15012 ( .B1(n13307), .B2(n13306), .A(n13305), .ZN(n13315) );
  NOR2_X1 U15013 ( .A1(n14141), .A2(n13354), .ZN(n13311) );
  NOR2_X1 U15014 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8546), .ZN(n13599) );
  AOI21_X1 U15015 ( .B1(n13959), .B2(n13346), .A(n13599), .ZN(n13308) );
  OAI21_X1 U15016 ( .B1(n13309), .B2(n13349), .A(n13308), .ZN(n13310) );
  AOI211_X1 U15017 ( .C1(n13312), .C2(n13351), .A(n13311), .B(n13310), .ZN(
        n13313) );
  OAI21_X1 U15018 ( .B1(n13315), .B2(n13314), .A(n13313), .ZN(P3_U3174) );
  XNOR2_X1 U15019 ( .A(n13316), .B(n13846), .ZN(n13317) );
  NAND2_X1 U15020 ( .A1(n13317), .A2(n13343), .ZN(n13322) );
  AOI22_X1 U15021 ( .A1(n13318), .A2(n13857), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13319) );
  OAI21_X1 U15022 ( .B1(n13826), .B2(n13335), .A(n13319), .ZN(n13320) );
  AOI21_X1 U15023 ( .B1(n13860), .B2(n13351), .A(n13320), .ZN(n13321) );
  OAI211_X1 U15024 ( .C1(n13862), .C2(n13354), .A(n13322), .B(n13321), .ZN(
        P3_U3175) );
  INV_X1 U15025 ( .A(n14054), .ZN(n13330) );
  OAI211_X1 U15026 ( .C1(n13325), .C2(n13324), .A(n13323), .B(n13343), .ZN(
        n13329) );
  NAND2_X1 U15027 ( .A1(n13346), .A2(n13915), .ZN(n13326) );
  NAND2_X1 U15028 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13731)
         );
  OAI211_X1 U15029 ( .C1(n13349), .C2(n13943), .A(n13326), .B(n13731), .ZN(
        n13327) );
  AOI21_X1 U15030 ( .B1(n13908), .B2(n13351), .A(n13327), .ZN(n13328) );
  OAI211_X1 U15031 ( .C1(n13330), .C2(n13354), .A(n13329), .B(n13328), .ZN(
        P3_U3178) );
  XNOR2_X1 U15032 ( .A(n13332), .B(n13331), .ZN(n13333) );
  NAND2_X1 U15033 ( .A1(n13333), .A2(n13343), .ZN(n13339) );
  OAI22_X1 U15034 ( .A1(n12951), .A2(n13335), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13334), .ZN(n13337) );
  NOR2_X1 U15035 ( .A1(n13349), .A2(n13827), .ZN(n13336) );
  AOI211_X1 U15036 ( .C1(n13804), .C2(n13351), .A(n13337), .B(n13336), .ZN(
        n13338) );
  OAI211_X1 U15037 ( .C1(n14100), .C2(n13354), .A(n13339), .B(n13338), .ZN(
        P3_U3180) );
  AND2_X1 U15038 ( .A1(n13341), .A2(n13340), .ZN(n13345) );
  OAI211_X1 U15039 ( .C1(n13345), .C2(n13344), .A(n13343), .B(n13342), .ZN(
        n13353) );
  NAND2_X1 U15040 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(P3_U3151), .ZN(n13650)
         );
  NAND2_X1 U15041 ( .A1(n13346), .A2(n13958), .ZN(n13347) );
  OAI211_X1 U15042 ( .C1(n13349), .C2(n13348), .A(n13650), .B(n13347), .ZN(
        n13350) );
  AOI21_X1 U15043 ( .B1(n13962), .B2(n13351), .A(n13350), .ZN(n13352) );
  OAI211_X1 U15044 ( .C1(n13354), .C2(n14133), .A(n13353), .B(n13352), .ZN(
        P3_U3181) );
  NAND2_X1 U15045 ( .A1(n13356), .A2(n13355), .ZN(n13359) );
  NAND2_X1 U15046 ( .A1(n13357), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13358) );
  NAND2_X1 U15047 ( .A1(n13359), .A2(n13358), .ZN(n13361) );
  XNOR2_X1 U15048 ( .A(n14854), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n13360) );
  XNOR2_X1 U15049 ( .A(n13361), .B(n13360), .ZN(n14149) );
  NAND2_X1 U15050 ( .A1(n14149), .A2(n13370), .ZN(n13363) );
  OR2_X1 U15051 ( .A1(n12960), .A2(n14145), .ZN(n13362) );
  NAND2_X1 U15052 ( .A1(n13363), .A2(n13362), .ZN(n13555) );
  NAND2_X1 U15053 ( .A1(n13364), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13368) );
  NAND2_X1 U15054 ( .A1(n13365), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13367) );
  NAND2_X1 U15055 ( .A1(n7238), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13366) );
  OR2_X1 U15056 ( .A1(n13555), .A2(n13760), .ZN(n13519) );
  NAND2_X1 U15057 ( .A1(n13371), .A2(n13370), .ZN(n13374) );
  OR2_X1 U15058 ( .A1(n12960), .A2(n13372), .ZN(n13373) );
  NAND2_X1 U15059 ( .A1(n13374), .A2(n13373), .ZN(n13513) );
  AOI22_X1 U15060 ( .A1(n13555), .A2(n13760), .B1(n14089), .B2(n13571), .ZN(
        n13556) );
  INV_X1 U15061 ( .A(n13556), .ZN(n13518) );
  NAND2_X1 U15062 ( .A1(n13375), .A2(n7308), .ZN(n13377) );
  AND2_X1 U15063 ( .A1(n13377), .A2(n13376), .ZN(n13482) );
  NAND2_X1 U15064 ( .A1(n13482), .A2(n13474), .ZN(n13481) );
  OAI211_X1 U15065 ( .C1(n13912), .C2(n13379), .A(n13521), .B(n13378), .ZN(
        n13466) );
  NAND2_X1 U15066 ( .A1(n13586), .A2(n13380), .ZN(n13381) );
  NAND2_X1 U15067 ( .A1(n13382), .A2(n13381), .ZN(n13389) );
  NAND2_X1 U15068 ( .A1(n13389), .A2(n13383), .ZN(n13385) );
  OAI211_X1 U15069 ( .C1(n13386), .C2(n13385), .A(n13384), .B(n13395), .ZN(
        n13387) );
  NAND2_X1 U15070 ( .A1(n13387), .A2(n13393), .ZN(n13398) );
  NOR2_X1 U15071 ( .A1(n13389), .A2(n13388), .ZN(n13390) );
  OAI21_X1 U15072 ( .B1(n13391), .B2(n13390), .A(n13523), .ZN(n13394) );
  NAND3_X1 U15073 ( .A1(n13394), .A2(n13393), .A3(n13392), .ZN(n13396) );
  NAND2_X1 U15074 ( .A1(n13396), .A2(n13395), .ZN(n13397) );
  MUX2_X1 U15075 ( .A(n13398), .B(n13397), .S(n13474), .Z(n13399) );
  NAND3_X1 U15076 ( .A1(n13399), .A2(n13528), .A3(n13533), .ZN(n13410) );
  MUX2_X1 U15077 ( .A(n13401), .B(n13400), .S(n13509), .Z(n13407) );
  INV_X1 U15078 ( .A(n13533), .ZN(n13406) );
  NAND2_X1 U15079 ( .A1(n13582), .A2(n13402), .ZN(n13404) );
  MUX2_X1 U15080 ( .A(n13404), .B(n13403), .S(n13509), .Z(n13405) );
  OAI21_X1 U15081 ( .B1(n13407), .B2(n13406), .A(n13405), .ZN(n13408) );
  INV_X1 U15082 ( .A(n13408), .ZN(n13409) );
  NAND2_X1 U15083 ( .A1(n13410), .A2(n13409), .ZN(n13417) );
  MUX2_X1 U15084 ( .A(n13412), .B(n13411), .S(n13474), .Z(n13413) );
  OAI21_X1 U15085 ( .B1(n13417), .B2(n13414), .A(n13413), .ZN(n13419) );
  INV_X1 U15086 ( .A(n13415), .ZN(n13416) );
  NAND2_X1 U15087 ( .A1(n13417), .A2(n13416), .ZN(n13418) );
  AOI21_X1 U15088 ( .B1(n13419), .B2(n13418), .A(n13529), .ZN(n13425) );
  NAND2_X1 U15089 ( .A1(n13580), .A2(n13420), .ZN(n13422) );
  MUX2_X1 U15090 ( .A(n13422), .B(n13421), .S(n13509), .Z(n13423) );
  NAND2_X1 U15091 ( .A1(n13423), .A2(n13527), .ZN(n13424) );
  OR2_X1 U15092 ( .A1(n13425), .A2(n13424), .ZN(n13434) );
  NOR2_X1 U15093 ( .A1(n13522), .A2(n7854), .ZN(n13427) );
  AOI21_X1 U15094 ( .B1(n13434), .B2(n13427), .A(n7244), .ZN(n13429) );
  OAI21_X1 U15095 ( .B1(n13429), .B2(n12207), .A(n13428), .ZN(n13438) );
  INV_X1 U15096 ( .A(n13430), .ZN(n13431) );
  NOR2_X1 U15097 ( .A1(n13522), .A2(n13431), .ZN(n13433) );
  AOI21_X1 U15098 ( .B1(n13434), .B2(n13433), .A(n13432), .ZN(n13436) );
  OAI21_X1 U15099 ( .B1(n13436), .B2(n12207), .A(n13435), .ZN(n13437) );
  MUX2_X1 U15100 ( .A(n13438), .B(n13437), .S(n13509), .Z(n13442) );
  AND2_X1 U15101 ( .A1(n13448), .A2(n13439), .ZN(n13440) );
  OAI22_X1 U15102 ( .A1(n13442), .A2(n13441), .B1(n13509), .B2(n13440), .ZN(
        n13446) );
  AOI21_X1 U15103 ( .B1(n13443), .B2(n13445), .A(n13474), .ZN(n13444) );
  AOI21_X1 U15104 ( .B1(n13446), .B2(n13445), .A(n13444), .ZN(n13453) );
  OAI21_X1 U15105 ( .B1(n13448), .B2(n13474), .A(n13447), .ZN(n13452) );
  MUX2_X1 U15106 ( .A(n13450), .B(n13449), .S(n13509), .Z(n13451) );
  OAI211_X1 U15107 ( .C1(n13453), .C2(n13452), .A(n13977), .B(n13451), .ZN(
        n13457) );
  MUX2_X1 U15108 ( .A(n13455), .B(n13454), .S(n13509), .Z(n13456) );
  NAND3_X1 U15109 ( .A1(n13457), .A2(n13953), .A3(n13456), .ZN(n13461) );
  MUX2_X1 U15110 ( .A(n13459), .B(n13458), .S(n13509), .Z(n13460) );
  NAND3_X1 U15111 ( .A1(n13461), .A2(n13941), .A3(n13460), .ZN(n13464) );
  INV_X1 U15112 ( .A(n13930), .ZN(n13462) );
  NOR2_X1 U15113 ( .A1(n13912), .A2(n13462), .ZN(n13463) );
  NAND2_X1 U15114 ( .A1(n13464), .A2(n13463), .ZN(n13470) );
  OAI211_X1 U15115 ( .C1(n13470), .C2(n14129), .A(n13893), .B(n8229), .ZN(
        n13465) );
  MUX2_X1 U15116 ( .A(n13466), .B(n13465), .S(n13474), .Z(n13473) );
  MUX2_X1 U15117 ( .A(n13474), .B(n13468), .S(n13467), .Z(n13469) );
  NOR2_X1 U15118 ( .A1(n13470), .A2(n13469), .ZN(n13472) );
  MUX2_X1 U15119 ( .A(n13521), .B(n8229), .S(n13509), .Z(n13471) );
  OAI211_X1 U15120 ( .C1(n13473), .C2(n13472), .A(n13878), .B(n13471), .ZN(
        n13478) );
  MUX2_X1 U15121 ( .A(n13476), .B(n13475), .S(n13474), .Z(n13477) );
  NAND2_X1 U15122 ( .A1(n13478), .A2(n13477), .ZN(n13480) );
  NOR2_X1 U15123 ( .A1(n13855), .A2(n13867), .ZN(n13542) );
  MUX2_X1 U15124 ( .A(n13481), .B(n13480), .S(n13542), .Z(n13486) );
  INV_X1 U15125 ( .A(n13841), .ZN(n13485) );
  INV_X1 U15126 ( .A(n13482), .ZN(n13483) );
  NAND2_X1 U15127 ( .A1(n13483), .A2(n13509), .ZN(n13484) );
  NAND3_X1 U15128 ( .A1(n13486), .A2(n13485), .A3(n13484), .ZN(n13490) );
  NAND2_X1 U15129 ( .A1(n14035), .A2(n13826), .ZN(n13488) );
  MUX2_X1 U15130 ( .A(n13488), .B(n13487), .S(n13509), .Z(n13489) );
  INV_X1 U15131 ( .A(n13785), .ZN(n13501) );
  NAND2_X1 U15132 ( .A1(n13491), .A2(n13499), .ZN(n13492) );
  NAND2_X1 U15133 ( .A1(n13494), .A2(n13813), .ZN(n13495) );
  NAND2_X1 U15134 ( .A1(n13496), .A2(n13495), .ZN(n13498) );
  NAND4_X1 U15135 ( .A1(n13501), .A2(n13811), .A3(n13825), .A4(n13798), .ZN(
        n13544) );
  NAND2_X1 U15136 ( .A1(n13502), .A2(n13509), .ZN(n13503) );
  AND2_X1 U15137 ( .A1(n13503), .A2(n13765), .ZN(n13504) );
  NAND2_X1 U15138 ( .A1(n13505), .A2(n13504), .ZN(n13508) );
  NAND2_X1 U15139 ( .A1(n13508), .A2(n13506), .ZN(n13511) );
  AND2_X1 U15140 ( .A1(n13508), .A2(n13507), .ZN(n13510) );
  INV_X1 U15141 ( .A(n13571), .ZN(n13512) );
  NAND2_X1 U15142 ( .A1(n13513), .A2(n13512), .ZN(n13514) );
  NAND2_X1 U15143 ( .A1(n13519), .A2(n13514), .ZN(n13520) );
  INV_X1 U15144 ( .A(n13515), .ZN(n13516) );
  INV_X1 U15145 ( .A(n13520), .ZN(n13547) );
  NAND2_X1 U15146 ( .A1(n8229), .A2(n13521), .ZN(n13897) );
  INV_X1 U15147 ( .A(n13522), .ZN(n13525) );
  NAND3_X1 U15148 ( .A1(n13525), .A2(n13524), .A3(n13523), .ZN(n13531) );
  NAND4_X1 U15149 ( .A1(n8243), .A2(n13528), .A3(n13527), .A4(n13526), .ZN(
        n13530) );
  NOR4_X1 U15150 ( .A1(n13531), .A2(n13530), .A3(n12207), .A4(n13529), .ZN(
        n13534) );
  NAND4_X1 U15151 ( .A1(n13533), .A2(n13534), .A3(n13532), .A4(n11263), .ZN(
        n13537) );
  INV_X1 U15152 ( .A(n13992), .ZN(n13536) );
  NOR4_X1 U15153 ( .A1(n13537), .A2(n13536), .A3(n13535), .A4(n13972), .ZN(
        n13538) );
  NAND4_X1 U15154 ( .A1(n13538), .A2(n13953), .A3(n13930), .A4(n13941), .ZN(
        n13539) );
  NOR4_X1 U15155 ( .A1(n13540), .A2(n13912), .A3(n13897), .A4(n13539), .ZN(
        n13541) );
  NAND2_X1 U15156 ( .A1(n13542), .A2(n13541), .ZN(n13543) );
  NOR4_X1 U15157 ( .A1(n13771), .A2(n13544), .A3(n13841), .A4(n13543), .ZN(
        n13545) );
  NAND4_X1 U15158 ( .A1(n13547), .A2(n13556), .A3(n13546), .A4(n13545), .ZN(
        n13548) );
  INV_X1 U15159 ( .A(n13551), .ZN(n13552) );
  INV_X1 U15160 ( .A(n13760), .ZN(n13570) );
  OAI21_X1 U15161 ( .B1(n14089), .B2(n13570), .A(n13554), .ZN(n13557) );
  OAI22_X1 U15162 ( .A1(n13558), .A2(n13557), .B1(n14086), .B2(n13556), .ZN(
        n13559) );
  XNOR2_X1 U15163 ( .A(n13559), .B(n13743), .ZN(n13561) );
  NOR2_X1 U15164 ( .A1(n13561), .A2(n13560), .ZN(n13562) );
  NOR3_X1 U15165 ( .A1(n13564), .A2(n13603), .A3(n8827), .ZN(n13567) );
  OAI21_X1 U15166 ( .B1(n13568), .B2(n13565), .A(P3_B_REG_SCAN_IN), .ZN(n13566) );
  OAI22_X1 U15167 ( .A1(n13569), .A2(n13568), .B1(n13567), .B2(n13566), .ZN(
        P3_U3296) );
  MUX2_X1 U15168 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13570), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15169 ( .A(n13571), .B(P3_DATAO_REG_30__SCAN_IN), .S(n13587), .Z(
        P3_U3521) );
  MUX2_X1 U15170 ( .A(n13572), .B(P3_DATAO_REG_29__SCAN_IN), .S(n13587), .Z(
        P3_U3520) );
  MUX2_X1 U15171 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13573), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15172 ( .A(n13574), .B(P3_DATAO_REG_27__SCAN_IN), .S(n13587), .Z(
        P3_U3518) );
  MUX2_X1 U15173 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13575), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15174 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13843), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15175 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12946), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U15176 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n7492), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15177 ( .A(n13857), .B(P3_DATAO_REG_21__SCAN_IN), .S(n13587), .Z(
        P3_U3512) );
  MUX2_X1 U15178 ( .A(n13866), .B(P3_DATAO_REG_20__SCAN_IN), .S(n13587), .Z(
        P3_U3511) );
  MUX2_X1 U15179 ( .A(n13915), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13587), .Z(
        P3_U3510) );
  MUX2_X1 U15180 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13924), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15181 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13914), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15182 ( .A(n13958), .B(P3_DATAO_REG_16__SCAN_IN), .S(n13587), .Z(
        P3_U3507) );
  MUX2_X1 U15183 ( .A(n13974), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13587), .Z(
        P3_U3506) );
  MUX2_X1 U15184 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13959), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15185 ( .A(n13995), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13587), .Z(
        P3_U3504) );
  MUX2_X1 U15186 ( .A(n13576), .B(P3_DATAO_REG_12__SCAN_IN), .S(n13587), .Z(
        P3_U3503) );
  MUX2_X1 U15187 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13998), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15188 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13577), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15189 ( .A(n13578), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13587), .Z(
        P3_U3500) );
  MUX2_X1 U15190 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13579), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15191 ( .A(n13580), .B(P3_DATAO_REG_7__SCAN_IN), .S(n13587), .Z(
        P3_U3498) );
  MUX2_X1 U15192 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13581), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15193 ( .A(n13582), .B(P3_DATAO_REG_5__SCAN_IN), .S(n13587), .Z(
        P3_U3496) );
  MUX2_X1 U15194 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13583), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15195 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13584), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15196 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13585), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15197 ( .A(n13586), .B(P3_DATAO_REG_1__SCAN_IN), .S(n13587), .Z(
        P3_U3492) );
  MUX2_X1 U15198 ( .A(n13588), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13587), .Z(
        P3_U3491) );
  INV_X1 U15199 ( .A(n13624), .ZN(n13591) );
  OAI21_X1 U15200 ( .B1(n13592), .B2(n13608), .A(n13591), .ZN(n13594) );
  INV_X1 U15201 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13593) );
  AOI21_X1 U15202 ( .B1(n13594), .B2(n13593), .A(n13623), .ZN(n13615) );
  INV_X1 U15203 ( .A(n13608), .ZN(n13617) );
  INV_X1 U15204 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n13602) );
  INV_X1 U15205 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14081) );
  INV_X1 U15206 ( .A(n13604), .ZN(n13596) );
  NOR2_X1 U15207 ( .A1(n7279), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n13598) );
  OAI21_X1 U15208 ( .B1(n13632), .B2(n13598), .A(n13722), .ZN(n13601) );
  INV_X1 U15209 ( .A(n13599), .ZN(n13600) );
  OAI211_X1 U15210 ( .C1(n13602), .C2(n15853), .A(n13601), .B(n13600), .ZN(
        n13613) );
  MUX2_X1 U15211 ( .A(n13605), .B(n13604), .S(n10630), .Z(n13606) );
  NAND2_X1 U15212 ( .A1(n13607), .A2(n13606), .ZN(n13610) );
  MUX2_X1 U15213 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n10630), .Z(n13616) );
  XNOR2_X1 U15214 ( .A(n13616), .B(n13608), .ZN(n13609) );
  NAND2_X1 U15215 ( .A1(n13610), .A2(n13609), .ZN(n13611) );
  AOI21_X1 U15216 ( .B1(n13622), .B2(n13611), .A(n15843), .ZN(n13612) );
  AOI211_X1 U15217 ( .C1(n13754), .C2(n13617), .A(n13613), .B(n13612), .ZN(
        n13614) );
  OAI21_X1 U15218 ( .B1(n13615), .B2(n15872), .A(n13614), .ZN(P3_U3195) );
  INV_X1 U15219 ( .A(n13616), .ZN(n13618) );
  NAND2_X1 U15220 ( .A1(n13618), .A2(n13617), .ZN(n13619) );
  MUX2_X1 U15221 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n10630), .Z(n13653) );
  XNOR2_X1 U15222 ( .A(n13653), .B(n13656), .ZN(n13620) );
  AOI21_X1 U15223 ( .B1(n13622), .B2(n13619), .A(n13620), .ZN(n13641) );
  AND2_X1 U15224 ( .A1(n13620), .A2(n13619), .ZN(n13621) );
  NAND2_X1 U15225 ( .A1(n13622), .A2(n13621), .ZN(n13654) );
  NAND2_X1 U15226 ( .A1(n13654), .A2(n15863), .ZN(n13640) );
  INV_X1 U15227 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13625) );
  AOI22_X1 U15228 ( .A1(n13656), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n13625), 
        .B2(n13634), .ZN(n13626) );
  AOI21_X1 U15229 ( .B1(n13627), .B2(n13626), .A(n13642), .ZN(n13629) );
  AOI22_X1 U15230 ( .A1(n13754), .A2(n13656), .B1(n15521), .B2(
        P3_ADDR_REG_14__SCAN_IN), .ZN(n13628) );
  OAI21_X1 U15231 ( .B1(n15872), .B2(n13629), .A(n13628), .ZN(n13630) );
  NOR2_X1 U15232 ( .A1(n13631), .A2(n13630), .ZN(n13639) );
  INV_X1 U15233 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14076) );
  AOI22_X1 U15234 ( .A1(n13656), .A2(P3_REG1_REG_14__SCAN_IN), .B1(n14076), 
        .B2(n13634), .ZN(n13635) );
  AOI21_X1 U15235 ( .B1(n13636), .B2(n13635), .A(n13647), .ZN(n13637) );
  OR2_X1 U15236 ( .A1(n13637), .A2(n15866), .ZN(n13638) );
  OAI211_X1 U15237 ( .C1(n13641), .C2(n13640), .A(n13639), .B(n13638), .ZN(
        P3_U3196) );
  OAI21_X1 U15238 ( .B1(n13643), .B2(n13657), .A(n13671), .ZN(n13645) );
  INV_X1 U15239 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13644) );
  AOI21_X1 U15240 ( .B1(n13645), .B2(n13644), .A(n13672), .ZN(n13665) );
  NOR2_X1 U15241 ( .A1(n13656), .A2(n14076), .ZN(n13646) );
  OR2_X2 U15242 ( .A1(n13647), .A2(n13646), .ZN(n13648) );
  INV_X1 U15243 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14071) );
  AOI21_X1 U15244 ( .B1(n13649), .B2(n14071), .A(n13667), .ZN(n13662) );
  INV_X1 U15245 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n13651) );
  OAI21_X1 U15246 ( .B1(n15853), .B2(n13651), .A(n13650), .ZN(n13652) );
  AOI21_X1 U15247 ( .B1(n7458), .B2(n13754), .A(n13652), .ZN(n13661) );
  INV_X1 U15248 ( .A(n13653), .ZN(n13655) );
  MUX2_X1 U15249 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n10630), .Z(n13658) );
  NAND2_X1 U15250 ( .A1(n13659), .A2(n13658), .ZN(n13680) );
  OAI211_X1 U15251 ( .C1(n13659), .C2(n13658), .A(n13680), .B(n15863), .ZN(
        n13660) );
  OAI211_X1 U15252 ( .C1(n13662), .C2(n15866), .A(n13661), .B(n13660), .ZN(
        n13663) );
  INV_X1 U15253 ( .A(n13663), .ZN(n13664) );
  OAI21_X1 U15254 ( .B1(n13665), .B2(n15872), .A(n13664), .ZN(P3_U3197) );
  INV_X1 U15255 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n14067) );
  AOI22_X1 U15256 ( .A1(n13688), .A2(P3_REG1_REG_16__SCAN_IN), .B1(n14067), 
        .B2(n13695), .ZN(n13668) );
  AOI21_X1 U15257 ( .B1(n13669), .B2(n13668), .A(n13691), .ZN(n13690) );
  INV_X1 U15258 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13670) );
  AOI22_X1 U15259 ( .A1(n13688), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n13670), 
        .B2(n13695), .ZN(n13675) );
  INV_X1 U15260 ( .A(n13671), .ZN(n13673) );
  NOR2_X1 U15261 ( .A1(n13673), .A2(n13672), .ZN(n13674) );
  AOI21_X1 U15262 ( .B1(n13675), .B2(n13674), .A(n13694), .ZN(n13678) );
  NAND2_X1 U15263 ( .A1(n15521), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n13676) );
  OAI211_X1 U15264 ( .C1(n15872), .C2(n13678), .A(n13677), .B(n13676), .ZN(
        n13687) );
  INV_X1 U15265 ( .A(n13679), .ZN(n13681) );
  OAI21_X1 U15266 ( .B1(n7458), .B2(n13681), .A(n13680), .ZN(n13702) );
  MUX2_X1 U15267 ( .A(n13670), .B(n14067), .S(n10630), .Z(n13682) );
  NOR2_X1 U15268 ( .A1(n13682), .A2(n13688), .ZN(n13700) );
  NAND2_X1 U15269 ( .A1(n13682), .A2(n13688), .ZN(n13701) );
  INV_X1 U15270 ( .A(n13701), .ZN(n13683) );
  NOR2_X1 U15271 ( .A1(n13700), .A2(n13683), .ZN(n13684) );
  XNOR2_X1 U15272 ( .A(n13702), .B(n13684), .ZN(n13685) );
  NOR2_X1 U15273 ( .A1(n13685), .A2(n15843), .ZN(n13686) );
  AOI211_X1 U15274 ( .C1(n13754), .C2(n13688), .A(n13687), .B(n13686), .ZN(
        n13689) );
  OAI21_X1 U15275 ( .B1(n13690), .B2(n15866), .A(n13689), .ZN(P3_U3198) );
  INV_X1 U15276 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13693) );
  AOI21_X1 U15277 ( .B1(n13693), .B2(n13692), .A(n13714), .ZN(n13708) );
  INV_X1 U15278 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15810) );
  INV_X1 U15279 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13696) );
  OAI211_X1 U15280 ( .C1(n15853), .C2(n15810), .A(n13699), .B(n13698), .ZN(
        n13706) );
  MUX2_X1 U15281 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n10630), .Z(n13711) );
  XNOR2_X1 U15282 ( .A(n13711), .B(n13710), .ZN(n13703) );
  NOR2_X1 U15283 ( .A1(n13704), .A2(n13703), .ZN(n13709) );
  AOI211_X1 U15284 ( .C1(n13704), .C2(n13703), .A(n15843), .B(n13709), .ZN(
        n13705) );
  OAI21_X1 U15285 ( .B1(n13708), .B2(n15866), .A(n13707), .ZN(P3_U3199) );
  MUX2_X1 U15286 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n10630), .Z(n13713) );
  AOI21_X1 U15287 ( .B1(n13711), .B2(n13710), .A(n13709), .ZN(n13750) );
  XNOR2_X1 U15288 ( .A(n13750), .B(n13749), .ZN(n13712) );
  NOR2_X1 U15289 ( .A1(n13712), .A2(n13713), .ZN(n13748) );
  AOI21_X1 U15290 ( .B1(n13713), .B2(n13712), .A(n13748), .ZN(n13736) );
  OR2_X1 U15291 ( .A1(n13715), .A2(n13727), .ZN(n13720) );
  NAND2_X1 U15292 ( .A1(n13716), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13737) );
  INV_X1 U15293 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13717) );
  NAND2_X1 U15294 ( .A1(n13749), .A2(n13717), .ZN(n13718) );
  NAND2_X1 U15295 ( .A1(n13737), .A2(n13718), .ZN(n13719) );
  AND3_X1 U15296 ( .A1(n13721), .A2(n13720), .A3(n13719), .ZN(n13723) );
  OAI21_X1 U15297 ( .B1(n13739), .B2(n13723), .A(n13722), .ZN(n13735) );
  INV_X1 U15298 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15818) );
  INV_X1 U15299 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13910) );
  NOR2_X1 U15300 ( .A1(n13749), .A2(n13910), .ZN(n13740) );
  AOI21_X1 U15301 ( .B1(n13749), .B2(n13910), .A(n13740), .ZN(n13729) );
  NAND2_X1 U15302 ( .A1(n13729), .A2(n13728), .ZN(n13742) );
  OAI21_X1 U15303 ( .B1(n13729), .B2(n13728), .A(n13742), .ZN(n13730) );
  NAND2_X1 U15304 ( .A1(n7465), .A2(n13730), .ZN(n13732) );
  OAI211_X1 U15305 ( .C1(n15853), .C2(n15818), .A(n13732), .B(n13731), .ZN(
        n13733) );
  AOI21_X1 U15306 ( .B1(n13749), .B2(n13754), .A(n13733), .ZN(n13734) );
  OAI211_X1 U15307 ( .C1(n13736), .C2(n15843), .A(n13735), .B(n13734), .ZN(
        P3_U3200) );
  XNOR2_X1 U15308 ( .A(n13743), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13746) );
  INV_X1 U15309 ( .A(n13737), .ZN(n13738) );
  INV_X1 U15310 ( .A(n13740), .ZN(n13741) );
  XNOR2_X1 U15311 ( .A(n13743), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13747) );
  AOI21_X1 U15312 ( .B1(n15521), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n13744), 
        .ZN(n13745) );
  MUX2_X1 U15313 ( .A(n13747), .B(n13746), .S(n10630), .Z(n13751) );
  NOR2_X1 U15314 ( .A1(n13752), .A2(n15843), .ZN(n13753) );
  OAI21_X1 U15315 ( .B1(n13756), .B2(n15866), .A(n7291), .ZN(P3_U3201) );
  NAND2_X1 U15316 ( .A1(n13757), .A2(n14004), .ZN(n13761) );
  INV_X1 U15317 ( .A(n13758), .ZN(n13759) );
  NAND3_X1 U15318 ( .A1(n13966), .A2(n13761), .A3(n14084), .ZN(n13763) );
  OAI21_X1 U15319 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n13966), .A(n13763), 
        .ZN(n13762) );
  OAI21_X1 U15320 ( .B1(n14086), .B2(n14006), .A(n13762), .ZN(P3_U3202) );
  OAI21_X1 U15321 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n13966), .A(n13763), 
        .ZN(n13764) );
  OAI21_X1 U15322 ( .B1(n14089), .B2(n14006), .A(n13764), .ZN(P3_U3203) );
  AOI21_X1 U15323 ( .B1(n13766), .B2(n13765), .A(n14002), .ZN(n13769) );
  OAI22_X1 U15324 ( .A1(n13767), .A2(n13944), .B1(n12951), .B2(n13946), .ZN(
        n13768) );
  INV_X1 U15325 ( .A(n13783), .ZN(n13773) );
  OAI21_X1 U15326 ( .B1(n13773), .B2(n13772), .A(n13771), .ZN(n13775) );
  NAND2_X1 U15327 ( .A1(n13775), .A2(n13774), .ZN(n14015) );
  INV_X1 U15328 ( .A(n14015), .ZN(n13779) );
  AOI22_X1 U15329 ( .A1(n13963), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n14004), 
        .B2(n13776), .ZN(n13777) );
  OAI21_X1 U15330 ( .B1(n14017), .B2(n14006), .A(n13777), .ZN(n13778) );
  AOI21_X1 U15331 ( .B1(n13779), .B2(n13981), .A(n13778), .ZN(n13780) );
  OAI21_X1 U15332 ( .B1(n14014), .B2(n13963), .A(n13780), .ZN(P3_U3205) );
  NAND2_X1 U15333 ( .A1(n13781), .A2(n13785), .ZN(n13782) );
  OAI21_X1 U15334 ( .B1(n13786), .B2(n13785), .A(n13784), .ZN(n13789) );
  OAI22_X1 U15335 ( .A1(n13813), .A2(n13946), .B1(n13787), .B2(n13944), .ZN(
        n13788) );
  INV_X1 U15336 ( .A(n14018), .ZN(n13796) );
  AOI22_X1 U15337 ( .A1(n13963), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n14004), 
        .B2(n13792), .ZN(n13793) );
  OAI21_X1 U15338 ( .B1(n14096), .B2(n14006), .A(n13793), .ZN(n13794) );
  AOI21_X1 U15339 ( .B1(n14019), .B2(n14008), .A(n13794), .ZN(n13795) );
  OAI21_X1 U15340 ( .B1(n13796), .B2(n13963), .A(n13795), .ZN(P3_U3206) );
  XNOR2_X1 U15341 ( .A(n13797), .B(n13798), .ZN(n13803) );
  XNOR2_X1 U15342 ( .A(n13799), .B(n13798), .ZN(n13801) );
  OAI22_X1 U15343 ( .A1(n13827), .A2(n13946), .B1(n12951), .B2(n13944), .ZN(
        n13800) );
  AOI21_X1 U15344 ( .B1(n13801), .B2(n13970), .A(n13800), .ZN(n13802) );
  OAI21_X1 U15345 ( .B1(n13885), .B2(n13803), .A(n13802), .ZN(n14022) );
  INV_X1 U15346 ( .A(n14022), .ZN(n13808) );
  INV_X1 U15347 ( .A(n13803), .ZN(n14023) );
  AOI22_X1 U15348 ( .A1(n13963), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n14004), 
        .B2(n13804), .ZN(n13805) );
  OAI21_X1 U15349 ( .B1(n14100), .B2(n14006), .A(n13805), .ZN(n13806) );
  AOI21_X1 U15350 ( .B1(n14023), .B2(n14008), .A(n13806), .ZN(n13807) );
  OAI21_X1 U15351 ( .B1(n13808), .B2(n13963), .A(n13807), .ZN(P3_U3207) );
  XNOR2_X1 U15352 ( .A(n13809), .B(n13811), .ZN(n13817) );
  XOR2_X1 U15353 ( .A(n13811), .B(n7225), .Z(n13815) );
  OAI22_X1 U15354 ( .A1(n13813), .A2(n13944), .B1(n13812), .B2(n13946), .ZN(
        n13814) );
  AOI21_X1 U15355 ( .B1(n13815), .B2(n13970), .A(n13814), .ZN(n13816) );
  OAI21_X1 U15356 ( .B1(n13885), .B2(n13817), .A(n13816), .ZN(n14026) );
  INV_X1 U15357 ( .A(n14026), .ZN(n13822) );
  INV_X1 U15358 ( .A(n13817), .ZN(n14027) );
  AOI22_X1 U15359 ( .A1(n13963), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n14004), 
        .B2(n13818), .ZN(n13819) );
  OAI21_X1 U15360 ( .B1(n14104), .B2(n14006), .A(n13819), .ZN(n13820) );
  AOI21_X1 U15361 ( .B1(n14027), .B2(n14008), .A(n13820), .ZN(n13821) );
  OAI21_X1 U15362 ( .B1(n13822), .B2(n13963), .A(n13821), .ZN(P3_U3208) );
  XNOR2_X1 U15363 ( .A(n13823), .B(n13825), .ZN(n13831) );
  XNOR2_X1 U15364 ( .A(n13824), .B(n13825), .ZN(n13829) );
  OAI22_X1 U15365 ( .A1(n13827), .A2(n13944), .B1(n13826), .B2(n13946), .ZN(
        n13828) );
  AOI21_X1 U15366 ( .B1(n13829), .B2(n13970), .A(n13828), .ZN(n13830) );
  OAI21_X1 U15367 ( .B1(n13885), .B2(n13831), .A(n13830), .ZN(n14030) );
  INV_X1 U15368 ( .A(n14030), .ZN(n13836) );
  INV_X1 U15369 ( .A(n13831), .ZN(n14031) );
  AOI22_X1 U15370 ( .A1(n13963), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n14004), 
        .B2(n13832), .ZN(n13833) );
  OAI21_X1 U15371 ( .B1(n14108), .B2(n14006), .A(n13833), .ZN(n13834) );
  AOI21_X1 U15372 ( .B1(n14031), .B2(n14008), .A(n13834), .ZN(n13835) );
  OAI21_X1 U15373 ( .B1(n13836), .B2(n13963), .A(n13835), .ZN(P3_U3209) );
  NAND2_X1 U15374 ( .A1(n13837), .A2(n13841), .ZN(n13838) );
  NAND2_X1 U15375 ( .A1(n13839), .A2(n13838), .ZN(n14037) );
  OAI211_X1 U15376 ( .C1(n13842), .C2(n13841), .A(n13840), .B(n13970), .ZN(
        n13845) );
  NAND2_X1 U15377 ( .A1(n13843), .A2(n13996), .ZN(n13844) );
  OAI211_X1 U15378 ( .C1(n13846), .C2(n13946), .A(n13845), .B(n13844), .ZN(
        n14034) );
  NAND2_X1 U15379 ( .A1(n14034), .A2(n13966), .ZN(n13852) );
  INV_X1 U15380 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n13849) );
  INV_X1 U15381 ( .A(n13847), .ZN(n13848) );
  OAI22_X1 U15382 ( .A1(n13966), .A2(n13849), .B1(n13848), .B2(n13983), .ZN(
        n13850) );
  AOI21_X1 U15383 ( .B1(n14035), .B2(n13986), .A(n13850), .ZN(n13851) );
  OAI211_X1 U15384 ( .C1(n13968), .C2(n14037), .A(n13852), .B(n13851), .ZN(
        P3_U3210) );
  XNOR2_X1 U15385 ( .A(n13853), .B(n13855), .ZN(n14041) );
  OAI211_X1 U15386 ( .C1(n7226), .C2(n13855), .A(n13854), .B(n13970), .ZN(
        n13859) );
  AOI22_X1 U15387 ( .A1(n12946), .A2(n13996), .B1(n13997), .B2(n13857), .ZN(
        n13858) );
  NAND2_X1 U15388 ( .A1(n13859), .A2(n13858), .ZN(n14038) );
  AOI22_X1 U15389 ( .A1(n13963), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n14004), 
        .B2(n13860), .ZN(n13861) );
  OAI21_X1 U15390 ( .B1(n13862), .B2(n14006), .A(n13861), .ZN(n13863) );
  AOI21_X1 U15391 ( .B1(n14038), .B2(n13966), .A(n13863), .ZN(n13864) );
  OAI21_X1 U15392 ( .B1(n13968), .B2(n14041), .A(n13864), .ZN(P3_U3211) );
  XOR2_X1 U15393 ( .A(n13867), .B(n13865), .Z(n13871) );
  AOI22_X1 U15394 ( .A1(n7492), .A2(n13996), .B1(n13997), .B2(n13866), .ZN(
        n13870) );
  XNOR2_X1 U15395 ( .A(n13868), .B(n13867), .ZN(n14043) );
  NAND2_X1 U15396 ( .A1(n14043), .A2(n13994), .ZN(n13869) );
  OAI211_X1 U15397 ( .C1(n13871), .C2(n14002), .A(n13870), .B(n13869), .ZN(
        n14042) );
  INV_X1 U15398 ( .A(n14042), .ZN(n13876) );
  AOI22_X1 U15399 ( .A1(n13963), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n14004), 
        .B2(n13872), .ZN(n13873) );
  OAI21_X1 U15400 ( .B1(n14114), .B2(n14006), .A(n13873), .ZN(n13874) );
  AOI21_X1 U15401 ( .B1(n14043), .B2(n14008), .A(n13874), .ZN(n13875) );
  OAI21_X1 U15402 ( .B1(n13876), .B2(n13963), .A(n13875), .ZN(P3_U3212) );
  XNOR2_X1 U15403 ( .A(n13877), .B(n13878), .ZN(n13886) );
  XNOR2_X1 U15404 ( .A(n13879), .B(n13878), .ZN(n13883) );
  OAI22_X1 U15405 ( .A1(n13881), .A2(n13946), .B1(n13880), .B2(n13944), .ZN(
        n13882) );
  AOI21_X1 U15406 ( .B1(n13883), .B2(n13970), .A(n13882), .ZN(n13884) );
  OAI21_X1 U15407 ( .B1(n13885), .B2(n13886), .A(n13884), .ZN(n14046) );
  INV_X1 U15408 ( .A(n14046), .ZN(n13891) );
  INV_X1 U15409 ( .A(n13886), .ZN(n14047) );
  AOI22_X1 U15410 ( .A1(n13963), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n14004), 
        .B2(n13887), .ZN(n13888) );
  OAI21_X1 U15411 ( .B1(n14118), .B2(n14006), .A(n13888), .ZN(n13889) );
  AOI21_X1 U15412 ( .B1(n14047), .B2(n14008), .A(n13889), .ZN(n13890) );
  OAI21_X1 U15413 ( .B1(n13891), .B2(n13963), .A(n13890), .ZN(P3_U3213) );
  OR2_X1 U15414 ( .A1(n13933), .A2(n13892), .ZN(n13894) );
  NAND2_X1 U15415 ( .A1(n13894), .A2(n13893), .ZN(n13895) );
  XNOR2_X1 U15416 ( .A(n13895), .B(n13897), .ZN(n14053) );
  XOR2_X1 U15417 ( .A(n13896), .B(n13897), .Z(n13898) );
  OAI222_X1 U15418 ( .A1(n13944), .A2(n13900), .B1(n13946), .B2(n13899), .C1(
        n14002), .C2(n13898), .ZN(n14050) );
  AOI22_X1 U15419 ( .A1(n13963), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n14004), 
        .B2(n13901), .ZN(n13902) );
  OAI21_X1 U15420 ( .B1(n13903), .B2(n14006), .A(n13902), .ZN(n13904) );
  AOI21_X1 U15421 ( .B1(n14050), .B2(n13966), .A(n13904), .ZN(n13905) );
  OAI21_X1 U15422 ( .B1(n13968), .B2(n14053), .A(n13905), .ZN(P3_U3214) );
  NAND2_X1 U15423 ( .A1(n13933), .A2(n13906), .ZN(n13907) );
  XNOR2_X1 U15424 ( .A(n13907), .B(n13912), .ZN(n14057) );
  INV_X1 U15425 ( .A(n13908), .ZN(n13909) );
  OAI22_X1 U15426 ( .A1(n13966), .A2(n13910), .B1(n13909), .B2(n13983), .ZN(
        n13918) );
  OAI21_X1 U15427 ( .B1(n7222), .B2(n13912), .A(n13911), .ZN(n13916) );
  AOI222_X1 U15428 ( .A1(n13970), .A2(n13916), .B1(n13915), .B2(n13996), .C1(
        n13914), .C2(n13997), .ZN(n14056) );
  NOR2_X1 U15429 ( .A1(n14056), .A2(n13963), .ZN(n13917) );
  AOI211_X1 U15430 ( .C1(n13986), .C2(n14054), .A(n13918), .B(n13917), .ZN(
        n13919) );
  OAI21_X1 U15431 ( .B1(n13968), .B2(n14057), .A(n13919), .ZN(P3_U3215) );
  NAND2_X1 U15432 ( .A1(n13920), .A2(n13930), .ZN(n13921) );
  NAND2_X1 U15433 ( .A1(n13921), .A2(n13970), .ZN(n13922) );
  OR2_X1 U15434 ( .A1(n13923), .A2(n13922), .ZN(n13926) );
  AOI22_X1 U15435 ( .A1(n13924), .A2(n13996), .B1(n13997), .B2(n13958), .ZN(
        n13925) );
  INV_X1 U15436 ( .A(n13927), .ZN(n13928) );
  OAI22_X1 U15437 ( .A1(n13966), .A2(n13696), .B1(n13928), .B2(n13983), .ZN(
        n13929) );
  AOI21_X1 U15438 ( .B1(n14123), .B2(n13986), .A(n13929), .ZN(n13935) );
  OR2_X1 U15439 ( .A1(n13931), .A2(n13930), .ZN(n13932) );
  NAND2_X1 U15440 ( .A1(n13933), .A2(n13932), .ZN(n14059) );
  NAND2_X1 U15441 ( .A1(n14059), .A2(n13981), .ZN(n13934) );
  OAI211_X1 U15442 ( .C1(n14061), .C2(n13963), .A(n13935), .B(n13934), .ZN(
        P3_U3216) );
  OAI21_X1 U15443 ( .B1(n13937), .B2(n13941), .A(n13936), .ZN(n14066) );
  INV_X1 U15444 ( .A(n14066), .ZN(n13951) );
  INV_X1 U15445 ( .A(n13938), .ZN(n13939) );
  AOI21_X1 U15446 ( .B1(n13941), .B2(n13940), .A(n13939), .ZN(n13942) );
  OAI222_X1 U15447 ( .A1(n13946), .A2(n13945), .B1(n13944), .B2(n13943), .C1(
        n14002), .C2(n13942), .ZN(n14065) );
  AOI22_X1 U15448 ( .A1(n13963), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n14004), 
        .B2(n13947), .ZN(n13948) );
  OAI21_X1 U15449 ( .B1(n14129), .B2(n14006), .A(n13948), .ZN(n13949) );
  AOI21_X1 U15450 ( .B1(n14065), .B2(n13966), .A(n13949), .ZN(n13950) );
  OAI21_X1 U15451 ( .B1(n13968), .B2(n13951), .A(n13950), .ZN(P3_U3217) );
  OAI21_X1 U15452 ( .B1(n13954), .B2(n13953), .A(n13952), .ZN(n14070) );
  INV_X1 U15453 ( .A(n14070), .ZN(n13969) );
  OAI211_X1 U15454 ( .C1(n13957), .C2(n13956), .A(n13955), .B(n13970), .ZN(
        n13961) );
  AOI22_X1 U15455 ( .A1(n13959), .A2(n13997), .B1(n13996), .B2(n13958), .ZN(
        n13960) );
  NAND2_X1 U15456 ( .A1(n13961), .A2(n13960), .ZN(n14069) );
  AOI22_X1 U15457 ( .A1(n13963), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n14004), 
        .B2(n13962), .ZN(n13964) );
  OAI21_X1 U15458 ( .B1(n14133), .B2(n14006), .A(n13964), .ZN(n13965) );
  AOI21_X1 U15459 ( .B1(n14069), .B2(n13966), .A(n13965), .ZN(n13967) );
  OAI21_X1 U15460 ( .B1(n13969), .B2(n13968), .A(n13967), .ZN(P3_U3218) );
  OAI211_X1 U15461 ( .C1(n13973), .C2(n13972), .A(n13971), .B(n13970), .ZN(
        n13976) );
  AOI22_X1 U15462 ( .A1(n13997), .A2(n13995), .B1(n13974), .B2(n13996), .ZN(
        n13975) );
  AND2_X1 U15463 ( .A1(n13976), .A2(n13975), .ZN(n14074) );
  OR2_X1 U15464 ( .A1(n13978), .A2(n13977), .ZN(n13979) );
  NAND2_X1 U15465 ( .A1(n13980), .A2(n13979), .ZN(n14073) );
  NAND2_X1 U15466 ( .A1(n14073), .A2(n13981), .ZN(n13989) );
  INV_X1 U15467 ( .A(n13982), .ZN(n13984) );
  OAI22_X1 U15468 ( .A1(n13966), .A2(n13625), .B1(n13984), .B2(n13983), .ZN(
        n13985) );
  AOI21_X1 U15469 ( .B1(n13987), .B2(n13986), .A(n13985), .ZN(n13988) );
  OAI211_X1 U15470 ( .C1(n14074), .C2(n13963), .A(n13989), .B(n13988), .ZN(
        P3_U3219) );
  XNOR2_X1 U15471 ( .A(n7224), .B(n13992), .ZN(n14001) );
  OAI21_X1 U15472 ( .B1(n13993), .B2(n13992), .A(n13991), .ZN(n16058) );
  NAND2_X1 U15473 ( .A1(n16058), .A2(n13994), .ZN(n14000) );
  AOI22_X1 U15474 ( .A1(n13998), .A2(n13997), .B1(n13996), .B2(n13995), .ZN(
        n13999) );
  OAI211_X1 U15475 ( .C1(n14002), .C2(n14001), .A(n14000), .B(n13999), .ZN(
        n16056) );
  INV_X1 U15476 ( .A(n16056), .ZN(n14010) );
  AOI22_X1 U15477 ( .A1(n13963), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n14004), 
        .B2(n14003), .ZN(n14005) );
  OAI21_X1 U15478 ( .B1(n16055), .B2(n14006), .A(n14005), .ZN(n14007) );
  AOI21_X1 U15479 ( .B1(n16058), .B2(n14008), .A(n14007), .ZN(n14009) );
  OAI21_X1 U15480 ( .B1(n14010), .B2(n13963), .A(n14009), .ZN(P3_U3221) );
  NOR2_X1 U15481 ( .A1(n12991), .A2(n14084), .ZN(n14012) );
  AOI21_X1 U15482 ( .B1(n12991), .B2(P3_REG1_REG_31__SCAN_IN), .A(n14012), 
        .ZN(n14011) );
  OAI21_X1 U15483 ( .B1(n14086), .B2(n14083), .A(n14011), .ZN(P3_U3490) );
  AOI21_X1 U15484 ( .B1(n12991), .B2(P3_REG1_REG_30__SCAN_IN), .A(n14012), 
        .ZN(n14013) );
  OAI21_X1 U15485 ( .B1(n14089), .B2(n14083), .A(n14013), .ZN(P3_U3489) );
  OAI21_X1 U15486 ( .B1(n14058), .B2(n14015), .A(n14014), .ZN(n14090) );
  OAI21_X1 U15487 ( .B1(n14017), .B2(n14083), .A(n14016), .ZN(P3_U3487) );
  INV_X1 U15488 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n14020) );
  MUX2_X1 U15489 ( .A(n14020), .B(n14093), .S(n16061), .Z(n14021) );
  INV_X1 U15490 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n14024) );
  AOI21_X1 U15491 ( .B1(n16059), .B2(n14023), .A(n14022), .ZN(n14097) );
  MUX2_X1 U15492 ( .A(n14024), .B(n14097), .S(n16061), .Z(n14025) );
  OAI21_X1 U15493 ( .B1(n14100), .B2(n14083), .A(n14025), .ZN(P3_U3485) );
  INV_X1 U15494 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n14028) );
  AOI21_X1 U15495 ( .B1(n16059), .B2(n14027), .A(n14026), .ZN(n14101) );
  MUX2_X1 U15496 ( .A(n14028), .B(n14101), .S(n16061), .Z(n14029) );
  OAI21_X1 U15497 ( .B1(n14104), .B2(n14083), .A(n14029), .ZN(P3_U3484) );
  INV_X1 U15498 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n14032) );
  AOI21_X1 U15499 ( .B1(n16059), .B2(n14031), .A(n14030), .ZN(n14105) );
  MUX2_X1 U15500 ( .A(n14032), .B(n14105), .S(n16061), .Z(n14033) );
  OAI21_X1 U15501 ( .B1(n14108), .B2(n14083), .A(n14033), .ZN(P3_U3483) );
  AOI21_X1 U15502 ( .B1(n15940), .B2(n14035), .A(n14034), .ZN(n14036) );
  OAI21_X1 U15503 ( .B1(n14058), .B2(n14037), .A(n14036), .ZN(n14109) );
  MUX2_X1 U15504 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n14109), .S(n16061), .Z(
        P3_U3482) );
  AOI21_X1 U15505 ( .B1(n15940), .B2(n14039), .A(n14038), .ZN(n14040) );
  OAI21_X1 U15506 ( .B1(n14058), .B2(n14041), .A(n14040), .ZN(n14110) );
  MUX2_X1 U15507 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n14110), .S(n16061), .Z(
        P3_U3481) );
  INV_X1 U15508 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n14044) );
  AOI21_X1 U15509 ( .B1(n16059), .B2(n14043), .A(n14042), .ZN(n14111) );
  MUX2_X1 U15510 ( .A(n14044), .B(n14111), .S(n16061), .Z(n14045) );
  OAI21_X1 U15511 ( .B1(n14114), .B2(n14083), .A(n14045), .ZN(P3_U3480) );
  INV_X1 U15512 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n14048) );
  AOI21_X1 U15513 ( .B1(n16059), .B2(n14047), .A(n14046), .ZN(n14115) );
  MUX2_X1 U15514 ( .A(n14048), .B(n14115), .S(n16061), .Z(n14049) );
  OAI21_X1 U15515 ( .B1(n14118), .B2(n14083), .A(n14049), .ZN(P3_U3479) );
  AOI21_X1 U15516 ( .B1(n15940), .B2(n14051), .A(n14050), .ZN(n14052) );
  OAI21_X1 U15517 ( .B1(n14058), .B2(n14053), .A(n14052), .ZN(n14119) );
  MUX2_X1 U15518 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n14119), .S(n16061), .Z(
        P3_U3478) );
  NAND2_X1 U15519 ( .A1(n14054), .A2(n15940), .ZN(n14055) );
  OAI211_X1 U15520 ( .C1(n14058), .C2(n14057), .A(n14056), .B(n14055), .ZN(
        n14120) );
  MUX2_X1 U15521 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n14120), .S(n16061), .Z(
        P3_U3477) );
  NAND2_X1 U15522 ( .A1(n14059), .A2(n14080), .ZN(n14060) );
  NAND2_X1 U15523 ( .A1(n14061), .A2(n14060), .ZN(n14121) );
  MUX2_X1 U15524 ( .A(n14121), .B(P3_REG1_REG_17__SCAN_IN), .S(n12991), .Z(
        n14062) );
  AOI21_X1 U15525 ( .B1(n14063), .B2(n14123), .A(n14062), .ZN(n14064) );
  INV_X1 U15526 ( .A(n14064), .ZN(P3_U3476) );
  AOI21_X1 U15527 ( .B1(n14080), .B2(n14066), .A(n14065), .ZN(n14126) );
  MUX2_X1 U15528 ( .A(n14067), .B(n14126), .S(n16061), .Z(n14068) );
  OAI21_X1 U15529 ( .B1(n14129), .B2(n14083), .A(n14068), .ZN(P3_U3475) );
  AOI21_X1 U15530 ( .B1(n14070), .B2(n14080), .A(n14069), .ZN(n14130) );
  MUX2_X1 U15531 ( .A(n14071), .B(n14130), .S(n16061), .Z(n14072) );
  OAI21_X1 U15532 ( .B1(n14083), .B2(n14133), .A(n14072), .ZN(P3_U3474) );
  NAND2_X1 U15533 ( .A1(n14073), .A2(n14080), .ZN(n14075) );
  MUX2_X1 U15534 ( .A(n14076), .B(n14134), .S(n16061), .Z(n14077) );
  OAI21_X1 U15535 ( .B1(n14137), .B2(n14083), .A(n14077), .ZN(P3_U3473) );
  AOI21_X1 U15536 ( .B1(n14080), .B2(n14079), .A(n14078), .ZN(n14138) );
  MUX2_X1 U15537 ( .A(n14081), .B(n14138), .S(n16061), .Z(n14082) );
  OAI21_X1 U15538 ( .B1(n14083), .B2(n14141), .A(n14082), .ZN(P3_U3472) );
  NOR2_X1 U15539 ( .A1(n14084), .A2(n16062), .ZN(n14087) );
  AOI21_X1 U15540 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n16062), .A(n14087), 
        .ZN(n14085) );
  OAI21_X1 U15541 ( .B1(n14086), .B2(n14142), .A(n14085), .ZN(P3_U3458) );
  AOI21_X1 U15542 ( .B1(n16062), .B2(P3_REG0_REG_30__SCAN_IN), .A(n14087), 
        .ZN(n14088) );
  OAI21_X1 U15543 ( .B1(n14089), .B2(n14142), .A(n14088), .ZN(P3_U3457) );
  INV_X1 U15544 ( .A(n14092), .ZN(P3_U3455) );
  INV_X1 U15545 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n14094) );
  MUX2_X1 U15546 ( .A(n14094), .B(n14093), .S(n16065), .Z(n14095) );
  INV_X1 U15547 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n14098) );
  MUX2_X1 U15548 ( .A(n14098), .B(n14097), .S(n16065), .Z(n14099) );
  OAI21_X1 U15549 ( .B1(n14100), .B2(n14142), .A(n14099), .ZN(P3_U3453) );
  INV_X1 U15550 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n14102) );
  MUX2_X1 U15551 ( .A(n14102), .B(n14101), .S(n16065), .Z(n14103) );
  OAI21_X1 U15552 ( .B1(n14104), .B2(n14142), .A(n14103), .ZN(P3_U3452) );
  INV_X1 U15553 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n14106) );
  MUX2_X1 U15554 ( .A(n14106), .B(n14105), .S(n16065), .Z(n14107) );
  OAI21_X1 U15555 ( .B1(n14108), .B2(n14142), .A(n14107), .ZN(P3_U3451) );
  MUX2_X1 U15556 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n14109), .S(n16065), .Z(
        P3_U3450) );
  MUX2_X1 U15557 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n14110), .S(n16065), .Z(
        P3_U3449) );
  INV_X1 U15558 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n14112) );
  MUX2_X1 U15559 ( .A(n14112), .B(n14111), .S(n16065), .Z(n14113) );
  OAI21_X1 U15560 ( .B1(n14114), .B2(n14142), .A(n14113), .ZN(P3_U3448) );
  INV_X1 U15561 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n14116) );
  MUX2_X1 U15562 ( .A(n14116), .B(n14115), .S(n16065), .Z(n14117) );
  OAI21_X1 U15563 ( .B1(n14118), .B2(n14142), .A(n14117), .ZN(P3_U3447) );
  MUX2_X1 U15564 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n14119), .S(n16065), .Z(
        P3_U3446) );
  MUX2_X1 U15565 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n14120), .S(n16065), .Z(
        P3_U3444) );
  MUX2_X1 U15566 ( .A(n14121), .B(P3_REG0_REG_17__SCAN_IN), .S(n16062), .Z(
        n14122) );
  AOI21_X1 U15567 ( .B1(n14124), .B2(n14123), .A(n14122), .ZN(n14125) );
  INV_X1 U15568 ( .A(n14125), .ZN(P3_U3441) );
  INV_X1 U15569 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n14127) );
  MUX2_X1 U15570 ( .A(n14127), .B(n14126), .S(n16065), .Z(n14128) );
  OAI21_X1 U15571 ( .B1(n14129), .B2(n14142), .A(n14128), .ZN(P3_U3438) );
  INV_X1 U15572 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n14131) );
  MUX2_X1 U15573 ( .A(n14131), .B(n14130), .S(n16065), .Z(n14132) );
  OAI21_X1 U15574 ( .B1(n14142), .B2(n14133), .A(n14132), .ZN(P3_U3435) );
  INV_X1 U15575 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14135) );
  MUX2_X1 U15576 ( .A(n14135), .B(n14134), .S(n16065), .Z(n14136) );
  OAI21_X1 U15577 ( .B1(n14137), .B2(n14142), .A(n14136), .ZN(P3_U3432) );
  INV_X1 U15578 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14139) );
  MUX2_X1 U15579 ( .A(n14139), .B(n14138), .S(n16065), .Z(n14140) );
  OAI21_X1 U15580 ( .B1(n14142), .B2(n14141), .A(n14140), .ZN(P3_U3429) );
  MUX2_X1 U15581 ( .A(P3_D_REG_0__SCAN_IN), .B(n7567), .S(n14143), .Z(P3_U3376) );
  INV_X1 U15582 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n14144) );
  NAND3_X1 U15583 ( .A1(n14144), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n14146) );
  OAI22_X1 U15584 ( .A1(n8268), .A2(n14146), .B1(n14145), .B2(n14155), .ZN(
        n14147) );
  AOI21_X1 U15585 ( .B1(n14149), .B2(n14148), .A(n14147), .ZN(n14150) );
  INV_X1 U15586 ( .A(n14150), .ZN(P3_U3264) );
  INV_X1 U15587 ( .A(n14154), .ZN(n14157) );
  INV_X1 U15588 ( .A(n14563), .ZN(n14748) );
  NOR2_X1 U15589 ( .A1(n14484), .A2(n14716), .ZN(n14199) );
  XNOR2_X1 U15590 ( .A(n14573), .B(n10662), .ZN(n14197) );
  XNOR2_X1 U15591 ( .A(n14784), .B(n14188), .ZN(n14182) );
  NAND2_X1 U15592 ( .A1(n14507), .A2(n14633), .ZN(n14181) );
  NAND2_X1 U15593 ( .A1(n14466), .A2(n14633), .ZN(n14162) );
  INV_X1 U15594 ( .A(n14162), .ZN(n14166) );
  XNOR2_X1 U15595 ( .A(n14723), .B(n10662), .ZN(n14165) );
  INV_X1 U15596 ( .A(n14281), .ZN(n14161) );
  INV_X1 U15597 ( .A(n14159), .ZN(n14160) );
  NOR2_X1 U15598 ( .A1(n14161), .A2(n14160), .ZN(n14163) );
  XNOR2_X1 U15599 ( .A(n14165), .B(n14162), .ZN(n14280) );
  XNOR2_X1 U15600 ( .A(n14698), .B(n14229), .ZN(n14217) );
  AND2_X1 U15601 ( .A1(n14497), .A2(n14633), .ZN(n14167) );
  NAND2_X1 U15602 ( .A1(n14217), .A2(n14167), .ZN(n14168) );
  OAI21_X1 U15603 ( .B1(n14217), .B2(n14167), .A(n14168), .ZN(n14325) );
  INV_X1 U15604 ( .A(n14168), .ZN(n14173) );
  XNOR2_X1 U15605 ( .A(n14686), .B(n14229), .ZN(n14169) );
  AND2_X1 U15606 ( .A1(n14470), .A2(n14633), .ZN(n14170) );
  NAND2_X1 U15607 ( .A1(n14169), .A2(n14170), .ZN(n14178) );
  INV_X1 U15608 ( .A(n14169), .ZN(n14297) );
  INV_X1 U15609 ( .A(n14170), .ZN(n14171) );
  NAND2_X1 U15610 ( .A1(n14297), .A2(n14171), .ZN(n14172) );
  XNOR2_X1 U15611 ( .A(n14789), .B(n10662), .ZN(n14174) );
  AND2_X1 U15612 ( .A1(n14474), .A2(n14633), .ZN(n14175) );
  NAND2_X1 U15613 ( .A1(n14174), .A2(n14175), .ZN(n14179) );
  INV_X1 U15614 ( .A(n14174), .ZN(n14241) );
  INV_X1 U15615 ( .A(n14175), .ZN(n14176) );
  NAND2_X1 U15616 ( .A1(n14241), .A2(n14176), .ZN(n14177) );
  NAND2_X1 U15617 ( .A1(n14179), .A2(n14177), .ZN(n14298) );
  INV_X1 U15618 ( .A(n14179), .ZN(n14180) );
  XNOR2_X1 U15619 ( .A(n14182), .B(n14181), .ZN(n14243) );
  XOR2_X1 U15620 ( .A(n10662), .B(n14778), .Z(n14184) );
  XNOR2_X1 U15621 ( .A(n14183), .B(n14184), .ZN(n14312) );
  INV_X1 U15622 ( .A(n14183), .ZN(n14185) );
  XNOR2_X1 U15623 ( .A(n14609), .B(n14188), .ZN(n14253) );
  NAND2_X1 U15624 ( .A1(n14480), .A2(n14633), .ZN(n14189) );
  NOR2_X1 U15625 ( .A1(n14253), .A2(n14189), .ZN(n14190) );
  AOI21_X1 U15626 ( .B1(n14253), .B2(n14189), .A(n14190), .ZN(n14289) );
  INV_X1 U15627 ( .A(n14190), .ZN(n14191) );
  NAND2_X1 U15628 ( .A1(n14288), .A2(n14191), .ZN(n14196) );
  XNOR2_X1 U15629 ( .A(n14759), .B(n10662), .ZN(n14331) );
  AND2_X1 U15630 ( .A1(n14482), .A2(n14633), .ZN(n14192) );
  NAND2_X1 U15631 ( .A1(n14331), .A2(n14192), .ZN(n14198) );
  INV_X1 U15632 ( .A(n14331), .ZN(n14194) );
  INV_X1 U15633 ( .A(n14192), .ZN(n14193) );
  NAND2_X1 U15634 ( .A1(n14194), .A2(n14193), .ZN(n14195) );
  AND2_X1 U15635 ( .A1(n14198), .A2(n14195), .ZN(n14251) );
  XNOR2_X1 U15636 ( .A(n14197), .B(n14199), .ZN(n14334) );
  XNOR2_X1 U15637 ( .A(n14563), .B(n10662), .ZN(n14227) );
  AND2_X1 U15638 ( .A1(n14520), .A2(n14633), .ZN(n14200) );
  NAND2_X1 U15639 ( .A1(n14227), .A2(n14200), .ZN(n14237) );
  OAI21_X1 U15640 ( .B1(n14227), .B2(n14200), .A(n14237), .ZN(n14202) );
  NAND2_X1 U15641 ( .A1(n14526), .A2(n14338), .ZN(n14204) );
  OR2_X1 U15642 ( .A1(n14484), .A2(n14313), .ZN(n14203) );
  NAND2_X1 U15643 ( .A1(n14204), .A2(n14203), .ZN(n14550) );
  INV_X1 U15644 ( .A(n14205), .ZN(n14557) );
  OAI22_X1 U15645 ( .A1(n14557), .A2(n14351), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14206), .ZN(n14207) );
  AOI21_X1 U15646 ( .B1(n14550), .B2(n14348), .A(n14207), .ZN(n14208) );
  AOI22_X1 U15647 ( .A1(n14209), .A2(n14311), .B1(n14330), .B2(n14478), .ZN(
        n14215) );
  INV_X1 U15648 ( .A(n14210), .ZN(n14214) );
  INV_X1 U15649 ( .A(n14476), .ZN(n14509) );
  OAI22_X1 U15650 ( .A1(n14515), .A2(n14453), .B1(n14509), .B2(n14313), .ZN(
        n14615) );
  AOI22_X1 U15651 ( .A1(n14615), .A2(n14348), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14211) );
  OAI21_X1 U15652 ( .B1(n14621), .B2(n14351), .A(n14211), .ZN(n14212) );
  AOI21_X1 U15653 ( .B1(n14769), .B2(n14358), .A(n14212), .ZN(n14213) );
  OAI21_X1 U15654 ( .B1(n14215), .B2(n14214), .A(n14213), .ZN(P2_U3188) );
  INV_X1 U15655 ( .A(n14686), .ZN(n14793) );
  OAI21_X1 U15656 ( .B1(n14324), .B2(n14216), .A(n14311), .ZN(n14219) );
  NAND3_X1 U15657 ( .A1(n14217), .A2(n14330), .A3(n14497), .ZN(n14218) );
  NAND2_X1 U15658 ( .A1(n14219), .A2(n14218), .ZN(n14220) );
  NAND2_X1 U15659 ( .A1(n14299), .A2(n14220), .ZN(n14226) );
  INV_X1 U15660 ( .A(n14683), .ZN(n14224) );
  AND2_X1 U15661 ( .A1(n14497), .A2(n14525), .ZN(n14221) );
  AOI21_X1 U15662 ( .B1(n14474), .B2(n14338), .A(n14221), .ZN(n14678) );
  OAI21_X1 U15663 ( .B1(n14341), .B2(n14678), .A(n14222), .ZN(n14223) );
  AOI21_X1 U15664 ( .B1(n14224), .B2(n14339), .A(n14223), .ZN(n14225) );
  OAI211_X1 U15665 ( .C1(n14793), .C2(n14309), .A(n14226), .B(n14225), .ZN(
        P2_U3191) );
  NAND3_X1 U15666 ( .A1(n14227), .A2(n14330), .A3(n14520), .ZN(n14228) );
  MUX2_X1 U15667 ( .A(n14486), .B(n14741), .S(n14716), .Z(n14230) );
  XNOR2_X1 U15668 ( .A(n14230), .B(n10662), .ZN(n14235) );
  NAND2_X1 U15669 ( .A1(n14231), .A2(n14235), .ZN(n14240) );
  AOI22_X1 U15670 ( .A1(n14520), .A2(n14525), .B1(n14361), .B2(n14338), .ZN(
        n14539) );
  INV_X1 U15671 ( .A(n14543), .ZN(n14232) );
  AOI22_X1 U15672 ( .A1(n14232), .A2(n14339), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14233) );
  OAI21_X1 U15673 ( .B1(n14539), .B2(n14341), .A(n14233), .ZN(n14234) );
  AOI21_X1 U15674 ( .B1(n14545), .B2(n14358), .A(n14234), .ZN(n14239) );
  INV_X1 U15675 ( .A(n14235), .ZN(n14236) );
  NOR3_X1 U15676 ( .A1(n14241), .A2(n14505), .A3(n14296), .ZN(n14242) );
  AOI21_X1 U15677 ( .B1(n14300), .B2(n14311), .A(n14242), .ZN(n14250) );
  INV_X1 U15678 ( .A(n14243), .ZN(n14249) );
  INV_X1 U15679 ( .A(n14784), .ZN(n14656) );
  AOI22_X1 U15680 ( .A1(n14476), .A2(n14338), .B1(n14525), .B2(n14474), .ZN(
        n14648) );
  OAI22_X1 U15681 ( .A1(n14648), .A2(n14341), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14244), .ZN(n14245) );
  AOI21_X1 U15682 ( .B1(n14653), .B2(n14339), .A(n14245), .ZN(n14246) );
  OAI21_X1 U15683 ( .B1(n14656), .B2(n14309), .A(n14246), .ZN(n14247) );
  AOI21_X1 U15684 ( .B1(n7362), .B2(n14311), .A(n14247), .ZN(n14248) );
  OAI21_X1 U15685 ( .B1(n14250), .B2(n14249), .A(n14248), .ZN(P2_U3195) );
  INV_X1 U15686 ( .A(n14759), .ZN(n14262) );
  INV_X1 U15687 ( .A(n14251), .ZN(n14252) );
  AOI21_X1 U15688 ( .B1(n14288), .B2(n14252), .A(n14353), .ZN(n14255) );
  NOR3_X1 U15689 ( .A1(n14253), .A2(n14515), .A3(n14296), .ZN(n14254) );
  OAI21_X1 U15690 ( .B1(n14255), .B2(n14254), .A(n14333), .ZN(n14261) );
  OR2_X1 U15691 ( .A1(n14484), .A2(n14453), .ZN(n14257) );
  NAND2_X1 U15692 ( .A1(n14480), .A2(n14525), .ZN(n14256) );
  NAND2_X1 U15693 ( .A1(n14257), .A2(n14256), .ZN(n14583) );
  OAI22_X1 U15694 ( .A1(n14589), .A2(n14351), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14258), .ZN(n14259) );
  AOI21_X1 U15695 ( .B1(n14583), .B2(n14348), .A(n14259), .ZN(n14260) );
  OAI211_X1 U15696 ( .C1(n14262), .C2(n14309), .A(n14261), .B(n14260), .ZN(
        P2_U3197) );
  OAI21_X1 U15697 ( .B1(n14265), .B2(n14264), .A(n14263), .ZN(n14266) );
  NAND2_X1 U15698 ( .A1(n14266), .A2(n14311), .ZN(n14275) );
  NAND2_X1 U15699 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n15575) );
  INV_X1 U15700 ( .A(n15575), .ZN(n14267) );
  AOI21_X1 U15701 ( .B1(n14348), .B2(n14268), .A(n14267), .ZN(n14274) );
  NAND2_X1 U15702 ( .A1(n14358), .A2(n14269), .ZN(n14273) );
  INV_X1 U15703 ( .A(n14270), .ZN(n14271) );
  NAND2_X1 U15704 ( .A1(n14339), .A2(n14271), .ZN(n14272) );
  NAND4_X1 U15705 ( .A1(n14275), .A2(n14274), .A3(n14273), .A4(n14272), .ZN(
        P2_U3199) );
  AND2_X1 U15706 ( .A1(n14463), .A2(n14525), .ZN(n14276) );
  AOI21_X1 U15707 ( .B1(n14497), .B2(n14338), .A(n14276), .ZN(n14712) );
  INV_X1 U15708 ( .A(n14712), .ZN(n14277) );
  AOI22_X1 U15709 ( .A1(n14348), .A2(n14277), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14278) );
  OAI21_X1 U15710 ( .B1(n14351), .B2(n14719), .A(n14278), .ZN(n14279) );
  AOI21_X1 U15711 ( .B1(n14723), .B2(n14358), .A(n14279), .ZN(n14286) );
  INV_X1 U15712 ( .A(n14280), .ZN(n14283) );
  INV_X1 U15713 ( .A(n14463), .ZN(n14492) );
  OAI22_X1 U15714 ( .A1(n14281), .A2(n14353), .B1(n14492), .B2(n14296), .ZN(
        n14282) );
  NAND3_X1 U15715 ( .A1(n14284), .A2(n14283), .A3(n14282), .ZN(n14285) );
  OAI211_X1 U15716 ( .C1(n14287), .C2(n14353), .A(n14286), .B(n14285), .ZN(
        P2_U3200) );
  OAI211_X1 U15717 ( .C1(n14290), .C2(n14289), .A(n14288), .B(n14311), .ZN(
        n14295) );
  INV_X1 U15718 ( .A(n14482), .ZN(n14516) );
  OAI22_X1 U15719 ( .A1(n14516), .A2(n14453), .B1(n14512), .B2(n14313), .ZN(
        n14599) );
  INV_X1 U15720 ( .A(n14608), .ZN(n14292) );
  OAI22_X1 U15721 ( .A1(n14351), .A2(n14292), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14291), .ZN(n14293) );
  AOI21_X1 U15722 ( .B1(n14599), .B2(n14348), .A(n14293), .ZN(n14294) );
  OAI211_X1 U15723 ( .C1(n7706), .C2(n14309), .A(n14295), .B(n14294), .ZN(
        P2_U3201) );
  INV_X1 U15724 ( .A(n14789), .ZN(n14662) );
  INV_X1 U15725 ( .A(n14470), .ZN(n14501) );
  NOR3_X1 U15726 ( .A1(n14297), .A2(n14501), .A3(n14296), .ZN(n14303) );
  AOI21_X1 U15727 ( .B1(n14299), .B2(n14298), .A(n14353), .ZN(n14302) );
  INV_X1 U15728 ( .A(n14300), .ZN(n14301) );
  OAI21_X1 U15729 ( .B1(n14303), .B2(n14302), .A(n14301), .ZN(n14308) );
  INV_X1 U15730 ( .A(n14663), .ZN(n14306) );
  AOI22_X1 U15731 ( .A1(n14507), .A2(n14338), .B1(n14525), .B2(n14470), .ZN(
        n14670) );
  OAI22_X1 U15732 ( .A1(n14670), .A2(n14341), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14304), .ZN(n14305) );
  AOI21_X1 U15733 ( .B1(n14306), .B2(n14339), .A(n14305), .ZN(n14307) );
  OAI211_X1 U15734 ( .C1(n14662), .C2(n14309), .A(n14308), .B(n14307), .ZN(
        P2_U3205) );
  INV_X1 U15735 ( .A(n14310), .ZN(n14319) );
  AOI22_X1 U15736 ( .A1(n14312), .A2(n14311), .B1(n14330), .B2(n14476), .ZN(
        n14318) );
  OAI22_X1 U15737 ( .A1(n14512), .A2(n14453), .B1(n14314), .B2(n14313), .ZN(
        n14628) );
  AOI22_X1 U15738 ( .A1(n14628), .A2(n14348), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14315) );
  OAI21_X1 U15739 ( .B1(n14636), .B2(n14351), .A(n14315), .ZN(n14316) );
  AOI21_X1 U15740 ( .B1(n14778), .B2(n14358), .A(n14316), .ZN(n14317) );
  OAI21_X1 U15741 ( .B1(n14319), .B2(n14318), .A(n14317), .ZN(P2_U3207) );
  INV_X1 U15742 ( .A(n14696), .ZN(n14323) );
  NAND2_X1 U15743 ( .A1(n14470), .A2(n14338), .ZN(n14321) );
  NAND2_X1 U15744 ( .A1(n14466), .A2(n14525), .ZN(n14320) );
  NAND2_X1 U15745 ( .A1(n14321), .A2(n14320), .ZN(n14693) );
  AOI22_X1 U15746 ( .A1(n14348), .A2(n14693), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14322) );
  OAI21_X1 U15747 ( .B1(n14351), .B2(n14323), .A(n14322), .ZN(n14328) );
  AOI211_X1 U15748 ( .C1(n14326), .C2(n14325), .A(n14353), .B(n14324), .ZN(
        n14327) );
  AOI211_X1 U15749 ( .C1(n14698), .C2(n14358), .A(n14328), .B(n14327), .ZN(
        n14329) );
  INV_X1 U15750 ( .A(n14329), .ZN(P2_U3210) );
  NAND3_X1 U15751 ( .A1(n14331), .A2(n14330), .A3(n14482), .ZN(n14332) );
  OAI21_X1 U15752 ( .B1(n14333), .B2(n14353), .A(n14332), .ZN(n14336) );
  INV_X1 U15753 ( .A(n14334), .ZN(n14335) );
  NAND2_X1 U15754 ( .A1(n14336), .A2(n14335), .ZN(n14344) );
  AND2_X1 U15755 ( .A1(n14482), .A2(n14525), .ZN(n14337) );
  AOI21_X1 U15756 ( .B1(n14520), .B2(n14338), .A(n14337), .ZN(n14577) );
  AOI22_X1 U15757 ( .A1(n14571), .A2(n14339), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14340) );
  OAI21_X1 U15758 ( .B1(n14577), .B2(n14341), .A(n14340), .ZN(n14342) );
  AOI21_X1 U15759 ( .B1(n14755), .B2(n14358), .A(n14342), .ZN(n14343) );
  OAI211_X1 U15760 ( .C1(n14345), .C2(n14353), .A(n14344), .B(n14343), .ZN(
        P2_U3212) );
  INV_X1 U15761 ( .A(n14346), .ZN(n14347) );
  AOI22_X1 U15762 ( .A1(n14348), .A2(n14347), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14349) );
  OAI21_X1 U15763 ( .B1(n14351), .B2(n14350), .A(n14349), .ZN(n14357) );
  AOI211_X1 U15764 ( .C1(n14355), .C2(n14354), .A(n14353), .B(n14352), .ZN(
        n14356) );
  AOI211_X1 U15765 ( .C1(n14359), .C2(n14358), .A(n14357), .B(n14356), .ZN(
        n14360) );
  INV_X1 U15766 ( .A(n14360), .ZN(P2_U3213) );
  MUX2_X1 U15767 ( .A(n14454), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14376), .Z(
        P2_U3562) );
  MUX2_X1 U15768 ( .A(n14528), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14376), .Z(
        P2_U3561) );
  MUX2_X1 U15769 ( .A(n14361), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14376), .Z(
        P2_U3560) );
  MUX2_X1 U15770 ( .A(n14526), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14376), .Z(
        P2_U3559) );
  MUX2_X1 U15771 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n14520), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15772 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n14517), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15773 ( .A(n14482), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14376), .Z(
        P2_U3556) );
  MUX2_X1 U15774 ( .A(n14480), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14376), .Z(
        P2_U3555) );
  MUX2_X1 U15775 ( .A(n14478), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14376), .Z(
        P2_U3554) );
  MUX2_X1 U15776 ( .A(n14476), .B(P2_DATAO_REG_22__SCAN_IN), .S(n14376), .Z(
        P2_U3553) );
  MUX2_X1 U15777 ( .A(n14507), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14376), .Z(
        P2_U3552) );
  MUX2_X1 U15778 ( .A(n14474), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14376), .Z(
        P2_U3551) );
  MUX2_X1 U15779 ( .A(n14470), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14376), .Z(
        P2_U3550) );
  MUX2_X1 U15780 ( .A(n14497), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14376), .Z(
        P2_U3549) );
  MUX2_X1 U15781 ( .A(n14466), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14376), .Z(
        P2_U3548) );
  MUX2_X1 U15782 ( .A(n14463), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14376), .Z(
        P2_U3547) );
  MUX2_X1 U15783 ( .A(n14362), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14376), .Z(
        P2_U3546) );
  MUX2_X1 U15784 ( .A(n14363), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14376), .Z(
        P2_U3545) );
  MUX2_X1 U15785 ( .A(n14364), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14376), .Z(
        P2_U3544) );
  MUX2_X1 U15786 ( .A(n14365), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14376), .Z(
        P2_U3543) );
  MUX2_X1 U15787 ( .A(n14366), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14376), .Z(
        P2_U3542) );
  MUX2_X1 U15788 ( .A(n14367), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14376), .Z(
        P2_U3541) );
  MUX2_X1 U15789 ( .A(n14368), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14376), .Z(
        P2_U3540) );
  MUX2_X1 U15790 ( .A(n14369), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14376), .Z(
        P2_U3539) );
  MUX2_X1 U15791 ( .A(n14370), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14376), .Z(
        P2_U3538) );
  MUX2_X1 U15792 ( .A(n14371), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14376), .Z(
        P2_U3537) );
  MUX2_X1 U15793 ( .A(n14372), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14376), .Z(
        P2_U3536) );
  MUX2_X1 U15794 ( .A(n14373), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14376), .Z(
        P2_U3535) );
  MUX2_X1 U15795 ( .A(n14374), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14376), .Z(
        P2_U3534) );
  MUX2_X1 U15796 ( .A(n14375), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14376), .Z(
        P2_U3533) );
  MUX2_X1 U15797 ( .A(n14377), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14376), .Z(
        P2_U3532) );
  OAI211_X1 U15798 ( .C1(n14380), .C2(n14379), .A(n15602), .B(n14378), .ZN(
        n14391) );
  MUX2_X1 U15799 ( .A(n10525), .B(P2_REG2_REG_3__SCAN_IN), .S(n14387), .Z(
        n14381) );
  NAND3_X1 U15800 ( .A1(n15547), .A2(n14382), .A3(n14381), .ZN(n14383) );
  NAND3_X1 U15801 ( .A1(n15611), .A2(n14384), .A3(n14383), .ZN(n14390) );
  NOR2_X1 U15802 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14385), .ZN(n14386) );
  AOI21_X1 U15803 ( .B1(n15627), .B2(n14387), .A(n14386), .ZN(n14389) );
  NAND2_X1 U15804 ( .A1(n15619), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n14388) );
  NAND4_X1 U15805 ( .A1(n14391), .A2(n14390), .A3(n14389), .A4(n14388), .ZN(
        P2_U3217) );
  OAI211_X1 U15806 ( .C1(n14394), .C2(n14393), .A(n15602), .B(n14392), .ZN(
        n14404) );
  MUX2_X1 U15807 ( .A(n11805), .B(P2_REG2_REG_7__SCAN_IN), .S(n14400), .Z(
        n14395) );
  NAND3_X1 U15808 ( .A1(n15583), .A2(n14396), .A3(n14395), .ZN(n14397) );
  NAND3_X1 U15809 ( .A1(n15611), .A2(n14410), .A3(n14397), .ZN(n14403) );
  INV_X1 U15810 ( .A(n14398), .ZN(n14399) );
  AOI21_X1 U15811 ( .B1(n15627), .B2(n14400), .A(n14399), .ZN(n14402) );
  NAND2_X1 U15812 ( .A1(n15619), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n14401) );
  NAND4_X1 U15813 ( .A1(n14404), .A2(n14403), .A3(n14402), .A4(n14401), .ZN(
        P2_U3221) );
  OAI211_X1 U15814 ( .C1(n14407), .C2(n14406), .A(n15602), .B(n14405), .ZN(
        n14419) );
  MUX2_X1 U15815 ( .A(n11756), .B(P2_REG2_REG_8__SCAN_IN), .S(n14415), .Z(
        n14408) );
  NAND3_X1 U15816 ( .A1(n14410), .A2(n14409), .A3(n14408), .ZN(n14411) );
  NAND3_X1 U15817 ( .A1(n15611), .A2(n14412), .A3(n14411), .ZN(n14418) );
  INV_X1 U15818 ( .A(n14413), .ZN(n14414) );
  AOI21_X1 U15819 ( .B1(n15627), .B2(n14415), .A(n14414), .ZN(n14417) );
  NAND2_X1 U15820 ( .A1(n15619), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n14416) );
  NAND4_X1 U15821 ( .A1(n14419), .A2(n14418), .A3(n14417), .A4(n14416), .ZN(
        P2_U3222) );
  NOR2_X1 U15822 ( .A1(n15543), .A2(n14420), .ZN(n14421) );
  AOI211_X1 U15823 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n15619), .A(n14422), 
        .B(n14421), .ZN(n14435) );
  AOI21_X1 U15824 ( .B1(n14424), .B2(n14423), .A(n15622), .ZN(n14426) );
  NAND2_X1 U15825 ( .A1(n14426), .A2(n14425), .ZN(n14434) );
  INV_X1 U15826 ( .A(n14427), .ZN(n14432) );
  MUX2_X1 U15827 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n14429), .S(n14428), .Z(
        n14431) );
  OAI211_X1 U15828 ( .C1(n14432), .C2(n14431), .A(n15611), .B(n14430), .ZN(
        n14433) );
  NAND3_X1 U15829 ( .A1(n14435), .A2(n14434), .A3(n14433), .ZN(P2_U3224) );
  AOI211_X1 U15830 ( .C1(n14438), .C2(n14437), .A(n15622), .B(n14436), .ZN(
        n14439) );
  INV_X1 U15831 ( .A(n14439), .ZN(n14448) );
  AND2_X1 U15832 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14442) );
  NOR2_X1 U15833 ( .A1(n15543), .A2(n14440), .ZN(n14441) );
  AOI211_X1 U15834 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n15619), .A(n14442), 
        .B(n14441), .ZN(n14447) );
  OAI211_X1 U15835 ( .C1(n14445), .C2(n14444), .A(n14443), .B(n15611), .ZN(
        n14446) );
  NAND3_X1 U15836 ( .A1(n14448), .A2(n14447), .A3(n14446), .ZN(P2_U3231) );
  INV_X1 U15837 ( .A(n14698), .ZN(n14801) );
  NAND2_X1 U15838 ( .A1(n14801), .A2(n14715), .ZN(n14695) );
  NAND2_X1 U15839 ( .A1(n14660), .A2(n14656), .ZN(n14650) );
  NAND2_X1 U15840 ( .A1(n14449), .A2(n14716), .ZN(n14731) );
  NOR2_X1 U15841 ( .A1(n12155), .A2(n14450), .ZN(n14455) );
  INV_X1 U15842 ( .A(P2_B_REG_SCAN_IN), .ZN(n14451) );
  NOR2_X1 U15843 ( .A1(n14868), .A2(n14451), .ZN(n14452) );
  NOR2_X1 U15844 ( .A1(n14453), .A2(n14452), .ZN(n14527) );
  NAND2_X1 U15845 ( .A1(n14454), .A2(n14527), .ZN(n14732) );
  NOR2_X1 U15846 ( .A1(n15891), .A2(n14732), .ZN(n14459) );
  AOI211_X1 U15847 ( .C1(n14730), .C2(n14722), .A(n14455), .B(n14459), .ZN(
        n14456) );
  OAI21_X1 U15848 ( .B1(n14731), .B2(n14725), .A(n14456), .ZN(P2_U3234) );
  OAI211_X1 U15849 ( .C1(n14487), .C2(n14734), .A(n14457), .B(n14716), .ZN(
        n14733) );
  NOR2_X1 U15850 ( .A1(n12155), .A2(n14458), .ZN(n14460) );
  AOI211_X1 U15851 ( .C1(n14461), .C2(n14722), .A(n14460), .B(n14459), .ZN(
        n14462) );
  OAI21_X1 U15852 ( .B1(n14733), .B2(n14725), .A(n14462), .ZN(P2_U3235) );
  NAND2_X1 U15853 ( .A1(n14808), .A2(n14463), .ZN(n14464) );
  OR2_X1 U15854 ( .A1(n14723), .A2(n14466), .ZN(n14467) );
  OR2_X1 U15855 ( .A1(n14698), .A2(n14497), .ZN(n14469) );
  INV_X1 U15856 ( .A(n14676), .ZN(n14674) );
  OR2_X1 U15857 ( .A1(n14686), .A2(n14470), .ZN(n14471) );
  NAND2_X1 U15858 ( .A1(n14472), .A2(n14471), .ZN(n14659) );
  NOR2_X1 U15859 ( .A1(n14789), .A2(n14474), .ZN(n14473) );
  NAND2_X1 U15860 ( .A1(n14789), .A2(n14474), .ZN(n14475) );
  NAND2_X1 U15861 ( .A1(n14778), .A2(n14476), .ZN(n14477) );
  OR2_X1 U15862 ( .A1(n14769), .A2(n14478), .ZN(n14479) );
  NAND2_X1 U15863 ( .A1(n14601), .A2(n14514), .ZN(n14604) );
  NAND2_X1 U15864 ( .A1(n14609), .A2(n14480), .ZN(n14481) );
  INV_X1 U15865 ( .A(n14581), .ZN(n14586) );
  NAND2_X1 U15866 ( .A1(n14587), .A2(n14586), .ZN(n14585) );
  NAND2_X1 U15867 ( .A1(n14759), .A2(n14482), .ZN(n14483) );
  NAND2_X1 U15868 ( .A1(n14585), .A2(n14483), .ZN(n14568) );
  OR2_X2 U15869 ( .A1(n14568), .A2(n14576), .ZN(n14566) );
  NAND2_X1 U15870 ( .A1(n14573), .A2(n14484), .ZN(n14485) );
  AOI211_X1 U15871 ( .C1(n14736), .C2(n14541), .A(n14633), .B(n14487), .ZN(
        n14735) );
  INV_X1 U15872 ( .A(n14736), .ZN(n14491) );
  INV_X1 U15873 ( .A(n14488), .ZN(n14489) );
  AOI22_X1 U15874 ( .A1(n14489), .A2(n15884), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14697), .ZN(n14490) );
  OAI21_X1 U15875 ( .B1(n14491), .B2(n14661), .A(n14490), .ZN(n14531) );
  OR2_X1 U15876 ( .A1(n14808), .A2(n14492), .ZN(n14706) );
  NAND2_X1 U15877 ( .A1(n14494), .A2(n14493), .ZN(n14711) );
  OR2_X1 U15878 ( .A1(n14723), .A2(n14495), .ZN(n14496) );
  INV_X1 U15879 ( .A(n14497), .ZN(n14499) );
  NAND2_X1 U15880 ( .A1(n14698), .A2(n14499), .ZN(n14498) );
  OR2_X1 U15881 ( .A1(n14698), .A2(n14499), .ZN(n14500) );
  NAND2_X1 U15882 ( .A1(n14686), .A2(n14501), .ZN(n14502) );
  AND2_X1 U15883 ( .A1(n14789), .A2(n14505), .ZN(n14504) );
  OR2_X1 U15884 ( .A1(n14789), .A2(n14505), .ZN(n14506) );
  NOR2_X1 U15885 ( .A1(n14778), .A2(n14509), .ZN(n14508) );
  NAND2_X1 U15886 ( .A1(n14778), .A2(n14509), .ZN(n14510) );
  NAND2_X1 U15887 ( .A1(n14769), .A2(n14512), .ZN(n14513) );
  INV_X1 U15888 ( .A(n14514), .ZN(n14602) );
  OR2_X1 U15889 ( .A1(n14573), .A2(n14517), .ZN(n14518) );
  INV_X1 U15890 ( .A(n14520), .ZN(n14521) );
  NAND2_X1 U15891 ( .A1(n14538), .A2(n14522), .ZN(n14523) );
  NAND2_X1 U15892 ( .A1(n14526), .A2(n14525), .ZN(n14530) );
  OAI21_X1 U15893 ( .B1(n14728), .B2(n14739), .A(n14532), .ZN(P2_U3236) );
  OAI21_X1 U15894 ( .B1(n14534), .B2(n14535), .A(n14533), .ZN(n14744) );
  INV_X1 U15895 ( .A(n14744), .ZN(n14822) );
  NAND2_X1 U15896 ( .A1(n14536), .A2(n14535), .ZN(n14537) );
  NAND3_X1 U15897 ( .A1(n14538), .A2(n14710), .A3(n14537), .ZN(n14540) );
  OAI211_X1 U15898 ( .C1(n14741), .C2(n14558), .A(n14716), .B(n14541), .ZN(
        n14740) );
  OAI22_X1 U15899 ( .A1(n14543), .A2(n14718), .B1(n14542), .B2(n12155), .ZN(
        n14544) );
  AOI21_X1 U15900 ( .B1(n14545), .B2(n14722), .A(n14544), .ZN(n14546) );
  OAI21_X1 U15901 ( .B1(n14740), .B2(n14725), .A(n14546), .ZN(n14547) );
  AOI21_X1 U15902 ( .B1(n14743), .B2(n12155), .A(n14547), .ZN(n14548) );
  OAI21_X1 U15903 ( .B1(n14822), .B2(n14728), .A(n14548), .ZN(P2_U3237) );
  XNOR2_X1 U15904 ( .A(n14549), .B(n14552), .ZN(n14551) );
  AND2_X1 U15905 ( .A1(n14553), .A2(n14552), .ZN(n14554) );
  NOR2_X1 U15906 ( .A1(n14555), .A2(n14554), .ZN(n14750) );
  NAND2_X1 U15907 ( .A1(n14750), .A2(n14642), .ZN(n14565) );
  OAI22_X1 U15908 ( .A1(n14557), .A2(n14718), .B1(n14556), .B2(n12155), .ZN(
        n14562) );
  INV_X1 U15909 ( .A(n14570), .ZN(n14560) );
  INV_X1 U15910 ( .A(n14558), .ZN(n14559) );
  OAI211_X1 U15911 ( .C1(n14748), .C2(n14560), .A(n14559), .B(n14716), .ZN(
        n14746) );
  NOR2_X1 U15912 ( .A1(n14746), .A2(n14725), .ZN(n14561) );
  AOI211_X1 U15913 ( .C1(n14722), .C2(n14563), .A(n14562), .B(n14561), .ZN(
        n14564) );
  OAI211_X1 U15914 ( .C1(n15891), .C2(n14747), .A(n14565), .B(n14564), .ZN(
        P2_U3238) );
  INV_X1 U15915 ( .A(n14566), .ZN(n14567) );
  AOI21_X1 U15916 ( .B1(n14576), .B2(n14568), .A(n14567), .ZN(n14757) );
  OR2_X1 U15917 ( .A1(n14573), .A2(n14593), .ZN(n14569) );
  AND3_X1 U15918 ( .A1(n14570), .A2(n14569), .A3(n14716), .ZN(n14754) );
  AOI22_X1 U15919 ( .A1(n14571), .A2(n15884), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n15891), .ZN(n14572) );
  OAI21_X1 U15920 ( .B1(n14573), .B2(n14661), .A(n14572), .ZN(n14574) );
  AOI21_X1 U15921 ( .B1(n14754), .B2(n14667), .A(n14574), .ZN(n14580) );
  XOR2_X1 U15922 ( .A(n14576), .B(n14575), .Z(n14578) );
  OAI21_X1 U15923 ( .B1(n14578), .B2(n14679), .A(n14577), .ZN(n14753) );
  NAND2_X1 U15924 ( .A1(n14753), .A2(n12155), .ZN(n14579) );
  OAI211_X1 U15925 ( .C1(n14757), .C2(n14728), .A(n14580), .B(n14579), .ZN(
        P2_U3239) );
  XNOR2_X1 U15926 ( .A(n14582), .B(n14581), .ZN(n14584) );
  AOI21_X1 U15927 ( .B1(n14584), .B2(n14710), .A(n14583), .ZN(n14761) );
  OAI21_X1 U15928 ( .B1(n14587), .B2(n14586), .A(n14585), .ZN(n14762) );
  OAI22_X1 U15929 ( .A1(n14589), .A2(n14718), .B1(n14588), .B2(n12155), .ZN(
        n14590) );
  AOI21_X1 U15930 ( .B1(n14759), .B2(n14722), .A(n14590), .ZN(n14595) );
  NAND2_X1 U15931 ( .A1(n14759), .A2(n14606), .ZN(n14591) );
  NAND2_X1 U15932 ( .A1(n14591), .A2(n14716), .ZN(n14592) );
  NOR2_X1 U15933 ( .A1(n14593), .A2(n14592), .ZN(n14758) );
  NAND2_X1 U15934 ( .A1(n14758), .A2(n14667), .ZN(n14594) );
  OAI211_X1 U15935 ( .C1(n14762), .C2(n14728), .A(n14595), .B(n14594), .ZN(
        n14596) );
  INV_X1 U15936 ( .A(n14596), .ZN(n14597) );
  OAI21_X1 U15937 ( .B1(n14697), .B2(n14761), .A(n14597), .ZN(P2_U3240) );
  XNOR2_X1 U15938 ( .A(n14598), .B(n14602), .ZN(n14600) );
  AOI21_X1 U15939 ( .B1(n14600), .B2(n14710), .A(n14599), .ZN(n14764) );
  INV_X1 U15940 ( .A(n14601), .ZN(n14603) );
  NAND2_X1 U15941 ( .A1(n14603), .A2(n14602), .ZN(n14605) );
  AND2_X1 U15942 ( .A1(n14605), .A2(n14604), .ZN(n14766) );
  AOI21_X1 U15943 ( .B1(n14609), .B2(n14619), .A(n14633), .ZN(n14607) );
  NAND2_X1 U15944 ( .A1(n14607), .A2(n14606), .ZN(n14763) );
  AOI22_X1 U15945 ( .A1(n14608), .A2(n15884), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14697), .ZN(n14611) );
  NAND2_X1 U15946 ( .A1(n14609), .A2(n14722), .ZN(n14610) );
  OAI211_X1 U15947 ( .C1(n14763), .C2(n14725), .A(n14611), .B(n14610), .ZN(
        n14612) );
  AOI21_X1 U15948 ( .B1(n14766), .B2(n14642), .A(n14612), .ZN(n14613) );
  OAI21_X1 U15949 ( .B1(n14697), .B2(n14764), .A(n14613), .ZN(P2_U3241) );
  XNOR2_X1 U15950 ( .A(n14614), .B(n14617), .ZN(n14616) );
  AOI21_X1 U15951 ( .B1(n14616), .B2(n14710), .A(n14615), .ZN(n14771) );
  OAI21_X1 U15952 ( .B1(n7295), .B2(n7690), .A(n14618), .ZN(n14774) );
  AOI21_X1 U15953 ( .B1(n14769), .B2(n14634), .A(n14633), .ZN(n14620) );
  NAND2_X1 U15954 ( .A1(n14620), .A2(n14619), .ZN(n14770) );
  INV_X1 U15955 ( .A(n14621), .ZN(n14622) );
  AOI22_X1 U15956 ( .A1(n14622), .A2(n15884), .B1(n14697), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n14624) );
  NAND2_X1 U15957 ( .A1(n14769), .A2(n14722), .ZN(n14623) );
  OAI211_X1 U15958 ( .C1(n14770), .C2(n14725), .A(n14624), .B(n14623), .ZN(
        n14625) );
  AOI21_X1 U15959 ( .B1(n14774), .B2(n14642), .A(n14625), .ZN(n14626) );
  OAI21_X1 U15960 ( .B1(n14697), .B2(n14771), .A(n14626), .ZN(P2_U3242) );
  XOR2_X1 U15961 ( .A(n14630), .B(n14627), .Z(n14629) );
  AOI21_X1 U15962 ( .B1(n14629), .B2(n14710), .A(n14628), .ZN(n14780) );
  INV_X1 U15963 ( .A(n14630), .ZN(n14632) );
  OAI21_X1 U15964 ( .B1(n7298), .B2(n14632), .A(n14631), .ZN(n14781) );
  INV_X1 U15965 ( .A(n14781), .ZN(n14643) );
  INV_X1 U15966 ( .A(n14778), .ZN(n14640) );
  AOI21_X1 U15967 ( .B1(n14650), .B2(n14778), .A(n14633), .ZN(n14635) );
  AND2_X1 U15968 ( .A1(n14635), .A2(n14634), .ZN(n14777) );
  NAND2_X1 U15969 ( .A1(n14777), .A2(n14667), .ZN(n14639) );
  INV_X1 U15970 ( .A(n14636), .ZN(n14637) );
  AOI22_X1 U15971 ( .A1(n14697), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14637), 
        .B2(n15884), .ZN(n14638) );
  OAI211_X1 U15972 ( .C1(n14640), .C2(n14661), .A(n14639), .B(n14638), .ZN(
        n14641) );
  AOI21_X1 U15973 ( .B1(n14643), .B2(n14642), .A(n14641), .ZN(n14644) );
  OAI21_X1 U15974 ( .B1(n15891), .B2(n14780), .A(n14644), .ZN(P2_U3243) );
  XOR2_X1 U15975 ( .A(n14646), .B(n14645), .Z(n14786) );
  XNOR2_X1 U15976 ( .A(n14647), .B(n14646), .ZN(n14649) );
  OAI21_X1 U15977 ( .B1(n14649), .B2(n14679), .A(n14648), .ZN(n14782) );
  INV_X1 U15978 ( .A(n14660), .ZN(n14652) );
  INV_X1 U15979 ( .A(n14650), .ZN(n14651) );
  AOI211_X1 U15980 ( .C1(n14784), .C2(n14652), .A(n14633), .B(n14651), .ZN(
        n14783) );
  NAND2_X1 U15981 ( .A1(n14783), .A2(n14667), .ZN(n14655) );
  AOI22_X1 U15982 ( .A1(n14697), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14653), 
        .B2(n15884), .ZN(n14654) );
  OAI211_X1 U15983 ( .C1(n14656), .C2(n14661), .A(n14655), .B(n14654), .ZN(
        n14657) );
  AOI21_X1 U15984 ( .B1(n14782), .B2(n12155), .A(n14657), .ZN(n14658) );
  OAI21_X1 U15985 ( .B1(n14786), .B2(n14728), .A(n14658), .ZN(P2_U3244) );
  XNOR2_X1 U15986 ( .A(n14659), .B(n14669), .ZN(n14791) );
  AOI211_X1 U15987 ( .C1(n14789), .C2(n14681), .A(n14633), .B(n14660), .ZN(
        n14788) );
  NOR2_X1 U15988 ( .A1(n14662), .A2(n14661), .ZN(n14666) );
  OAI22_X1 U15989 ( .A1(n12155), .A2(n14664), .B1(n14663), .B2(n14718), .ZN(
        n14665) );
  AOI211_X1 U15990 ( .C1(n14788), .C2(n14667), .A(n14666), .B(n14665), .ZN(
        n14673) );
  XOR2_X1 U15991 ( .A(n14669), .B(n14668), .Z(n14671) );
  OAI21_X1 U15992 ( .B1(n14671), .B2(n14679), .A(n14670), .ZN(n14787) );
  NAND2_X1 U15993 ( .A1(n14787), .A2(n12155), .ZN(n14672) );
  OAI211_X1 U15994 ( .C1(n14791), .C2(n14728), .A(n14673), .B(n14672), .ZN(
        P2_U3245) );
  XNOR2_X1 U15995 ( .A(n14675), .B(n14674), .ZN(n14796) );
  INV_X1 U15996 ( .A(n14796), .ZN(n14842) );
  XNOR2_X1 U15997 ( .A(n14677), .B(n14676), .ZN(n14680) );
  OAI21_X1 U15998 ( .B1(n14680), .B2(n14679), .A(n14678), .ZN(n14795) );
  INV_X1 U15999 ( .A(n14695), .ZN(n14682) );
  OAI211_X1 U16000 ( .C1(n14682), .C2(n14793), .A(n14716), .B(n14681), .ZN(
        n14792) );
  OAI22_X1 U16001 ( .A1(n12155), .A2(n14684), .B1(n14683), .B2(n14718), .ZN(
        n14685) );
  AOI21_X1 U16002 ( .B1(n14686), .B2(n14722), .A(n14685), .ZN(n14687) );
  OAI21_X1 U16003 ( .B1(n14792), .B2(n14725), .A(n14687), .ZN(n14688) );
  AOI21_X1 U16004 ( .B1(n14795), .B2(n12155), .A(n14688), .ZN(n14689) );
  OAI21_X1 U16005 ( .B1(n14842), .B2(n14728), .A(n14689), .ZN(P2_U3246) );
  XNOR2_X1 U16006 ( .A(n14690), .B(n14691), .ZN(n14804) );
  INV_X1 U16007 ( .A(n14804), .ZN(n14846) );
  XNOR2_X1 U16008 ( .A(n14692), .B(n14691), .ZN(n14694) );
  AOI21_X1 U16009 ( .B1(n14694), .B2(n14710), .A(n14693), .ZN(n14800) );
  INV_X1 U16010 ( .A(n14800), .ZN(n14702) );
  OAI211_X1 U16011 ( .C1(n14801), .C2(n14715), .A(n14716), .B(n14695), .ZN(
        n14799) );
  AOI22_X1 U16012 ( .A1(n14697), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14696), 
        .B2(n15884), .ZN(n14700) );
  NAND2_X1 U16013 ( .A1(n14698), .A2(n14722), .ZN(n14699) );
  OAI211_X1 U16014 ( .C1(n14799), .C2(n14725), .A(n14700), .B(n14699), .ZN(
        n14701) );
  AOI21_X1 U16015 ( .B1(n14702), .B2(n12155), .A(n14701), .ZN(n14703) );
  OAI21_X1 U16016 ( .B1(n14846), .B2(n14728), .A(n14703), .ZN(P2_U3247) );
  OAI21_X1 U16017 ( .B1(n14705), .B2(n14707), .A(n14704), .ZN(n16154) );
  INV_X1 U16018 ( .A(n16154), .ZN(n14729) );
  NAND3_X1 U16019 ( .A1(n14708), .A2(n14707), .A3(n14706), .ZN(n14709) );
  NAND3_X1 U16020 ( .A1(n14711), .A2(n14710), .A3(n14709), .ZN(n14713) );
  NAND2_X1 U16021 ( .A1(n14713), .A2(n14712), .ZN(n16152) );
  INV_X1 U16022 ( .A(n14723), .ZN(n16150) );
  INV_X1 U16023 ( .A(n14715), .ZN(n14717) );
  OAI211_X1 U16024 ( .C1(n16150), .C2(n7703), .A(n14717), .B(n14716), .ZN(
        n16148) );
  OAI22_X1 U16025 ( .A1(n12155), .A2(n14720), .B1(n14719), .B2(n14718), .ZN(
        n14721) );
  AOI21_X1 U16026 ( .B1(n14723), .B2(n14722), .A(n14721), .ZN(n14724) );
  OAI21_X1 U16027 ( .B1(n16148), .B2(n14725), .A(n14724), .ZN(n14726) );
  AOI21_X1 U16028 ( .B1(n16152), .B2(n12155), .A(n14726), .ZN(n14727) );
  OAI21_X1 U16029 ( .B1(n14729), .B2(n14728), .A(n14727), .ZN(P2_U3248) );
  OAI211_X1 U16030 ( .C1(n7702), .C2(n16149), .A(n14731), .B(n14732), .ZN(
        n14817) );
  MUX2_X1 U16031 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14817), .S(n16156), .Z(
        P2_U3530) );
  OAI211_X1 U16032 ( .C1(n14734), .C2(n16149), .A(n14733), .B(n14732), .ZN(
        n14818) );
  MUX2_X1 U16033 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14818), .S(n16156), .Z(
        P2_U3529) );
  AOI21_X1 U16034 ( .B1(n16112), .B2(n14736), .A(n14735), .ZN(n14737) );
  MUX2_X1 U16035 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14819), .S(n16156), .Z(
        P2_U3528) );
  INV_X1 U16036 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n14745) );
  OAI21_X1 U16037 ( .B1(n14741), .B2(n16149), .A(n14740), .ZN(n14742) );
  INV_X1 U16038 ( .A(n14750), .ZN(n14825) );
  INV_X1 U16039 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n14751) );
  AOI21_X1 U16040 ( .B1(n14750), .B2(n14803), .A(n14749), .ZN(n14823) );
  MUX2_X1 U16041 ( .A(n14751), .B(n14823), .S(n16156), .Z(n14752) );
  OAI21_X1 U16042 ( .B1(n14825), .B2(n14816), .A(n14752), .ZN(P2_U3526) );
  AOI211_X1 U16043 ( .C1(n16112), .C2(n14755), .A(n14754), .B(n14753), .ZN(
        n14756) );
  OAI21_X1 U16044 ( .B1(n14757), .B2(n16006), .A(n14756), .ZN(n14826) );
  MUX2_X1 U16045 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14826), .S(n16156), .Z(
        P2_U3525) );
  AOI21_X1 U16046 ( .B1(n16112), .B2(n14759), .A(n14758), .ZN(n14760) );
  OAI211_X1 U16047 ( .C1(n14762), .C2(n16006), .A(n14761), .B(n14760), .ZN(
        n14827) );
  MUX2_X1 U16048 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14827), .S(n16156), .Z(
        P2_U3524) );
  OAI211_X1 U16049 ( .C1(n7706), .C2(n16149), .A(n14764), .B(n14763), .ZN(
        n14765) );
  AOI21_X1 U16050 ( .B1(n14766), .B2(n14803), .A(n14765), .ZN(n14829) );
  INV_X1 U16051 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n14767) );
  MUX2_X1 U16052 ( .A(n14829), .B(n14767), .S(n16155), .Z(n14768) );
  OAI21_X1 U16053 ( .B1(n14831), .B2(n14816), .A(n14768), .ZN(P2_U3523) );
  INV_X1 U16054 ( .A(n14774), .ZN(n14835) );
  INV_X1 U16055 ( .A(n14769), .ZN(n14772) );
  OAI211_X1 U16056 ( .C1(n14772), .C2(n16149), .A(n14771), .B(n14770), .ZN(
        n14773) );
  AOI21_X1 U16057 ( .B1(n14774), .B2(n14803), .A(n14773), .ZN(n14833) );
  INV_X1 U16058 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14775) );
  MUX2_X1 U16059 ( .A(n14833), .B(n14775), .S(n16155), .Z(n14776) );
  OAI21_X1 U16060 ( .B1(n14835), .B2(n14816), .A(n14776), .ZN(P2_U3522) );
  AOI21_X1 U16061 ( .B1(n16112), .B2(n14778), .A(n14777), .ZN(n14779) );
  OAI211_X1 U16062 ( .C1(n14781), .C2(n16006), .A(n14780), .B(n14779), .ZN(
        n14836) );
  MUX2_X1 U16063 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14836), .S(n16156), .Z(
        P2_U3521) );
  AOI211_X1 U16064 ( .C1(n16112), .C2(n14784), .A(n14783), .B(n14782), .ZN(
        n14785) );
  OAI21_X1 U16065 ( .B1(n14786), .B2(n16006), .A(n14785), .ZN(n14837) );
  MUX2_X1 U16066 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14837), .S(n16156), .Z(
        P2_U3520) );
  AOI211_X1 U16067 ( .C1(n16112), .C2(n14789), .A(n14788), .B(n14787), .ZN(
        n14790) );
  OAI21_X1 U16068 ( .B1(n16006), .B2(n14791), .A(n14790), .ZN(n14838) );
  MUX2_X1 U16069 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14838), .S(n16156), .Z(
        P2_U3519) );
  OAI21_X1 U16070 ( .B1(n14793), .B2(n16149), .A(n14792), .ZN(n14794) );
  AOI211_X1 U16071 ( .C1(n14796), .C2(n14803), .A(n14795), .B(n14794), .ZN(
        n14839) );
  MUX2_X1 U16072 ( .A(n14797), .B(n14839), .S(n16156), .Z(n14798) );
  OAI21_X1 U16073 ( .B1(n14842), .B2(n14816), .A(n14798), .ZN(P2_U3518) );
  INV_X1 U16074 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14805) );
  OAI211_X1 U16075 ( .C1(n14801), .C2(n16149), .A(n14800), .B(n14799), .ZN(
        n14802) );
  AOI21_X1 U16076 ( .B1(n14804), .B2(n14803), .A(n14802), .ZN(n14843) );
  MUX2_X1 U16077 ( .A(n14805), .B(n14843), .S(n16156), .Z(n14806) );
  OAI21_X1 U16078 ( .B1(n14846), .B2(n14816), .A(n14806), .ZN(P2_U3517) );
  OR2_X1 U16079 ( .A1(n14850), .A2(n14807), .ZN(n14814) );
  INV_X1 U16080 ( .A(n14808), .ZN(n14810) );
  OAI21_X1 U16081 ( .B1(n14810), .B2(n16149), .A(n14809), .ZN(n14811) );
  NOR2_X1 U16082 ( .A1(n14812), .A2(n14811), .ZN(n14813) );
  MUX2_X1 U16083 ( .A(n8248), .B(n12333), .S(n16155), .Z(n14815) );
  OAI21_X1 U16084 ( .B1(n14850), .B2(n14816), .A(n14815), .ZN(P2_U3515) );
  MUX2_X1 U16085 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n14817), .S(n16117), .Z(
        P2_U3498) );
  MUX2_X1 U16086 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14818), .S(n16117), .Z(
        P2_U3497) );
  MUX2_X1 U16087 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14819), .S(n16117), .Z(
        P2_U3496) );
  INV_X1 U16088 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n14821) );
  INV_X1 U16089 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n14824) );
  MUX2_X1 U16090 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14826), .S(n16117), .Z(
        P2_U3493) );
  MUX2_X1 U16091 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14827), .S(n16117), .Z(
        P2_U3492) );
  INV_X1 U16092 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n14828) );
  MUX2_X1 U16093 ( .A(n14829), .B(n14828), .S(n16157), .Z(n14830) );
  OAI21_X1 U16094 ( .B1(n14831), .B2(n14849), .A(n14830), .ZN(P2_U3491) );
  INV_X1 U16095 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14832) );
  MUX2_X1 U16096 ( .A(n14833), .B(n14832), .S(n16157), .Z(n14834) );
  OAI21_X1 U16097 ( .B1(n14835), .B2(n14849), .A(n14834), .ZN(P2_U3490) );
  MUX2_X1 U16098 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14836), .S(n16117), .Z(
        P2_U3489) );
  MUX2_X1 U16099 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14837), .S(n16117), .Z(
        P2_U3488) );
  MUX2_X1 U16100 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14838), .S(n16117), .Z(
        P2_U3487) );
  INV_X1 U16101 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14840) );
  MUX2_X1 U16102 ( .A(n14840), .B(n14839), .S(n16117), .Z(n14841) );
  OAI21_X1 U16103 ( .B1(n14842), .B2(n14849), .A(n14841), .ZN(P2_U3486) );
  INV_X1 U16104 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14844) );
  MUX2_X1 U16105 ( .A(n14844), .B(n14843), .S(n16117), .Z(n14845) );
  OAI21_X1 U16106 ( .B1(n14846), .B2(n14849), .A(n14845), .ZN(P2_U3484) );
  INV_X1 U16107 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n14847) );
  MUX2_X1 U16108 ( .A(n8248), .B(n14847), .S(n16157), .Z(n14848) );
  OAI21_X1 U16109 ( .B1(n14850), .B2(n14849), .A(n14848), .ZN(P2_U3478) );
  INV_X1 U16110 ( .A(n14851), .ZN(n15505) );
  NAND3_X1 U16111 ( .A1(n14853), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14855) );
  OAI22_X1 U16112 ( .A1(n14852), .A2(n14855), .B1(n14854), .B2(n14871), .ZN(
        n14856) );
  INV_X1 U16113 ( .A(n14856), .ZN(n14857) );
  OAI21_X1 U16114 ( .B1(n15505), .B2(n14869), .A(n14857), .ZN(P2_U3296) );
  OAI222_X1 U16115 ( .A1(n14860), .A2(P2_U3088), .B1(n14869), .B2(n14859), 
        .C1(n14858), .C2(n14871), .ZN(P2_U3297) );
  NAND2_X1 U16116 ( .A1(n14862), .A2(n14861), .ZN(n14864) );
  OAI211_X1 U16117 ( .C1(n14866), .C2(n14865), .A(n14864), .B(n14863), .ZN(
        P2_U3299) );
  INV_X1 U16118 ( .A(n14867), .ZN(n15509) );
  OAI222_X1 U16119 ( .A1(n14871), .A2(n14870), .B1(n14869), .B2(n15509), .C1(
        P2_U3088), .C2(n14868), .ZN(P2_U3300) );
  INV_X1 U16120 ( .A(n14872), .ZN(n14873) );
  MUX2_X1 U16121 ( .A(n14873), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U16122 ( .A1(n15413), .A2(n14905), .ZN(n14875) );
  NAND2_X1 U16123 ( .A1(n15056), .A2(n7404), .ZN(n14874) );
  NAND2_X1 U16124 ( .A1(n14875), .A2(n14874), .ZN(n14876) );
  XNOR2_X1 U16125 ( .A(n14876), .B(n14954), .ZN(n14880) );
  NAND2_X1 U16126 ( .A1(n15413), .A2(n7404), .ZN(n14878) );
  NAND2_X1 U16127 ( .A1(n15056), .A2(n14953), .ZN(n14877) );
  NAND2_X1 U16128 ( .A1(n14878), .A2(n14877), .ZN(n14879) );
  NOR2_X1 U16129 ( .A1(n14880), .A2(n14879), .ZN(n14951) );
  AOI22_X1 U16130 ( .A1(n15429), .A2(n9798), .B1(n14953), .B2(n15059), .ZN(
        n14895) );
  INV_X1 U16131 ( .A(n14895), .ZN(n14897) );
  NAND2_X1 U16132 ( .A1(n15429), .A2(n14905), .ZN(n14882) );
  NAND2_X1 U16133 ( .A1(n15059), .A2(n9798), .ZN(n14881) );
  NAND2_X1 U16134 ( .A1(n14882), .A2(n14881), .ZN(n14883) );
  XNOR2_X1 U16135 ( .A(n14883), .B(n14954), .ZN(n14896) );
  NAND2_X1 U16136 ( .A1(n15433), .A2(n14905), .ZN(n14889) );
  NAND2_X1 U16137 ( .A1(n15257), .A2(n7404), .ZN(n14888) );
  NAND2_X1 U16138 ( .A1(n14889), .A2(n14888), .ZN(n14890) );
  XNOR2_X1 U16139 ( .A(n14890), .B(n14954), .ZN(n14893) );
  AOI22_X1 U16140 ( .A1(n15433), .A2(n9798), .B1(n14953), .B2(n15257), .ZN(
        n14891) );
  XNOR2_X1 U16141 ( .A(n14893), .B(n14891), .ZN(n14927) );
  INV_X1 U16142 ( .A(n14891), .ZN(n14892) );
  XNOR2_X1 U16143 ( .A(n14896), .B(n14895), .ZN(n15003) );
  NAND2_X1 U16144 ( .A1(n15425), .A2(n14905), .ZN(n14899) );
  NAND2_X1 U16145 ( .A1(n15058), .A2(n7404), .ZN(n14898) );
  NAND2_X1 U16146 ( .A1(n14899), .A2(n14898), .ZN(n14900) );
  XNOR2_X1 U16147 ( .A(n14900), .B(n14954), .ZN(n14901) );
  AOI22_X1 U16148 ( .A1(n15425), .A2(n7404), .B1(n14953), .B2(n15058), .ZN(
        n14902) );
  XNOR2_X1 U16149 ( .A(n14901), .B(n14902), .ZN(n14977) );
  INV_X1 U16150 ( .A(n14901), .ZN(n14903) );
  NAND2_X1 U16151 ( .A1(n14903), .A2(n14902), .ZN(n14904) );
  NAND2_X1 U16152 ( .A1(n15420), .A2(n14905), .ZN(n14907) );
  NAND2_X1 U16153 ( .A1(n15057), .A2(n7404), .ZN(n14906) );
  NAND2_X1 U16154 ( .A1(n14907), .A2(n14906), .ZN(n14908) );
  XNOR2_X1 U16155 ( .A(n14908), .B(n14954), .ZN(n14911) );
  NAND2_X1 U16156 ( .A1(n15420), .A2(n7404), .ZN(n14910) );
  NAND2_X1 U16157 ( .A1(n15057), .A2(n14953), .ZN(n14909) );
  NAND2_X1 U16158 ( .A1(n14910), .A2(n14909), .ZN(n14912) );
  INV_X1 U16159 ( .A(n14911), .ZN(n14914) );
  INV_X1 U16160 ( .A(n14912), .ZN(n14913) );
  NAND2_X1 U16161 ( .A1(n14914), .A2(n14913), .ZN(n15033) );
  OAI21_X1 U16162 ( .B1(n14916), .B2(n14915), .A(n14952), .ZN(n14917) );
  NOR2_X1 U16163 ( .A1(n14918), .A2(n15049), .ZN(n14921) );
  OAI22_X1 U16164 ( .A1(n15177), .A2(n15036), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14919), .ZN(n14920) );
  AOI211_X1 U16165 ( .C1(n14987), .C2(n14922), .A(n14921), .B(n14920), .ZN(
        n14923) );
  INV_X1 U16166 ( .A(n15433), .ZN(n14935) );
  OAI21_X1 U16167 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n14928) );
  NAND2_X1 U16168 ( .A1(n14928), .A2(n16093), .ZN(n14934) );
  OAI22_X1 U16169 ( .A1(n14969), .A2(n15357), .B1(n14929), .B2(n15359), .ZN(
        n15236) );
  INV_X1 U16170 ( .A(n14930), .ZN(n15238) );
  OAI22_X1 U16171 ( .A1(n16098), .A2(n15238), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14931), .ZN(n14932) );
  AOI21_X1 U16172 ( .B1(n15236), .B2(n15020), .A(n14932), .ZN(n14933) );
  OAI211_X1 U16173 ( .C1(n14935), .C2(n16091), .A(n14934), .B(n14933), .ZN(
        P1_U3216) );
  OAI211_X1 U16174 ( .C1(n14938), .C2(n14937), .A(n14936), .B(n16093), .ZN(
        n14942) );
  AOI22_X1 U16175 ( .A1(n16089), .A2(n15072), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14941) );
  AOI22_X1 U16176 ( .A1(n9912), .A2(n14987), .B1(n16087), .B2(n15074), .ZN(
        n14940) );
  NAND2_X1 U16177 ( .A1(n15040), .A2(n15906), .ZN(n14939) );
  NAND4_X1 U16178 ( .A1(n14942), .A2(n14941), .A3(n14940), .A4(n14939), .ZN(
        P1_U3218) );
  NOR2_X1 U16179 ( .A1(n14944), .A2(n8045), .ZN(n14945) );
  XNOR2_X1 U16180 ( .A(n14946), .B(n14945), .ZN(n14950) );
  NAND2_X1 U16181 ( .A1(n7201), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15152) );
  OAI21_X1 U16182 ( .B1(n15341), .B2(n15049), .A(n15152), .ZN(n14948) );
  OAI22_X1 U16183 ( .A1(n15310), .A2(n15036), .B1(n15311), .B2(n16098), .ZN(
        n14947) );
  AOI211_X1 U16184 ( .C1(n15460), .C2(n15040), .A(n14948), .B(n14947), .ZN(
        n14949) );
  OAI21_X1 U16185 ( .B1(n14950), .B2(n15042), .A(n14949), .ZN(P1_U3219) );
  AOI22_X1 U16186 ( .A1(n15408), .A2(n14905), .B1(n9798), .B2(n15401), .ZN(
        n14957) );
  AOI22_X1 U16187 ( .A1(n15408), .A2(n9798), .B1(n14953), .B2(n15401), .ZN(
        n14955) );
  XNOR2_X1 U16188 ( .A(n14955), .B(n14954), .ZN(n14956) );
  OAI22_X1 U16189 ( .A1(n15190), .A2(n15049), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14959), .ZN(n14964) );
  INV_X1 U16190 ( .A(n14960), .ZN(n14961) );
  OAI22_X1 U16191 ( .A1(n14962), .A2(n15036), .B1(n16098), .B2(n14961), .ZN(
        n14963) );
  AOI211_X1 U16192 ( .C1(n15408), .C2(n15040), .A(n14964), .B(n14963), .ZN(
        n14965) );
  OAI21_X1 U16193 ( .B1(n14967), .B2(n7324), .A(n14966), .ZN(n14968) );
  NAND2_X1 U16194 ( .A1(n14968), .A2(n16093), .ZN(n14975) );
  OR2_X1 U16195 ( .A1(n14969), .A2(n15359), .ZN(n14971) );
  NAND2_X1 U16196 ( .A1(n15061), .A2(n16030), .ZN(n14970) );
  NAND2_X1 U16197 ( .A1(n14971), .A2(n14970), .ZN(n15277) );
  INV_X1 U16198 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14972) );
  OAI22_X1 U16199 ( .A1(n15270), .A2(n16098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14972), .ZN(n14973) );
  AOI21_X1 U16200 ( .B1(n15277), .B2(n15020), .A(n14973), .ZN(n14974) );
  OAI211_X1 U16201 ( .C1(n15273), .C2(n16091), .A(n14975), .B(n14974), .ZN(
        P1_U3223) );
  XOR2_X1 U16202 ( .A(n14977), .B(n14976), .Z(n14983) );
  NAND2_X1 U16203 ( .A1(n15059), .A2(n16030), .ZN(n14979) );
  NAND2_X1 U16204 ( .A1(n15057), .A2(n15376), .ZN(n14978) );
  AND2_X1 U16205 ( .A1(n14979), .A2(n14978), .ZN(n15204) );
  AOI22_X1 U16206 ( .A1(n14987), .A2(n15212), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14980) );
  OAI21_X1 U16207 ( .B1(n15204), .B2(n15026), .A(n14980), .ZN(n14981) );
  AOI21_X1 U16208 ( .B1(n15425), .B2(n15040), .A(n14981), .ZN(n14982) );
  OAI21_X1 U16209 ( .B1(n14983), .B2(n15042), .A(n14982), .ZN(P1_U3225) );
  AOI21_X1 U16210 ( .B1(n14986), .B2(n14984), .A(n14985), .ZN(n14992) );
  AOI22_X1 U16211 ( .A1(n14987), .A2(n15361), .B1(n16087), .B2(n16088), .ZN(
        n14989) );
  OAI211_X1 U16212 ( .C1(n15360), .C2(n15036), .A(n14989), .B(n14988), .ZN(
        n14990) );
  AOI21_X1 U16213 ( .B1(n16133), .B2(n15040), .A(n14990), .ZN(n14991) );
  OAI21_X1 U16214 ( .B1(n14992), .B2(n15042), .A(n14991), .ZN(P1_U3226) );
  XNOR2_X1 U16215 ( .A(n14994), .B(n14993), .ZN(n14995) );
  XNOR2_X1 U16216 ( .A(n14996), .B(n14995), .ZN(n15000) );
  NAND2_X1 U16217 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15114)
         );
  OAI21_X1 U16218 ( .B1(n15340), .B2(n15049), .A(n15114), .ZN(n14998) );
  OAI22_X1 U16219 ( .A1(n15341), .A2(n15036), .B1(n15342), .B2(n16098), .ZN(
        n14997) );
  AOI211_X1 U16220 ( .C1(n15474), .C2(n15040), .A(n14998), .B(n14997), .ZN(
        n14999) );
  OAI21_X1 U16221 ( .B1(n15000), .B2(n15042), .A(n14999), .ZN(P1_U3228) );
  INV_X1 U16222 ( .A(n15429), .ZN(n15232) );
  OAI21_X1 U16223 ( .B1(n15003), .B2(n15002), .A(n15001), .ZN(n15004) );
  NAND2_X1 U16224 ( .A1(n15004), .A2(n16093), .ZN(n15011) );
  NAND2_X1 U16225 ( .A1(n15257), .A2(n16030), .ZN(n15006) );
  NAND2_X1 U16226 ( .A1(n15058), .A2(n15376), .ZN(n15005) );
  NAND2_X1 U16227 ( .A1(n15006), .A2(n15005), .ZN(n15225) );
  INV_X1 U16228 ( .A(n15229), .ZN(n15008) );
  OAI22_X1 U16229 ( .A1(n16098), .A2(n15008), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15007), .ZN(n15009) );
  AOI21_X1 U16230 ( .B1(n15020), .B2(n15225), .A(n15009), .ZN(n15010) );
  OAI211_X1 U16231 ( .C1(n15232), .C2(n16091), .A(n15011), .B(n15010), .ZN(
        P1_U3229) );
  AOI211_X1 U16232 ( .C1(n15014), .C2(n15013), .A(n15042), .B(n15012), .ZN(
        n15015) );
  INV_X1 U16233 ( .A(n15015), .ZN(n15022) );
  NAND2_X1 U16234 ( .A1(n15259), .A2(n15376), .ZN(n15017) );
  NAND2_X1 U16235 ( .A1(n15062), .A2(n16030), .ZN(n15016) );
  NAND2_X1 U16236 ( .A1(n15017), .A2(n15016), .ZN(n15287) );
  OAI22_X1 U16237 ( .A1(n15295), .A2(n16098), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15018), .ZN(n15019) );
  AOI21_X1 U16238 ( .B1(n15287), .B2(n15020), .A(n15019), .ZN(n15021) );
  OAI211_X1 U16239 ( .C1(n15452), .C2(n16091), .A(n15022), .B(n15021), .ZN(
        P1_U3233) );
  AOI21_X1 U16240 ( .B1(n15025), .B2(n15024), .A(n15023), .ZN(n15030) );
  AOI22_X1 U16241 ( .A1(n15062), .A2(n15376), .B1(n16030), .B2(n15064), .ZN(
        n15324) );
  NOR2_X1 U16242 ( .A1(n15324), .A2(n15026), .ZN(n15028) );
  NAND2_X1 U16243 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15128)
         );
  OAI21_X1 U16244 ( .B1(n16098), .B2(n15328), .A(n15128), .ZN(n15027) );
  AOI211_X1 U16245 ( .C1(n15466), .C2(n15040), .A(n15028), .B(n15027), .ZN(
        n15029) );
  OAI21_X1 U16246 ( .B1(n15030), .B2(n15042), .A(n15029), .ZN(P1_U3238) );
  NAND2_X1 U16247 ( .A1(n15033), .A2(n15032), .ZN(n15034) );
  XNOR2_X1 U16248 ( .A(n15031), .B(n15034), .ZN(n15043) );
  OAI22_X1 U16249 ( .A1(n15190), .A2(n15036), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15035), .ZN(n15039) );
  INV_X1 U16250 ( .A(n15195), .ZN(n15037) );
  OAI22_X1 U16251 ( .A1(n15191), .A2(n15049), .B1(n16098), .B2(n15037), .ZN(
        n15038) );
  AOI211_X1 U16252 ( .C1(n15420), .C2(n15040), .A(n15039), .B(n15038), .ZN(
        n15041) );
  OAI21_X1 U16253 ( .B1(n15043), .B2(n15042), .A(n15041), .ZN(P1_U3240) );
  OAI211_X1 U16254 ( .C1(n15045), .C2(n15047), .A(n15046), .B(n16093), .ZN(
        n15054) );
  NAND2_X1 U16255 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15654)
         );
  INV_X1 U16256 ( .A(n15654), .ZN(n15052) );
  INV_X1 U16257 ( .A(n15048), .ZN(n15378) );
  OAI22_X1 U16258 ( .A1(n15050), .A2(n15049), .B1(n16098), .B2(n15378), .ZN(
        n15051) );
  AOI211_X1 U16259 ( .C1(n16089), .C2(n15375), .A(n15052), .B(n15051), .ZN(
        n15053) );
  OAI211_X1 U16260 ( .C1(n16124), .C2(n16091), .A(n15054), .B(n15053), .ZN(
        P1_U3241) );
  MUX2_X1 U16261 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n15155), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16262 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15400), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16263 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n15055), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16264 ( .A(n15401), .B(P1_DATAO_REG_28__SCAN_IN), .S(n15076), .Z(
        P1_U3588) );
  MUX2_X1 U16265 ( .A(n15056), .B(P1_DATAO_REG_27__SCAN_IN), .S(n15076), .Z(
        P1_U3587) );
  MUX2_X1 U16266 ( .A(n15057), .B(P1_DATAO_REG_26__SCAN_IN), .S(n15076), .Z(
        P1_U3586) );
  MUX2_X1 U16267 ( .A(n15058), .B(P1_DATAO_REG_25__SCAN_IN), .S(n15076), .Z(
        P1_U3585) );
  MUX2_X1 U16268 ( .A(n15059), .B(P1_DATAO_REG_24__SCAN_IN), .S(n15076), .Z(
        P1_U3584) );
  MUX2_X1 U16269 ( .A(n15257), .B(P1_DATAO_REG_23__SCAN_IN), .S(n15076), .Z(
        P1_U3583) );
  MUX2_X1 U16270 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15060), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16271 ( .A(n15259), .B(P1_DATAO_REG_21__SCAN_IN), .S(n15076), .Z(
        P1_U3581) );
  MUX2_X1 U16272 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15061), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16273 ( .A(n15062), .B(P1_DATAO_REG_19__SCAN_IN), .S(n15076), .Z(
        P1_U3579) );
  MUX2_X1 U16274 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15063), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16275 ( .A(n15064), .B(P1_DATAO_REG_17__SCAN_IN), .S(n15076), .Z(
        P1_U3577) );
  MUX2_X1 U16276 ( .A(n15375), .B(P1_DATAO_REG_16__SCAN_IN), .S(n15076), .Z(
        P1_U3576) );
  MUX2_X1 U16277 ( .A(n16088), .B(P1_DATAO_REG_15__SCAN_IN), .S(n15076), .Z(
        P1_U3575) );
  MUX2_X1 U16278 ( .A(n15374), .B(P1_DATAO_REG_14__SCAN_IN), .S(n15076), .Z(
        P1_U3574) );
  MUX2_X1 U16279 ( .A(n16086), .B(P1_DATAO_REG_13__SCAN_IN), .S(n15076), .Z(
        P1_U3573) );
  MUX2_X1 U16280 ( .A(n15065), .B(P1_DATAO_REG_12__SCAN_IN), .S(n15076), .Z(
        P1_U3572) );
  MUX2_X1 U16281 ( .A(n15066), .B(P1_DATAO_REG_11__SCAN_IN), .S(n15076), .Z(
        P1_U3571) );
  MUX2_X1 U16282 ( .A(n15067), .B(P1_DATAO_REG_10__SCAN_IN), .S(n15076), .Z(
        P1_U3570) );
  MUX2_X1 U16283 ( .A(n16029), .B(P1_DATAO_REG_9__SCAN_IN), .S(n15076), .Z(
        P1_U3569) );
  MUX2_X1 U16284 ( .A(n15068), .B(P1_DATAO_REG_8__SCAN_IN), .S(n15076), .Z(
        P1_U3568) );
  MUX2_X1 U16285 ( .A(n15069), .B(P1_DATAO_REG_7__SCAN_IN), .S(n15076), .Z(
        P1_U3567) );
  MUX2_X1 U16286 ( .A(n15070), .B(P1_DATAO_REG_6__SCAN_IN), .S(n15076), .Z(
        P1_U3566) );
  MUX2_X1 U16287 ( .A(n15071), .B(P1_DATAO_REG_5__SCAN_IN), .S(n15076), .Z(
        P1_U3565) );
  MUX2_X1 U16288 ( .A(n15072), .B(P1_DATAO_REG_4__SCAN_IN), .S(n15076), .Z(
        P1_U3564) );
  MUX2_X1 U16289 ( .A(n15073), .B(P1_DATAO_REG_3__SCAN_IN), .S(n15076), .Z(
        P1_U3563) );
  MUX2_X1 U16290 ( .A(n15074), .B(P1_DATAO_REG_2__SCAN_IN), .S(n15076), .Z(
        P1_U3562) );
  MUX2_X1 U16291 ( .A(n15075), .B(P1_DATAO_REG_1__SCAN_IN), .S(n15076), .Z(
        P1_U3561) );
  MUX2_X1 U16292 ( .A(n10907), .B(P1_DATAO_REG_0__SCAN_IN), .S(n15076), .Z(
        P1_U3560) );
  OAI21_X1 U16293 ( .B1(n15079), .B2(n15078), .A(n15077), .ZN(n15080) );
  NAND2_X1 U16294 ( .A1(n15080), .A2(n15652), .ZN(n15092) );
  AOI21_X1 U16295 ( .B1(n15639), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n15081), .ZN(
        n15091) );
  INV_X1 U16296 ( .A(n15082), .ZN(n15084) );
  MUX2_X1 U16297 ( .A(n11936), .B(P1_REG2_REG_9__SCAN_IN), .S(n15088), .Z(
        n15083) );
  NAND2_X1 U16298 ( .A1(n15084), .A2(n15083), .ZN(n15086) );
  OAI211_X1 U16299 ( .C1(n15087), .C2(n15086), .A(n15085), .B(n15143), .ZN(
        n15090) );
  NAND2_X1 U16300 ( .A1(n15147), .A2(n15088), .ZN(n15089) );
  NAND4_X1 U16301 ( .A1(n15092), .A2(n15091), .A3(n15090), .A4(n15089), .ZN(
        P1_U3252) );
  OAI211_X1 U16302 ( .C1(n15095), .C2(n15094), .A(n15093), .B(n15652), .ZN(
        n15104) );
  NOR2_X1 U16303 ( .A1(n15647), .A2(n15096), .ZN(n15097) );
  AOI211_X1 U16304 ( .C1(n15639), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n15098), 
        .B(n15097), .ZN(n15103) );
  OAI211_X1 U16305 ( .C1(n15101), .C2(n15100), .A(n15099), .B(n15143), .ZN(
        n15102) );
  NAND3_X1 U16306 ( .A1(n15104), .A2(n15103), .A3(n15102), .ZN(P1_U3256) );
  AOI21_X1 U16307 ( .B1(n15106), .B2(P1_REG1_REG_16__SCAN_IN), .A(n15105), 
        .ZN(n15108) );
  XNOR2_X1 U16308 ( .A(n15124), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n15107) );
  AOI211_X1 U16309 ( .C1(n15108), .C2(n15107), .A(n15145), .B(n15123), .ZN(
        n15119) );
  OAI21_X1 U16310 ( .B1(n15110), .B2(n12491), .A(n15109), .ZN(n15113) );
  INV_X1 U16311 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15121) );
  NOR2_X1 U16312 ( .A1(n15122), .A2(n15121), .ZN(n15111) );
  AOI21_X1 U16313 ( .B1(n15121), .B2(n15122), .A(n15111), .ZN(n15112) );
  NAND2_X1 U16314 ( .A1(n15112), .A2(n15113), .ZN(n15120) );
  OAI211_X1 U16315 ( .C1(n15113), .C2(n15112), .A(n15120), .B(n15143), .ZN(
        n15117) );
  INV_X1 U16316 ( .A(n15114), .ZN(n15115) );
  AOI21_X1 U16317 ( .B1(n15639), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n15115), 
        .ZN(n15116) );
  OAI211_X1 U16318 ( .C1(n15647), .C2(n15122), .A(n15117), .B(n15116), .ZN(
        n15118) );
  OR2_X1 U16319 ( .A1(n15119), .A2(n15118), .ZN(P1_U3260) );
  OAI21_X1 U16320 ( .B1(n15122), .B2(n15121), .A(n15120), .ZN(n15139) );
  XNOR2_X1 U16321 ( .A(n15139), .B(n15125), .ZN(n15137) );
  XNOR2_X1 U16322 ( .A(n15137), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n15133) );
  AND2_X1 U16323 ( .A1(n15127), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n15135) );
  INV_X1 U16324 ( .A(n15135), .ZN(n15126) );
  OAI211_X1 U16325 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n15127), .A(n15126), 
        .B(n15652), .ZN(n15132) );
  INV_X1 U16326 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15129) );
  OAI21_X1 U16327 ( .B1(n15656), .B2(n15129), .A(n15128), .ZN(n15130) );
  AOI21_X1 U16328 ( .B1(n15138), .B2(n15147), .A(n15130), .ZN(n15131) );
  OAI211_X1 U16329 ( .C1(n15133), .C2(n15649), .A(n15132), .B(n15131), .ZN(
        P1_U3261) );
  NOR2_X1 U16330 ( .A1(n15135), .A2(n15134), .ZN(n15136) );
  XNOR2_X1 U16331 ( .A(n15136), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n15146) );
  NAND2_X1 U16332 ( .A1(n15137), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n15141) );
  NAND2_X1 U16333 ( .A1(n15139), .A2(n15138), .ZN(n15140) );
  NAND2_X1 U16334 ( .A1(n15141), .A2(n15140), .ZN(n15142) );
  XOR2_X1 U16335 ( .A(n15142), .B(P1_REG2_REG_19__SCAN_IN), .Z(n15144) );
  AOI22_X1 U16336 ( .A1(n15146), .A2(n15652), .B1(n15143), .B2(n15144), .ZN(
        n15151) );
  INV_X1 U16337 ( .A(n15144), .ZN(n15148) );
  NAND2_X1 U16338 ( .A1(n15633), .A2(P1_B_REG_SCAN_IN), .ZN(n15154) );
  AND2_X1 U16339 ( .A1(n15376), .A2(n15154), .ZN(n15399) );
  NAND2_X1 U16340 ( .A1(n15155), .A2(n15399), .ZN(n15395) );
  NOR2_X1 U16341 ( .A1(n15395), .A2(n16001), .ZN(n15161) );
  NOR2_X1 U16342 ( .A1(n7734), .A2(n15365), .ZN(n15157) );
  AOI211_X1 U16343 ( .C1(n16001), .C2(P1_REG2_REG_31__SCAN_IN), .A(n15161), 
        .B(n15157), .ZN(n15158) );
  OAI21_X1 U16344 ( .B1(n15993), .B2(n15394), .A(n15158), .ZN(P1_U3263) );
  OAI211_X1 U16345 ( .C1(n15165), .C2(n15397), .A(n15445), .B(n15159), .ZN(
        n15396) );
  NOR2_X1 U16346 ( .A1(n15397), .A2(n15365), .ZN(n15160) );
  AOI211_X1 U16347 ( .C1(n16001), .C2(P1_REG2_REG_30__SCAN_IN), .A(n15161), 
        .B(n15160), .ZN(n15162) );
  OAI21_X1 U16348 ( .B1(n15993), .B2(n15396), .A(n15162), .ZN(P1_U3264) );
  NAND2_X1 U16349 ( .A1(n15408), .A2(n15401), .ZN(n15163) );
  AOI211_X1 U16350 ( .C1(n15167), .C2(n15166), .A(n15974), .B(n15165), .ZN(
        n15405) );
  NOR2_X1 U16351 ( .A1(n15403), .A2(n15365), .ZN(n15175) );
  AOI22_X1 U16352 ( .A1(n16001), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n15168), 
        .B2(n15990), .ZN(n15172) );
  INV_X1 U16353 ( .A(n15169), .ZN(n15170) );
  NAND3_X1 U16354 ( .A1(n15400), .A2(n15399), .A3(n15170), .ZN(n15171) );
  OAI211_X1 U16355 ( .C1(n15173), .C2(n15177), .A(n15172), .B(n15171), .ZN(
        n15174) );
  AOI211_X1 U16356 ( .C1(n15405), .C2(n15368), .A(n15175), .B(n15174), .ZN(
        n15185) );
  NAND2_X1 U16357 ( .A1(n15408), .A2(n15177), .ZN(n15178) );
  NAND2_X1 U16358 ( .A1(n15179), .A2(n15178), .ZN(n15181) );
  NAND2_X1 U16359 ( .A1(n15181), .A2(n15180), .ZN(n15183) );
  NAND2_X1 U16360 ( .A1(n15398), .A2(n15389), .ZN(n15184) );
  OAI211_X1 U16361 ( .C1(n15407), .C2(n15392), .A(n15185), .B(n15184), .ZN(
        P1_U3356) );
  XNOR2_X1 U16362 ( .A(n15186), .B(n15187), .ZN(n15421) );
  XNOR2_X1 U16363 ( .A(n15188), .B(n15187), .ZN(n15189) );
  OAI222_X1 U16364 ( .A1(n15357), .A2(n15191), .B1(n15359), .B2(n15190), .C1(
        n16136), .C2(n15189), .ZN(n15418) );
  INV_X1 U16365 ( .A(n15211), .ZN(n15194) );
  INV_X1 U16366 ( .A(n15192), .ZN(n15193) );
  AOI211_X1 U16367 ( .C1(n15420), .C2(n15194), .A(n15974), .B(n15193), .ZN(
        n15419) );
  NAND2_X1 U16368 ( .A1(n15419), .A2(n15368), .ZN(n15197) );
  AOI22_X1 U16369 ( .A1(n16001), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n15195), 
        .B2(n15990), .ZN(n15196) );
  OAI211_X1 U16370 ( .C1(n15198), .C2(n15365), .A(n15197), .B(n15196), .ZN(
        n15199) );
  AOI21_X1 U16371 ( .B1(n15418), .B2(n7218), .A(n15199), .ZN(n15200) );
  OAI21_X1 U16372 ( .B1(n15421), .B2(n15392), .A(n15200), .ZN(P1_U3267) );
  OAI21_X1 U16373 ( .B1(n15205), .B2(n16136), .A(n15204), .ZN(n15423) );
  INV_X1 U16374 ( .A(n15423), .ZN(n15218) );
  AOI21_X1 U16375 ( .B1(n15208), .B2(n15207), .A(n15206), .ZN(n15422) );
  INV_X1 U16376 ( .A(n15425), .ZN(n15215) );
  NAND2_X1 U16377 ( .A1(n15425), .A2(n15228), .ZN(n15209) );
  NAND2_X1 U16378 ( .A1(n15209), .A2(n15445), .ZN(n15210) );
  NOR2_X1 U16379 ( .A1(n15211), .A2(n15210), .ZN(n15424) );
  NAND2_X1 U16380 ( .A1(n15424), .A2(n15368), .ZN(n15214) );
  AOI22_X1 U16381 ( .A1(n16001), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n15212), 
        .B2(n15990), .ZN(n15213) );
  OAI211_X1 U16382 ( .C1(n15215), .C2(n15365), .A(n15214), .B(n15213), .ZN(
        n15216) );
  AOI21_X1 U16383 ( .B1(n15422), .B2(n15355), .A(n15216), .ZN(n15217) );
  OAI21_X1 U16384 ( .B1(n15218), .B2(n16001), .A(n15217), .ZN(P1_U3268) );
  OAI21_X1 U16385 ( .B1(n7346), .B2(n15220), .A(n15219), .ZN(n15221) );
  INV_X1 U16386 ( .A(n15221), .ZN(n15431) );
  OAI211_X1 U16387 ( .C1(n15224), .C2(n15223), .A(n15222), .B(n16119), .ZN(
        n15227) );
  INV_X1 U16388 ( .A(n15225), .ZN(n15226) );
  NAND2_X1 U16389 ( .A1(n15227), .A2(n15226), .ZN(n15427) );
  AOI211_X1 U16390 ( .C1(n15429), .C2(n15242), .A(n15974), .B(n7735), .ZN(
        n15428) );
  NAND2_X1 U16391 ( .A1(n15428), .A2(n15368), .ZN(n15231) );
  AOI22_X1 U16392 ( .A1(n16001), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n15229), 
        .B2(n15990), .ZN(n15230) );
  OAI211_X1 U16393 ( .C1(n15232), .C2(n15365), .A(n15231), .B(n15230), .ZN(
        n15233) );
  AOI21_X1 U16394 ( .B1(n15427), .B2(n7218), .A(n15233), .ZN(n15234) );
  OAI21_X1 U16395 ( .B1(n15431), .B2(n15392), .A(n15234), .ZN(P1_U3269) );
  XNOR2_X1 U16396 ( .A(n15235), .B(n7923), .ZN(n15237) );
  AOI21_X1 U16397 ( .B1(n15237), .B2(n16119), .A(n15236), .ZN(n15435) );
  OAI21_X1 U16398 ( .B1(n15238), .B2(n15377), .A(n15435), .ZN(n15247) );
  AOI21_X1 U16399 ( .B1(n7923), .B2(n15240), .A(n15239), .ZN(n15241) );
  INV_X1 U16400 ( .A(n15241), .ZN(n15436) );
  AOI22_X1 U16401 ( .A1(n15433), .A2(n15991), .B1(n16001), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n15245) );
  AOI21_X1 U16402 ( .B1(n15433), .B2(n15256), .A(n15974), .ZN(n15243) );
  AND2_X1 U16403 ( .A1(n15243), .A2(n15242), .ZN(n15432) );
  NAND2_X1 U16404 ( .A1(n15432), .A2(n15368), .ZN(n15244) );
  OAI211_X1 U16405 ( .C1(n15436), .C2(n15392), .A(n15245), .B(n15244), .ZN(
        n15246) );
  AOI21_X1 U16406 ( .B1(n7218), .B2(n15247), .A(n15246), .ZN(n15248) );
  INV_X1 U16407 ( .A(n15248), .ZN(P1_U3270) );
  OAI21_X1 U16408 ( .B1(n15251), .B2(n15250), .A(n15249), .ZN(n15252) );
  INV_X1 U16409 ( .A(n15252), .ZN(n15443) );
  OAI21_X1 U16410 ( .B1(n15255), .B2(n15254), .A(n15253), .ZN(n15441) );
  OAI211_X1 U16411 ( .C1(n15439), .C2(n15269), .A(n15445), .B(n15256), .ZN(
        n15438) );
  NOR2_X1 U16412 ( .A1(n15438), .A2(n15993), .ZN(n15266) );
  AND2_X1 U16413 ( .A1(n15257), .A2(n15376), .ZN(n15258) );
  AOI21_X1 U16414 ( .B1(n15259), .B2(n16030), .A(n15258), .ZN(n15437) );
  INV_X1 U16415 ( .A(n15437), .ZN(n15263) );
  INV_X1 U16416 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n15260) );
  OAI22_X1 U16417 ( .A1(n15261), .A2(n15377), .B1(n15260), .B2(n7218), .ZN(
        n15262) );
  AOI21_X1 U16418 ( .B1(n15263), .B2(n7218), .A(n15262), .ZN(n15264) );
  OAI21_X1 U16419 ( .B1(n15439), .B2(n15365), .A(n15264), .ZN(n15265) );
  AOI211_X1 U16420 ( .C1(n15441), .C2(n15389), .A(n15266), .B(n15265), .ZN(
        n15267) );
  OAI21_X1 U16421 ( .B1(n15443), .B2(n15392), .A(n15267), .ZN(P1_U3271) );
  XNOR2_X1 U16422 ( .A(n15268), .B(n15276), .ZN(n15449) );
  AOI21_X1 U16423 ( .B1(n15444), .B2(n7357), .A(n15269), .ZN(n15446) );
  INV_X1 U16424 ( .A(n15270), .ZN(n15271) );
  AOI22_X1 U16425 ( .A1(n15271), .A2(n15990), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n16001), .ZN(n15272) );
  OAI21_X1 U16426 ( .B1(n15273), .B2(n15365), .A(n15272), .ZN(n15280) );
  AOI211_X1 U16427 ( .C1(n15276), .C2(n15275), .A(n16136), .B(n15274), .ZN(
        n15278) );
  NOR2_X1 U16428 ( .A1(n15278), .A2(n15277), .ZN(n15448) );
  NOR2_X1 U16429 ( .A1(n15448), .A2(n16001), .ZN(n15279) );
  AOI211_X1 U16430 ( .C1(n15446), .C2(n15347), .A(n15280), .B(n15279), .ZN(
        n15281) );
  OAI21_X1 U16431 ( .B1(n15449), .B2(n15392), .A(n15281), .ZN(P1_U3272) );
  NAND2_X1 U16432 ( .A1(n15283), .A2(n15282), .ZN(n15284) );
  NAND2_X1 U16433 ( .A1(n15284), .A2(n16119), .ZN(n15285) );
  OR2_X1 U16434 ( .A1(n15286), .A2(n15285), .ZN(n15289) );
  INV_X1 U16435 ( .A(n15287), .ZN(n15288) );
  NAND2_X1 U16436 ( .A1(n15291), .A2(n15290), .ZN(n15292) );
  AND2_X1 U16437 ( .A1(n15293), .A2(n15292), .ZN(n15454) );
  NAND2_X1 U16438 ( .A1(n15454), .A2(n15355), .ZN(n15301) );
  INV_X1 U16439 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n15294) );
  OAI22_X1 U16440 ( .A1(n15295), .A2(n15377), .B1(n15294), .B2(n7218), .ZN(
        n15298) );
  AOI21_X1 U16441 ( .B1(n15309), .B2(n15299), .A(n15974), .ZN(n15296) );
  NAND2_X1 U16442 ( .A1(n7357), .A2(n15296), .ZN(n15450) );
  NOR2_X1 U16443 ( .A1(n15450), .A2(n15993), .ZN(n15297) );
  AOI211_X1 U16444 ( .C1(n15991), .C2(n15299), .A(n15298), .B(n15297), .ZN(
        n15300) );
  OAI211_X1 U16445 ( .C1(n16001), .C2(n15451), .A(n15301), .B(n15300), .ZN(
        P1_U3273) );
  OAI21_X1 U16446 ( .B1(n15304), .B2(n15303), .A(n15302), .ZN(n15305) );
  INV_X1 U16447 ( .A(n15305), .ZN(n15463) );
  OAI21_X1 U16448 ( .B1(n15308), .B2(n15307), .A(n15306), .ZN(n15457) );
  NAND2_X1 U16449 ( .A1(n15457), .A2(n15355), .ZN(n15318) );
  AOI211_X1 U16450 ( .C1(n15460), .C2(n15326), .A(n15974), .B(n7743), .ZN(
        n15458) );
  INV_X1 U16451 ( .A(n15460), .ZN(n15315) );
  OAI22_X1 U16452 ( .A1(n15310), .A2(n15359), .B1(n15341), .B2(n15357), .ZN(
        n15459) );
  OAI22_X1 U16453 ( .A1(n15312), .A2(n7218), .B1(n15311), .B2(n15377), .ZN(
        n15313) );
  AOI21_X1 U16454 ( .B1(n15459), .B2(n7218), .A(n15313), .ZN(n15314) );
  OAI21_X1 U16455 ( .B1(n15315), .B2(n15365), .A(n15314), .ZN(n15316) );
  AOI21_X1 U16456 ( .B1(n15458), .B2(n15368), .A(n15316), .ZN(n15317) );
  OAI211_X1 U16457 ( .C1(n15463), .C2(n15371), .A(n15318), .B(n15317), .ZN(
        P1_U3274) );
  XNOR2_X1 U16458 ( .A(n15320), .B(n15319), .ZN(n15468) );
  OAI211_X1 U16459 ( .C1(n15323), .C2(n15322), .A(n16119), .B(n15321), .ZN(
        n15325) );
  NAND2_X1 U16460 ( .A1(n15325), .A2(n15324), .ZN(n15464) );
  INV_X1 U16461 ( .A(n15466), .ZN(n15332) );
  INV_X1 U16462 ( .A(n15326), .ZN(n15327) );
  AOI211_X1 U16463 ( .C1(n15466), .C2(n15339), .A(n15974), .B(n15327), .ZN(
        n15465) );
  NAND2_X1 U16464 ( .A1(n15465), .A2(n15368), .ZN(n15331) );
  INV_X1 U16465 ( .A(n15328), .ZN(n15329) );
  AOI22_X1 U16466 ( .A1(n15329), .A2(n15990), .B1(n16001), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n15330) );
  OAI211_X1 U16467 ( .C1(n15332), .C2(n15365), .A(n15331), .B(n15330), .ZN(
        n15333) );
  AOI21_X1 U16468 ( .B1(n15464), .B2(n7218), .A(n15333), .ZN(n15334) );
  OAI21_X1 U16469 ( .B1(n15468), .B2(n15392), .A(n15334), .ZN(P1_U3275) );
  XOR2_X1 U16470 ( .A(n15335), .B(n15338), .Z(n15477) );
  NAND2_X1 U16471 ( .A1(n15337), .A2(n15338), .ZN(n15470) );
  NAND3_X1 U16472 ( .A1(n15336), .A2(n15470), .A3(n15355), .ZN(n15350) );
  OAI21_X1 U16473 ( .B1(n7271), .B2(n15345), .A(n15339), .ZN(n15471) );
  INV_X1 U16474 ( .A(n15471), .ZN(n15348) );
  OAI22_X1 U16475 ( .A1(n15341), .A2(n15359), .B1(n15340), .B2(n15357), .ZN(
        n15473) );
  OAI22_X1 U16476 ( .A1(n7218), .A2(n15121), .B1(n15342), .B2(n15377), .ZN(
        n15343) );
  AOI21_X1 U16477 ( .B1(n15473), .B2(n7218), .A(n15343), .ZN(n15344) );
  OAI21_X1 U16478 ( .B1(n15345), .B2(n15365), .A(n15344), .ZN(n15346) );
  AOI21_X1 U16479 ( .B1(n15348), .B2(n15347), .A(n15346), .ZN(n15349) );
  OAI211_X1 U16480 ( .C1(n15477), .C2(n15371), .A(n15350), .B(n15349), .ZN(
        P1_U3276) );
  XNOR2_X1 U16481 ( .A(n15352), .B(n15351), .ZN(n16137) );
  XNOR2_X1 U16482 ( .A(n15354), .B(n15353), .ZN(n16140) );
  NAND2_X1 U16483 ( .A1(n16140), .A2(n15355), .ZN(n15370) );
  OAI21_X1 U16484 ( .B1(n15382), .B2(n15366), .A(n15445), .ZN(n15356) );
  NOR2_X1 U16485 ( .A1(n15356), .A2(n7271), .ZN(n16131) );
  OAI22_X1 U16486 ( .A1(n15360), .A2(n15359), .B1(n15358), .B2(n15357), .ZN(
        n16132) );
  AOI21_X1 U16487 ( .B1(n15361), .B2(n15990), .A(n16132), .ZN(n15362) );
  NOR2_X1 U16488 ( .A1(n15362), .A2(n16001), .ZN(n15363) );
  AOI21_X1 U16489 ( .B1(n16001), .B2(P1_REG2_REG_16__SCAN_IN), .A(n15363), 
        .ZN(n15364) );
  OAI21_X1 U16490 ( .B1(n15366), .B2(n15365), .A(n15364), .ZN(n15367) );
  AOI21_X1 U16491 ( .B1(n16131), .B2(n15368), .A(n15367), .ZN(n15369) );
  OAI211_X1 U16492 ( .C1(n16137), .C2(n15371), .A(n15370), .B(n15369), .ZN(
        P1_U3277) );
  OAI21_X1 U16493 ( .B1(n15373), .B2(n15387), .A(n15372), .ZN(n16127) );
  INV_X1 U16494 ( .A(n16127), .ZN(n15393) );
  AOI22_X1 U16495 ( .A1(n15376), .A2(n15375), .B1(n15374), .B2(n16030), .ZN(
        n16121) );
  OAI21_X1 U16496 ( .B1(n15378), .B2(n15377), .A(n16121), .ZN(n15379) );
  MUX2_X1 U16497 ( .A(P1_REG2_REG_15__SCAN_IN), .B(n15379), .S(n7218), .Z(
        n15385) );
  NAND2_X1 U16498 ( .A1(n15386), .A2(n15380), .ZN(n15381) );
  NAND2_X1 U16499 ( .A1(n15381), .A2(n15445), .ZN(n15383) );
  OR2_X1 U16500 ( .A1(n15383), .A2(n15382), .ZN(n16122) );
  NOR2_X1 U16501 ( .A1(n16122), .A2(n15993), .ZN(n15384) );
  AOI211_X1 U16502 ( .C1(n15991), .C2(n15386), .A(n15385), .B(n15384), .ZN(
        n15391) );
  NAND2_X1 U16503 ( .A1(n15388), .A2(n15387), .ZN(n16118) );
  NAND3_X1 U16504 ( .A1(n16120), .A2(n16118), .A3(n15389), .ZN(n15390) );
  OAI211_X1 U16505 ( .C1(n15393), .C2(n15392), .A(n15391), .B(n15390), .ZN(
        P1_U3278) );
  OAI211_X1 U16506 ( .C1(n7734), .C2(n16123), .A(n15394), .B(n15395), .ZN(
        n15478) );
  MUX2_X1 U16507 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15478), .S(n16143), .Z(
        P1_U3559) );
  OAI211_X1 U16508 ( .C1(n15397), .C2(n16123), .A(n15396), .B(n15395), .ZN(
        n15479) );
  MUX2_X1 U16509 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15479), .S(n16143), .Z(
        P1_U3558) );
  AOI22_X1 U16510 ( .A1(n16030), .A2(n15401), .B1(n15400), .B2(n15399), .ZN(
        n15402) );
  OAI21_X1 U16511 ( .B1(n15403), .B2(n16123), .A(n15402), .ZN(n15404) );
  MUX2_X1 U16512 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15480), .S(n16143), .Z(
        P1_U3557) );
  AOI22_X1 U16513 ( .A1(n15409), .A2(n15445), .B1(n16134), .B2(n15408), .ZN(
        n15410) );
  OAI211_X1 U16514 ( .C1(n15469), .C2(n15412), .A(n15411), .B(n15410), .ZN(
        n15481) );
  MUX2_X1 U16515 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15481), .S(n16143), .Z(
        P1_U3556) );
  AOI22_X1 U16516 ( .A1(n15414), .A2(n15445), .B1(n16134), .B2(n15413), .ZN(
        n15415) );
  OAI211_X1 U16517 ( .C1(n15417), .C2(n16021), .A(n15416), .B(n15415), .ZN(
        n15482) );
  MUX2_X1 U16518 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15482), .S(n16143), .Z(
        P1_U3555) );
  MUX2_X1 U16519 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15483), .S(n16143), .Z(
        P1_U3554) );
  INV_X1 U16520 ( .A(n15422), .ZN(n15426) );
  MUX2_X1 U16521 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n7333), .S(n16143), .Z(
        P1_U3553) );
  AOI211_X1 U16522 ( .C1(n16134), .C2(n15429), .A(n15428), .B(n15427), .ZN(
        n15430) );
  OAI21_X1 U16523 ( .B1(n15469), .B2(n15431), .A(n15430), .ZN(n15484) );
  MUX2_X1 U16524 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15484), .S(n16143), .Z(
        P1_U3552) );
  AOI21_X1 U16525 ( .B1(n16134), .B2(n15433), .A(n15432), .ZN(n15434) );
  OAI211_X1 U16526 ( .C1(n15436), .C2(n15469), .A(n15435), .B(n15434), .ZN(
        n15485) );
  MUX2_X1 U16527 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15485), .S(n16143), .Z(
        P1_U3551) );
  OAI211_X1 U16528 ( .C1(n16123), .C2(n15439), .A(n15438), .B(n15437), .ZN(
        n15440) );
  AOI21_X1 U16529 ( .B1(n15441), .B2(n16119), .A(n15440), .ZN(n15442) );
  OAI21_X1 U16530 ( .B1(n15469), .B2(n15443), .A(n15442), .ZN(n15486) );
  MUX2_X1 U16531 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15486), .S(n16143), .Z(
        P1_U3550) );
  AOI22_X1 U16532 ( .A1(n15446), .A2(n15445), .B1(n16134), .B2(n15444), .ZN(
        n15447) );
  OAI211_X1 U16533 ( .C1(n15469), .C2(n15449), .A(n15448), .B(n15447), .ZN(
        n15487) );
  MUX2_X1 U16534 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15487), .S(n16143), .Z(
        P1_U3549) );
  INV_X1 U16535 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n15455) );
  OAI211_X1 U16536 ( .C1(n15452), .C2(n16123), .A(n15451), .B(n15450), .ZN(
        n15453) );
  AOI21_X1 U16537 ( .B1(n15454), .B2(n16139), .A(n15453), .ZN(n15488) );
  MUX2_X1 U16538 ( .A(n15455), .B(n15488), .S(n16143), .Z(n15456) );
  INV_X1 U16539 ( .A(n15456), .ZN(P1_U3548) );
  NAND2_X1 U16540 ( .A1(n15457), .A2(n16139), .ZN(n15462) );
  AOI211_X1 U16541 ( .C1(n16134), .C2(n15460), .A(n15459), .B(n15458), .ZN(
        n15461) );
  OAI211_X1 U16542 ( .C1(n16136), .C2(n15463), .A(n15462), .B(n15461), .ZN(
        n15491) );
  MUX2_X1 U16543 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15491), .S(n16143), .Z(
        P1_U3547) );
  AOI211_X1 U16544 ( .C1(n16134), .C2(n15466), .A(n15465), .B(n15464), .ZN(
        n15467) );
  OAI21_X1 U16545 ( .B1(n15469), .B2(n15468), .A(n15467), .ZN(n15492) );
  MUX2_X1 U16546 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15492), .S(n16143), .Z(
        P1_U3546) );
  NAND3_X1 U16547 ( .A1(n15336), .A2(n16139), .A3(n15470), .ZN(n15476) );
  NOR2_X1 U16548 ( .A1(n15471), .A2(n15974), .ZN(n15472) );
  AOI211_X1 U16549 ( .C1(n16134), .C2(n15474), .A(n15473), .B(n15472), .ZN(
        n15475) );
  OAI211_X1 U16550 ( .C1(n16136), .C2(n15477), .A(n15476), .B(n15475), .ZN(
        n15493) );
  MUX2_X1 U16551 ( .A(n15493), .B(P1_REG1_REG_17__SCAN_IN), .S(n16141), .Z(
        P1_U3545) );
  MUX2_X1 U16552 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15478), .S(n16147), .Z(
        P1_U3527) );
  MUX2_X1 U16553 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15479), .S(n16147), .Z(
        P1_U3526) );
  MUX2_X1 U16554 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15480), .S(n16147), .Z(
        P1_U3525) );
  MUX2_X1 U16555 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15481), .S(n16147), .Z(
        P1_U3524) );
  MUX2_X1 U16556 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15482), .S(n16147), .Z(
        P1_U3523) );
  MUX2_X1 U16557 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15483), .S(n16147), .Z(
        P1_U3522) );
  MUX2_X1 U16558 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n7333), .S(n16147), .Z(
        P1_U3521) );
  MUX2_X1 U16559 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15484), .S(n16147), .Z(
        P1_U3520) );
  MUX2_X1 U16560 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15485), .S(n16147), .Z(
        P1_U3519) );
  MUX2_X1 U16561 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15486), .S(n16147), .Z(
        P1_U3518) );
  MUX2_X1 U16562 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15487), .S(n16147), .Z(
        P1_U3517) );
  INV_X1 U16563 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15489) );
  MUX2_X1 U16564 ( .A(n15489), .B(n15488), .S(n16147), .Z(n15490) );
  INV_X1 U16565 ( .A(n15490), .ZN(P1_U3516) );
  MUX2_X1 U16566 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15491), .S(n16147), .Z(
        P1_U3515) );
  MUX2_X1 U16567 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15492), .S(n16147), .Z(
        P1_U3513) );
  MUX2_X1 U16568 ( .A(n15493), .B(P1_REG0_REG_17__SCAN_IN), .S(n16144), .Z(
        P1_U3510) );
  MUX2_X1 U16570 ( .A(n15496), .B(P1_D_REG_1__SCAN_IN), .S(n7198), .Z(P1_U3446) );
  MUX2_X1 U16571 ( .A(n15497), .B(P1_D_REG_0__SCAN_IN), .S(n7198), .Z(P1_U3445) );
  INV_X1 U16572 ( .A(n15498), .ZN(n15499) );
  NOR4_X1 U16573 ( .A1(n15499), .A2(P1_IR_REG_30__SCAN_IN), .A3(n15501), .A4(
        P1_U3086), .ZN(n15502) );
  AOI21_X1 U16574 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n15503), .A(n15502), 
        .ZN(n15504) );
  OAI21_X1 U16575 ( .B1(n15505), .B2(n15510), .A(n15504), .ZN(P1_U3324) );
  OAI222_X1 U16576 ( .A1(n15512), .A2(n15507), .B1(n7201), .B2(n9771), .C1(
        n15510), .C2(n15506), .ZN(P1_U3326) );
  OAI222_X1 U16577 ( .A1(n15512), .A2(n15511), .B1(n15510), .B2(n15509), .C1(
        n15508), .C2(P1_U3086), .ZN(P1_U3328) );
  MUX2_X1 U16578 ( .A(n15514), .B(n15513), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16579 ( .A(n15515), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U16580 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n7198), .ZN(P1_U3323) );
  AND2_X1 U16581 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n7198), .ZN(P1_U3322) );
  AND2_X1 U16582 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n7198), .ZN(P1_U3321) );
  AND2_X1 U16583 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n7198), .ZN(P1_U3320) );
  AND2_X1 U16584 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n7198), .ZN(P1_U3319) );
  AND2_X1 U16585 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n7198), .ZN(P1_U3318) );
  AND2_X1 U16586 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n7198), .ZN(P1_U3317) );
  AND2_X1 U16587 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n7198), .ZN(P1_U3316) );
  AND2_X1 U16588 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n7198), .ZN(P1_U3315) );
  AND2_X1 U16589 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n7198), .ZN(P1_U3314) );
  AND2_X1 U16590 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n7198), .ZN(P1_U3313) );
  AND2_X1 U16591 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n7198), .ZN(P1_U3312) );
  AND2_X1 U16592 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n7198), .ZN(P1_U3311) );
  AND2_X1 U16593 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n7198), .ZN(P1_U3310) );
  AND2_X1 U16594 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n7198), .ZN(P1_U3309) );
  AND2_X1 U16595 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n7198), .ZN(P1_U3308) );
  AND2_X1 U16596 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n7198), .ZN(P1_U3307) );
  AND2_X1 U16597 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n7198), .ZN(P1_U3306) );
  AND2_X1 U16598 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n7198), .ZN(P1_U3305) );
  AND2_X1 U16599 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n7198), .ZN(P1_U3304) );
  AND2_X1 U16600 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n7198), .ZN(P1_U3303) );
  AND2_X1 U16601 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n7198), .ZN(P1_U3302) );
  AND2_X1 U16602 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n7198), .ZN(P1_U3301) );
  AND2_X1 U16603 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n7198), .ZN(P1_U3300) );
  AND2_X1 U16604 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n7198), .ZN(P1_U3299) );
  AND2_X1 U16605 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n7198), .ZN(P1_U3298) );
  AND2_X1 U16606 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n7198), .ZN(P1_U3297) );
  AND2_X1 U16607 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n7198), .ZN(P1_U3296) );
  AND2_X1 U16608 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n7198), .ZN(P1_U3295) );
  AND2_X1 U16609 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n7198), .ZN(P1_U3294) );
  INV_X1 U16610 ( .A(n15525), .ZN(n15522) );
  AOI21_X1 U16611 ( .B1(n15518), .B2(n15522), .A(n15517), .ZN(P2_U3417) );
  AND2_X1 U16612 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15520), .ZN(P2_U3295) );
  AND2_X1 U16613 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15520), .ZN(P2_U3294) );
  AND2_X1 U16614 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15520), .ZN(P2_U3293) );
  AND2_X1 U16615 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15520), .ZN(P2_U3292) );
  AND2_X1 U16616 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15520), .ZN(P2_U3291) );
  AND2_X1 U16617 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15520), .ZN(P2_U3290) );
  AND2_X1 U16618 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15520), .ZN(P2_U3289) );
  AND2_X1 U16619 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15520), .ZN(P2_U3288) );
  AND2_X1 U16620 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15520), .ZN(P2_U3287) );
  AND2_X1 U16621 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15520), .ZN(P2_U3286) );
  AND2_X1 U16622 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15520), .ZN(P2_U3285) );
  AND2_X1 U16623 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15520), .ZN(P2_U3284) );
  AND2_X1 U16624 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15520), .ZN(P2_U3283) );
  AND2_X1 U16625 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15520), .ZN(P2_U3282) );
  AND2_X1 U16626 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15520), .ZN(P2_U3281) );
  AND2_X1 U16627 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15520), .ZN(P2_U3280) );
  AND2_X1 U16628 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15520), .ZN(P2_U3279) );
  AND2_X1 U16629 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15520), .ZN(P2_U3278) );
  AND2_X1 U16630 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15520), .ZN(P2_U3277) );
  AND2_X1 U16631 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15520), .ZN(P2_U3276) );
  AND2_X1 U16632 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15520), .ZN(P2_U3275) );
  AND2_X1 U16633 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15520), .ZN(P2_U3274) );
  AND2_X1 U16634 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15520), .ZN(P2_U3273) );
  AND2_X1 U16635 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15520), .ZN(P2_U3272) );
  AND2_X1 U16636 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15520), .ZN(P2_U3271) );
  AND2_X1 U16637 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15520), .ZN(P2_U3270) );
  AND2_X1 U16638 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15520), .ZN(P2_U3269) );
  AND2_X1 U16639 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15520), .ZN(P2_U3268) );
  AND2_X1 U16640 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15520), .ZN(P2_U3267) );
  AND2_X1 U16641 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15520), .ZN(P2_U3266) );
  NOR2_X1 U16642 ( .A1(n15619), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16643 ( .A1(P3_U3897), .A2(n15521), .ZN(P3_U3150) );
  AOI22_X1 U16644 ( .A1(n15525), .A2(n15524), .B1(n15523), .B2(n15522), .ZN(
        P2_U3416) );
  AOI22_X1 U16645 ( .A1(n15619), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n15539) );
  OAI21_X1 U16646 ( .B1(n15528), .B2(n15527), .A(n15526), .ZN(n15532) );
  NAND3_X1 U16647 ( .A1(n15530), .A2(n15529), .A3(n9707), .ZN(n15531) );
  OAI21_X1 U16648 ( .B1(n15622), .B2(n15532), .A(n15531), .ZN(n15533) );
  INV_X1 U16649 ( .A(n15533), .ZN(n15538) );
  OAI211_X1 U16650 ( .C1(n15536), .C2(n15535), .A(n15611), .B(n15534), .ZN(
        n15537) );
  NAND3_X1 U16651 ( .A1(n15539), .A2(n15538), .A3(n15537), .ZN(P2_U3215) );
  AOI22_X1 U16652 ( .A1(n15619), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15552) );
  OAI21_X1 U16653 ( .B1(n15542), .B2(n15541), .A(n15540), .ZN(n15545) );
  OAI22_X1 U16654 ( .A1(n15622), .A2(n15545), .B1(n15544), .B2(n15543), .ZN(
        n15546) );
  INV_X1 U16655 ( .A(n15546), .ZN(n15551) );
  OAI211_X1 U16656 ( .C1(n15549), .C2(n15548), .A(n15611), .B(n15547), .ZN(
        n15550) );
  NAND3_X1 U16657 ( .A1(n15552), .A2(n15551), .A3(n15550), .ZN(P2_U3216) );
  AOI22_X1 U16658 ( .A1(n15619), .A2(P2_ADDR_REG_4__SCAN_IN), .B1(n15627), 
        .B2(n15553), .ZN(n15558) );
  OAI211_X1 U16659 ( .C1(n15556), .C2(n15555), .A(n15602), .B(n15554), .ZN(
        n15557) );
  AND2_X1 U16660 ( .A1(n15558), .A2(n15557), .ZN(n15564) );
  NAND2_X1 U16661 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n15563) );
  OAI211_X1 U16662 ( .C1(n15561), .C2(n15560), .A(n15611), .B(n15559), .ZN(
        n15562) );
  NAND3_X1 U16663 ( .A1(n15564), .A2(n15563), .A3(n15562), .ZN(P2_U3218) );
  AOI22_X1 U16664 ( .A1(n15619), .A2(P2_ADDR_REG_5__SCAN_IN), .B1(n15627), 
        .B2(n15565), .ZN(n15570) );
  OAI211_X1 U16665 ( .C1(n15568), .C2(n15567), .A(n15602), .B(n15566), .ZN(
        n15569) );
  AND2_X1 U16666 ( .A1(n15570), .A2(n15569), .ZN(n15576) );
  OAI211_X1 U16667 ( .C1(n15573), .C2(n15572), .A(n15611), .B(n15571), .ZN(
        n15574) );
  NAND3_X1 U16668 ( .A1(n15576), .A2(n15575), .A3(n15574), .ZN(P2_U3219) );
  AOI22_X1 U16669 ( .A1(n15619), .A2(P2_ADDR_REG_6__SCAN_IN), .B1(n15627), 
        .B2(n15577), .ZN(n15582) );
  OAI211_X1 U16670 ( .C1(n15580), .C2(n15579), .A(n15602), .B(n15578), .ZN(
        n15581) );
  AND2_X1 U16671 ( .A1(n15582), .A2(n15581), .ZN(n15588) );
  OAI211_X1 U16672 ( .C1(n15585), .C2(n15584), .A(n15611), .B(n15583), .ZN(
        n15586) );
  NAND3_X1 U16673 ( .A1(n15588), .A2(n15587), .A3(n15586), .ZN(P2_U3220) );
  INV_X1 U16674 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15601) );
  NOR2_X1 U16675 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15589), .ZN(n15594) );
  AOI211_X1 U16676 ( .C1(n15592), .C2(n15591), .A(n15622), .B(n15590), .ZN(
        n15593) );
  AOI211_X1 U16677 ( .C1(n15627), .C2(n15595), .A(n15594), .B(n15593), .ZN(
        n15600) );
  OAI211_X1 U16678 ( .C1(n15598), .C2(n15597), .A(n15611), .B(n15596), .ZN(
        n15599) );
  OAI211_X1 U16679 ( .C1(n15616), .C2(n15601), .A(n15600), .B(n15599), .ZN(
        P2_U3230) );
  INV_X1 U16680 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15767) );
  AND2_X1 U16681 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n15608) );
  OAI211_X1 U16682 ( .C1(n15605), .C2(n15604), .A(n15603), .B(n15602), .ZN(
        n15606) );
  INV_X1 U16683 ( .A(n15606), .ZN(n15607) );
  AOI211_X1 U16684 ( .C1(n15627), .C2(n15609), .A(n15608), .B(n15607), .ZN(
        n15615) );
  OAI211_X1 U16685 ( .C1(n15613), .C2(n15612), .A(n15611), .B(n15610), .ZN(
        n15614) );
  OAI211_X1 U16686 ( .C1(n15616), .C2(n15767), .A(n15615), .B(n15614), .ZN(
        P2_U3227) );
  AOI21_X1 U16687 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n15618), .A(n15617), 
        .ZN(n15631) );
  AOI22_X1 U16688 ( .A1(n15619), .A2(P2_ADDR_REG_12__SCAN_IN), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(P2_U3088), .ZN(n15629) );
  NAND2_X1 U16689 ( .A1(n15621), .A2(n15620), .ZN(n15623) );
  AOI21_X1 U16690 ( .B1(n15624), .B2(n15623), .A(n15622), .ZN(n15625) );
  AOI21_X1 U16691 ( .B1(n15627), .B2(n15626), .A(n15625), .ZN(n15628) );
  OAI211_X1 U16692 ( .C1(n15631), .C2(n15630), .A(n15629), .B(n15628), .ZN(
        P2_U3226) );
  NOR2_X1 U16693 ( .A1(n15632), .A2(n15880), .ZN(n15636) );
  NOR2_X1 U16694 ( .A1(n15633), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n15635) );
  MUX2_X1 U16695 ( .A(n15636), .B(n15635), .S(n15634), .Z(n15637) );
  OR2_X1 U16696 ( .A1(n15638), .A2(n15637), .ZN(n15642) );
  AOI22_X1 U16697 ( .A1(n15639), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n7201), .ZN(n15640) );
  OAI21_X1 U16698 ( .B1(n15642), .B2(n15641), .A(n15640), .ZN(P1_U3243) );
  INV_X1 U16699 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15790) );
  OAI21_X1 U16700 ( .B1(n15644), .B2(n16128), .A(n15643), .ZN(n15653) );
  AOI21_X1 U16701 ( .B1(n15646), .B2(P1_REG2_REG_15__SCAN_IN), .A(n15645), 
        .ZN(n15650) );
  OAI22_X1 U16702 ( .A1(n15650), .A2(n15649), .B1(n15648), .B2(n15647), .ZN(
        n15651) );
  AOI21_X1 U16703 ( .B1(n15653), .B2(n15652), .A(n15651), .ZN(n15655) );
  OAI211_X1 U16704 ( .C1(n15790), .C2(n15656), .A(n15655), .B(n15654), .ZN(
        P1_U3258) );
  NAND2_X1 U16705 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n15657), .ZN(n15663) );
  OAI21_X1 U16706 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n15657), .A(n15663), .ZN(
        n15658) );
  XOR2_X1 U16707 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15658), .Z(SUB_1596_U53) );
  INV_X1 U16708 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n15660) );
  NOR2_X1 U16709 ( .A1(n15659), .A2(n15660), .ZN(n15661) );
  NAND2_X1 U16710 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15658), .ZN(n15830) );
  XNOR2_X1 U16711 ( .A(n15660), .B(n15659), .ZN(n15829) );
  NOR2_X1 U16712 ( .A1(n15830), .A2(n15829), .ZN(n15828) );
  XOR2_X1 U16713 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n15672), .Z(n15666) );
  NAND2_X1 U16714 ( .A1(n15667), .A2(n15666), .ZN(n15668) );
  OAI21_X1 U16715 ( .B1(n15667), .B2(n15666), .A(n15668), .ZN(n15665) );
  XNOR2_X1 U16716 ( .A(n15665), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  NOR2_X1 U16717 ( .A1(n15667), .A2(n15666), .ZN(n15669) );
  NOR2_X1 U16718 ( .A1(n15671), .A2(n15670), .ZN(n15674) );
  NOR2_X1 U16719 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n15672), .ZN(n15673) );
  INV_X1 U16720 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15675) );
  OAI21_X1 U16721 ( .B1(n15676), .B2(n15675), .A(n15685), .ZN(SUB_1596_U60) );
  NOR2_X1 U16722 ( .A1(n15678), .A2(n15677), .ZN(n15681) );
  NOR2_X1 U16723 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n15679), .ZN(n15680) );
  XOR2_X1 U16724 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P3_ADDR_REG_4__SCAN_IN), .Z(
        n15682) );
  XNOR2_X1 U16725 ( .A(n15689), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15688) );
  NAND2_X1 U16726 ( .A1(n15684), .A2(n15683), .ZN(n15686) );
  NOR2_X1 U16727 ( .A1(n15688), .A2(n15687), .ZN(n15690) );
  AOI21_X1 U16728 ( .B1(n15688), .B2(n15687), .A(n15690), .ZN(SUB_1596_U59) );
  AND2_X1 U16729 ( .A1(n15689), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n15691) );
  XNOR2_X1 U16730 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n15694) );
  XOR2_X1 U16731 ( .A(n15694), .B(n15702), .Z(n15696) );
  NOR2_X1 U16732 ( .A1(n15697), .A2(n15696), .ZN(n15698) );
  AOI21_X1 U16733 ( .B1(n15697), .B2(n15696), .A(n15698), .ZN(n15695) );
  XOR2_X1 U16734 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15695), .Z(SUB_1596_U58) );
  NAND2_X1 U16735 ( .A1(n15697), .A2(n15696), .ZN(n15699) );
  XNOR2_X1 U16736 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n15703) );
  AND2_X1 U16737 ( .A1(n15700), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n15701) );
  XNOR2_X1 U16738 ( .A(n15703), .B(n15705), .ZN(n15825) );
  NAND2_X1 U16739 ( .A1(n15826), .A2(n15825), .ZN(n15704) );
  NOR2_X1 U16740 ( .A1(n15826), .A2(n15825), .ZN(n15824) );
  XOR2_X1 U16741 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n15710), .Z(n15712) );
  XNOR2_X1 U16742 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n15712), .ZN(n15708) );
  OAI21_X1 U16743 ( .B1(n15709), .B2(n15708), .A(n15716), .ZN(SUB_1596_U56) );
  INV_X1 U16744 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15722) );
  INV_X1 U16745 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15726) );
  XNOR2_X1 U16746 ( .A(n15726), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n15724) );
  NAND2_X1 U16747 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n15710), .ZN(n15714) );
  INV_X1 U16748 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15711) );
  NAND2_X1 U16749 ( .A1(n15712), .A2(n15711), .ZN(n15713) );
  NAND2_X1 U16750 ( .A1(n15714), .A2(n15713), .ZN(n15723) );
  XOR2_X1 U16751 ( .A(n15724), .B(n15723), .Z(n15719) );
  NAND2_X1 U16752 ( .A1(n15715), .A2(n7711), .ZN(n15717) );
  NAND2_X1 U16753 ( .A1(n15719), .A2(n15718), .ZN(n15721) );
  INV_X1 U16754 ( .A(n15720), .ZN(n15728) );
  NAND2_X1 U16755 ( .A1(n15722), .A2(n15721), .ZN(n15727) );
  OAI222_X1 U16756 ( .A1(n15722), .A2(n15721), .B1(n15722), .B2(n15728), .C1(
        n15720), .C2(n15727), .ZN(SUB_1596_U55) );
  XOR2_X1 U16757 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Z(
        n15735) );
  XNOR2_X1 U16758 ( .A(n15736), .B(n15735), .ZN(n15731) );
  NAND2_X1 U16759 ( .A1(n15731), .A2(n15730), .ZN(n15732) );
  OAI21_X1 U16760 ( .B1(n15731), .B2(n15730), .A(n15732), .ZN(n15729) );
  XNOR2_X1 U16761 ( .A(n15729), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  INV_X1 U16762 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15743) );
  NOR2_X1 U16763 ( .A1(n15731), .A2(n15730), .ZN(n15733) );
  OAI21_X1 U16764 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(n15733), .A(n15732), .ZN(
        n15734) );
  INV_X1 U16765 ( .A(n15734), .ZN(n15739) );
  INV_X1 U16766 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15738) );
  XNOR2_X1 U16767 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n15744) );
  XNOR2_X1 U16768 ( .A(n15745), .B(n15744), .ZN(n15740) );
  OAI222_X1 U16769 ( .A1(n15743), .A2(n15742), .B1(n15743), .B2(n15749), .C1(
        n15741), .C2(n15748), .ZN(SUB_1596_U70) );
  XNOR2_X1 U16770 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n15747) );
  INV_X1 U16771 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15833) );
  NAND2_X1 U16772 ( .A1(n15745), .A2(n15744), .ZN(n15746) );
  XOR2_X1 U16773 ( .A(n15747), .B(n15756), .Z(n15752) );
  AOI21_X1 U16774 ( .B1(n15752), .B2(n15751), .A(n15753), .ZN(n15750) );
  XOR2_X1 U16775 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15750), .Z(SUB_1596_U69)
         );
  NAND2_X1 U16776 ( .A1(n15752), .A2(n15751), .ZN(n15754) );
  XNOR2_X1 U16777 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n11465), .ZN(n15765) );
  INV_X1 U16778 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15854) );
  NOR2_X1 U16779 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n15854), .ZN(n15757) );
  INV_X1 U16780 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15755) );
  XOR2_X1 U16781 ( .A(n15765), .B(n15764), .Z(n15760) );
  INV_X1 U16782 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15758) );
  OAI21_X1 U16783 ( .B1(n15759), .B2(n15758), .A(n15762), .ZN(SUB_1596_U68) );
  NAND2_X1 U16784 ( .A1(n15761), .A2(n15760), .ZN(n15763) );
  XNOR2_X1 U16785 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n15770) );
  XNOR2_X1 U16786 ( .A(n15770), .B(n15769), .ZN(n15773) );
  NAND2_X1 U16787 ( .A1(n15768), .A2(n15767), .ZN(n15775) );
  OAI21_X1 U16788 ( .B1(n15768), .B2(n15767), .A(n15775), .ZN(SUB_1596_U67) );
  INV_X1 U16789 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15772) );
  NAND2_X1 U16790 ( .A1(n15770), .A2(n15769), .ZN(n15771) );
  XNOR2_X1 U16791 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n15779) );
  XNOR2_X1 U16792 ( .A(n15778), .B(n15779), .ZN(n15783) );
  NAND2_X1 U16793 ( .A1(n15774), .A2(n15773), .ZN(n15776) );
  OAI21_X1 U16794 ( .B1(n15783), .B2(n15782), .A(n15784), .ZN(n15777) );
  XNOR2_X1 U16795 ( .A(n15777), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  XNOR2_X1 U16796 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(n15790), .ZN(n15788) );
  INV_X1 U16797 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15781) );
  NAND2_X1 U16798 ( .A1(n15779), .A2(n15778), .ZN(n15780) );
  XOR2_X1 U16799 ( .A(n15788), .B(n15787), .Z(n15792) );
  AOI21_X1 U16800 ( .B1(n15792), .B2(n15791), .A(n15793), .ZN(n15786) );
  XOR2_X1 U16801 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15786), .Z(SUB_1596_U65)
         );
  NOR2_X1 U16802 ( .A1(n15788), .A2(n15787), .ZN(n15789) );
  AOI21_X1 U16803 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n15790), .A(n15789), 
        .ZN(n15799) );
  XNOR2_X1 U16804 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n15799), .ZN(n15800) );
  XNOR2_X1 U16805 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n15800), .ZN(n15795) );
  NAND2_X1 U16806 ( .A1(n15796), .A2(n15795), .ZN(n15797) );
  OAI21_X1 U16807 ( .B1(n15795), .B2(n15796), .A(n15797), .ZN(n15794) );
  XNOR2_X1 U16808 ( .A(n15794), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  NAND2_X1 U16809 ( .A1(n15799), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n15802) );
  NAND2_X1 U16810 ( .A1(n15802), .A2(n15801), .ZN(n15809) );
  XOR2_X1 U16811 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n15809), .Z(n15811) );
  XOR2_X1 U16812 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n15811), .Z(n15806) );
  INV_X1 U16813 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15805) );
  XNOR2_X1 U16814 ( .A(n15806), .B(n15805), .ZN(n15803) );
  NOR2_X1 U16815 ( .A1(n15804), .A2(n15803), .ZN(n15807) );
  AOI21_X1 U16816 ( .B1(n15804), .B2(n15803), .A(n15807), .ZN(SUB_1596_U63) );
  NOR2_X1 U16817 ( .A1(n15806), .A2(n15805), .ZN(n15808) );
  NAND2_X1 U16818 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15809), .ZN(n15813) );
  NAND2_X1 U16819 ( .A1(n15811), .A2(n15810), .ZN(n15812) );
  NAND2_X1 U16820 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15818), .ZN(n15814) );
  OAI21_X1 U16821 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15818), .A(n15814), 
        .ZN(n15815) );
  XNOR2_X1 U16822 ( .A(n15816), .B(n15815), .ZN(n15821) );
  NOR2_X1 U16823 ( .A1(n15816), .A2(n15815), .ZN(n15817) );
  AOI21_X1 U16824 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15818), .A(n15817), 
        .ZN(n15820) );
  XNOR2_X1 U16825 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n15819) );
  XNOR2_X1 U16826 ( .A(n15820), .B(n15819), .ZN(n15823) );
  AOI21_X1 U16827 ( .B1(n15826), .B2(n15825), .A(n15824), .ZN(n15827) );
  XOR2_X1 U16828 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n15827), .Z(SUB_1596_U57) );
  AOI21_X1 U16829 ( .B1(n15830), .B2(n15829), .A(n15828), .ZN(SUB_1596_U5) );
  AOI21_X1 U16830 ( .B1(n7375), .B2(n15832), .A(n15831), .ZN(n15849) );
  OAI22_X1 U16831 ( .A1(n15856), .A2(n15834), .B1(n15833), .B2(n15853), .ZN(
        n15846) );
  INV_X1 U16832 ( .A(n15835), .ZN(n15836) );
  AOI21_X1 U16833 ( .B1(n15838), .B2(n15837), .A(n15836), .ZN(n15844) );
  AOI21_X1 U16834 ( .B1(n15841), .B2(n15840), .A(n15839), .ZN(n15842) );
  OAI22_X1 U16835 ( .A1(n15844), .A2(n15843), .B1(n15842), .B2(n15866), .ZN(
        n15845) );
  NOR3_X1 U16836 ( .A1(n15847), .A2(n15846), .A3(n15845), .ZN(n15848) );
  OAI21_X1 U16837 ( .B1(n15849), .B2(n15872), .A(n15848), .ZN(P3_U3192) );
  AOI21_X1 U16838 ( .B1(n15852), .B2(n15851), .A(n15850), .ZN(n15873) );
  OAI22_X1 U16839 ( .A1(n15856), .A2(n15855), .B1(n15854), .B2(n15853), .ZN(
        n15869) );
  AOI21_X1 U16840 ( .B1(n15859), .B2(n15858), .A(n15857), .ZN(n15867) );
  OAI21_X1 U16841 ( .B1(n15862), .B2(n15861), .A(n15860), .ZN(n15864) );
  NAND2_X1 U16842 ( .A1(n15864), .A2(n15863), .ZN(n15865) );
  OAI21_X1 U16843 ( .B1(n15867), .B2(n15866), .A(n15865), .ZN(n15868) );
  NOR3_X1 U16844 ( .A1(n15870), .A2(n15869), .A3(n15868), .ZN(n15871) );
  OAI21_X1 U16845 ( .B1(n15873), .B2(n15872), .A(n15871), .ZN(P3_U3193) );
  OAI221_X1 U16846 ( .B1(P1_RD_REG_SCAN_IN), .B2(P2_RD_REG_SCAN_IN), .C1(n7989), .C2(n7987), .A(n15874), .ZN(U29) );
  NOR2_X1 U16847 ( .A1(n15875), .A2(n16021), .ZN(n15876) );
  AOI211_X1 U16848 ( .C1(n15879), .C2(n15878), .A(n15877), .B(n15876), .ZN(
        n15882) );
  AOI22_X1 U16849 ( .A1(n16143), .A2(n15882), .B1(n15880), .B2(n16141), .ZN(
        P1_U3528) );
  INV_X1 U16850 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15881) );
  AOI22_X1 U16851 ( .A1(n16147), .A2(n15882), .B1(n15881), .B2(n16144), .ZN(
        P1_U3459) );
  AOI21_X1 U16852 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n15884), .A(n15883), .ZN(
        n15890) );
  NAND2_X1 U16853 ( .A1(n16006), .A2(n15885), .ZN(n15889) );
  AOI22_X1 U16854 ( .A1(n15887), .A2(n15886), .B1(P2_REG2_REG_0__SCAN_IN), 
        .B2(n15891), .ZN(n15888) );
  OAI221_X1 U16855 ( .B1(n15891), .B2(n15890), .C1(n15891), .C2(n15889), .A(
        n15888), .ZN(P2_U3265) );
  INV_X1 U16856 ( .A(n15892), .ZN(n15894) );
  AOI211_X1 U16857 ( .C1(n16059), .C2(n15895), .A(n15894), .B(n15893), .ZN(
        n15898) );
  AOI22_X1 U16858 ( .A1(n16061), .A2(n15898), .B1(n15896), .B2(n12991), .ZN(
        P3_U3461) );
  INV_X1 U16859 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15897) );
  AOI22_X1 U16860 ( .A1(n16065), .A2(n15898), .B1(n15897), .B2(n16062), .ZN(
        P3_U3396) );
  NOR2_X1 U16861 ( .A1(n15899), .A2(n16054), .ZN(n15901) );
  AOI211_X1 U16862 ( .C1(n16059), .C2(n15902), .A(n15901), .B(n15900), .ZN(
        n15904) );
  AOI22_X1 U16863 ( .A1(n16061), .A2(n15904), .B1(n10860), .B2(n12991), .ZN(
        P3_U3462) );
  INV_X1 U16864 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15903) );
  AOI22_X1 U16865 ( .A1(n16065), .A2(n15904), .B1(n15903), .B2(n16062), .ZN(
        P3_U3399) );
  AOI21_X1 U16866 ( .B1(n16026), .B2(n15911), .A(n15905), .ZN(n15913) );
  AOI22_X1 U16867 ( .A1(n16001), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n15990), 
        .B2(n9912), .ZN(n15908) );
  NAND2_X1 U16868 ( .A1(n15991), .A2(n15906), .ZN(n15907) );
  OAI211_X1 U16869 ( .C1(n15909), .C2(n15993), .A(n15908), .B(n15907), .ZN(
        n15910) );
  AOI21_X1 U16870 ( .B1(n15911), .B2(n15996), .A(n15910), .ZN(n15912) );
  OAI21_X1 U16871 ( .B1(n16001), .B2(n15913), .A(n15912), .ZN(P1_U3290) );
  NOR2_X1 U16872 ( .A1(n15914), .A2(n16054), .ZN(n15916) );
  AOI211_X1 U16873 ( .C1(n16059), .C2(n15917), .A(n15916), .B(n15915), .ZN(
        n15919) );
  AOI22_X1 U16874 ( .A1(n16061), .A2(n15919), .B1(n10881), .B2(n12991), .ZN(
        P3_U3463) );
  INV_X1 U16875 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15918) );
  AOI22_X1 U16876 ( .A1(n16065), .A2(n15919), .B1(n15918), .B2(n16062), .ZN(
        P3_U3402) );
  INV_X1 U16877 ( .A(n15920), .ZN(n15921) );
  NAND3_X1 U16878 ( .A1(n15923), .A2(n15922), .A3(n15921), .ZN(n15926) );
  INV_X1 U16879 ( .A(n15924), .ZN(n15925) );
  AOI211_X1 U16880 ( .C1(n16139), .C2(n15927), .A(n15926), .B(n15925), .ZN(
        n15930) );
  INV_X1 U16881 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15928) );
  AOI22_X1 U16882 ( .A1(n16143), .A2(n15930), .B1(n15928), .B2(n16141), .ZN(
        P1_U3532) );
  INV_X1 U16883 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15929) );
  AOI22_X1 U16884 ( .A1(n16147), .A2(n15930), .B1(n15929), .B2(n16144), .ZN(
        P1_U3471) );
  INV_X1 U16885 ( .A(n16021), .ZN(n16066) );
  INV_X1 U16886 ( .A(n15931), .ZN(n15932) );
  NAND2_X1 U16887 ( .A1(n15933), .A2(n15932), .ZN(n15935) );
  AOI211_X1 U16888 ( .C1(n16066), .C2(n15936), .A(n15935), .B(n15934), .ZN(
        n15938) );
  AOI22_X1 U16889 ( .A1(n16143), .A2(n15938), .B1(n10340), .B2(n16141), .ZN(
        P1_U3533) );
  INV_X1 U16890 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15937) );
  AOI22_X1 U16891 ( .A1(n16147), .A2(n15938), .B1(n15937), .B2(n16144), .ZN(
        P1_U3474) );
  AOI22_X1 U16892 ( .A1(n15941), .A2(n16059), .B1(n15940), .B2(n15939), .ZN(
        n15942) );
  AND2_X1 U16893 ( .A1(n15943), .A2(n15942), .ZN(n15946) );
  AOI22_X1 U16894 ( .A1(n16061), .A2(n15946), .B1(n15944), .B2(n12991), .ZN(
        P3_U3465) );
  INV_X1 U16895 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15945) );
  AOI22_X1 U16896 ( .A1(n16065), .A2(n15946), .B1(n15945), .B2(n16062), .ZN(
        P3_U3408) );
  OAI21_X1 U16897 ( .B1(n15948), .B2(n16123), .A(n15947), .ZN(n15950) );
  AOI211_X1 U16898 ( .C1(n16066), .C2(n15951), .A(n15950), .B(n15949), .ZN(
        n15954) );
  INV_X1 U16899 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n15952) );
  AOI22_X1 U16900 ( .A1(n16143), .A2(n15954), .B1(n15952), .B2(n16141), .ZN(
        P1_U3534) );
  INV_X1 U16901 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15953) );
  AOI22_X1 U16902 ( .A1(n16147), .A2(n15954), .B1(n15953), .B2(n16144), .ZN(
        P1_U3477) );
  INV_X1 U16903 ( .A(n15958), .ZN(n15961) );
  OAI211_X1 U16904 ( .C1(n15957), .C2(n16123), .A(n15956), .B(n15955), .ZN(
        n15960) );
  NOR2_X1 U16905 ( .A1(n15958), .A2(n16021), .ZN(n15959) );
  AOI211_X1 U16906 ( .C1(n15961), .C2(n16026), .A(n15960), .B(n15959), .ZN(
        n15963) );
  AOI22_X1 U16907 ( .A1(n16143), .A2(n15963), .B1(n10403), .B2(n16141), .ZN(
        P1_U3535) );
  INV_X1 U16908 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15962) );
  AOI22_X1 U16909 ( .A1(n16147), .A2(n15963), .B1(n15962), .B2(n16144), .ZN(
        P1_U3480) );
  OAI22_X1 U16910 ( .A1(n15965), .A2(n16011), .B1(n15964), .B2(n16054), .ZN(
        n15967) );
  NOR2_X1 U16911 ( .A1(n15967), .A2(n15966), .ZN(n15970) );
  INV_X1 U16912 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15968) );
  AOI22_X1 U16913 ( .A1(n16061), .A2(n15970), .B1(n15968), .B2(n12991), .ZN(
        P3_U3467) );
  INV_X1 U16914 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15969) );
  AOI22_X1 U16915 ( .A1(n16065), .A2(n15970), .B1(n15969), .B2(n16062), .ZN(
        P3_U3414) );
  NAND2_X1 U16916 ( .A1(n15971), .A2(n11930), .ZN(n15972) );
  INV_X1 U16917 ( .A(n15992), .ZN(n15978) );
  AOI21_X1 U16918 ( .B1(n15975), .B2(n15992), .A(n15974), .ZN(n15977) );
  NAND2_X1 U16919 ( .A1(n15977), .A2(n15976), .ZN(n15994) );
  OAI21_X1 U16920 ( .B1(n15978), .B2(n16123), .A(n15994), .ZN(n15987) );
  INV_X1 U16921 ( .A(n15979), .ZN(n15985) );
  INV_X1 U16922 ( .A(n15980), .ZN(n15981) );
  AOI211_X1 U16923 ( .C1(n15983), .C2(n15982), .A(n16136), .B(n15981), .ZN(
        n15984) );
  AOI211_X1 U16924 ( .C1(n16026), .C2(n15997), .A(n15985), .B(n15984), .ZN(
        n16000) );
  INV_X1 U16925 ( .A(n16000), .ZN(n15986) );
  AOI211_X1 U16926 ( .C1(n16066), .C2(n15997), .A(n15987), .B(n15986), .ZN(
        n15989) );
  AOI22_X1 U16927 ( .A1(n16143), .A2(n15989), .B1(n10615), .B2(n16141), .ZN(
        P1_U3536) );
  INV_X1 U16928 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15988) );
  AOI22_X1 U16929 ( .A1(n16147), .A2(n15989), .B1(n15988), .B2(n16144), .ZN(
        P1_U3483) );
  AOI222_X1 U16930 ( .A1(n15992), .A2(n15991), .B1(n7252), .B2(n15990), .C1(
        P1_REG2_REG_8__SCAN_IN), .C2(n16001), .ZN(n15999) );
  NOR2_X1 U16931 ( .A1(n15994), .A2(n15993), .ZN(n15995) );
  AOI21_X1 U16932 ( .B1(n15997), .B2(n15996), .A(n15995), .ZN(n15998) );
  OAI211_X1 U16933 ( .C1(n16001), .C2(n16000), .A(n15999), .B(n15998), .ZN(
        P1_U3285) );
  AOI21_X1 U16934 ( .B1(n16112), .B2(n16003), .A(n16002), .ZN(n16004) );
  OAI211_X1 U16935 ( .C1(n16007), .C2(n16006), .A(n16005), .B(n16004), .ZN(
        n16008) );
  INV_X1 U16936 ( .A(n16008), .ZN(n16009) );
  AOI22_X1 U16937 ( .A1(n16156), .A2(n16009), .B1(n10514), .B2(n16155), .ZN(
        P2_U3507) );
  AOI22_X1 U16938 ( .A1(n16117), .A2(n16009), .B1(n9067), .B2(n16157), .ZN(
        P2_U3454) );
  OAI22_X1 U16939 ( .A1(n16012), .A2(n16011), .B1(n16010), .B2(n16054), .ZN(
        n16013) );
  NOR2_X1 U16940 ( .A1(n16014), .A2(n16013), .ZN(n16017) );
  AOI22_X1 U16941 ( .A1(n16061), .A2(n16017), .B1(n16015), .B2(n12991), .ZN(
        P3_U3468) );
  INV_X1 U16942 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n16016) );
  AOI22_X1 U16943 ( .A1(n16065), .A2(n16017), .B1(n16016), .B2(n16062), .ZN(
        P3_U3417) );
  INV_X1 U16944 ( .A(n16022), .ZN(n16025) );
  AOI21_X1 U16945 ( .B1(n16134), .B2(n16019), .A(n16018), .ZN(n16020) );
  OAI21_X1 U16946 ( .B1(n16022), .B2(n16021), .A(n16020), .ZN(n16023) );
  AOI211_X1 U16947 ( .C1(n16026), .C2(n16025), .A(n16024), .B(n16023), .ZN(
        n16028) );
  AOI22_X1 U16948 ( .A1(n16143), .A2(n16028), .B1(n11160), .B2(n16141), .ZN(
        P1_U3537) );
  INV_X1 U16949 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n16027) );
  AOI22_X1 U16950 ( .A1(n16147), .A2(n16028), .B1(n16027), .B2(n16144), .ZN(
        P1_U3486) );
  AOI22_X1 U16951 ( .A1(n16031), .A2(n16134), .B1(n16030), .B2(n16029), .ZN(
        n16032) );
  OAI211_X1 U16952 ( .C1(n16034), .C2(n16136), .A(n16033), .B(n16032), .ZN(
        n16035) );
  AOI21_X1 U16953 ( .B1(n16036), .B2(n16139), .A(n16035), .ZN(n16038) );
  AOI22_X1 U16954 ( .A1(n16143), .A2(n16038), .B1(n11157), .B2(n16141), .ZN(
        P1_U3538) );
  INV_X1 U16955 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n16037) );
  AOI22_X1 U16956 ( .A1(n16147), .A2(n16038), .B1(n16037), .B2(n16144), .ZN(
        P1_U3489) );
  OAI21_X1 U16957 ( .B1(n7708), .B2(n16149), .A(n16039), .ZN(n16040) );
  AOI21_X1 U16958 ( .B1(n16042), .B2(n16041), .A(n16040), .ZN(n16043) );
  AND2_X1 U16959 ( .A1(n16044), .A2(n16043), .ZN(n16045) );
  AOI22_X1 U16960 ( .A1(n16156), .A2(n16045), .B1(n10579), .B2(n16155), .ZN(
        P2_U3509) );
  AOI22_X1 U16961 ( .A1(n16160), .A2(n16045), .B1(n9119), .B2(n16157), .ZN(
        P2_U3460) );
  NAND3_X1 U16962 ( .A1(n12302), .A2(n16046), .A3(n16139), .ZN(n16048) );
  OAI211_X1 U16963 ( .C1(n16049), .C2(n16123), .A(n16048), .B(n16047), .ZN(
        n16051) );
  NOR2_X1 U16964 ( .A1(n16051), .A2(n16050), .ZN(n16053) );
  AOI22_X1 U16965 ( .A1(n16143), .A2(n16053), .B1(n11237), .B2(n16141), .ZN(
        P1_U3539) );
  INV_X1 U16966 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n16052) );
  AOI22_X1 U16967 ( .A1(n16147), .A2(n16053), .B1(n16052), .B2(n16144), .ZN(
        P1_U3492) );
  NOR2_X1 U16968 ( .A1(n16055), .A2(n16054), .ZN(n16057) );
  AOI211_X1 U16969 ( .C1(n16059), .C2(n16058), .A(n16057), .B(n16056), .ZN(
        n16064) );
  INV_X1 U16970 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n16060) );
  AOI22_X1 U16971 ( .A1(n16061), .A2(n16064), .B1(n16060), .B2(n12991), .ZN(
        P3_U3471) );
  INV_X1 U16972 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n16063) );
  AOI22_X1 U16973 ( .A1(n16065), .A2(n16064), .B1(n16063), .B2(n16062), .ZN(
        P3_U3426) );
  NAND2_X1 U16974 ( .A1(n16067), .A2(n16066), .ZN(n16069) );
  OAI211_X1 U16975 ( .C1(n16070), .C2(n16123), .A(n16069), .B(n16068), .ZN(
        n16071) );
  NOR2_X1 U16976 ( .A1(n16072), .A2(n16071), .ZN(n16075) );
  AOI22_X1 U16977 ( .A1(n16143), .A2(n16075), .B1(n16073), .B2(n16141), .ZN(
        P1_U3540) );
  INV_X1 U16978 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n16074) );
  AOI22_X1 U16979 ( .A1(n16147), .A2(n16075), .B1(n16074), .B2(n16144), .ZN(
        P1_U3495) );
  OAI211_X1 U16980 ( .C1(n16078), .C2(n16123), .A(n16077), .B(n16076), .ZN(
        n16079) );
  AOI21_X1 U16981 ( .B1(n16080), .B2(n16139), .A(n16079), .ZN(n16082) );
  AOI22_X1 U16982 ( .A1(n16143), .A2(n16082), .B1(n11838), .B2(n16141), .ZN(
        P1_U3541) );
  INV_X1 U16983 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n16081) );
  AOI22_X1 U16984 ( .A1(n16147), .A2(n16082), .B1(n16081), .B2(n16144), .ZN(
        P1_U3498) );
  OAI21_X1 U16985 ( .B1(n16085), .B2(n16084), .A(n16083), .ZN(n16094) );
  AOI22_X1 U16986 ( .A1(n16089), .A2(n16088), .B1(n16087), .B2(n16086), .ZN(
        n16090) );
  OAI21_X1 U16987 ( .B1(n7737), .B2(n16091), .A(n16090), .ZN(n16092) );
  AOI21_X1 U16988 ( .B1(n16094), .B2(n16093), .A(n16092), .ZN(n16096) );
  OAI211_X1 U16989 ( .C1(n16098), .C2(n16097), .A(n16096), .B(n16095), .ZN(
        P1_U3215) );
  OAI211_X1 U16990 ( .C1(n7737), .C2(n16123), .A(n16100), .B(n16099), .ZN(
        n16103) );
  AND3_X1 U16991 ( .A1(n7359), .A2(n16139), .A3(n16101), .ZN(n16102) );
  AOI211_X1 U16992 ( .C1(n16104), .C2(n16119), .A(n16103), .B(n16102), .ZN(
        n16107) );
  AOI22_X1 U16993 ( .A1(n16143), .A2(n16107), .B1(n16105), .B2(n16141), .ZN(
        P1_U3542) );
  INV_X1 U16994 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n16106) );
  AOI22_X1 U16995 ( .A1(n16147), .A2(n16107), .B1(n16106), .B2(n16144), .ZN(
        P1_U3501) );
  NAND3_X1 U16996 ( .A1(n16109), .A2(n16108), .A3(n16153), .ZN(n16115) );
  AOI21_X1 U16997 ( .B1(n16112), .B2(n16111), .A(n16110), .ZN(n16113) );
  AOI22_X1 U16998 ( .A1(n16156), .A2(n16116), .B1(n11086), .B2(n16155), .ZN(
        P2_U3513) );
  AOI22_X1 U16999 ( .A1(n16117), .A2(n16116), .B1(n9232), .B2(n16157), .ZN(
        P2_U3472) );
  AND3_X1 U17000 ( .A1(n16120), .A2(n16119), .A3(n16118), .ZN(n16126) );
  OAI211_X1 U17001 ( .C1(n16124), .C2(n16123), .A(n16122), .B(n16121), .ZN(
        n16125) );
  AOI211_X1 U17002 ( .C1(n16127), .C2(n16139), .A(n16126), .B(n16125), .ZN(
        n16130) );
  AOI22_X1 U17003 ( .A1(n16143), .A2(n16130), .B1(n16128), .B2(n16141), .ZN(
        P1_U3543) );
  INV_X1 U17004 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n16129) );
  AOI22_X1 U17005 ( .A1(n16147), .A2(n16130), .B1(n16129), .B2(n16144), .ZN(
        P1_U3504) );
  AOI211_X1 U17006 ( .C1(n16134), .C2(n16133), .A(n16132), .B(n16131), .ZN(
        n16135) );
  OAI21_X1 U17007 ( .B1(n16137), .B2(n16136), .A(n16135), .ZN(n16138) );
  AOI21_X1 U17008 ( .B1(n16140), .B2(n16139), .A(n16138), .ZN(n16146) );
  AOI22_X1 U17009 ( .A1(n16143), .A2(n16146), .B1(n16142), .B2(n16141), .ZN(
        P1_U3544) );
  INV_X1 U17010 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n16145) );
  AOI22_X1 U17011 ( .A1(n16147), .A2(n16146), .B1(n16145), .B2(n16144), .ZN(
        P1_U3507) );
  OAI21_X1 U17012 ( .B1(n16150), .B2(n16149), .A(n16148), .ZN(n16151) );
  AOI211_X1 U17013 ( .C1(n16154), .C2(n16153), .A(n16152), .B(n16151), .ZN(
        n16159) );
  AOI22_X1 U17014 ( .A1(n16156), .A2(n16159), .B1(n12335), .B2(n16155), .ZN(
        P2_U3516) );
  INV_X1 U17015 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n16158) );
  AOI22_X1 U17016 ( .A1(n16160), .A2(n16159), .B1(n16158), .B2(n16157), .ZN(
        P2_U3481) );
  AOI21_X1 U17017 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16161) );
  OAI21_X1 U17018 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16161), 
        .ZN(U28) );
  NAND2_X1 U7369 ( .A1(n8267), .A2(n8268), .ZN(n14153) );
  CLKBUF_X2 U7307 ( .A(n12702), .Z(n12743) );
  CLKBUF_X1 U7314 ( .A(n12885), .Z(n7227) );
  CLKBUF_X1 U7331 ( .A(n9871), .Z(n9894) );
  CLKBUF_X1 U7367 ( .A(n8182), .Z(n7508) );
  CLKBUF_X2 U7388 ( .A(n9887), .Z(n14953) );
  CLKBUF_X1 U7498 ( .A(n7231), .Z(n8823) );
  CLKBUF_X1 U7606 ( .A(n9606), .Z(n7207) );
  AND2_X1 U7698 ( .A1(n15495), .A2(n15494), .ZN(n16168) );
endmodule

